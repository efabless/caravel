magic
tech sky130A
magscale 1 2
timestamp 1665749829
<< viali >>
rect 581 10761 615 10795
rect 5273 10761 5307 10795
rect 8861 10761 8895 10795
rect 11897 10761 11931 10795
rect 12817 10761 12851 10795
rect 17969 10761 18003 10795
rect 18245 10761 18279 10795
rect 2513 10693 2547 10727
rect 6561 10693 6595 10727
rect 9689 10693 9723 10727
rect 11805 10693 11839 10727
rect 14381 10693 14415 10727
rect 17233 10693 17267 10727
rect 17693 10693 17727 10727
rect 1133 10625 1167 10659
rect 1961 10625 1995 10659
rect 2053 10625 2087 10659
rect 3065 10625 3099 10659
rect 3249 10625 3283 10659
rect 4813 10625 4847 10659
rect 5917 10625 5951 10659
rect 6469 10625 6503 10659
rect 7113 10625 7147 10659
rect 8033 10625 8067 10659
rect 9965 10625 9999 10659
rect 10609 10625 10643 10659
rect 11161 10625 11195 10659
rect 12541 10625 12575 10659
rect 12725 10625 12759 10659
rect 13829 10625 13863 10659
rect 14933 10625 14967 10659
rect 16773 10625 16807 10659
rect 765 10557 799 10591
rect 857 10557 891 10591
rect 1685 10557 1719 10591
rect 2881 10557 2915 10591
rect 3341 10557 3375 10591
rect 4537 10557 4571 10591
rect 4629 10557 4663 10591
rect 5733 10557 5767 10591
rect 6929 10557 6963 10591
rect 7849 10557 7883 10591
rect 8769 10557 8803 10591
rect 9045 10557 9079 10591
rect 9229 10557 9263 10591
rect 11897 10557 11931 10591
rect 12081 10557 12115 10591
rect 12265 10557 12299 10591
rect 12633 10557 12667 10591
rect 13001 10557 13035 10591
rect 13553 10557 13587 10591
rect 14657 10557 14691 10591
rect 16681 10557 16715 10591
rect 17877 10557 17911 10591
rect 18061 10557 18095 10591
rect 18429 10557 18463 10591
rect 1593 10489 1627 10523
rect 10517 10489 10551 10523
rect 11437 10489 11471 10523
rect 12449 10489 12483 10523
rect 13921 10489 13955 10523
rect 15117 10489 15151 10523
rect 16037 10489 16071 10523
rect 16405 10489 16439 10523
rect 17601 10489 17635 10523
rect 2145 10421 2179 10455
rect 2697 10421 2731 10455
rect 3709 10421 3743 10455
rect 4077 10421 4111 10455
rect 4169 10421 4203 10455
rect 5365 10421 5399 10455
rect 5825 10421 5859 10455
rect 7021 10421 7055 10455
rect 7481 10421 7515 10455
rect 7941 10421 7975 10455
rect 8401 10421 8435 10455
rect 9137 10421 9171 10455
rect 9505 10421 9539 10455
rect 10057 10421 10091 10455
rect 10425 10421 10459 10455
rect 11345 10421 11379 10455
rect 13001 10421 13035 10455
rect 14013 10421 14047 10455
rect 15209 10421 15243 10455
rect 15577 10421 15611 10455
rect 15945 10421 15979 10455
rect 16129 10421 16163 10455
rect 16221 10421 16255 10455
rect 16497 10421 16531 10455
rect 17141 10421 17175 10455
rect 6009 10217 6043 10251
rect 17417 10217 17451 10251
rect 17509 10217 17543 10251
rect 17877 10217 17911 10251
rect 1317 10149 1351 10183
rect 5181 10149 5215 10183
rect 5457 10149 5491 10183
rect 12035 10149 12069 10183
rect 16405 10149 16439 10183
rect 16589 10149 16623 10183
rect 18153 10149 18187 10183
rect 673 10081 707 10115
rect 2145 10081 2179 10115
rect 4905 10081 4939 10115
rect 7297 10081 7331 10115
rect 9873 10081 9907 10115
rect 9965 10081 9999 10115
rect 10241 10081 10275 10115
rect 16681 10081 16715 10115
rect 16865 10081 16899 10115
rect 18061 10081 18095 10115
rect 18245 10081 18279 10115
rect 18337 10081 18371 10115
rect 949 10013 983 10047
rect 1869 10013 1903 10047
rect 2053 10013 2087 10047
rect 4169 10013 4203 10047
rect 4537 10013 4571 10047
rect 4629 10013 4663 10047
rect 7481 10013 7515 10047
rect 7849 10013 7883 10047
rect 10149 10013 10183 10047
rect 10609 10013 10643 10047
rect 12633 10013 12667 10047
rect 13001 10013 13035 10047
rect 17693 10013 17727 10047
rect 581 9945 615 9979
rect 2513 9945 2547 9979
rect 4721 9945 4755 9979
rect 9275 9945 9309 9979
rect 12449 9945 12483 9979
rect 1593 9877 1627 9911
rect 2743 9877 2777 9911
rect 4813 9877 4847 9911
rect 9505 9877 9539 9911
rect 9597 9877 9631 9911
rect 10057 9877 10091 9911
rect 12265 9877 12299 9911
rect 14427 9877 14461 9911
rect 15117 9877 15151 9911
rect 16773 9877 16807 9911
rect 17049 9877 17083 9911
rect 3985 9673 4019 9707
rect 4353 9673 4387 9707
rect 5837 9673 5871 9707
rect 6285 9673 6319 9707
rect 15945 9673 15979 9707
rect 18429 9673 18463 9707
rect 3617 9605 3651 9639
rect 8447 9605 8481 9639
rect 8677 9605 8711 9639
rect 10609 9605 10643 9639
rect 10793 9605 10827 9639
rect 13139 9605 13173 9639
rect 15393 9605 15427 9639
rect 18337 9605 18371 9639
rect 765 9537 799 9571
rect 3893 9537 3927 9571
rect 6101 9537 6135 9571
rect 8861 9537 8895 9571
rect 9137 9537 9171 9571
rect 11713 9537 11747 9571
rect 16221 9537 16255 9571
rect 16589 9537 16623 9571
rect 18015 9537 18049 9571
rect 18245 9537 18279 9571
rect 489 9469 523 9503
rect 581 9469 615 9503
rect 1041 9469 1075 9503
rect 1133 9463 1167 9497
rect 1261 9469 1295 9503
rect 1501 9469 1535 9503
rect 3617 9469 3651 9503
rect 4077 9469 4111 9503
rect 4169 9469 4203 9503
rect 6653 9469 6687 9503
rect 7021 9469 7055 9503
rect 10885 9469 10919 9503
rect 11345 9469 11379 9503
rect 13461 9469 13495 9503
rect 15485 9469 15519 9503
rect 16129 9469 16163 9503
rect 18521 9469 18555 9503
rect 765 9401 799 9435
rect 1777 9401 1811 9435
rect 857 9333 891 9367
rect 3249 9333 3283 9367
rect 6561 9333 6595 9367
rect 11161 9333 11195 9367
rect 14749 9333 14783 9367
rect 15669 9333 15703 9367
rect 1777 9129 1811 9163
rect 5089 9129 5123 9163
rect 11805 9129 11839 9163
rect 13553 9129 13587 9163
rect 1041 9061 1075 9095
rect 2789 9061 2823 9095
rect 7481 9061 7515 9095
rect 9689 9061 9723 9095
rect 12265 9061 12299 9095
rect 637 8993 671 9027
rect 765 8993 799 9027
rect 857 8993 891 9027
rect 1225 8993 1259 9027
rect 2145 8993 2179 9027
rect 2237 8993 2271 9027
rect 4445 8993 4479 9027
rect 4721 8993 4755 9027
rect 4905 8993 4939 9027
rect 7021 8993 7055 9027
rect 7297 8993 7331 9027
rect 7849 8993 7883 9027
rect 9873 8993 9907 9027
rect 12081 8993 12115 9027
rect 14473 8993 14507 9027
rect 17049 8993 17083 9027
rect 2329 8925 2363 8959
rect 7941 8925 7975 8959
rect 10241 8925 10275 8959
rect 11667 8925 11701 8959
rect 11805 8925 11839 8959
rect 14841 8925 14875 8959
rect 15209 8925 15243 8959
rect 17509 8925 17543 8959
rect 1593 8857 1627 8891
rect 4813 8857 4847 8891
rect 14197 8857 14231 8891
rect 16589 8857 16623 8891
rect 4537 8789 4571 8823
rect 5733 8789 5767 8823
rect 11989 8789 12023 8823
rect 14749 8789 14783 8823
rect 16773 8789 16807 8823
rect 3433 8585 3467 8619
rect 3709 8585 3743 8619
rect 3985 8585 4019 8619
rect 4261 8585 4295 8619
rect 6561 8585 6595 8619
rect 9965 8585 9999 8619
rect 10701 8585 10735 8619
rect 14749 8585 14783 8619
rect 15393 8585 15427 8619
rect 18337 8585 18371 8619
rect 1317 8517 1351 8551
rect 10517 8517 10551 8551
rect 17877 8517 17911 8551
rect 1041 8449 1075 8483
rect 8493 8449 8527 8483
rect 11069 8449 11103 8483
rect 17785 8449 17819 8483
rect 673 8381 707 8415
rect 949 8381 983 8415
rect 1501 8381 1535 8415
rect 3341 8381 3375 8415
rect 3525 8381 3559 8415
rect 3893 8381 3927 8415
rect 4353 8381 4387 8415
rect 6561 8381 6595 8415
rect 6745 8381 6779 8415
rect 10701 8381 10735 8415
rect 10885 8381 10919 8415
rect 11437 8381 11471 8415
rect 13001 8381 13035 8415
rect 13185 8381 13219 8415
rect 13461 8381 13495 8415
rect 15301 8381 15335 8415
rect 15485 8381 15519 8415
rect 15669 8381 15703 8415
rect 18061 8381 18095 8415
rect 1777 8313 1811 8347
rect 6101 8313 6135 8347
rect 8677 8313 8711 8347
rect 12863 8313 12897 8347
rect 15853 8313 15887 8347
rect 17693 8313 17727 8347
rect 18429 8313 18463 8347
rect 581 8245 615 8279
rect 3249 8245 3283 8279
rect 13093 8245 13127 8279
rect 17141 8245 17175 8279
rect 17969 8245 18003 8279
rect 3065 8041 3099 8075
rect 4905 8041 4939 8075
rect 7205 8041 7239 8075
rect 8309 8041 8343 8075
rect 18337 8041 18371 8075
rect 673 7973 707 8007
rect 857 7973 891 8007
rect 2145 7973 2179 8007
rect 3770 7973 3804 8007
rect 10149 7973 10183 8007
rect 11989 7973 12023 8007
rect 14105 7973 14139 8007
rect 14473 7973 14507 8007
rect 18061 7973 18095 8007
rect 489 7905 523 7939
rect 1317 7905 1351 7939
rect 5181 7905 5215 7939
rect 5457 7905 5491 7939
rect 6101 7905 6135 7939
rect 6285 7905 6319 7939
rect 6837 7905 6871 7939
rect 7021 7905 7055 7939
rect 7573 7905 7607 7939
rect 7757 7905 7791 7939
rect 9597 7905 9631 7939
rect 11805 7905 11839 7939
rect 12081 7905 12115 7939
rect 12265 7905 12299 7939
rect 14289 7905 14323 7939
rect 14932 7905 14966 7939
rect 15025 7905 15059 7939
rect 16865 7905 16899 7939
rect 17049 7905 17083 7939
rect 17233 7905 17267 7939
rect 18245 7905 18279 7939
rect 18429 7905 18463 7939
rect 1041 7837 1075 7871
rect 1225 7837 1259 7871
rect 2237 7837 2271 7871
rect 2421 7837 2455 7871
rect 3157 7837 3191 7871
rect 3341 7837 3375 7871
rect 3525 7837 3559 7871
rect 5089 7837 5123 7871
rect 9873 7837 9907 7871
rect 16589 7837 16623 7871
rect 17509 7837 17543 7871
rect 1777 7769 1811 7803
rect 2697 7769 2731 7803
rect 11805 7769 11839 7803
rect 14657 7769 14691 7803
rect 1685 7701 1719 7735
rect 7665 7701 7699 7735
rect 11621 7701 11655 7735
rect 13737 7701 13771 7735
rect 15117 7701 15151 7735
rect 673 7497 707 7531
rect 8309 7497 8343 7531
rect 11345 7497 11379 7531
rect 13093 7497 13127 7531
rect 581 7429 615 7463
rect 3433 7429 3467 7463
rect 14749 7429 14783 7463
rect 18337 7429 18371 7463
rect 765 7361 799 7395
rect 1317 7361 1351 7395
rect 4169 7361 4203 7395
rect 4813 7361 4847 7395
rect 6285 7361 6319 7395
rect 8217 7361 8251 7395
rect 8401 7361 8435 7395
rect 9413 7361 9447 7395
rect 10333 7361 10367 7395
rect 489 7293 523 7327
rect 1041 7293 1075 7327
rect 1225 7293 1259 7327
rect 1501 7293 1535 7327
rect 3525 7293 3559 7327
rect 3709 7293 3743 7327
rect 4077 7293 4111 7327
rect 4353 7293 4387 7327
rect 4629 7293 4663 7327
rect 4997 7293 5031 7327
rect 5273 7293 5307 7327
rect 5549 7293 5583 7327
rect 6101 7293 6135 7327
rect 6653 7293 6687 7327
rect 8079 7293 8113 7327
rect 8493 7293 8527 7327
rect 9045 7293 9079 7327
rect 9597 7293 9631 7327
rect 10425 7293 10459 7327
rect 12817 7293 12851 7327
rect 13277 7293 13311 7327
rect 15301 7293 15335 7327
rect 15455 7293 15489 7327
rect 16067 7293 16101 7327
rect 16221 7293 16255 7327
rect 16313 7293 16347 7327
rect 18521 7293 18555 7327
rect 1777 7225 1811 7259
rect 5825 7225 5859 7259
rect 8677 7225 8711 7259
rect 9689 7225 9723 7259
rect 10517 7225 10551 7259
rect 13001 7225 13035 7259
rect 13185 7225 13219 7259
rect 13461 7225 13495 7259
rect 15853 7225 15887 7259
rect 16589 7225 16623 7259
rect 857 7157 891 7191
rect 3249 7157 3283 7191
rect 3617 7157 3651 7191
rect 3985 7157 4019 7191
rect 10057 7157 10091 7191
rect 10885 7157 10919 7191
rect 15669 7157 15703 7191
rect 18061 7157 18095 7191
rect 673 6953 707 6987
rect 1777 6953 1811 6987
rect 2421 6953 2455 6987
rect 3893 6953 3927 6987
rect 4813 6953 4847 6987
rect 8677 6953 8711 6987
rect 9137 6953 9171 6987
rect 16865 6953 16899 6987
rect 1317 6885 1351 6919
rect 3065 6885 3099 6919
rect 4353 6885 4387 6919
rect 7205 6885 7239 6919
rect 15393 6885 15427 6919
rect 765 6817 799 6851
rect 857 6817 891 6851
rect 1133 6817 1167 6851
rect 3157 6817 3191 6851
rect 4261 6817 4295 6851
rect 7021 6817 7055 6851
rect 7665 6817 7699 6851
rect 7849 6817 7883 6851
rect 7941 6817 7975 6851
rect 8125 6817 8159 6851
rect 8585 6817 8619 6851
rect 9137 6817 9171 6851
rect 9321 6817 9355 6851
rect 9505 6817 9539 6851
rect 9873 6817 9907 6851
rect 11621 6817 11655 6851
rect 11989 6817 12023 6851
rect 14197 6817 14231 6851
rect 14289 6817 14323 6851
rect 14473 6817 14507 6851
rect 14657 6817 14691 6851
rect 14811 6817 14845 6851
rect 17305 6817 17339 6851
rect 1501 6749 1535 6783
rect 1685 6749 1719 6783
rect 2329 6749 2363 6783
rect 3249 6749 3283 6783
rect 4537 6749 4571 6783
rect 7757 6749 7791 6783
rect 8769 6749 8803 6783
rect 11713 6749 11747 6783
rect 12449 6749 12483 6783
rect 13921 6749 13955 6783
rect 15117 6749 15151 6783
rect 17049 6749 17083 6783
rect 3801 6681 3835 6715
rect 5733 6681 5767 6715
rect 8217 6681 8251 6715
rect 12357 6681 12391 6715
rect 14289 6681 14323 6715
rect 15025 6681 15059 6715
rect 949 6613 983 6647
rect 2145 6613 2179 6647
rect 2697 6613 2731 6647
rect 3525 6613 3559 6647
rect 5181 6613 5215 6647
rect 11805 6613 11839 6647
rect 11897 6613 11931 6647
rect 18429 6613 18463 6647
rect 581 6409 615 6443
rect 4445 6409 4479 6443
rect 11326 6409 11360 6443
rect 15669 6409 15703 6443
rect 17693 6409 17727 6443
rect 18245 6409 18279 6443
rect 765 6341 799 6375
rect 3249 6341 3283 6375
rect 4261 6341 4295 6375
rect 13737 6341 13771 6375
rect 1869 6273 1903 6307
rect 5089 6273 5123 6307
rect 5917 6273 5951 6307
rect 8493 6273 8527 6307
rect 11069 6273 11103 6307
rect 13921 6273 13955 6307
rect 857 6205 891 6239
rect 1041 6205 1075 6239
rect 1317 6205 1351 6239
rect 1501 6205 1535 6239
rect 3525 6205 3559 6239
rect 3985 6205 4019 6239
rect 5733 6205 5767 6239
rect 6285 6205 6319 6239
rect 6377 6205 6411 6239
rect 6561 6205 6595 6239
rect 8677 6205 8711 6239
rect 8861 6205 8895 6239
rect 15853 6205 15887 6239
rect 17877 6205 17911 6239
rect 18429 6205 18463 6239
rect 4905 6137 4939 6171
rect 8217 6137 8251 6171
rect 9137 6137 9171 6171
rect 10701 6137 10735 6171
rect 13093 6137 13127 6171
rect 13277 6137 13311 6171
rect 14197 6137 14231 6171
rect 16129 6137 16163 6171
rect 18061 6137 18095 6171
rect 1225 6069 1259 6103
rect 3617 6069 3651 6103
rect 4813 6069 4847 6103
rect 5365 6069 5399 6103
rect 5825 6069 5859 6103
rect 6285 6069 6319 6103
rect 6745 6069 6779 6103
rect 8861 6069 8895 6103
rect 10885 6069 10919 6103
rect 13553 6069 13587 6103
rect 17601 6069 17635 6103
rect 1225 5865 1259 5899
rect 2513 5865 2547 5899
rect 2789 5865 2823 5899
rect 5733 5865 5767 5899
rect 9045 5865 9079 5899
rect 9873 5865 9907 5899
rect 14657 5865 14691 5899
rect 17877 5865 17911 5899
rect 1409 5797 1443 5831
rect 4077 5797 4111 5831
rect 4169 5797 4203 5831
rect 4629 5797 4663 5831
rect 7021 5797 7055 5831
rect 11345 5797 11379 5831
rect 12081 5797 12115 5831
rect 12725 5797 12759 5831
rect 16129 5797 16163 5831
rect 16865 5797 16899 5831
rect 1225 5729 1259 5763
rect 1593 5729 1627 5763
rect 1685 5729 1719 5763
rect 1777 5729 1811 5763
rect 2145 5729 2179 5763
rect 3157 5729 3191 5763
rect 7113 5729 7147 5763
rect 7297 5729 7331 5763
rect 7665 5729 7699 5763
rect 7941 5729 7975 5763
rect 8585 5729 8619 5763
rect 8677 5729 8711 5763
rect 9413 5729 9447 5763
rect 11713 5729 11747 5763
rect 11897 5729 11931 5763
rect 16497 5729 16531 5763
rect 16651 5729 16685 5763
rect 17417 5729 17451 5763
rect 18061 5729 18095 5763
rect 18337 5729 18371 5763
rect 2053 5661 2087 5695
rect 4353 5661 4387 5695
rect 5181 5661 5215 5695
rect 8769 5661 8803 5695
rect 9505 5661 9539 5695
rect 11621 5661 11655 5695
rect 12438 5661 12472 5695
rect 16405 5661 16439 5695
rect 17509 5661 17543 5695
rect 17601 5661 17635 5695
rect 18245 5661 18279 5695
rect 3709 5593 3743 5627
rect 7757 5593 7791 5627
rect 7849 5593 7883 5627
rect 8125 5593 8159 5627
rect 18153 5593 18187 5627
rect 765 5525 799 5559
rect 3525 5525 3559 5559
rect 4905 5525 4939 5559
rect 7297 5525 7331 5559
rect 8217 5525 8251 5559
rect 12265 5525 12299 5559
rect 14197 5525 14231 5559
rect 14381 5525 14415 5559
rect 17049 5525 17083 5559
rect 1501 5321 1535 5355
rect 5825 5321 5859 5355
rect 6469 5321 6503 5355
rect 7389 5321 7423 5355
rect 8861 5321 8895 5355
rect 15853 5321 15887 5355
rect 17417 5321 17451 5355
rect 17969 5321 18003 5355
rect 13093 5253 13127 5287
rect 15393 5253 15427 5287
rect 3249 5185 3283 5219
rect 3893 5185 3927 5219
rect 6745 5185 6779 5219
rect 8033 5185 8067 5219
rect 8769 5185 8803 5219
rect 8953 5185 8987 5219
rect 9413 5185 9447 5219
rect 16313 5185 16347 5219
rect 16405 5185 16439 5219
rect 16957 5185 16991 5219
rect 17785 5185 17819 5219
rect 4261 5117 4295 5151
rect 5825 5117 5859 5151
rect 6009 5117 6043 5151
rect 6837 5117 6871 5151
rect 6929 5117 6963 5151
rect 8309 5117 8343 5151
rect 8677 5117 8711 5151
rect 9045 5117 9079 5151
rect 12817 5117 12851 5151
rect 12909 5117 12943 5151
rect 13093 5117 13127 5151
rect 13461 5117 13495 5151
rect 15301 5117 15335 5151
rect 15577 5117 15611 5151
rect 16773 5117 16807 5151
rect 16865 5117 16899 5151
rect 17141 5117 17175 5151
rect 17233 5117 17267 5151
rect 17693 5117 17727 5151
rect 18245 5117 18279 5151
rect 2973 5049 3007 5083
rect 5733 5049 5767 5083
rect 7757 5049 7791 5083
rect 8217 5049 8251 5083
rect 13737 5049 13771 5083
rect 15485 5049 15519 5083
rect 16221 5049 16255 5083
rect 18337 5049 18371 5083
rect 18521 5049 18555 5083
rect 3709 4981 3743 5015
rect 7297 4981 7331 5015
rect 7849 4981 7883 5015
rect 10839 4981 10873 5015
rect 11529 4981 11563 5015
rect 13277 4981 13311 5015
rect 15209 4981 15243 5015
rect 16773 4981 16807 5015
rect 18429 4981 18463 5015
rect 2973 4777 3007 4811
rect 6377 4777 6411 4811
rect 6837 4777 6871 4811
rect 8217 4777 8251 4811
rect 9413 4777 9447 4811
rect 14657 4777 14691 4811
rect 16497 4777 16531 4811
rect 18429 4777 18463 4811
rect 5641 4709 5675 4743
rect 7481 4709 7515 4743
rect 7941 4709 7975 4743
rect 8033 4709 8067 4743
rect 15770 4709 15804 4743
rect 16129 4709 16163 4743
rect 3157 4641 3191 4675
rect 5181 4641 5215 4675
rect 5457 4641 5491 4675
rect 6101 4641 6135 4675
rect 6745 4641 6779 4675
rect 7757 4641 7791 4675
rect 7849 4641 7883 4675
rect 9321 4641 9355 4675
rect 9965 4641 9999 4675
rect 10241 4641 10275 4675
rect 12449 4641 12483 4675
rect 12633 4641 12667 4675
rect 12725 4641 12759 4675
rect 16405 4641 16439 4675
rect 17233 4641 17267 4675
rect 17877 4641 17911 4675
rect 18153 4641 18187 4675
rect 18337 4641 18371 4675
rect 3433 4573 3467 4607
rect 6009 4573 6043 4607
rect 7021 4573 7055 4607
rect 8309 4573 8343 4607
rect 9505 4573 9539 4607
rect 9873 4573 9907 4607
rect 10333 4573 10367 4607
rect 10609 4573 10643 4607
rect 12081 4573 12115 4607
rect 13001 4573 13035 4607
rect 16037 4573 16071 4607
rect 5273 4505 5307 4539
rect 5365 4505 5399 4539
rect 5733 4505 5767 4539
rect 8677 4505 8711 4539
rect 8953 4505 8987 4539
rect 10057 4505 10091 4539
rect 17969 4505 18003 4539
rect 18061 4505 18095 4539
rect 4905 4437 4939 4471
rect 7205 4437 7239 4471
rect 8769 4437 8803 4471
rect 10241 4437 10275 4471
rect 12265 4437 12299 4471
rect 14473 4437 14507 4471
rect 17325 4437 17359 4471
rect 17693 4437 17727 4471
rect 4077 4233 4111 4267
rect 16116 4233 16150 4267
rect 7113 4165 7147 4199
rect 15255 4165 15289 4199
rect 18061 4165 18095 4199
rect 3709 4097 3743 4131
rect 4261 4097 4295 4131
rect 4997 4097 5031 4131
rect 5825 4097 5859 4131
rect 6101 4097 6135 4131
rect 6469 4097 6503 4131
rect 6561 4097 6595 4131
rect 7389 4097 7423 4131
rect 10471 4097 10505 4131
rect 11437 4097 11471 4131
rect 13461 4097 13495 4131
rect 15853 4097 15887 4131
rect 18245 4097 18279 4131
rect 1961 4029 1995 4063
rect 7481 4029 7515 4063
rect 7757 4029 7791 4063
rect 7941 4029 7975 4063
rect 8033 4029 8067 4063
rect 8171 4029 8205 4063
rect 8309 4029 8343 4063
rect 8493 4029 8527 4063
rect 8677 4029 8711 4063
rect 9045 4029 9079 4063
rect 10793 4029 10827 4063
rect 11069 4029 11103 4063
rect 11253 4029 11287 4063
rect 11805 4029 11839 4063
rect 13231 4029 13265 4063
rect 13829 4029 13863 4063
rect 15485 4029 15519 4063
rect 17693 4029 17727 4063
rect 17786 4029 17820 4063
rect 18429 4029 18463 4063
rect 18521 4029 18555 4063
rect 2237 3961 2271 3995
rect 10701 3961 10735 3995
rect 4353 3893 4387 3927
rect 4721 3893 4755 3927
rect 4813 3893 4847 3927
rect 5181 3893 5215 3927
rect 5549 3893 5583 3927
rect 5641 3893 5675 3927
rect 6653 3893 6687 3927
rect 7021 3893 7055 3927
rect 7757 3893 7791 3927
rect 8401 3893 8435 3927
rect 11069 3893 11103 3927
rect 15577 3893 15611 3927
rect 17601 3893 17635 3927
rect 18245 3893 18279 3927
rect 2513 3689 2547 3723
rect 7297 3689 7331 3723
rect 9965 3689 9999 3723
rect 13369 3689 13403 3723
rect 13553 3689 13587 3723
rect 14289 3689 14323 3723
rect 14841 3689 14875 3723
rect 18337 3689 18371 3723
rect 2145 3621 2179 3655
rect 4721 3621 4755 3655
rect 6101 3621 6135 3655
rect 8769 3621 8803 3655
rect 10333 3621 10367 3655
rect 17049 3621 17083 3655
rect 2053 3553 2087 3587
rect 4905 3553 4939 3587
rect 5181 3553 5215 3587
rect 5719 3553 5753 3587
rect 6377 3553 6411 3587
rect 6469 3553 6503 3587
rect 6561 3553 6595 3587
rect 6837 3553 6871 3587
rect 7113 3553 7147 3587
rect 7757 3553 7791 3587
rect 7922 3553 7956 3587
rect 8033 3553 8067 3587
rect 8217 3553 8251 3587
rect 8677 3553 8711 3587
rect 8861 3553 8895 3587
rect 9229 3553 9263 3587
rect 9965 3553 9999 3587
rect 11897 3553 11931 3587
rect 13093 3553 13127 3587
rect 13277 3553 13311 3587
rect 13720 3553 13754 3587
rect 13829 3553 13863 3587
rect 14105 3553 14139 3587
rect 14197 3553 14231 3587
rect 14483 3553 14517 3587
rect 15954 3553 15988 3587
rect 16221 3553 16255 3587
rect 16497 3553 16531 3587
rect 16865 3553 16899 3587
rect 17325 3553 17359 3587
rect 17693 3553 17727 3587
rect 17969 3553 18003 3587
rect 18061 3553 18095 3587
rect 18521 3553 18555 3587
rect 1961 3485 1995 3519
rect 2697 3485 2731 3519
rect 2973 3485 3007 3519
rect 5549 3485 5583 3519
rect 7481 3485 7515 3519
rect 8401 3485 8435 3519
rect 9505 3485 9539 3519
rect 12265 3485 12299 3519
rect 12817 3485 12851 3519
rect 14657 3485 14691 3519
rect 17141 3485 17175 3519
rect 17233 3485 17267 3519
rect 17601 3485 17635 3519
rect 17785 3485 17819 3519
rect 4537 3417 4571 3451
rect 6745 3417 6779 3451
rect 14013 3417 14047 3451
rect 18245 3417 18279 3451
rect 4445 3349 4479 3383
rect 5273 3349 5307 3383
rect 5917 3349 5951 3383
rect 6929 3349 6963 3383
rect 7757 3349 7791 3383
rect 8033 3349 8067 3383
rect 8493 3349 8527 3383
rect 9137 3349 9171 3383
rect 14473 3349 14507 3383
rect 17509 3349 17543 3383
rect 3893 3145 3927 3179
rect 6285 3145 6319 3179
rect 7481 3145 7515 3179
rect 7757 3145 7791 3179
rect 11391 3145 11425 3179
rect 13553 3145 13587 3179
rect 18061 3145 18095 3179
rect 7389 3077 7423 3111
rect 8217 3077 8251 3111
rect 9505 3077 9539 3111
rect 18337 3077 18371 3111
rect 2237 3009 2271 3043
rect 4353 3009 4387 3043
rect 4537 3009 4571 3043
rect 5365 3009 5399 3043
rect 6837 3009 6871 3043
rect 7297 3009 7331 3043
rect 8769 3009 8803 3043
rect 9045 3009 9079 3043
rect 9137 3009 9171 3043
rect 9689 3009 9723 3043
rect 10885 3009 10919 3043
rect 13185 3009 13219 3043
rect 13737 3009 13771 3043
rect 15853 3009 15887 3043
rect 16129 3009 16163 3043
rect 1869 2941 1903 2975
rect 4261 2941 4295 2975
rect 5641 2941 5675 2975
rect 6653 2941 6687 2975
rect 6745 2941 6779 2975
rect 7389 2941 7423 2975
rect 7757 2941 7791 2975
rect 7941 2941 7975 2975
rect 8401 2941 8435 2975
rect 9229 2941 9263 2975
rect 9413 2941 9447 2975
rect 9781 2941 9815 2975
rect 10333 2941 10367 2975
rect 10701 2941 10735 2975
rect 12817 2941 12851 2975
rect 13461 2941 13495 2975
rect 13829 2941 13863 2975
rect 14197 2941 14231 2975
rect 17693 2941 17727 2975
rect 17877 2941 17911 2975
rect 18521 2941 18555 2975
rect 3709 2873 3743 2907
rect 6101 2873 6135 2907
rect 7113 2873 7147 2907
rect 8953 2873 8987 2907
rect 10499 2873 10533 2907
rect 13737 2873 13771 2907
rect 4721 2805 4755 2839
rect 5089 2805 5123 2839
rect 5181 2805 5215 2839
rect 8769 2805 8803 2839
rect 10609 2805 10643 2839
rect 11161 2805 11195 2839
rect 15623 2805 15657 2839
rect 17601 2805 17635 2839
rect 2881 2601 2915 2635
rect 3341 2601 3375 2635
rect 5181 2601 5215 2635
rect 9321 2601 9355 2635
rect 16313 2601 16347 2635
rect 1961 2533 1995 2567
rect 14657 2533 14691 2567
rect 16773 2533 16807 2567
rect 2329 2465 2363 2499
rect 3249 2465 3283 2499
rect 3893 2465 3927 2499
rect 4721 2465 4755 2499
rect 5089 2465 5123 2499
rect 5273 2465 5307 2499
rect 5733 2465 5767 2499
rect 6101 2465 6135 2499
rect 6469 2465 6503 2499
rect 6745 2465 6779 2499
rect 7297 2465 7331 2499
rect 9597 2465 9631 2499
rect 11621 2465 11655 2499
rect 12265 2465 12299 2499
rect 14197 2465 14231 2499
rect 14381 2465 14415 2499
rect 14933 2465 14967 2499
rect 15189 2465 15223 2499
rect 17417 2465 17451 2499
rect 18245 2465 18279 2499
rect 3433 2397 3467 2431
rect 3801 2397 3835 2431
rect 4445 2397 4479 2431
rect 7481 2397 7515 2431
rect 7757 2397 7791 2431
rect 9321 2397 9355 2431
rect 11345 2397 11379 2431
rect 12541 2397 12575 2431
rect 17141 2397 17175 2431
rect 17325 2397 17359 2431
rect 18153 2397 18187 2431
rect 4537 2329 4571 2363
rect 9505 2329 9539 2363
rect 14381 2329 14415 2363
rect 17877 2329 17911 2363
rect 4169 2261 4203 2295
rect 4905 2261 4939 2295
rect 5457 2261 5491 2295
rect 9229 2261 9263 2295
rect 9873 2261 9907 2295
rect 11897 2261 11931 2295
rect 11989 2261 12023 2295
rect 14013 2261 14047 2295
rect 16497 2261 16531 2295
rect 17785 2261 17819 2295
rect 4629 2057 4663 2091
rect 6009 2057 6043 2091
rect 7297 2057 7331 2091
rect 8309 2057 8343 2091
rect 9413 2057 9447 2091
rect 9781 2057 9815 2091
rect 10793 2057 10827 2091
rect 12265 2057 12299 2091
rect 12633 2057 12667 2091
rect 16773 2057 16807 2091
rect 16865 2057 16899 2091
rect 17049 2057 17083 2091
rect 18521 2057 18555 2091
rect 10609 1989 10643 2023
rect 17969 1989 18003 2023
rect 5825 1921 5859 1955
rect 6285 1921 6319 1955
rect 6469 1921 6503 1955
rect 6745 1921 6779 1955
rect 7113 1921 7147 1955
rect 7573 1921 7607 1955
rect 9317 1921 9351 1955
rect 10057 1921 10091 1955
rect 11621 1921 11655 1955
rect 12035 1921 12069 1955
rect 13277 1921 13311 1955
rect 13921 1921 13955 1955
rect 14105 1921 14139 1955
rect 14289 1921 14323 1955
rect 16497 1921 16531 1955
rect 16957 1921 16991 1955
rect 17601 1921 17635 1955
rect 3065 1853 3099 1887
rect 4261 1853 4295 1887
rect 4353 1853 4387 1887
rect 4445 1853 4479 1887
rect 4813 1853 4847 1887
rect 4997 1853 5031 1887
rect 5089 1853 5123 1887
rect 5273 1853 5307 1887
rect 5733 1853 5767 1887
rect 6101 1853 6135 1887
rect 7757 1853 7791 1887
rect 8217 1847 8251 1881
rect 8861 1853 8895 1887
rect 8953 1853 8987 1887
rect 9041 1853 9075 1887
rect 9229 1853 9263 1887
rect 9505 1853 9539 1887
rect 9597 1853 9631 1887
rect 10701 1853 10735 1887
rect 11897 1853 11931 1887
rect 12173 1853 12207 1887
rect 12357 1853 12391 1887
rect 12817 1853 12851 1887
rect 16681 1853 16715 1887
rect 17509 1853 17543 1887
rect 17877 1853 17911 1887
rect 18061 1853 18095 1887
rect 18337 1853 18371 1887
rect 18521 1853 18555 1887
rect 2973 1785 3007 1819
rect 10149 1785 10183 1819
rect 11529 1785 11563 1819
rect 14556 1785 14590 1819
rect 16313 1785 16347 1819
rect 17417 1785 17451 1819
rect 4077 1717 4111 1751
rect 5825 1717 5859 1751
rect 7113 1717 7147 1751
rect 7665 1717 7699 1751
rect 8125 1717 8159 1751
rect 10241 1717 10275 1751
rect 11069 1717 11103 1751
rect 11437 1717 11471 1751
rect 13461 1717 13495 1751
rect 13829 1717 13863 1751
rect 15669 1717 15703 1751
rect 15853 1717 15887 1751
rect 16221 1717 16255 1751
rect 4675 1513 4709 1547
rect 5181 1513 5215 1547
rect 6193 1513 6227 1547
rect 7481 1513 7515 1547
rect 7941 1513 7975 1547
rect 8769 1513 8803 1547
rect 10425 1513 10459 1547
rect 11437 1513 11471 1547
rect 11989 1513 12023 1547
rect 12541 1513 12575 1547
rect 12909 1513 12943 1547
rect 13737 1513 13771 1547
rect 14105 1513 14139 1547
rect 14473 1513 14507 1547
rect 16313 1513 16347 1547
rect 18061 1513 18095 1547
rect 11161 1445 11195 1479
rect 16773 1445 16807 1479
rect 17693 1445 17727 1479
rect 2881 1377 2915 1411
rect 5273 1377 5307 1411
rect 6101 1377 6135 1411
rect 7757 1377 7791 1411
rect 8309 1377 8343 1411
rect 9413 1377 9447 1411
rect 9873 1377 9907 1411
rect 10149 1377 10183 1411
rect 10701 1377 10735 1411
rect 11345 1377 11379 1411
rect 11529 1377 11563 1411
rect 12265 1377 12299 1411
rect 13185 1377 13219 1411
rect 13277 1377 13311 1411
rect 13645 1377 13679 1411
rect 14933 1377 14967 1411
rect 15200 1377 15234 1411
rect 17877 1377 17911 1411
rect 18153 1377 18187 1411
rect 18337 1377 18371 1411
rect 3249 1309 3283 1343
rect 6377 1309 6411 1343
rect 7481 1309 7515 1343
rect 8401 1309 8435 1343
rect 8493 1309 8527 1343
rect 9689 1309 9723 1343
rect 12541 1309 12575 1343
rect 13461 1309 13495 1343
rect 17049 1309 17083 1343
rect 17417 1309 17451 1343
rect 5733 1241 5767 1275
rect 9505 1241 9539 1275
rect 9597 1241 9631 1275
rect 12357 1241 12391 1275
rect 14289 1241 14323 1275
rect 16497 1241 16531 1275
rect 7665 1173 7699 1207
rect 10885 1173 10919 1207
rect 11897 1173 11931 1207
rect 12817 1173 12851 1207
rect 13277 1173 13311 1207
rect 14749 1173 14783 1207
rect 18429 1173 18463 1207
rect 7481 969 7515 1003
rect 8769 969 8803 1003
rect 9873 969 9907 1003
rect 10241 969 10275 1003
rect 13553 969 13587 1003
rect 15577 969 15611 1003
rect 16589 969 16623 1003
rect 17141 969 17175 1003
rect 17417 969 17451 1003
rect 18337 969 18371 1003
rect 14105 901 14139 935
rect 14197 901 14231 935
rect 14473 901 14507 935
rect 15485 901 15519 935
rect 6837 833 6871 867
rect 7941 833 7975 867
rect 8125 833 8159 867
rect 9965 833 9999 867
rect 12357 833 12391 867
rect 13277 833 13311 867
rect 16037 833 16071 867
rect 6929 765 6963 799
rect 8769 765 8803 799
rect 9873 765 9907 799
rect 12817 765 12851 799
rect 13001 765 13035 799
rect 13829 765 13863 799
rect 14013 765 14047 799
rect 14289 765 14323 799
rect 14841 765 14875 799
rect 15025 765 15059 799
rect 15209 765 15243 799
rect 17693 765 17727 799
rect 17877 765 17911 799
rect 18521 765 18555 799
rect 7849 697 7883 731
rect 16129 697 16163 731
rect 16221 697 16255 731
rect 16865 697 16899 731
rect 7297 629 7331 663
rect 12081 629 12115 663
rect 12541 629 12575 663
rect 12725 629 12759 663
rect 13093 629 13127 663
rect 15209 629 15243 663
rect 18061 629 18095 663
<< metal1 >>
rect 7282 11364 7288 11416
rect 7340 11404 7346 11416
rect 9674 11404 9680 11416
rect 7340 11376 9680 11404
rect 7340 11364 7346 11376
rect 9674 11364 9680 11376
rect 9732 11404 9738 11416
rect 17586 11404 17592 11416
rect 9732 11376 17592 11404
rect 9732 11364 9738 11376
rect 17586 11364 17592 11376
rect 17644 11364 17650 11416
rect 1302 11228 1308 11280
rect 1360 11268 1366 11280
rect 4522 11268 4528 11280
rect 1360 11240 4528 11268
rect 1360 11228 1366 11240
rect 4522 11228 4528 11240
rect 4580 11228 4586 11280
rect 4614 11228 4620 11280
rect 4672 11268 4678 11280
rect 6546 11268 6552 11280
rect 4672 11240 6552 11268
rect 4672 11228 4678 11240
rect 6546 11228 6552 11240
rect 6604 11268 6610 11280
rect 9766 11268 9772 11280
rect 6604 11240 9772 11268
rect 6604 11228 6610 11240
rect 9766 11228 9772 11240
rect 9824 11228 9830 11280
rect 4154 11160 4160 11212
rect 4212 11200 4218 11212
rect 4632 11200 4660 11228
rect 4212 11172 4660 11200
rect 4212 11160 4218 11172
rect 9122 11160 9128 11212
rect 9180 11200 9186 11212
rect 12250 11200 12256 11212
rect 9180 11172 12256 11200
rect 9180 11160 9186 11172
rect 12250 11160 12256 11172
rect 12308 11160 12314 11212
rect 1946 11092 1952 11144
rect 2004 11132 2010 11144
rect 8754 11132 8760 11144
rect 2004 11104 8760 11132
rect 2004 11092 2010 11104
rect 8754 11092 8760 11104
rect 8812 11092 8818 11144
rect 9214 11092 9220 11144
rect 9272 11132 9278 11144
rect 12158 11132 12164 11144
rect 9272 11104 12164 11132
rect 9272 11092 9278 11104
rect 12158 11092 12164 11104
rect 12216 11092 12222 11144
rect 16114 11092 16120 11144
rect 16172 11132 16178 11144
rect 17678 11132 17684 11144
rect 16172 11104 17684 11132
rect 16172 11092 16178 11104
rect 17678 11092 17684 11104
rect 17736 11092 17742 11144
rect 566 11024 572 11076
rect 624 11064 630 11076
rect 2866 11064 2872 11076
rect 624 11036 2872 11064
rect 624 11024 630 11036
rect 2866 11024 2872 11036
rect 2924 11024 2930 11076
rect 2958 11024 2964 11076
rect 3016 11064 3022 11076
rect 4982 11064 4988 11076
rect 3016 11036 4988 11064
rect 3016 11024 3022 11036
rect 4982 11024 4988 11036
rect 5040 11024 5046 11076
rect 6914 11064 6920 11076
rect 5184 11036 6920 11064
rect 1854 10956 1860 11008
rect 1912 10996 1918 11008
rect 5184 10996 5212 11036
rect 6914 11024 6920 11036
rect 6972 11024 6978 11076
rect 11882 11024 11888 11076
rect 11940 11064 11946 11076
rect 16574 11064 16580 11076
rect 11940 11036 16580 11064
rect 11940 11024 11946 11036
rect 16574 11024 16580 11036
rect 16632 11024 16638 11076
rect 1912 10968 5212 10996
rect 1912 10956 1918 10968
rect 5258 10956 5264 11008
rect 5316 10996 5322 11008
rect 7650 10996 7656 11008
rect 5316 10968 7656 10996
rect 5316 10956 5322 10968
rect 7650 10956 7656 10968
rect 7708 10956 7714 11008
rect 12066 10956 12072 11008
rect 12124 10996 12130 11008
rect 18230 10996 18236 11008
rect 12124 10968 18236 10996
rect 12124 10956 12130 10968
rect 18230 10956 18236 10968
rect 18288 10956 18294 11008
rect 184 10906 18924 10928
rect 184 10854 3110 10906
rect 3162 10854 3174 10906
rect 3226 10854 3238 10906
rect 3290 10854 3302 10906
rect 3354 10854 3366 10906
rect 3418 10854 6210 10906
rect 6262 10854 6274 10906
rect 6326 10854 6338 10906
rect 6390 10854 6402 10906
rect 6454 10854 6466 10906
rect 6518 10854 9310 10906
rect 9362 10854 9374 10906
rect 9426 10854 9438 10906
rect 9490 10854 9502 10906
rect 9554 10854 9566 10906
rect 9618 10854 12410 10906
rect 12462 10854 12474 10906
rect 12526 10854 12538 10906
rect 12590 10854 12602 10906
rect 12654 10854 12666 10906
rect 12718 10854 15510 10906
rect 15562 10854 15574 10906
rect 15626 10854 15638 10906
rect 15690 10854 15702 10906
rect 15754 10854 15766 10906
rect 15818 10854 18610 10906
rect 18662 10854 18674 10906
rect 18726 10854 18738 10906
rect 18790 10854 18802 10906
rect 18854 10854 18866 10906
rect 18918 10854 18924 10906
rect 184 10832 18924 10854
rect 566 10792 572 10804
rect 527 10764 572 10792
rect 566 10752 572 10764
rect 624 10752 630 10804
rect 4338 10792 4344 10804
rect 2056 10764 4344 10792
rect 1118 10656 1124 10668
rect 1079 10628 1124 10656
rect 1118 10616 1124 10628
rect 1176 10616 1182 10668
rect 1946 10656 1952 10668
rect 1907 10628 1952 10656
rect 1946 10616 1952 10628
rect 2004 10616 2010 10668
rect 2056 10665 2084 10764
rect 4338 10752 4344 10764
rect 4396 10752 4402 10804
rect 5258 10792 5264 10804
rect 5219 10764 5264 10792
rect 5258 10752 5264 10764
rect 5316 10752 5322 10804
rect 5810 10792 5816 10804
rect 5644 10764 5816 10792
rect 2498 10724 2504 10736
rect 2459 10696 2504 10724
rect 2498 10684 2504 10696
rect 2556 10684 2562 10736
rect 2041 10659 2099 10665
rect 2041 10625 2053 10659
rect 2087 10625 2099 10659
rect 2041 10619 2099 10625
rect 2958 10616 2964 10668
rect 3016 10656 3022 10668
rect 3053 10659 3111 10665
rect 3053 10656 3065 10659
rect 3016 10628 3065 10656
rect 3016 10616 3022 10628
rect 3053 10625 3065 10628
rect 3099 10625 3111 10659
rect 3053 10619 3111 10625
rect 3237 10659 3295 10665
rect 3237 10625 3249 10659
rect 3283 10656 3295 10659
rect 4062 10656 4068 10668
rect 3283 10628 4068 10656
rect 3283 10625 3295 10628
rect 3237 10619 3295 10625
rect 4062 10616 4068 10628
rect 4120 10616 4126 10668
rect 4801 10659 4859 10665
rect 4801 10625 4813 10659
rect 4847 10656 4859 10659
rect 5644 10656 5672 10764
rect 5810 10752 5816 10764
rect 5868 10792 5874 10804
rect 8849 10795 8907 10801
rect 5868 10764 6776 10792
rect 5868 10752 5874 10764
rect 6549 10727 6607 10733
rect 6549 10724 6561 10727
rect 4847 10628 5672 10656
rect 5736 10696 6561 10724
rect 4847 10625 4859 10628
rect 4801 10619 4859 10625
rect 750 10588 756 10600
rect 711 10560 756 10588
rect 750 10548 756 10560
rect 808 10548 814 10600
rect 845 10591 903 10597
rect 845 10557 857 10591
rect 891 10588 903 10591
rect 1394 10588 1400 10600
rect 891 10560 1400 10588
rect 891 10557 903 10560
rect 845 10551 903 10557
rect 1394 10548 1400 10560
rect 1452 10548 1458 10600
rect 1670 10588 1676 10600
rect 1631 10560 1676 10588
rect 1670 10548 1676 10560
rect 1728 10548 1734 10600
rect 2774 10548 2780 10600
rect 2832 10588 2838 10600
rect 2869 10591 2927 10597
rect 2869 10588 2881 10591
rect 2832 10560 2881 10588
rect 2832 10548 2838 10560
rect 2869 10557 2881 10560
rect 2915 10557 2927 10591
rect 2869 10551 2927 10557
rect 3329 10591 3387 10597
rect 3329 10557 3341 10591
rect 3375 10588 3387 10591
rect 4522 10588 4528 10600
rect 3375 10560 4200 10588
rect 4483 10560 4528 10588
rect 3375 10557 3387 10560
rect 3329 10551 3387 10557
rect 474 10480 480 10532
rect 532 10520 538 10532
rect 1581 10523 1639 10529
rect 1581 10520 1593 10523
rect 532 10492 1593 10520
rect 532 10480 538 10492
rect 1581 10489 1593 10492
rect 1627 10489 1639 10523
rect 1581 10483 1639 10489
rect 2130 10412 2136 10464
rect 2188 10452 2194 10464
rect 2682 10452 2688 10464
rect 2188 10424 2233 10452
rect 2643 10424 2688 10452
rect 2188 10412 2194 10424
rect 2682 10412 2688 10424
rect 2740 10412 2746 10464
rect 3697 10455 3755 10461
rect 3697 10421 3709 10455
rect 3743 10452 3755 10455
rect 3878 10452 3884 10464
rect 3743 10424 3884 10452
rect 3743 10421 3755 10424
rect 3697 10415 3755 10421
rect 3878 10412 3884 10424
rect 3936 10412 3942 10464
rect 4062 10452 4068 10464
rect 4023 10424 4068 10452
rect 4062 10412 4068 10424
rect 4120 10412 4126 10464
rect 4172 10461 4200 10560
rect 4522 10548 4528 10560
rect 4580 10548 4586 10600
rect 4614 10548 4620 10600
rect 4672 10588 4678 10600
rect 5736 10597 5764 10696
rect 6549 10693 6561 10696
rect 6595 10693 6607 10727
rect 6748 10724 6776 10764
rect 8849 10761 8861 10795
rect 8895 10792 8907 10795
rect 9766 10792 9772 10804
rect 8895 10764 9772 10792
rect 8895 10761 8907 10764
rect 8849 10755 8907 10761
rect 9766 10752 9772 10764
rect 9824 10792 9830 10804
rect 11882 10792 11888 10804
rect 9824 10764 9996 10792
rect 11843 10764 11888 10792
rect 9824 10752 9830 10764
rect 9214 10724 9220 10736
rect 6748 10696 9220 10724
rect 6549 10687 6607 10693
rect 5902 10656 5908 10668
rect 5863 10628 5908 10656
rect 5902 10616 5908 10628
rect 5960 10616 5966 10668
rect 6457 10659 6515 10665
rect 6457 10625 6469 10659
rect 6503 10656 6515 10659
rect 7006 10656 7012 10668
rect 6503 10628 7012 10656
rect 6503 10625 6515 10628
rect 6457 10619 6515 10625
rect 7006 10616 7012 10628
rect 7064 10616 7070 10668
rect 7116 10665 7144 10696
rect 9214 10684 9220 10696
rect 9272 10684 9278 10736
rect 9674 10724 9680 10736
rect 9635 10696 9680 10724
rect 9674 10684 9680 10696
rect 9732 10684 9738 10736
rect 7101 10659 7159 10665
rect 7101 10625 7113 10659
rect 7147 10625 7159 10659
rect 7101 10619 7159 10625
rect 7374 10616 7380 10668
rect 7432 10656 7438 10668
rect 8021 10659 8079 10665
rect 8021 10656 8033 10659
rect 7432 10628 8033 10656
rect 7432 10616 7438 10628
rect 8021 10625 8033 10628
rect 8067 10625 8079 10659
rect 9692 10656 9720 10684
rect 9968 10665 9996 10764
rect 11882 10752 11888 10764
rect 11940 10752 11946 10804
rect 11974 10752 11980 10804
rect 12032 10792 12038 10804
rect 12805 10795 12863 10801
rect 12805 10792 12817 10795
rect 12032 10764 12817 10792
rect 12032 10752 12038 10764
rect 12805 10761 12817 10764
rect 12851 10761 12863 10795
rect 12805 10755 12863 10761
rect 14918 10752 14924 10804
rect 14976 10792 14982 10804
rect 17954 10792 17960 10804
rect 14976 10764 17960 10792
rect 14976 10752 14982 10764
rect 17954 10752 17960 10764
rect 18012 10752 18018 10804
rect 18230 10792 18236 10804
rect 18191 10764 18236 10792
rect 18230 10752 18236 10764
rect 18288 10752 18294 10804
rect 11793 10727 11851 10733
rect 11793 10693 11805 10727
rect 11839 10724 11851 10727
rect 13446 10724 13452 10736
rect 11839 10696 13452 10724
rect 11839 10693 11851 10696
rect 11793 10687 11851 10693
rect 13446 10684 13452 10696
rect 13504 10684 13510 10736
rect 14369 10727 14427 10733
rect 14369 10693 14381 10727
rect 14415 10724 14427 10727
rect 17221 10727 17279 10733
rect 17221 10724 17233 10727
rect 14415 10696 17233 10724
rect 14415 10693 14427 10696
rect 14369 10687 14427 10693
rect 17221 10693 17233 10696
rect 17267 10693 17279 10727
rect 17678 10724 17684 10736
rect 17639 10696 17684 10724
rect 17221 10687 17279 10693
rect 17678 10684 17684 10696
rect 17736 10684 17742 10736
rect 8021 10619 8079 10625
rect 9048 10628 9720 10656
rect 9953 10659 10011 10665
rect 5721 10591 5779 10597
rect 4672 10560 4717 10588
rect 4672 10548 4678 10560
rect 5721 10557 5733 10591
rect 5767 10557 5779 10591
rect 5721 10551 5779 10557
rect 6917 10591 6975 10597
rect 6917 10557 6929 10591
rect 6963 10588 6975 10591
rect 7190 10588 7196 10600
rect 6963 10560 7196 10588
rect 6963 10557 6975 10560
rect 6917 10551 6975 10557
rect 7190 10548 7196 10560
rect 7248 10548 7254 10600
rect 7837 10591 7895 10597
rect 7837 10557 7849 10591
rect 7883 10588 7895 10591
rect 8110 10588 8116 10600
rect 7883 10560 8116 10588
rect 7883 10557 7895 10560
rect 7837 10551 7895 10557
rect 8110 10548 8116 10560
rect 8168 10548 8174 10600
rect 8202 10548 8208 10600
rect 8260 10588 8266 10600
rect 9048 10597 9076 10628
rect 9953 10625 9965 10659
rect 9999 10656 10011 10659
rect 10134 10656 10140 10668
rect 9999 10628 10140 10656
rect 9999 10625 10011 10628
rect 9953 10619 10011 10625
rect 10134 10616 10140 10628
rect 10192 10616 10198 10668
rect 10594 10656 10600 10668
rect 10555 10628 10600 10656
rect 10594 10616 10600 10628
rect 10652 10656 10658 10668
rect 11149 10659 11207 10665
rect 11149 10656 11161 10659
rect 10652 10628 11161 10656
rect 10652 10616 10658 10628
rect 11149 10625 11161 10628
rect 11195 10625 11207 10659
rect 11149 10619 11207 10625
rect 12158 10616 12164 10668
rect 12216 10656 12222 10668
rect 12529 10659 12587 10665
rect 12529 10656 12541 10659
rect 12216 10628 12541 10656
rect 12216 10616 12222 10628
rect 12529 10625 12541 10628
rect 12575 10625 12587 10659
rect 12529 10619 12587 10625
rect 12713 10659 12771 10665
rect 12713 10625 12725 10659
rect 12759 10656 12771 10659
rect 12894 10656 12900 10668
rect 12759 10628 12900 10656
rect 12759 10625 12771 10628
rect 12713 10619 12771 10625
rect 12894 10616 12900 10628
rect 12952 10616 12958 10668
rect 13817 10659 13875 10665
rect 13817 10625 13829 10659
rect 13863 10656 13875 10659
rect 14458 10656 14464 10668
rect 13863 10628 14464 10656
rect 13863 10625 13875 10628
rect 13817 10619 13875 10625
rect 14458 10616 14464 10628
rect 14516 10616 14522 10668
rect 14918 10656 14924 10668
rect 14879 10628 14924 10656
rect 14918 10616 14924 10628
rect 14976 10616 14982 10668
rect 16761 10659 16819 10665
rect 15028 10628 16712 10656
rect 8757 10591 8815 10597
rect 8757 10588 8769 10591
rect 8260 10560 8769 10588
rect 8260 10548 8266 10560
rect 8757 10557 8769 10560
rect 8803 10557 8815 10591
rect 8757 10551 8815 10557
rect 9033 10591 9091 10597
rect 9033 10557 9045 10591
rect 9079 10557 9091 10591
rect 9214 10588 9220 10600
rect 9175 10560 9220 10588
rect 9033 10551 9091 10557
rect 9214 10548 9220 10560
rect 9272 10548 9278 10600
rect 9306 10548 9312 10600
rect 9364 10588 9370 10600
rect 11514 10588 11520 10600
rect 9364 10560 11520 10588
rect 9364 10548 9370 10560
rect 11514 10548 11520 10560
rect 11572 10548 11578 10600
rect 11882 10588 11888 10600
rect 11843 10560 11888 10588
rect 11882 10548 11888 10560
rect 11940 10548 11946 10600
rect 12066 10588 12072 10600
rect 12027 10560 12072 10588
rect 12066 10548 12072 10560
rect 12124 10548 12130 10600
rect 12250 10588 12256 10600
rect 12211 10560 12256 10588
rect 12250 10548 12256 10560
rect 12308 10548 12314 10600
rect 12621 10591 12679 10597
rect 12621 10588 12633 10591
rect 12360 10560 12633 10588
rect 9766 10480 9772 10532
rect 9824 10520 9830 10532
rect 10505 10523 10563 10529
rect 10505 10520 10517 10523
rect 9824 10492 10517 10520
rect 9824 10480 9830 10492
rect 10505 10489 10517 10492
rect 10551 10489 10563 10523
rect 10505 10483 10563 10489
rect 11425 10523 11483 10529
rect 11425 10489 11437 10523
rect 11471 10520 11483 10523
rect 11471 10492 12112 10520
rect 11471 10489 11483 10492
rect 11425 10483 11483 10489
rect 4157 10455 4215 10461
rect 4157 10421 4169 10455
rect 4203 10421 4215 10455
rect 4157 10415 4215 10421
rect 5353 10455 5411 10461
rect 5353 10421 5365 10455
rect 5399 10452 5411 10455
rect 5442 10452 5448 10464
rect 5399 10424 5448 10452
rect 5399 10421 5411 10424
rect 5353 10415 5411 10421
rect 5442 10412 5448 10424
rect 5500 10412 5506 10464
rect 5534 10412 5540 10464
rect 5592 10452 5598 10464
rect 5813 10455 5871 10461
rect 5813 10452 5825 10455
rect 5592 10424 5825 10452
rect 5592 10412 5598 10424
rect 5813 10421 5825 10424
rect 5859 10452 5871 10455
rect 6086 10452 6092 10464
rect 5859 10424 6092 10452
rect 5859 10421 5871 10424
rect 5813 10415 5871 10421
rect 6086 10412 6092 10424
rect 6144 10452 6150 10464
rect 7009 10455 7067 10461
rect 7009 10452 7021 10455
rect 6144 10424 7021 10452
rect 6144 10412 6150 10424
rect 7009 10421 7021 10424
rect 7055 10452 7067 10455
rect 7282 10452 7288 10464
rect 7055 10424 7288 10452
rect 7055 10421 7067 10424
rect 7009 10415 7067 10421
rect 7282 10412 7288 10424
rect 7340 10412 7346 10464
rect 7469 10455 7527 10461
rect 7469 10421 7481 10455
rect 7515 10452 7527 10455
rect 7558 10452 7564 10464
rect 7515 10424 7564 10452
rect 7515 10421 7527 10424
rect 7469 10415 7527 10421
rect 7558 10412 7564 10424
rect 7616 10412 7622 10464
rect 7650 10412 7656 10464
rect 7708 10452 7714 10464
rect 7929 10455 7987 10461
rect 7929 10452 7941 10455
rect 7708 10424 7941 10452
rect 7708 10412 7714 10424
rect 7929 10421 7941 10424
rect 7975 10452 7987 10455
rect 8202 10452 8208 10464
rect 7975 10424 8208 10452
rect 7975 10421 7987 10424
rect 7929 10415 7987 10421
rect 8202 10412 8208 10424
rect 8260 10452 8266 10464
rect 8389 10455 8447 10461
rect 8389 10452 8401 10455
rect 8260 10424 8401 10452
rect 8260 10412 8266 10424
rect 8389 10421 8401 10424
rect 8435 10421 8447 10455
rect 8389 10415 8447 10421
rect 9122 10412 9128 10464
rect 9180 10452 9186 10464
rect 9490 10452 9496 10464
rect 9180 10424 9225 10452
rect 9451 10424 9496 10452
rect 9180 10412 9186 10424
rect 9490 10412 9496 10424
rect 9548 10412 9554 10464
rect 9950 10412 9956 10464
rect 10008 10452 10014 10464
rect 10045 10455 10103 10461
rect 10045 10452 10057 10455
rect 10008 10424 10057 10452
rect 10008 10412 10014 10424
rect 10045 10421 10057 10424
rect 10091 10421 10103 10455
rect 10045 10415 10103 10421
rect 10134 10412 10140 10464
rect 10192 10452 10198 10464
rect 10413 10455 10471 10461
rect 10413 10452 10425 10455
rect 10192 10424 10425 10452
rect 10192 10412 10198 10424
rect 10413 10421 10425 10424
rect 10459 10421 10471 10455
rect 11330 10452 11336 10464
rect 11291 10424 11336 10452
rect 10413 10415 10471 10421
rect 11330 10412 11336 10424
rect 11388 10412 11394 10464
rect 12084 10452 12112 10492
rect 12158 10480 12164 10532
rect 12216 10520 12222 10532
rect 12360 10520 12388 10560
rect 12621 10557 12633 10560
rect 12667 10557 12679 10591
rect 12621 10551 12679 10557
rect 12802 10548 12808 10600
rect 12860 10588 12866 10600
rect 12989 10591 13047 10597
rect 12989 10588 13001 10591
rect 12860 10560 13001 10588
rect 12860 10548 12866 10560
rect 12989 10557 13001 10560
rect 13035 10557 13047 10591
rect 12989 10551 13047 10557
rect 13541 10591 13599 10597
rect 13541 10557 13553 10591
rect 13587 10588 13599 10591
rect 14642 10588 14648 10600
rect 13587 10560 14648 10588
rect 13587 10557 13599 10560
rect 13541 10551 13599 10557
rect 14642 10548 14648 10560
rect 14700 10548 14706 10600
rect 12216 10492 12388 10520
rect 12216 10480 12222 10492
rect 12434 10480 12440 10532
rect 12492 10520 12498 10532
rect 13814 10520 13820 10532
rect 12492 10492 12537 10520
rect 12728 10492 13820 10520
rect 12492 10480 12498 10492
rect 12728 10452 12756 10492
rect 13814 10480 13820 10492
rect 13872 10480 13878 10532
rect 13909 10523 13967 10529
rect 13909 10489 13921 10523
rect 13955 10520 13967 10523
rect 14826 10520 14832 10532
rect 13955 10492 14832 10520
rect 13955 10489 13967 10492
rect 13909 10483 13967 10489
rect 14826 10480 14832 10492
rect 14884 10480 14890 10532
rect 12986 10452 12992 10464
rect 12084 10424 12756 10452
rect 12947 10424 12992 10452
rect 12986 10412 12992 10424
rect 13044 10412 13050 10464
rect 14001 10455 14059 10461
rect 14001 10421 14013 10455
rect 14047 10452 14059 10455
rect 15028 10452 15056 10628
rect 15654 10548 15660 10600
rect 15712 10588 15718 10600
rect 16684 10597 16712 10628
rect 16761 10625 16773 10659
rect 16807 10656 16819 10659
rect 18230 10656 18236 10668
rect 16807 10628 18236 10656
rect 16807 10625 16819 10628
rect 16761 10619 16819 10625
rect 18230 10616 18236 10628
rect 18288 10616 18294 10668
rect 16669 10591 16727 10597
rect 15712 10560 16252 10588
rect 15712 10548 15718 10560
rect 15105 10523 15163 10529
rect 15105 10489 15117 10523
rect 15151 10520 15163 10523
rect 15286 10520 15292 10532
rect 15151 10492 15292 10520
rect 15151 10489 15163 10492
rect 15105 10483 15163 10489
rect 15286 10480 15292 10492
rect 15344 10480 15350 10532
rect 16022 10520 16028 10532
rect 15983 10492 16028 10520
rect 16022 10480 16028 10492
rect 16080 10480 16086 10532
rect 15194 10452 15200 10464
rect 14047 10424 15056 10452
rect 15155 10424 15200 10452
rect 14047 10421 14059 10424
rect 14001 10415 14059 10421
rect 15194 10412 15200 10424
rect 15252 10412 15258 10464
rect 15562 10452 15568 10464
rect 15523 10424 15568 10452
rect 15562 10412 15568 10424
rect 15620 10412 15626 10464
rect 15930 10452 15936 10464
rect 15891 10424 15936 10452
rect 15930 10412 15936 10424
rect 15988 10412 15994 10464
rect 16114 10452 16120 10464
rect 16075 10424 16120 10452
rect 16114 10412 16120 10424
rect 16172 10412 16178 10464
rect 16224 10461 16252 10560
rect 16669 10557 16681 10591
rect 16715 10588 16727 10591
rect 17770 10588 17776 10600
rect 16715 10560 17776 10588
rect 16715 10557 16727 10560
rect 16669 10551 16727 10557
rect 17770 10548 17776 10560
rect 17828 10548 17834 10600
rect 17862 10548 17868 10600
rect 17920 10588 17926 10600
rect 18049 10591 18107 10597
rect 17920 10560 17965 10588
rect 17920 10548 17926 10560
rect 18049 10557 18061 10591
rect 18095 10588 18107 10591
rect 18138 10588 18144 10600
rect 18095 10560 18144 10588
rect 18095 10557 18107 10560
rect 18049 10551 18107 10557
rect 18138 10548 18144 10560
rect 18196 10548 18202 10600
rect 18414 10588 18420 10600
rect 18375 10560 18420 10588
rect 18414 10548 18420 10560
rect 18472 10548 18478 10600
rect 16393 10523 16451 10529
rect 16393 10489 16405 10523
rect 16439 10520 16451 10523
rect 17586 10520 17592 10532
rect 16439 10492 17172 10520
rect 17547 10492 17592 10520
rect 16439 10489 16451 10492
rect 16393 10483 16451 10489
rect 16209 10455 16267 10461
rect 16209 10421 16221 10455
rect 16255 10421 16267 10455
rect 16482 10452 16488 10464
rect 16443 10424 16488 10452
rect 16209 10415 16267 10421
rect 16482 10412 16488 10424
rect 16540 10412 16546 10464
rect 17144 10461 17172 10492
rect 17586 10480 17592 10492
rect 17644 10480 17650 10532
rect 17129 10455 17187 10461
rect 17129 10421 17141 10455
rect 17175 10421 17187 10455
rect 17129 10415 17187 10421
rect 184 10362 18860 10384
rect 184 10310 4660 10362
rect 4712 10310 4724 10362
rect 4776 10310 4788 10362
rect 4840 10310 4852 10362
rect 4904 10310 4916 10362
rect 4968 10310 7760 10362
rect 7812 10310 7824 10362
rect 7876 10310 7888 10362
rect 7940 10310 7952 10362
rect 8004 10310 8016 10362
rect 8068 10310 10860 10362
rect 10912 10310 10924 10362
rect 10976 10310 10988 10362
rect 11040 10310 11052 10362
rect 11104 10310 11116 10362
rect 11168 10310 13960 10362
rect 14012 10310 14024 10362
rect 14076 10310 14088 10362
rect 14140 10310 14152 10362
rect 14204 10310 14216 10362
rect 14268 10310 17060 10362
rect 17112 10310 17124 10362
rect 17176 10310 17188 10362
rect 17240 10310 17252 10362
rect 17304 10310 17316 10362
rect 17368 10310 18860 10362
rect 184 10288 18860 10310
rect 2130 10208 2136 10260
rect 2188 10248 2194 10260
rect 5997 10251 6055 10257
rect 2188 10220 5948 10248
rect 2188 10208 2194 10220
rect 750 10180 756 10192
rect 663 10152 756 10180
rect 676 10121 704 10152
rect 750 10140 756 10152
rect 808 10180 814 10192
rect 1305 10183 1363 10189
rect 1305 10180 1317 10183
rect 808 10152 1317 10180
rect 808 10140 814 10152
rect 1305 10149 1317 10152
rect 1351 10180 1363 10183
rect 2682 10180 2688 10192
rect 1351 10152 2688 10180
rect 1351 10149 1363 10152
rect 1305 10143 1363 10149
rect 2682 10140 2688 10152
rect 2740 10140 2746 10192
rect 2866 10140 2872 10192
rect 2924 10180 2930 10192
rect 2924 10152 3174 10180
rect 2924 10140 2930 10152
rect 4706 10140 4712 10192
rect 4764 10180 4770 10192
rect 4982 10180 4988 10192
rect 4764 10152 4988 10180
rect 4764 10140 4770 10152
rect 4982 10140 4988 10152
rect 5040 10180 5046 10192
rect 5169 10183 5227 10189
rect 5169 10180 5181 10183
rect 5040 10152 5181 10180
rect 5040 10140 5046 10152
rect 5169 10149 5181 10152
rect 5215 10149 5227 10183
rect 5169 10143 5227 10149
rect 5445 10183 5503 10189
rect 5445 10149 5457 10183
rect 5491 10180 5503 10183
rect 5534 10180 5540 10192
rect 5491 10152 5540 10180
rect 5491 10149 5503 10152
rect 5445 10143 5503 10149
rect 661 10115 719 10121
rect 661 10081 673 10115
rect 707 10081 719 10115
rect 661 10075 719 10081
rect 2133 10115 2191 10121
rect 2133 10081 2145 10115
rect 2179 10112 2191 10115
rect 4890 10112 4896 10124
rect 2179 10084 3464 10112
rect 4851 10084 4896 10112
rect 2179 10081 2191 10084
rect 2133 10075 2191 10081
rect 937 10047 995 10053
rect 937 10013 949 10047
rect 983 10044 995 10047
rect 1854 10044 1860 10056
rect 983 10016 1860 10044
rect 983 10013 995 10016
rect 937 10007 995 10013
rect 1854 10004 1860 10016
rect 1912 10004 1918 10056
rect 2038 10044 2044 10056
rect 1999 10016 2044 10044
rect 2038 10004 2044 10016
rect 2096 10004 2102 10056
rect 2148 10016 3096 10044
rect 569 9979 627 9985
rect 569 9945 581 9979
rect 615 9976 627 9979
rect 2148 9976 2176 10016
rect 3068 9988 3096 10016
rect 615 9948 2176 9976
rect 2501 9979 2559 9985
rect 615 9945 627 9948
rect 569 9939 627 9945
rect 2501 9945 2513 9979
rect 2547 9976 2559 9979
rect 2958 9976 2964 9988
rect 2547 9948 2964 9976
rect 2547 9945 2559 9948
rect 2501 9939 2559 9945
rect 2958 9936 2964 9948
rect 3016 9936 3022 9988
rect 3050 9936 3056 9988
rect 3108 9936 3114 9988
rect 1394 9868 1400 9920
rect 1452 9908 1458 9920
rect 1581 9911 1639 9917
rect 1581 9908 1593 9911
rect 1452 9880 1593 9908
rect 1452 9868 1458 9880
rect 1581 9877 1593 9880
rect 1627 9908 1639 9911
rect 1946 9908 1952 9920
rect 1627 9880 1952 9908
rect 1627 9877 1639 9880
rect 1581 9871 1639 9877
rect 1946 9868 1952 9880
rect 2004 9868 2010 9920
rect 2731 9911 2789 9917
rect 2731 9877 2743 9911
rect 2777 9908 2789 9911
rect 3142 9908 3148 9920
rect 2777 9880 3148 9908
rect 2777 9877 2789 9880
rect 2731 9871 2789 9877
rect 3142 9868 3148 9880
rect 3200 9868 3206 9920
rect 3436 9908 3464 10084
rect 4890 10072 4896 10084
rect 4948 10072 4954 10124
rect 5184 10112 5212 10143
rect 5534 10140 5540 10152
rect 5592 10140 5598 10192
rect 5920 10180 5948 10220
rect 5997 10217 6009 10251
rect 6043 10248 6055 10251
rect 10134 10248 10140 10260
rect 6043 10220 10140 10248
rect 6043 10217 6055 10220
rect 5997 10211 6055 10217
rect 10134 10208 10140 10220
rect 10192 10208 10198 10260
rect 12986 10248 12992 10260
rect 10244 10220 12992 10248
rect 5920 10152 7420 10180
rect 5902 10112 5908 10124
rect 5184 10084 5908 10112
rect 5902 10072 5908 10084
rect 5960 10072 5966 10124
rect 7282 10112 7288 10124
rect 7243 10084 7288 10112
rect 7282 10072 7288 10084
rect 7340 10072 7346 10124
rect 7392 10112 7420 10152
rect 8202 10140 8208 10192
rect 8260 10140 8266 10192
rect 9490 10140 9496 10192
rect 9548 10180 9554 10192
rect 9548 10152 9996 10180
rect 9548 10140 9554 10152
rect 9858 10112 9864 10124
rect 7392 10084 7972 10112
rect 9819 10084 9864 10112
rect 4154 10044 4160 10056
rect 4115 10016 4160 10044
rect 4154 10004 4160 10016
rect 4212 10004 4218 10056
rect 4522 10044 4528 10056
rect 4483 10016 4528 10044
rect 4522 10004 4528 10016
rect 4580 10004 4586 10056
rect 4617 10047 4675 10053
rect 4617 10013 4629 10047
rect 4663 10044 4675 10047
rect 5166 10044 5172 10056
rect 4663 10016 5172 10044
rect 4663 10013 4675 10016
rect 4617 10007 4675 10013
rect 5166 10004 5172 10016
rect 5224 10004 5230 10056
rect 7466 10044 7472 10056
rect 7427 10016 7472 10044
rect 7466 10004 7472 10016
rect 7524 10004 7530 10056
rect 7834 10044 7840 10056
rect 7795 10016 7840 10044
rect 7834 10004 7840 10016
rect 7892 10004 7898 10056
rect 7944 10044 7972 10084
rect 9858 10072 9864 10084
rect 9916 10072 9922 10124
rect 9968 10121 9996 10152
rect 10244 10121 10272 10220
rect 12986 10208 12992 10220
rect 13044 10208 13050 10260
rect 15562 10208 15568 10260
rect 15620 10248 15626 10260
rect 17405 10251 17463 10257
rect 17405 10248 17417 10251
rect 15620 10220 17417 10248
rect 15620 10208 15626 10220
rect 17405 10217 17417 10220
rect 17451 10217 17463 10251
rect 17405 10211 17463 10217
rect 17494 10208 17500 10260
rect 17552 10248 17558 10260
rect 17865 10251 17923 10257
rect 17552 10220 17597 10248
rect 17552 10208 17558 10220
rect 17865 10217 17877 10251
rect 17911 10217 17923 10251
rect 17865 10211 17923 10217
rect 9953 10115 10011 10121
rect 9953 10081 9965 10115
rect 9999 10081 10011 10115
rect 9953 10075 10011 10081
rect 10229 10115 10287 10121
rect 10229 10081 10241 10115
rect 10275 10081 10287 10115
rect 11624 10112 11652 10166
rect 11882 10140 11888 10192
rect 11940 10180 11946 10192
rect 12023 10183 12081 10189
rect 12023 10180 12035 10183
rect 11940 10152 12035 10180
rect 11940 10140 11946 10152
rect 12023 10149 12035 10152
rect 12069 10149 12081 10183
rect 14642 10180 14648 10192
rect 14030 10152 14648 10180
rect 12023 10143 12081 10149
rect 14642 10140 14648 10152
rect 14700 10140 14706 10192
rect 15930 10140 15936 10192
rect 15988 10180 15994 10192
rect 16393 10183 16451 10189
rect 16393 10180 16405 10183
rect 15988 10152 16405 10180
rect 15988 10140 15994 10152
rect 16393 10149 16405 10152
rect 16439 10149 16451 10183
rect 16393 10143 16451 10149
rect 16482 10140 16488 10192
rect 16540 10180 16546 10192
rect 16577 10183 16635 10189
rect 16577 10180 16589 10183
rect 16540 10152 16589 10180
rect 16540 10140 16546 10152
rect 16577 10149 16589 10152
rect 16623 10149 16635 10183
rect 17880 10180 17908 10211
rect 18138 10180 18144 10192
rect 16577 10143 16635 10149
rect 16868 10152 17908 10180
rect 18099 10152 18144 10180
rect 12250 10112 12256 10124
rect 11624 10084 12256 10112
rect 10229 10075 10287 10081
rect 12250 10072 12256 10084
rect 12308 10072 12314 10124
rect 12434 10072 12440 10124
rect 12492 10112 12498 10124
rect 12492 10084 13124 10112
rect 12492 10072 12498 10084
rect 9674 10044 9680 10056
rect 7944 10016 9680 10044
rect 9674 10004 9680 10016
rect 9732 10004 9738 10056
rect 10134 10044 10140 10056
rect 10095 10016 10140 10044
rect 10134 10004 10140 10016
rect 10192 10004 10198 10056
rect 10597 10047 10655 10053
rect 10597 10044 10609 10047
rect 10244 10016 10609 10044
rect 4709 9979 4767 9985
rect 4709 9945 4721 9979
rect 4755 9976 4767 9979
rect 4982 9976 4988 9988
rect 4755 9948 4988 9976
rect 4755 9945 4767 9948
rect 4709 9939 4767 9945
rect 4982 9936 4988 9948
rect 5040 9936 5046 9988
rect 9263 9979 9321 9985
rect 9263 9945 9275 9979
rect 9309 9976 9321 9979
rect 10244 9976 10272 10016
rect 10597 10013 10609 10016
rect 10643 10013 10655 10047
rect 10597 10007 10655 10013
rect 11330 10004 11336 10056
rect 11388 10044 11394 10056
rect 12621 10047 12679 10053
rect 12621 10044 12633 10047
rect 11388 10016 12633 10044
rect 11388 10004 11394 10016
rect 12621 10013 12633 10016
rect 12667 10013 12679 10047
rect 12986 10044 12992 10056
rect 12947 10016 12992 10044
rect 12621 10007 12679 10013
rect 12986 10004 12992 10016
rect 13044 10004 13050 10056
rect 13096 10044 13124 10084
rect 15010 10072 15016 10124
rect 15068 10112 15074 10124
rect 15654 10112 15660 10124
rect 15068 10084 15660 10112
rect 15068 10072 15074 10084
rect 15654 10072 15660 10084
rect 15712 10072 15718 10124
rect 16868 10121 16896 10152
rect 18138 10140 18144 10152
rect 18196 10140 18202 10192
rect 16669 10115 16727 10121
rect 16669 10081 16681 10115
rect 16715 10081 16727 10115
rect 16669 10075 16727 10081
rect 16853 10115 16911 10121
rect 16853 10081 16865 10115
rect 16899 10081 16911 10115
rect 16853 10075 16911 10081
rect 16206 10044 16212 10056
rect 13096 10016 16212 10044
rect 16206 10004 16212 10016
rect 16264 10004 16270 10056
rect 9309 9948 10272 9976
rect 9309 9945 9321 9948
rect 9263 9939 9321 9945
rect 11790 9936 11796 9988
rect 11848 9976 11854 9988
rect 12437 9979 12495 9985
rect 12437 9976 12449 9979
rect 11848 9948 12449 9976
rect 11848 9936 11854 9948
rect 12437 9945 12449 9948
rect 12483 9945 12495 9979
rect 16684 9976 16712 10075
rect 17494 10072 17500 10124
rect 17552 10112 17558 10124
rect 17862 10112 17868 10124
rect 17552 10084 17868 10112
rect 17552 10072 17558 10084
rect 17862 10072 17868 10084
rect 17920 10112 17926 10124
rect 18049 10115 18107 10121
rect 18049 10112 18061 10115
rect 17920 10084 18061 10112
rect 17920 10072 17926 10084
rect 18049 10081 18061 10084
rect 18095 10081 18107 10115
rect 18230 10112 18236 10124
rect 18191 10084 18236 10112
rect 18049 10075 18107 10081
rect 18230 10072 18236 10084
rect 18288 10072 18294 10124
rect 18322 10072 18328 10124
rect 18380 10112 18386 10124
rect 18380 10084 18425 10112
rect 18380 10072 18386 10084
rect 17681 10047 17739 10053
rect 17681 10013 17693 10047
rect 17727 10044 17739 10047
rect 17727 10016 18092 10044
rect 17727 10013 17739 10016
rect 17681 10007 17739 10013
rect 17862 9976 17868 9988
rect 16684 9948 17868 9976
rect 12437 9939 12495 9945
rect 17862 9936 17868 9948
rect 17920 9936 17926 9988
rect 18064 9976 18092 10016
rect 18322 9976 18328 9988
rect 18064 9948 18328 9976
rect 18322 9936 18328 9948
rect 18380 9936 18386 9988
rect 4614 9908 4620 9920
rect 3436 9880 4620 9908
rect 4614 9868 4620 9880
rect 4672 9868 4678 9920
rect 4801 9911 4859 9917
rect 4801 9877 4813 9911
rect 4847 9908 4859 9911
rect 5350 9908 5356 9920
rect 4847 9880 5356 9908
rect 4847 9877 4859 9880
rect 4801 9871 4859 9877
rect 5350 9868 5356 9880
rect 5408 9868 5414 9920
rect 7834 9868 7840 9920
rect 7892 9908 7898 9920
rect 8386 9908 8392 9920
rect 7892 9880 8392 9908
rect 7892 9868 7898 9880
rect 8386 9868 8392 9880
rect 8444 9868 8450 9920
rect 8662 9868 8668 9920
rect 8720 9908 8726 9920
rect 9493 9911 9551 9917
rect 9493 9908 9505 9911
rect 8720 9880 9505 9908
rect 8720 9868 8726 9880
rect 9493 9877 9505 9880
rect 9539 9908 9551 9911
rect 9582 9908 9588 9920
rect 9539 9880 9588 9908
rect 9539 9877 9551 9880
rect 9493 9871 9551 9877
rect 9582 9868 9588 9880
rect 9640 9868 9646 9920
rect 10045 9911 10103 9917
rect 10045 9877 10057 9911
rect 10091 9908 10103 9911
rect 10226 9908 10232 9920
rect 10091 9880 10232 9908
rect 10091 9877 10103 9880
rect 10045 9871 10103 9877
rect 10226 9868 10232 9880
rect 10284 9868 10290 9920
rect 10778 9868 10784 9920
rect 10836 9908 10842 9920
rect 12158 9908 12164 9920
rect 10836 9880 12164 9908
rect 10836 9868 10842 9880
rect 12158 9868 12164 9880
rect 12216 9868 12222 9920
rect 12250 9868 12256 9920
rect 12308 9908 12314 9920
rect 14415 9911 14473 9917
rect 12308 9880 12353 9908
rect 12308 9868 12314 9880
rect 14415 9877 14427 9911
rect 14461 9908 14473 9911
rect 14918 9908 14924 9920
rect 14461 9880 14924 9908
rect 14461 9877 14473 9880
rect 14415 9871 14473 9877
rect 14918 9868 14924 9880
rect 14976 9868 14982 9920
rect 15105 9911 15163 9917
rect 15105 9877 15117 9911
rect 15151 9908 15163 9911
rect 15838 9908 15844 9920
rect 15151 9880 15844 9908
rect 15151 9877 15163 9880
rect 15105 9871 15163 9877
rect 15838 9868 15844 9880
rect 15896 9868 15902 9920
rect 16758 9908 16764 9920
rect 16719 9880 16764 9908
rect 16758 9868 16764 9880
rect 16816 9868 16822 9920
rect 16850 9868 16856 9920
rect 16908 9908 16914 9920
rect 17037 9911 17095 9917
rect 17037 9908 17049 9911
rect 16908 9880 17049 9908
rect 16908 9868 16914 9880
rect 17037 9877 17049 9880
rect 17083 9877 17095 9911
rect 17037 9871 17095 9877
rect 17954 9868 17960 9920
rect 18012 9908 18018 9920
rect 18230 9908 18236 9920
rect 18012 9880 18236 9908
rect 18012 9868 18018 9880
rect 18230 9868 18236 9880
rect 18288 9868 18294 9920
rect 184 9818 18924 9840
rect 184 9766 3110 9818
rect 3162 9766 3174 9818
rect 3226 9766 3238 9818
rect 3290 9766 3302 9818
rect 3354 9766 3366 9818
rect 3418 9766 6210 9818
rect 6262 9766 6274 9818
rect 6326 9766 6338 9818
rect 6390 9766 6402 9818
rect 6454 9766 6466 9818
rect 6518 9766 9310 9818
rect 9362 9766 9374 9818
rect 9426 9766 9438 9818
rect 9490 9766 9502 9818
rect 9554 9766 9566 9818
rect 9618 9766 12410 9818
rect 12462 9766 12474 9818
rect 12526 9766 12538 9818
rect 12590 9766 12602 9818
rect 12654 9766 12666 9818
rect 12718 9766 15510 9818
rect 15562 9766 15574 9818
rect 15626 9766 15638 9818
rect 15690 9766 15702 9818
rect 15754 9766 15766 9818
rect 15818 9766 18610 9818
rect 18662 9766 18674 9818
rect 18726 9766 18738 9818
rect 18790 9766 18802 9818
rect 18854 9766 18866 9818
rect 18918 9766 18924 9818
rect 184 9744 18924 9766
rect 3973 9707 4031 9713
rect 3973 9673 3985 9707
rect 4019 9704 4031 9707
rect 4154 9704 4160 9716
rect 4019 9676 4160 9704
rect 4019 9673 4031 9676
rect 3973 9667 4031 9673
rect 4154 9664 4160 9676
rect 4212 9664 4218 9716
rect 4338 9704 4344 9716
rect 4299 9676 4344 9704
rect 4338 9664 4344 9676
rect 4396 9664 4402 9716
rect 4522 9664 4528 9716
rect 4580 9664 4586 9716
rect 4614 9664 4620 9716
rect 4672 9704 4678 9716
rect 5074 9704 5080 9716
rect 4672 9676 5080 9704
rect 4672 9664 4678 9676
rect 5074 9664 5080 9676
rect 5132 9704 5138 9716
rect 5825 9707 5883 9713
rect 5825 9704 5837 9707
rect 5132 9676 5837 9704
rect 5132 9664 5138 9676
rect 5825 9673 5837 9676
rect 5871 9673 5883 9707
rect 5825 9667 5883 9673
rect 6086 9664 6092 9716
rect 6144 9704 6150 9716
rect 6273 9707 6331 9713
rect 6273 9704 6285 9707
rect 6144 9676 6285 9704
rect 6144 9664 6150 9676
rect 6273 9673 6285 9676
rect 6319 9673 6331 9707
rect 6273 9667 6331 9673
rect 7282 9664 7288 9716
rect 7340 9704 7346 9716
rect 13538 9704 13544 9716
rect 7340 9676 13544 9704
rect 7340 9664 7346 9676
rect 13538 9664 13544 9676
rect 13596 9664 13602 9716
rect 15286 9664 15292 9716
rect 15344 9704 15350 9716
rect 15933 9707 15991 9713
rect 15933 9704 15945 9707
rect 15344 9676 15945 9704
rect 15344 9664 15350 9676
rect 15933 9673 15945 9676
rect 15979 9673 15991 9707
rect 16114 9704 16120 9716
rect 15933 9667 15991 9673
rect 16040 9676 16120 9704
rect 1486 9636 1492 9648
rect 768 9608 1492 9636
rect 768 9577 796 9608
rect 1486 9596 1492 9608
rect 1544 9596 1550 9648
rect 3605 9639 3663 9645
rect 3605 9605 3617 9639
rect 3651 9636 3663 9639
rect 4540 9636 4568 9664
rect 3651 9608 4568 9636
rect 3651 9605 3663 9608
rect 3605 9599 3663 9605
rect 8386 9596 8392 9648
rect 8444 9645 8450 9648
rect 8444 9639 8493 9645
rect 8444 9605 8447 9639
rect 8481 9605 8493 9639
rect 8662 9636 8668 9648
rect 8623 9608 8668 9636
rect 8444 9599 8493 9605
rect 8444 9596 8450 9599
rect 8662 9596 8668 9608
rect 8720 9596 8726 9648
rect 8754 9596 8760 9648
rect 8812 9636 8818 9648
rect 10594 9636 10600 9648
rect 8812 9608 8984 9636
rect 10555 9608 10600 9636
rect 8812 9596 8818 9608
rect 753 9571 811 9577
rect 753 9537 765 9571
rect 799 9537 811 9571
rect 753 9531 811 9537
rect 1504 9540 3648 9568
rect 474 9500 480 9512
rect 435 9472 480 9500
rect 474 9460 480 9472
rect 532 9460 538 9512
rect 569 9503 627 9509
rect 569 9469 581 9503
rect 615 9500 627 9503
rect 1026 9500 1032 9512
rect 615 9472 888 9500
rect 987 9472 1032 9500
rect 615 9469 627 9472
rect 569 9463 627 9469
rect 658 9392 664 9444
rect 716 9432 722 9444
rect 753 9435 811 9441
rect 753 9432 765 9435
rect 716 9404 765 9432
rect 716 9392 722 9404
rect 753 9401 765 9404
rect 799 9401 811 9435
rect 860 9432 888 9472
rect 1026 9460 1032 9472
rect 1084 9460 1090 9512
rect 1118 9460 1124 9512
rect 1176 9494 1182 9512
rect 1249 9503 1307 9509
rect 1249 9500 1261 9503
rect 1176 9466 1215 9494
rect 1246 9469 1261 9500
rect 1295 9469 1307 9503
rect 1176 9460 1182 9466
rect 1246 9463 1307 9469
rect 1121 9457 1179 9460
rect 860 9404 980 9432
rect 753 9395 811 9401
rect 952 9376 980 9404
rect 842 9364 848 9376
rect 803 9336 848 9364
rect 842 9324 848 9336
rect 900 9324 906 9376
rect 934 9324 940 9376
rect 992 9324 998 9376
rect 1246 9364 1274 9463
rect 1394 9460 1400 9512
rect 1452 9500 1458 9512
rect 1504 9509 1532 9540
rect 3620 9509 3648 9540
rect 3694 9528 3700 9580
rect 3752 9568 3758 9580
rect 3881 9571 3939 9577
rect 3881 9568 3893 9571
rect 3752 9540 3893 9568
rect 3752 9528 3758 9540
rect 3881 9537 3893 9540
rect 3927 9537 3939 9571
rect 5718 9568 5724 9580
rect 3881 9531 3939 9537
rect 3988 9540 5724 9568
rect 1489 9503 1547 9509
rect 1489 9500 1501 9503
rect 1452 9472 1501 9500
rect 1452 9460 1458 9472
rect 1489 9469 1501 9472
rect 1535 9469 1547 9503
rect 1489 9463 1547 9469
rect 3605 9503 3663 9509
rect 3605 9469 3617 9503
rect 3651 9500 3663 9503
rect 3988 9500 4016 9540
rect 5718 9528 5724 9540
rect 5776 9528 5782 9580
rect 6089 9571 6147 9577
rect 6089 9537 6101 9571
rect 6135 9568 6147 9571
rect 8202 9568 8208 9580
rect 6135 9540 8208 9568
rect 6135 9537 6147 9540
rect 6089 9531 6147 9537
rect 8202 9528 8208 9540
rect 8260 9568 8266 9580
rect 8849 9571 8907 9577
rect 8849 9568 8861 9571
rect 8260 9540 8861 9568
rect 8260 9528 8266 9540
rect 8849 9537 8861 9540
rect 8895 9537 8907 9571
rect 8956 9568 8984 9608
rect 10594 9596 10600 9608
rect 10652 9596 10658 9648
rect 10778 9636 10784 9648
rect 10739 9608 10784 9636
rect 10778 9596 10784 9608
rect 10836 9596 10842 9648
rect 12986 9596 12992 9648
rect 13044 9636 13050 9648
rect 13127 9639 13185 9645
rect 13127 9636 13139 9639
rect 13044 9608 13139 9636
rect 13044 9596 13050 9608
rect 13127 9605 13139 9608
rect 13173 9605 13185 9639
rect 13127 9599 13185 9605
rect 15381 9639 15439 9645
rect 15381 9605 15393 9639
rect 15427 9636 15439 9639
rect 16040 9636 16068 9676
rect 16114 9664 16120 9676
rect 16172 9704 16178 9716
rect 16482 9704 16488 9716
rect 16172 9676 16488 9704
rect 16172 9664 16178 9676
rect 16482 9664 16488 9676
rect 16540 9664 16546 9716
rect 18230 9664 18236 9716
rect 18288 9704 18294 9716
rect 18417 9707 18475 9713
rect 18417 9704 18429 9707
rect 18288 9676 18429 9704
rect 18288 9664 18294 9676
rect 18417 9673 18429 9676
rect 18463 9673 18475 9707
rect 18417 9667 18475 9673
rect 15427 9608 16068 9636
rect 15427 9605 15439 9608
rect 15381 9599 15439 9605
rect 17862 9596 17868 9648
rect 17920 9636 17926 9648
rect 18325 9639 18383 9645
rect 18325 9636 18337 9639
rect 17920 9608 18337 9636
rect 17920 9596 17926 9608
rect 18325 9605 18337 9608
rect 18371 9605 18383 9639
rect 18325 9599 18383 9605
rect 9125 9571 9183 9577
rect 9125 9568 9137 9571
rect 8956 9540 9137 9568
rect 8849 9531 8907 9537
rect 9125 9537 9137 9540
rect 9171 9568 9183 9571
rect 9490 9568 9496 9580
rect 9171 9540 9496 9568
rect 9171 9537 9183 9540
rect 9125 9531 9183 9537
rect 9490 9528 9496 9540
rect 9548 9528 9554 9580
rect 9858 9528 9864 9580
rect 9916 9568 9922 9580
rect 10796 9568 10824 9596
rect 9916 9540 10824 9568
rect 11701 9571 11759 9577
rect 9916 9528 9922 9540
rect 11701 9537 11713 9571
rect 11747 9568 11759 9571
rect 11747 9540 14780 9568
rect 11747 9537 11759 9540
rect 11701 9531 11759 9537
rect 3651 9472 4016 9500
rect 4065 9503 4123 9509
rect 3651 9469 3663 9472
rect 3605 9463 3663 9469
rect 4065 9469 4077 9503
rect 4111 9469 4123 9503
rect 4065 9463 4123 9469
rect 1762 9432 1768 9444
rect 1723 9404 1768 9432
rect 1762 9392 1768 9404
rect 1820 9392 1826 9444
rect 3050 9432 3056 9444
rect 2990 9404 3056 9432
rect 3050 9392 3056 9404
rect 3108 9392 3114 9444
rect 3786 9392 3792 9444
rect 3844 9432 3850 9444
rect 4080 9432 4108 9463
rect 4154 9460 4160 9512
rect 4212 9500 4218 9512
rect 4212 9472 4257 9500
rect 4212 9460 4218 9472
rect 6546 9460 6552 9512
rect 6604 9500 6610 9512
rect 6641 9503 6699 9509
rect 6641 9500 6653 9503
rect 6604 9472 6653 9500
rect 6604 9460 6610 9472
rect 6641 9469 6653 9472
rect 6687 9469 6699 9503
rect 7006 9500 7012 9512
rect 6967 9472 7012 9500
rect 6641 9463 6699 9469
rect 7006 9460 7012 9472
rect 7064 9460 7070 9512
rect 10873 9503 10931 9509
rect 10873 9469 10885 9503
rect 10919 9469 10931 9503
rect 11330 9500 11336 9512
rect 11291 9472 11336 9500
rect 10873 9463 10931 9469
rect 3844 9404 4108 9432
rect 3844 9392 3850 9404
rect 5258 9392 5264 9444
rect 5316 9392 5322 9444
rect 7374 9432 7380 9444
rect 7300 9404 7380 9432
rect 2130 9364 2136 9376
rect 1246 9336 2136 9364
rect 2130 9324 2136 9336
rect 2188 9324 2194 9376
rect 3237 9367 3295 9373
rect 3237 9333 3249 9367
rect 3283 9364 3295 9367
rect 3602 9364 3608 9376
rect 3283 9336 3608 9364
rect 3283 9333 3295 9336
rect 3237 9327 3295 9333
rect 3602 9324 3608 9336
rect 3660 9324 3666 9376
rect 6549 9367 6607 9373
rect 6549 9333 6561 9367
rect 6595 9364 6607 9367
rect 6638 9364 6644 9376
rect 6595 9336 6644 9364
rect 6595 9333 6607 9336
rect 6549 9327 6607 9333
rect 6638 9324 6644 9336
rect 6696 9324 6702 9376
rect 6914 9324 6920 9376
rect 6972 9364 6978 9376
rect 7300 9364 7328 9404
rect 7374 9392 7380 9404
rect 7432 9392 7438 9444
rect 10410 9432 10416 9444
rect 10323 9404 10416 9432
rect 10410 9392 10416 9404
rect 10468 9432 10474 9444
rect 10888 9432 10916 9463
rect 11330 9460 11336 9472
rect 11388 9460 11394 9512
rect 13446 9500 13452 9512
rect 13407 9472 13452 9500
rect 13446 9460 13452 9472
rect 13504 9460 13510 9512
rect 11238 9432 11244 9444
rect 10468 9404 10824 9432
rect 10888 9404 11244 9432
rect 10468 9392 10474 9404
rect 10796 9376 10824 9404
rect 11238 9392 11244 9404
rect 11296 9392 11302 9444
rect 14642 9432 14648 9444
rect 12742 9404 14648 9432
rect 8294 9364 8300 9376
rect 6972 9336 8300 9364
rect 6972 9324 6978 9336
rect 8294 9324 8300 9336
rect 8352 9324 8358 9376
rect 9490 9324 9496 9376
rect 9548 9364 9554 9376
rect 9858 9364 9864 9376
rect 9548 9336 9864 9364
rect 9548 9324 9554 9336
rect 9858 9324 9864 9336
rect 9916 9324 9922 9376
rect 10778 9324 10784 9376
rect 10836 9364 10842 9376
rect 11149 9367 11207 9373
rect 11149 9364 11161 9367
rect 10836 9336 11161 9364
rect 10836 9324 10842 9336
rect 11149 9333 11161 9336
rect 11195 9364 11207 9367
rect 12250 9364 12256 9376
rect 11195 9336 12256 9364
rect 11195 9333 11207 9336
rect 11149 9327 11207 9333
rect 12250 9324 12256 9336
rect 12308 9364 12314 9376
rect 12820 9364 12848 9404
rect 14642 9392 14648 9404
rect 14700 9392 14706 9444
rect 14752 9432 14780 9540
rect 14826 9528 14832 9580
rect 14884 9568 14890 9580
rect 16209 9571 16267 9577
rect 16209 9568 16221 9571
rect 14884 9540 16221 9568
rect 14884 9528 14890 9540
rect 16209 9537 16221 9540
rect 16255 9537 16267 9571
rect 16209 9531 16267 9537
rect 16577 9571 16635 9577
rect 16577 9537 16589 9571
rect 16623 9568 16635 9571
rect 16758 9568 16764 9580
rect 16623 9540 16764 9568
rect 16623 9537 16635 9540
rect 16577 9531 16635 9537
rect 16758 9528 16764 9540
rect 16816 9528 16822 9580
rect 17586 9528 17592 9580
rect 17644 9528 17650 9580
rect 17770 9528 17776 9580
rect 17828 9568 17834 9580
rect 18003 9571 18061 9577
rect 18003 9568 18015 9571
rect 17828 9540 18015 9568
rect 17828 9528 17834 9540
rect 18003 9537 18015 9540
rect 18049 9568 18061 9571
rect 18233 9571 18291 9577
rect 18233 9568 18245 9571
rect 18049 9540 18245 9568
rect 18049 9537 18061 9540
rect 18003 9531 18061 9537
rect 18233 9537 18245 9540
rect 18279 9537 18291 9571
rect 18233 9531 18291 9537
rect 15194 9460 15200 9512
rect 15252 9500 15258 9512
rect 15473 9503 15531 9509
rect 15473 9500 15485 9503
rect 15252 9472 15485 9500
rect 15252 9460 15258 9472
rect 15473 9469 15485 9472
rect 15519 9469 15531 9503
rect 15473 9463 15531 9469
rect 16117 9503 16175 9509
rect 16117 9469 16129 9503
rect 16163 9500 16175 9503
rect 16666 9500 16672 9512
rect 16163 9472 16672 9500
rect 16163 9469 16175 9472
rect 16117 9463 16175 9469
rect 16666 9460 16672 9472
rect 16724 9460 16730 9512
rect 17402 9460 17408 9512
rect 17460 9500 17466 9512
rect 17604 9500 17632 9528
rect 18509 9503 18567 9509
rect 18509 9500 18521 9503
rect 17460 9472 18521 9500
rect 17460 9460 17466 9472
rect 18509 9469 18521 9472
rect 18555 9469 18567 9503
rect 18509 9463 18567 9469
rect 17770 9432 17776 9444
rect 14752 9404 16344 9432
rect 17618 9404 17776 9432
rect 14734 9364 14740 9376
rect 12308 9336 12848 9364
rect 14695 9336 14740 9364
rect 12308 9324 12314 9336
rect 14734 9324 14740 9336
rect 14792 9324 14798 9376
rect 15657 9367 15715 9373
rect 15657 9333 15669 9367
rect 15703 9364 15715 9367
rect 16022 9364 16028 9376
rect 15703 9336 16028 9364
rect 15703 9333 15715 9336
rect 15657 9327 15715 9333
rect 16022 9324 16028 9336
rect 16080 9324 16086 9376
rect 16316 9364 16344 9404
rect 17770 9392 17776 9404
rect 17828 9392 17834 9444
rect 18046 9364 18052 9376
rect 16316 9336 18052 9364
rect 18046 9324 18052 9336
rect 18104 9324 18110 9376
rect 184 9274 18860 9296
rect 184 9222 4660 9274
rect 4712 9222 4724 9274
rect 4776 9222 4788 9274
rect 4840 9222 4852 9274
rect 4904 9222 4916 9274
rect 4968 9222 7760 9274
rect 7812 9222 7824 9274
rect 7876 9222 7888 9274
rect 7940 9222 7952 9274
rect 8004 9222 8016 9274
rect 8068 9222 10860 9274
rect 10912 9222 10924 9274
rect 10976 9222 10988 9274
rect 11040 9222 11052 9274
rect 11104 9222 11116 9274
rect 11168 9222 13960 9274
rect 14012 9222 14024 9274
rect 14076 9222 14088 9274
rect 14140 9222 14152 9274
rect 14204 9222 14216 9274
rect 14268 9222 17060 9274
rect 17112 9222 17124 9274
rect 17176 9222 17188 9274
rect 17240 9222 17252 9274
rect 17304 9222 17316 9274
rect 17368 9222 18860 9274
rect 184 9200 18860 9222
rect 1670 9120 1676 9172
rect 1728 9160 1734 9172
rect 1765 9163 1823 9169
rect 1765 9160 1777 9163
rect 1728 9132 1777 9160
rect 1728 9120 1734 9132
rect 1765 9129 1777 9132
rect 1811 9129 1823 9163
rect 3694 9160 3700 9172
rect 1765 9123 1823 9129
rect 1872 9132 3700 9160
rect 1029 9095 1087 9101
rect 1029 9061 1041 9095
rect 1075 9092 1087 9095
rect 1872 9092 1900 9132
rect 3694 9120 3700 9132
rect 3752 9120 3758 9172
rect 4430 9120 4436 9172
rect 4488 9160 4494 9172
rect 5077 9163 5135 9169
rect 5077 9160 5089 9163
rect 4488 9132 5089 9160
rect 4488 9120 4494 9132
rect 5077 9129 5089 9132
rect 5123 9160 5135 9163
rect 8662 9160 8668 9172
rect 5123 9132 8668 9160
rect 5123 9129 5135 9132
rect 5077 9123 5135 9129
rect 8662 9120 8668 9132
rect 8720 9120 8726 9172
rect 11422 9120 11428 9172
rect 11480 9160 11486 9172
rect 11793 9163 11851 9169
rect 11793 9160 11805 9163
rect 11480 9132 11805 9160
rect 11480 9120 11486 9132
rect 11793 9129 11805 9132
rect 11839 9129 11851 9163
rect 13538 9160 13544 9172
rect 13499 9132 13544 9160
rect 11793 9123 11851 9129
rect 13538 9120 13544 9132
rect 13596 9120 13602 9172
rect 14642 9120 14648 9172
rect 14700 9160 14706 9172
rect 14700 9132 16344 9160
rect 14700 9120 14706 9132
rect 1075 9064 1900 9092
rect 1075 9061 1087 9064
rect 1029 9055 1087 9061
rect 2038 9052 2044 9104
rect 2096 9092 2102 9104
rect 2777 9095 2835 9101
rect 2777 9092 2789 9095
rect 2096 9064 2789 9092
rect 2096 9052 2102 9064
rect 2777 9061 2789 9064
rect 2823 9061 2835 9095
rect 2777 9055 2835 9061
rect 2866 9052 2872 9104
rect 2924 9092 2930 9104
rect 3050 9092 3056 9104
rect 2924 9064 3056 9092
rect 2924 9052 2930 9064
rect 3050 9052 3056 9064
rect 3108 9092 3114 9104
rect 5258 9092 5264 9104
rect 3108 9064 5264 9092
rect 3108 9052 3114 9064
rect 5258 9052 5264 9064
rect 5316 9052 5322 9104
rect 6822 9052 6828 9104
rect 6880 9092 6886 9104
rect 7466 9092 7472 9104
rect 6880 9064 7328 9092
rect 7427 9064 7472 9092
rect 6880 9052 6886 9064
rect 566 8984 572 9036
rect 624 9033 630 9036
rect 624 9027 683 9033
rect 624 8993 637 9027
rect 671 8993 683 9027
rect 750 9024 756 9036
rect 711 8996 756 9024
rect 624 8987 683 8993
rect 624 8984 630 8987
rect 750 8984 756 8996
rect 808 8984 814 9036
rect 845 9027 903 9033
rect 845 8993 857 9027
rect 891 9024 903 9027
rect 1210 9024 1216 9036
rect 891 8996 1072 9024
rect 1171 8996 1216 9024
rect 891 8993 903 8996
rect 845 8987 903 8993
rect 1044 8968 1072 8996
rect 1210 8984 1216 8996
rect 1268 8984 1274 9036
rect 2130 9024 2136 9036
rect 2091 8996 2136 9024
rect 2130 8984 2136 8996
rect 2188 8984 2194 9036
rect 2225 9027 2283 9033
rect 2225 8993 2237 9027
rect 2271 9024 2283 9027
rect 2682 9024 2688 9036
rect 2271 8996 2688 9024
rect 2271 8993 2283 8996
rect 2225 8987 2283 8993
rect 2682 8984 2688 8996
rect 2740 8984 2746 9036
rect 4430 9024 4436 9036
rect 4391 8996 4436 9024
rect 4430 8984 4436 8996
rect 4488 8984 4494 9036
rect 4709 9027 4767 9033
rect 4709 8993 4721 9027
rect 4755 8993 4767 9027
rect 4709 8987 4767 8993
rect 4893 9027 4951 9033
rect 4893 8993 4905 9027
rect 4939 9024 4951 9027
rect 4982 9024 4988 9036
rect 4939 8996 4988 9024
rect 4939 8993 4951 8996
rect 4893 8987 4951 8993
rect 1026 8916 1032 8968
rect 1084 8916 1090 8968
rect 2314 8956 2320 8968
rect 2275 8928 2320 8956
rect 2314 8916 2320 8928
rect 2372 8916 2378 8968
rect 3694 8916 3700 8968
rect 3752 8956 3758 8968
rect 4724 8956 4752 8987
rect 4982 8984 4988 8996
rect 5040 8984 5046 9036
rect 7300 9033 7328 9064
rect 7466 9052 7472 9064
rect 7524 9052 7530 9104
rect 9677 9095 9735 9101
rect 9677 9061 9689 9095
rect 9723 9092 9735 9095
rect 9950 9092 9956 9104
rect 9723 9064 9956 9092
rect 9723 9061 9735 9064
rect 9677 9055 9735 9061
rect 9950 9052 9956 9064
rect 10008 9052 10014 9104
rect 10778 9052 10784 9104
rect 10836 9052 10842 9104
rect 11514 9052 11520 9104
rect 11572 9092 11578 9104
rect 12253 9095 12311 9101
rect 12253 9092 12265 9095
rect 11572 9064 12265 9092
rect 11572 9052 11578 9064
rect 12253 9061 12265 9064
rect 12299 9061 12311 9095
rect 16316 9092 16344 9132
rect 17770 9092 17776 9104
rect 16238 9064 17776 9092
rect 12253 9055 12311 9061
rect 17770 9052 17776 9064
rect 17828 9052 17834 9104
rect 7009 9027 7067 9033
rect 7009 8993 7021 9027
rect 7055 8993 7067 9027
rect 7009 8987 7067 8993
rect 7285 9027 7343 9033
rect 7285 8993 7297 9027
rect 7331 9024 7343 9027
rect 7650 9024 7656 9036
rect 7331 8996 7656 9024
rect 7331 8993 7343 8996
rect 7285 8987 7343 8993
rect 3752 8928 4752 8956
rect 3752 8916 3758 8928
rect 1581 8891 1639 8897
rect 1581 8857 1593 8891
rect 1627 8888 1639 8891
rect 4062 8888 4068 8900
rect 1627 8860 4068 8888
rect 1627 8857 1639 8860
rect 1581 8851 1639 8857
rect 4062 8848 4068 8860
rect 4120 8848 4126 8900
rect 4154 8848 4160 8900
rect 4212 8888 4218 8900
rect 4801 8891 4859 8897
rect 4801 8888 4813 8891
rect 4212 8860 4813 8888
rect 4212 8848 4218 8860
rect 4801 8857 4813 8860
rect 4847 8857 4859 8891
rect 7024 8888 7052 8987
rect 7650 8984 7656 8996
rect 7708 8984 7714 9036
rect 7834 9024 7840 9036
rect 7795 8996 7840 9024
rect 7834 8984 7840 8996
rect 7892 8984 7898 9036
rect 9861 9027 9919 9033
rect 9861 8993 9873 9027
rect 9907 9024 9919 9027
rect 9907 8996 10364 9024
rect 9907 8993 9919 8996
rect 9861 8987 9919 8993
rect 7926 8956 7932 8968
rect 7887 8928 7932 8956
rect 7926 8916 7932 8928
rect 7984 8916 7990 8968
rect 10226 8956 10232 8968
rect 10187 8928 10232 8956
rect 10226 8916 10232 8928
rect 10284 8916 10290 8968
rect 10336 8956 10364 8996
rect 11670 8996 12020 9024
rect 10336 8928 11192 8956
rect 11164 8888 11192 8928
rect 11238 8916 11244 8968
rect 11296 8956 11302 8968
rect 11670 8965 11698 8996
rect 11655 8959 11713 8965
rect 11655 8956 11667 8959
rect 11296 8928 11667 8956
rect 11296 8916 11302 8928
rect 11655 8925 11667 8928
rect 11701 8925 11713 8959
rect 11655 8919 11713 8925
rect 11793 8959 11851 8965
rect 11793 8925 11805 8959
rect 11839 8956 11851 8959
rect 11882 8956 11888 8968
rect 11839 8928 11888 8956
rect 11839 8925 11851 8928
rect 11793 8919 11851 8925
rect 11882 8916 11888 8928
rect 11940 8916 11946 8968
rect 11992 8956 12020 8996
rect 12066 8984 12072 9036
rect 12124 9024 12130 9036
rect 14461 9027 14519 9033
rect 12124 8996 12169 9024
rect 12124 8984 12130 8996
rect 14461 8993 14473 9027
rect 14507 8993 14519 9027
rect 14461 8987 14519 8993
rect 13722 8956 13728 8968
rect 11992 8928 13728 8956
rect 13722 8916 13728 8928
rect 13780 8916 13786 8968
rect 14476 8956 14504 8987
rect 16574 8984 16580 9036
rect 16632 9024 16638 9036
rect 17037 9027 17095 9033
rect 17037 9024 17049 9027
rect 16632 8996 17049 9024
rect 16632 8984 16638 8996
rect 17037 8993 17049 8996
rect 17083 8993 17095 9027
rect 17037 8987 17095 8993
rect 14826 8956 14832 8968
rect 14476 8928 14832 8956
rect 14826 8916 14832 8928
rect 14884 8916 14890 8968
rect 15197 8959 15255 8965
rect 15197 8925 15209 8959
rect 15243 8956 15255 8959
rect 16850 8956 16856 8968
rect 15243 8928 16856 8956
rect 15243 8925 15255 8928
rect 15197 8919 15255 8925
rect 16850 8916 16856 8928
rect 16908 8916 16914 8968
rect 17494 8956 17500 8968
rect 17455 8928 17500 8956
rect 17494 8916 17500 8928
rect 17552 8916 17558 8968
rect 14185 8891 14243 8897
rect 14185 8888 14197 8891
rect 7024 8860 9812 8888
rect 11164 8860 14197 8888
rect 4801 8851 4859 8857
rect 4338 8780 4344 8832
rect 4396 8820 4402 8832
rect 4525 8823 4583 8829
rect 4525 8820 4537 8823
rect 4396 8792 4537 8820
rect 4396 8780 4402 8792
rect 4525 8789 4537 8792
rect 4571 8789 4583 8823
rect 5718 8820 5724 8832
rect 5679 8792 5724 8820
rect 4525 8783 4583 8789
rect 5718 8780 5724 8792
rect 5776 8780 5782 8832
rect 9784 8820 9812 8860
rect 14185 8857 14197 8860
rect 14231 8857 14243 8891
rect 14185 8851 14243 8857
rect 16577 8891 16635 8897
rect 16577 8857 16589 8891
rect 16623 8888 16635 8891
rect 16666 8888 16672 8900
rect 16623 8860 16672 8888
rect 16623 8857 16635 8860
rect 16577 8851 16635 8857
rect 16666 8848 16672 8860
rect 16724 8888 16730 8900
rect 17586 8888 17592 8900
rect 16724 8860 17592 8888
rect 16724 8848 16730 8860
rect 17586 8848 17592 8860
rect 17644 8848 17650 8900
rect 9858 8820 9864 8832
rect 9784 8792 9864 8820
rect 9858 8780 9864 8792
rect 9916 8780 9922 8832
rect 11974 8820 11980 8832
rect 11935 8792 11980 8820
rect 11974 8780 11980 8792
rect 12032 8780 12038 8832
rect 14737 8823 14795 8829
rect 14737 8789 14749 8823
rect 14783 8820 14795 8823
rect 15102 8820 15108 8832
rect 14783 8792 15108 8820
rect 14783 8789 14795 8792
rect 14737 8783 14795 8789
rect 15102 8780 15108 8792
rect 15160 8780 15166 8832
rect 16758 8820 16764 8832
rect 16719 8792 16764 8820
rect 16758 8780 16764 8792
rect 16816 8780 16822 8832
rect 184 8730 18924 8752
rect 184 8678 3110 8730
rect 3162 8678 3174 8730
rect 3226 8678 3238 8730
rect 3290 8678 3302 8730
rect 3354 8678 3366 8730
rect 3418 8678 6210 8730
rect 6262 8678 6274 8730
rect 6326 8678 6338 8730
rect 6390 8678 6402 8730
rect 6454 8678 6466 8730
rect 6518 8678 9310 8730
rect 9362 8678 9374 8730
rect 9426 8678 9438 8730
rect 9490 8678 9502 8730
rect 9554 8678 9566 8730
rect 9618 8678 12410 8730
rect 12462 8678 12474 8730
rect 12526 8678 12538 8730
rect 12590 8678 12602 8730
rect 12654 8678 12666 8730
rect 12718 8678 15510 8730
rect 15562 8678 15574 8730
rect 15626 8678 15638 8730
rect 15690 8678 15702 8730
rect 15754 8678 15766 8730
rect 15818 8678 18610 8730
rect 18662 8678 18674 8730
rect 18726 8678 18738 8730
rect 18790 8678 18802 8730
rect 18854 8678 18866 8730
rect 18918 8678 18924 8730
rect 184 8656 18924 8678
rect 750 8576 756 8628
rect 808 8616 814 8628
rect 3418 8616 3424 8628
rect 808 8588 2820 8616
rect 3379 8588 3424 8616
rect 808 8576 814 8588
rect 566 8372 572 8424
rect 624 8412 630 8424
rect 952 8421 980 8588
rect 1302 8548 1308 8560
rect 1263 8520 1308 8548
rect 1302 8508 1308 8520
rect 1360 8508 1366 8560
rect 2792 8548 2820 8588
rect 3418 8576 3424 8588
rect 3476 8576 3482 8628
rect 3694 8616 3700 8628
rect 3655 8588 3700 8616
rect 3694 8576 3700 8588
rect 3752 8576 3758 8628
rect 3970 8616 3976 8628
rect 3931 8588 3976 8616
rect 3970 8576 3976 8588
rect 4028 8576 4034 8628
rect 4246 8616 4252 8628
rect 4207 8588 4252 8616
rect 4246 8576 4252 8588
rect 4304 8576 4310 8628
rect 6546 8616 6552 8628
rect 6507 8588 6552 8616
rect 6546 8576 6552 8588
rect 6604 8576 6610 8628
rect 9674 8576 9680 8628
rect 9732 8616 9738 8628
rect 9953 8619 10011 8625
rect 9953 8616 9965 8619
rect 9732 8588 9965 8616
rect 9732 8576 9738 8588
rect 9953 8585 9965 8588
rect 9999 8585 10011 8619
rect 9953 8579 10011 8585
rect 10594 8576 10600 8628
rect 10652 8616 10658 8628
rect 10689 8619 10747 8625
rect 10689 8616 10701 8619
rect 10652 8588 10701 8616
rect 10652 8576 10658 8588
rect 10689 8585 10701 8588
rect 10735 8585 10747 8619
rect 10689 8579 10747 8585
rect 11072 8588 13768 8616
rect 3510 8548 3516 8560
rect 2792 8520 3516 8548
rect 3510 8508 3516 8520
rect 3568 8508 3574 8560
rect 3602 8508 3608 8560
rect 3660 8548 3666 8560
rect 3660 8520 3740 8548
rect 3660 8508 3666 8520
rect 1029 8483 1087 8489
rect 1029 8449 1041 8483
rect 1075 8480 1087 8483
rect 1118 8480 1124 8492
rect 1075 8452 1124 8480
rect 1075 8449 1087 8452
rect 1029 8443 1087 8449
rect 1118 8440 1124 8452
rect 1176 8480 1182 8492
rect 3418 8480 3424 8492
rect 1176 8452 3424 8480
rect 1176 8440 1182 8452
rect 3418 8440 3424 8452
rect 3476 8440 3482 8492
rect 3712 8480 3740 8520
rect 8294 8508 8300 8560
rect 8352 8548 8358 8560
rect 10505 8551 10563 8557
rect 10505 8548 10517 8551
rect 8352 8520 10517 8548
rect 8352 8508 8358 8520
rect 10505 8517 10517 8520
rect 10551 8517 10563 8551
rect 10505 8511 10563 8517
rect 5166 8480 5172 8492
rect 3712 8452 5172 8480
rect 661 8415 719 8421
rect 661 8412 673 8415
rect 624 8384 673 8412
rect 624 8372 630 8384
rect 661 8381 673 8384
rect 707 8381 719 8415
rect 661 8375 719 8381
rect 937 8415 995 8421
rect 937 8381 949 8415
rect 983 8381 995 8415
rect 937 8375 995 8381
rect 1394 8372 1400 8424
rect 1452 8412 1458 8424
rect 1489 8415 1547 8421
rect 1489 8412 1501 8415
rect 1452 8384 1501 8412
rect 1452 8372 1458 8384
rect 1489 8381 1501 8384
rect 1535 8381 1547 8415
rect 1489 8375 1547 8381
rect 2866 8372 2872 8424
rect 2924 8412 2930 8424
rect 3050 8412 3056 8424
rect 2924 8384 3056 8412
rect 2924 8372 2930 8384
rect 3050 8372 3056 8384
rect 3108 8372 3114 8424
rect 3329 8415 3387 8421
rect 3329 8381 3341 8415
rect 3375 8381 3387 8415
rect 3510 8412 3516 8424
rect 3471 8384 3516 8412
rect 3329 8375 3387 8381
rect 750 8304 756 8356
rect 808 8344 814 8356
rect 1765 8347 1823 8353
rect 1765 8344 1777 8347
rect 808 8316 1777 8344
rect 808 8304 814 8316
rect 1765 8313 1777 8316
rect 1811 8313 1823 8347
rect 3344 8344 3372 8375
rect 3510 8372 3516 8384
rect 3568 8372 3574 8424
rect 3712 8344 3740 8452
rect 5166 8440 5172 8452
rect 5224 8480 5230 8492
rect 5534 8480 5540 8492
rect 5224 8452 5540 8480
rect 5224 8440 5230 8452
rect 5534 8440 5540 8452
rect 5592 8440 5598 8492
rect 7098 8480 7104 8492
rect 6564 8452 7104 8480
rect 3878 8412 3884 8424
rect 3839 8384 3884 8412
rect 3878 8372 3884 8384
rect 3936 8372 3942 8424
rect 4246 8372 4252 8424
rect 4304 8412 4310 8424
rect 6564 8421 6592 8452
rect 7098 8440 7104 8452
rect 7156 8440 7162 8492
rect 7834 8440 7840 8492
rect 7892 8480 7898 8492
rect 11072 8489 11100 8588
rect 12250 8508 12256 8560
rect 12308 8548 12314 8560
rect 13740 8548 13768 8588
rect 13814 8576 13820 8628
rect 13872 8616 13878 8628
rect 14737 8619 14795 8625
rect 14737 8616 14749 8619
rect 13872 8588 14749 8616
rect 13872 8576 13878 8588
rect 14737 8585 14749 8588
rect 14783 8585 14795 8619
rect 14737 8579 14795 8585
rect 15381 8619 15439 8625
rect 15381 8585 15393 8619
rect 15427 8616 15439 8619
rect 15930 8616 15936 8628
rect 15427 8588 15936 8616
rect 15427 8585 15439 8588
rect 15381 8579 15439 8585
rect 15930 8576 15936 8588
rect 15988 8576 15994 8628
rect 18322 8616 18328 8628
rect 18283 8588 18328 8616
rect 18322 8576 18328 8588
rect 18380 8576 18386 8628
rect 12308 8520 13216 8548
rect 13740 8520 13860 8548
rect 12308 8508 12314 8520
rect 8481 8483 8539 8489
rect 8481 8480 8493 8483
rect 7892 8452 8493 8480
rect 7892 8440 7898 8452
rect 8481 8449 8493 8452
rect 8527 8480 8539 8483
rect 11057 8483 11115 8489
rect 8527 8452 11008 8480
rect 8527 8449 8539 8452
rect 8481 8443 8539 8449
rect 4341 8415 4399 8421
rect 4341 8412 4353 8415
rect 4304 8384 4353 8412
rect 4304 8372 4310 8384
rect 4341 8381 4353 8384
rect 4387 8381 4399 8415
rect 4341 8375 4399 8381
rect 6549 8415 6607 8421
rect 6549 8381 6561 8415
rect 6595 8381 6607 8415
rect 6549 8375 6607 8381
rect 6733 8415 6791 8421
rect 6733 8381 6745 8415
rect 6779 8412 6791 8415
rect 6914 8412 6920 8424
rect 6779 8384 6920 8412
rect 6779 8381 6791 8384
rect 6733 8375 6791 8381
rect 6914 8372 6920 8384
rect 6972 8412 6978 8424
rect 7926 8412 7932 8424
rect 6972 8384 7932 8412
rect 6972 8372 6978 8384
rect 7926 8372 7932 8384
rect 7984 8372 7990 8424
rect 9030 8372 9036 8424
rect 9088 8412 9094 8424
rect 10594 8412 10600 8424
rect 9088 8384 10600 8412
rect 9088 8372 9094 8384
rect 10594 8372 10600 8384
rect 10652 8372 10658 8424
rect 10689 8415 10747 8421
rect 10689 8381 10701 8415
rect 10735 8381 10747 8415
rect 10689 8375 10747 8381
rect 10873 8415 10931 8421
rect 10873 8381 10885 8415
rect 10919 8381 10931 8415
rect 10980 8412 11008 8452
rect 11057 8449 11069 8483
rect 11103 8449 11115 8483
rect 12802 8480 12808 8492
rect 11057 8443 11115 8449
rect 11164 8452 12808 8480
rect 11164 8412 11192 8452
rect 12802 8440 12808 8452
rect 12860 8440 12866 8492
rect 11422 8412 11428 8424
rect 10980 8384 11192 8412
rect 11383 8384 11428 8412
rect 10873 8375 10931 8381
rect 1765 8307 1823 8313
rect 3068 8316 3740 8344
rect 566 8276 572 8288
rect 527 8248 572 8276
rect 566 8236 572 8248
rect 624 8236 630 8288
rect 2590 8236 2596 8288
rect 2648 8276 2654 8288
rect 3068 8276 3096 8316
rect 4430 8304 4436 8356
rect 4488 8344 4494 8356
rect 6089 8347 6147 8353
rect 6089 8344 6101 8347
rect 4488 8316 6101 8344
rect 4488 8304 4494 8316
rect 6089 8313 6101 8316
rect 6135 8344 6147 8347
rect 8665 8347 8723 8353
rect 8665 8344 8677 8347
rect 6135 8316 8677 8344
rect 6135 8313 6147 8316
rect 6089 8307 6147 8313
rect 8665 8313 8677 8316
rect 8711 8313 8723 8347
rect 8665 8307 8723 8313
rect 8846 8304 8852 8356
rect 8904 8344 8910 8356
rect 10704 8344 10732 8375
rect 10778 8344 10784 8356
rect 8904 8316 10784 8344
rect 8904 8304 8910 8316
rect 10778 8304 10784 8316
rect 10836 8304 10842 8356
rect 2648 8248 3096 8276
rect 3237 8279 3295 8285
rect 2648 8236 2654 8248
rect 3237 8245 3249 8279
rect 3283 8276 3295 8279
rect 3418 8276 3424 8288
rect 3283 8248 3424 8276
rect 3283 8245 3295 8248
rect 3237 8239 3295 8245
rect 3418 8236 3424 8248
rect 3476 8276 3482 8288
rect 5350 8276 5356 8288
rect 3476 8248 5356 8276
rect 3476 8236 3482 8248
rect 5350 8236 5356 8248
rect 5408 8236 5414 8288
rect 10134 8236 10140 8288
rect 10192 8276 10198 8288
rect 10888 8276 10916 8375
rect 11422 8372 11428 8384
rect 11480 8372 11486 8424
rect 12342 8372 12348 8424
rect 12400 8412 12406 8424
rect 13188 8421 13216 8520
rect 13832 8492 13860 8520
rect 17586 8508 17592 8560
rect 17644 8548 17650 8560
rect 17865 8551 17923 8557
rect 17865 8548 17877 8551
rect 17644 8520 17877 8548
rect 17644 8508 17650 8520
rect 17865 8517 17877 8520
rect 17911 8517 17923 8551
rect 17865 8511 17923 8517
rect 13814 8440 13820 8492
rect 13872 8440 13878 8492
rect 14292 8452 15516 8480
rect 12989 8415 13047 8421
rect 12989 8412 13001 8415
rect 12400 8384 13001 8412
rect 12400 8372 12406 8384
rect 12989 8381 13001 8384
rect 13035 8381 13047 8415
rect 12989 8375 13047 8381
rect 13173 8415 13231 8421
rect 13173 8381 13185 8415
rect 13219 8381 13231 8415
rect 13173 8375 13231 8381
rect 13449 8415 13507 8421
rect 13449 8381 13461 8415
rect 13495 8412 13507 8415
rect 13538 8412 13544 8424
rect 13495 8384 13544 8412
rect 13495 8381 13507 8384
rect 13449 8375 13507 8381
rect 13538 8372 13544 8384
rect 13596 8372 13602 8424
rect 13722 8372 13728 8424
rect 13780 8412 13786 8424
rect 14292 8412 14320 8452
rect 13780 8384 14320 8412
rect 13780 8372 13786 8384
rect 14366 8372 14372 8424
rect 14424 8412 14430 8424
rect 15488 8421 15516 8452
rect 17678 8440 17684 8492
rect 17736 8480 17742 8492
rect 17773 8483 17831 8489
rect 17773 8480 17785 8483
rect 17736 8452 17785 8480
rect 17736 8440 17742 8452
rect 17773 8449 17785 8452
rect 17819 8449 17831 8483
rect 17773 8443 17831 8449
rect 15289 8415 15347 8421
rect 15289 8412 15301 8415
rect 14424 8384 15301 8412
rect 14424 8372 14430 8384
rect 15289 8381 15301 8384
rect 15335 8381 15347 8415
rect 15289 8375 15347 8381
rect 15473 8415 15531 8421
rect 15473 8381 15485 8415
rect 15519 8381 15531 8415
rect 15473 8375 15531 8381
rect 15657 8415 15715 8421
rect 15657 8381 15669 8415
rect 15703 8412 15715 8415
rect 16758 8412 16764 8424
rect 15703 8384 16764 8412
rect 15703 8381 15715 8384
rect 15657 8375 15715 8381
rect 16758 8372 16764 8384
rect 16816 8372 16822 8424
rect 16942 8372 16948 8424
rect 17000 8412 17006 8424
rect 18049 8415 18107 8421
rect 17000 8384 17816 8412
rect 17000 8372 17006 8384
rect 12158 8304 12164 8356
rect 12216 8304 12222 8356
rect 12851 8347 12909 8353
rect 12851 8313 12863 8347
rect 12897 8344 12909 8347
rect 14384 8344 14412 8372
rect 15838 8344 15844 8356
rect 12897 8316 14412 8344
rect 15488 8316 15700 8344
rect 15799 8316 15844 8344
rect 12897 8313 12909 8316
rect 12851 8307 12909 8313
rect 11514 8276 11520 8288
rect 10192 8248 11520 8276
rect 10192 8236 10198 8248
rect 11514 8236 11520 8248
rect 11572 8236 11578 8288
rect 12066 8236 12072 8288
rect 12124 8276 12130 8288
rect 12866 8276 12894 8307
rect 13078 8276 13084 8288
rect 12124 8248 12894 8276
rect 13039 8248 13084 8276
rect 12124 8236 12130 8248
rect 13078 8236 13084 8248
rect 13136 8236 13142 8288
rect 13170 8236 13176 8288
rect 13228 8276 13234 8288
rect 15488 8276 15516 8316
rect 13228 8248 15516 8276
rect 15672 8276 15700 8316
rect 15838 8304 15844 8316
rect 15896 8304 15902 8356
rect 17494 8344 17500 8356
rect 16776 8316 17500 8344
rect 16776 8276 16804 8316
rect 17494 8304 17500 8316
rect 17552 8304 17558 8356
rect 17681 8347 17739 8353
rect 17681 8313 17693 8347
rect 17727 8313 17739 8347
rect 17788 8344 17816 8384
rect 18049 8381 18061 8415
rect 18095 8412 18107 8415
rect 18322 8412 18328 8424
rect 18095 8384 18328 8412
rect 18095 8381 18107 8384
rect 18049 8375 18107 8381
rect 18322 8372 18328 8384
rect 18380 8372 18386 8424
rect 18417 8347 18475 8353
rect 18417 8344 18429 8347
rect 17788 8316 18429 8344
rect 17681 8307 17739 8313
rect 18417 8313 18429 8316
rect 18463 8313 18475 8347
rect 18417 8307 18475 8313
rect 15672 8248 16804 8276
rect 13228 8236 13234 8248
rect 16850 8236 16856 8288
rect 16908 8276 16914 8288
rect 17129 8279 17187 8285
rect 17129 8276 17141 8279
rect 16908 8248 17141 8276
rect 16908 8236 16914 8248
rect 17129 8245 17141 8248
rect 17175 8245 17187 8279
rect 17129 8239 17187 8245
rect 17402 8236 17408 8288
rect 17460 8276 17466 8288
rect 17696 8276 17724 8307
rect 17954 8276 17960 8288
rect 17460 8248 17724 8276
rect 17915 8248 17960 8276
rect 17460 8236 17466 8248
rect 17954 8236 17960 8248
rect 18012 8236 18018 8288
rect 184 8186 18860 8208
rect 184 8134 4660 8186
rect 4712 8134 4724 8186
rect 4776 8134 4788 8186
rect 4840 8134 4852 8186
rect 4904 8134 4916 8186
rect 4968 8134 7760 8186
rect 7812 8134 7824 8186
rect 7876 8134 7888 8186
rect 7940 8134 7952 8186
rect 8004 8134 8016 8186
rect 8068 8134 10860 8186
rect 10912 8134 10924 8186
rect 10976 8134 10988 8186
rect 11040 8134 11052 8186
rect 11104 8134 11116 8186
rect 11168 8134 13960 8186
rect 14012 8134 14024 8186
rect 14076 8134 14088 8186
rect 14140 8134 14152 8186
rect 14204 8134 14216 8186
rect 14268 8134 17060 8186
rect 17112 8134 17124 8186
rect 17176 8134 17188 8186
rect 17240 8134 17252 8186
rect 17304 8134 17316 8186
rect 17368 8134 18860 8186
rect 184 8112 18860 8134
rect 566 8032 572 8084
rect 624 8072 630 8084
rect 2406 8072 2412 8084
rect 624 8044 2412 8072
rect 624 8032 630 8044
rect 2406 8032 2412 8044
rect 2464 8032 2470 8084
rect 3053 8075 3111 8081
rect 3053 8041 3065 8075
rect 3099 8072 3111 8075
rect 4154 8072 4160 8084
rect 3099 8044 4160 8072
rect 3099 8041 3111 8044
rect 3053 8035 3111 8041
rect 4154 8032 4160 8044
rect 4212 8032 4218 8084
rect 4893 8075 4951 8081
rect 4893 8041 4905 8075
rect 4939 8072 4951 8075
rect 5074 8072 5080 8084
rect 4939 8044 5080 8072
rect 4939 8041 4951 8044
rect 4893 8035 4951 8041
rect 5074 8032 5080 8044
rect 5132 8032 5138 8084
rect 7190 8072 7196 8084
rect 7151 8044 7196 8072
rect 7190 8032 7196 8044
rect 7248 8032 7254 8084
rect 8297 8075 8355 8081
rect 8297 8041 8309 8075
rect 8343 8072 8355 8075
rect 9766 8072 9772 8084
rect 8343 8044 9772 8072
rect 8343 8041 8355 8044
rect 8297 8035 8355 8041
rect 9766 8032 9772 8044
rect 9824 8032 9830 8084
rect 10042 8032 10048 8084
rect 10100 8072 10106 8084
rect 14734 8072 14740 8084
rect 10100 8044 14740 8072
rect 10100 8032 10106 8044
rect 14734 8032 14740 8044
rect 14792 8032 14798 8084
rect 15010 8032 15016 8084
rect 15068 8032 15074 8084
rect 16206 8032 16212 8084
rect 16264 8072 16270 8084
rect 16264 8044 17172 8072
rect 16264 8032 16270 8044
rect 658 8004 664 8016
rect 619 7976 664 8004
rect 658 7964 664 7976
rect 716 7964 722 8016
rect 845 8007 903 8013
rect 845 7973 857 8007
rect 891 8004 903 8007
rect 2133 8007 2191 8013
rect 2133 8004 2145 8007
rect 891 7976 2145 8004
rect 891 7973 903 7976
rect 845 7967 903 7973
rect 2133 7973 2145 7976
rect 2179 7973 2191 8007
rect 2133 7967 2191 7973
rect 2958 7964 2964 8016
rect 3016 8004 3022 8016
rect 3758 8007 3816 8013
rect 3758 8004 3770 8007
rect 3016 7976 3770 8004
rect 3016 7964 3022 7976
rect 3758 7973 3770 7976
rect 3804 7973 3816 8007
rect 3758 7967 3816 7973
rect 3878 7964 3884 8016
rect 3936 7964 3942 8016
rect 4430 7964 4436 8016
rect 4488 8004 4494 8016
rect 4488 7976 5488 8004
rect 4488 7964 4494 7976
rect 477 7939 535 7945
rect 477 7905 489 7939
rect 523 7936 535 7939
rect 566 7936 572 7948
rect 523 7908 572 7936
rect 523 7905 535 7908
rect 477 7899 535 7905
rect 566 7896 572 7908
rect 624 7896 630 7948
rect 1118 7896 1124 7948
rect 1176 7936 1182 7948
rect 1305 7939 1363 7945
rect 1305 7936 1317 7939
rect 1176 7908 1317 7936
rect 1176 7896 1182 7908
rect 1305 7905 1317 7908
rect 1351 7905 1363 7939
rect 3896 7936 3924 7964
rect 1305 7899 1363 7905
rect 3344 7908 3924 7936
rect 1029 7871 1087 7877
rect 1029 7837 1041 7871
rect 1075 7837 1087 7871
rect 1210 7868 1216 7880
rect 1171 7840 1216 7868
rect 1029 7831 1087 7837
rect 1044 7800 1072 7831
rect 1210 7828 1216 7840
rect 1268 7828 1274 7880
rect 2222 7868 2228 7880
rect 2183 7840 2228 7868
rect 2222 7828 2228 7840
rect 2280 7828 2286 7880
rect 2406 7868 2412 7880
rect 2367 7840 2412 7868
rect 2406 7828 2412 7840
rect 2464 7828 2470 7880
rect 2774 7828 2780 7880
rect 2832 7868 2838 7880
rect 3344 7877 3372 7908
rect 4062 7896 4068 7948
rect 4120 7936 4126 7948
rect 5460 7945 5488 7976
rect 8386 7964 8392 8016
rect 8444 8004 8450 8016
rect 10137 8007 10195 8013
rect 10137 8004 10149 8007
rect 8444 7976 10149 8004
rect 8444 7964 8450 7976
rect 10137 7973 10149 7976
rect 10183 7973 10195 8007
rect 11698 8004 11704 8016
rect 11362 7976 11704 8004
rect 10137 7967 10195 7973
rect 11698 7964 11704 7976
rect 11756 7964 11762 8016
rect 11974 8004 11980 8016
rect 11935 7976 11980 8004
rect 11974 7964 11980 7976
rect 12032 8004 12038 8016
rect 14093 8007 14151 8013
rect 12032 7976 12434 8004
rect 12032 7964 12038 7976
rect 5169 7939 5227 7945
rect 5169 7936 5181 7939
rect 4120 7908 5181 7936
rect 4120 7896 4126 7908
rect 5169 7905 5181 7908
rect 5215 7905 5227 7939
rect 5169 7899 5227 7905
rect 5445 7939 5503 7945
rect 5445 7905 5457 7939
rect 5491 7905 5503 7939
rect 6086 7936 6092 7948
rect 6047 7908 6092 7936
rect 5445 7899 5503 7905
rect 6086 7896 6092 7908
rect 6144 7896 6150 7948
rect 6178 7896 6184 7948
rect 6236 7936 6242 7948
rect 6273 7939 6331 7945
rect 6273 7936 6285 7939
rect 6236 7908 6285 7936
rect 6236 7896 6242 7908
rect 6273 7905 6285 7908
rect 6319 7936 6331 7939
rect 6638 7936 6644 7948
rect 6319 7908 6644 7936
rect 6319 7905 6331 7908
rect 6273 7899 6331 7905
rect 6638 7896 6644 7908
rect 6696 7896 6702 7948
rect 6822 7936 6828 7948
rect 6783 7908 6828 7936
rect 6822 7896 6828 7908
rect 6880 7896 6886 7948
rect 7006 7936 7012 7948
rect 6967 7908 7012 7936
rect 7006 7896 7012 7908
rect 7064 7896 7070 7948
rect 7561 7939 7619 7945
rect 7561 7905 7573 7939
rect 7607 7936 7619 7939
rect 7650 7936 7656 7948
rect 7607 7908 7656 7936
rect 7607 7905 7619 7908
rect 7561 7899 7619 7905
rect 7650 7896 7656 7908
rect 7708 7896 7714 7948
rect 7745 7939 7803 7945
rect 7745 7905 7757 7939
rect 7791 7936 7803 7939
rect 8294 7936 8300 7948
rect 7791 7908 8300 7936
rect 7791 7905 7803 7908
rect 7745 7899 7803 7905
rect 8294 7896 8300 7908
rect 8352 7896 8358 7948
rect 9585 7939 9643 7945
rect 9585 7905 9597 7939
rect 9631 7936 9643 7939
rect 9766 7936 9772 7948
rect 9631 7908 9772 7936
rect 9631 7905 9643 7908
rect 9585 7899 9643 7905
rect 9766 7896 9772 7908
rect 9824 7896 9830 7948
rect 11790 7936 11796 7948
rect 11751 7908 11796 7936
rect 11790 7896 11796 7908
rect 11848 7896 11854 7948
rect 12066 7936 12072 7948
rect 12027 7908 12072 7936
rect 12066 7896 12072 7908
rect 12124 7896 12130 7948
rect 12253 7939 12311 7945
rect 12253 7905 12265 7939
rect 12299 7905 12311 7939
rect 12253 7899 12311 7905
rect 3145 7871 3203 7877
rect 3145 7868 3157 7871
rect 2832 7840 3157 7868
rect 2832 7828 2838 7840
rect 3145 7837 3157 7840
rect 3191 7837 3203 7871
rect 3145 7831 3203 7837
rect 3329 7871 3387 7877
rect 3329 7837 3341 7871
rect 3375 7837 3387 7871
rect 3510 7868 3516 7880
rect 3471 7840 3516 7868
rect 3329 7831 3387 7837
rect 3510 7828 3516 7840
rect 3568 7828 3574 7880
rect 4982 7828 4988 7880
rect 5040 7868 5046 7880
rect 5077 7871 5135 7877
rect 5077 7868 5089 7871
rect 5040 7840 5089 7868
rect 5040 7828 5046 7840
rect 5077 7837 5089 7840
rect 5123 7837 5135 7871
rect 5077 7831 5135 7837
rect 5718 7828 5724 7880
rect 5776 7868 5782 7880
rect 6546 7868 6552 7880
rect 5776 7840 6552 7868
rect 5776 7828 5782 7840
rect 6546 7828 6552 7840
rect 6604 7868 6610 7880
rect 9861 7871 9919 7877
rect 9861 7868 9873 7871
rect 6604 7840 9873 7868
rect 6604 7828 6610 7840
rect 9861 7837 9873 7840
rect 9907 7837 9919 7871
rect 12268 7868 12296 7899
rect 9861 7831 9919 7837
rect 11440 7840 12296 7868
rect 12406 7868 12434 7976
rect 14093 7973 14105 8007
rect 14139 8004 14151 8007
rect 14366 8004 14372 8016
rect 14139 7976 14372 8004
rect 14139 7973 14151 7976
rect 14093 7967 14151 7973
rect 14366 7964 14372 7976
rect 14424 7964 14430 8016
rect 14461 8007 14519 8013
rect 14461 7973 14473 8007
rect 14507 8004 14519 8007
rect 15028 8004 15056 8032
rect 14507 7976 15056 8004
rect 14507 7973 14519 7976
rect 14461 7967 14519 7973
rect 16114 7964 16120 8016
rect 16172 8004 16178 8016
rect 16482 8004 16488 8016
rect 16172 7976 16488 8004
rect 16172 7964 16178 7976
rect 16482 7964 16488 7976
rect 16540 7964 16546 8016
rect 16666 7964 16672 8016
rect 16724 8004 16730 8016
rect 17144 8004 17172 8044
rect 17310 8032 17316 8084
rect 17368 8072 17374 8084
rect 17402 8072 17408 8084
rect 17368 8044 17408 8072
rect 17368 8032 17374 8044
rect 17402 8032 17408 8044
rect 17460 8032 17466 8084
rect 18138 8032 18144 8084
rect 18196 8072 18202 8084
rect 18325 8075 18383 8081
rect 18325 8072 18337 8075
rect 18196 8044 18337 8072
rect 18196 8032 18202 8044
rect 18325 8041 18337 8044
rect 18371 8041 18383 8075
rect 18325 8035 18383 8041
rect 18049 8007 18107 8013
rect 18049 8004 18061 8007
rect 16724 7976 17080 8004
rect 17144 7976 18061 8004
rect 16724 7964 16730 7976
rect 13722 7896 13728 7948
rect 13780 7936 13786 7948
rect 14277 7939 14335 7945
rect 14277 7936 14289 7939
rect 13780 7908 14289 7936
rect 13780 7896 13786 7908
rect 14277 7905 14289 7908
rect 14323 7905 14335 7939
rect 14277 7899 14335 7905
rect 14920 7939 14978 7945
rect 14920 7905 14932 7939
rect 14966 7905 14978 7939
rect 14920 7899 14978 7905
rect 14936 7868 14964 7899
rect 15010 7896 15016 7948
rect 15068 7936 15074 7948
rect 15068 7908 15113 7936
rect 15068 7896 15074 7908
rect 16850 7896 16856 7948
rect 16908 7936 16914 7948
rect 17052 7945 17080 7976
rect 18049 7973 18061 7976
rect 18095 7973 18107 8007
rect 18049 7967 18107 7973
rect 17037 7939 17095 7945
rect 16908 7908 16953 7936
rect 16908 7896 16914 7908
rect 17037 7905 17049 7939
rect 17083 7905 17095 7939
rect 17037 7899 17095 7905
rect 17218 7896 17224 7948
rect 17276 7936 17282 7948
rect 17402 7936 17408 7948
rect 17276 7908 17408 7936
rect 17276 7896 17282 7908
rect 17402 7896 17408 7908
rect 17460 7896 17466 7948
rect 17678 7896 17684 7948
rect 17736 7936 17742 7948
rect 18233 7939 18291 7945
rect 18233 7936 18245 7939
rect 17736 7908 18245 7936
rect 17736 7896 17742 7908
rect 18233 7905 18245 7908
rect 18279 7905 18291 7939
rect 18414 7936 18420 7948
rect 18375 7908 18420 7936
rect 18233 7899 18291 7905
rect 18414 7896 18420 7908
rect 18472 7896 18478 7948
rect 16114 7868 16120 7880
rect 12406 7840 14780 7868
rect 14936 7840 16120 7868
rect 1486 7800 1492 7812
rect 1044 7772 1492 7800
rect 1486 7760 1492 7772
rect 1544 7800 1550 7812
rect 1765 7803 1823 7809
rect 1765 7800 1777 7803
rect 1544 7772 1777 7800
rect 1544 7760 1550 7772
rect 1765 7769 1777 7772
rect 1811 7769 1823 7803
rect 1765 7763 1823 7769
rect 2130 7760 2136 7812
rect 2188 7800 2194 7812
rect 2685 7803 2743 7809
rect 2685 7800 2697 7803
rect 2188 7772 2697 7800
rect 2188 7760 2194 7772
rect 2685 7769 2697 7772
rect 2731 7769 2743 7803
rect 2685 7763 2743 7769
rect 5166 7760 5172 7812
rect 5224 7800 5230 7812
rect 9122 7800 9128 7812
rect 5224 7772 9128 7800
rect 5224 7760 5230 7772
rect 9122 7760 9128 7772
rect 9180 7760 9186 7812
rect 1670 7732 1676 7744
rect 1631 7704 1676 7732
rect 1670 7692 1676 7704
rect 1728 7692 1734 7744
rect 2866 7692 2872 7744
rect 2924 7732 2930 7744
rect 3050 7732 3056 7744
rect 2924 7704 3056 7732
rect 2924 7692 2930 7704
rect 3050 7692 3056 7704
rect 3108 7732 3114 7744
rect 3694 7732 3700 7744
rect 3108 7704 3700 7732
rect 3108 7692 3114 7704
rect 3694 7692 3700 7704
rect 3752 7692 3758 7744
rect 3878 7692 3884 7744
rect 3936 7732 3942 7744
rect 5810 7732 5816 7744
rect 3936 7704 5816 7732
rect 3936 7692 3942 7704
rect 5810 7692 5816 7704
rect 5868 7692 5874 7744
rect 7653 7735 7711 7741
rect 7653 7701 7665 7735
rect 7699 7732 7711 7735
rect 8478 7732 8484 7744
rect 7699 7704 8484 7732
rect 7699 7701 7711 7704
rect 7653 7695 7711 7701
rect 8478 7692 8484 7704
rect 8536 7692 8542 7744
rect 9858 7692 9864 7744
rect 9916 7732 9922 7744
rect 11440 7732 11468 7840
rect 11793 7803 11851 7809
rect 11793 7769 11805 7803
rect 11839 7800 11851 7803
rect 11882 7800 11888 7812
rect 11839 7772 11888 7800
rect 11839 7769 11851 7772
rect 11793 7763 11851 7769
rect 11882 7760 11888 7772
rect 11940 7760 11946 7812
rect 13262 7760 13268 7812
rect 13320 7800 13326 7812
rect 14645 7803 14703 7809
rect 14645 7800 14657 7803
rect 13320 7772 14657 7800
rect 13320 7760 13326 7772
rect 14645 7769 14657 7772
rect 14691 7769 14703 7803
rect 14752 7800 14780 7840
rect 16114 7828 16120 7840
rect 16172 7828 16178 7880
rect 16577 7871 16635 7877
rect 16577 7837 16589 7871
rect 16623 7868 16635 7871
rect 16623 7840 16988 7868
rect 16623 7837 16635 7840
rect 16577 7831 16635 7837
rect 16960 7800 16988 7840
rect 17310 7828 17316 7880
rect 17368 7868 17374 7880
rect 17497 7871 17555 7877
rect 17497 7868 17509 7871
rect 17368 7840 17509 7868
rect 17368 7828 17374 7840
rect 17497 7837 17509 7840
rect 17543 7868 17555 7871
rect 17862 7868 17868 7880
rect 17543 7840 17868 7868
rect 17543 7837 17555 7840
rect 17497 7831 17555 7837
rect 17862 7828 17868 7840
rect 17920 7828 17926 7880
rect 18322 7800 18328 7812
rect 14752 7772 15424 7800
rect 16960 7772 18328 7800
rect 14645 7763 14703 7769
rect 9916 7704 11468 7732
rect 9916 7692 9922 7704
rect 11514 7692 11520 7744
rect 11572 7732 11578 7744
rect 11609 7735 11667 7741
rect 11609 7732 11621 7735
rect 11572 7704 11621 7732
rect 11572 7692 11578 7704
rect 11609 7701 11621 7704
rect 11655 7732 11667 7735
rect 12250 7732 12256 7744
rect 11655 7704 12256 7732
rect 11655 7701 11667 7704
rect 11609 7695 11667 7701
rect 12250 7692 12256 7704
rect 12308 7692 12314 7744
rect 13725 7735 13783 7741
rect 13725 7701 13737 7735
rect 13771 7732 13783 7735
rect 13814 7732 13820 7744
rect 13771 7704 13820 7732
rect 13771 7701 13783 7704
rect 13725 7695 13783 7701
rect 13814 7692 13820 7704
rect 13872 7692 13878 7744
rect 15105 7735 15163 7741
rect 15105 7701 15117 7735
rect 15151 7732 15163 7735
rect 15286 7732 15292 7744
rect 15151 7704 15292 7732
rect 15151 7701 15163 7704
rect 15105 7695 15163 7701
rect 15286 7692 15292 7704
rect 15344 7692 15350 7744
rect 15396 7732 15424 7772
rect 18322 7760 18328 7772
rect 18380 7760 18386 7812
rect 17402 7732 17408 7744
rect 15396 7704 17408 7732
rect 17402 7692 17408 7704
rect 17460 7692 17466 7744
rect 184 7642 18924 7664
rect 184 7590 3110 7642
rect 3162 7590 3174 7642
rect 3226 7590 3238 7642
rect 3290 7590 3302 7642
rect 3354 7590 3366 7642
rect 3418 7590 6210 7642
rect 6262 7590 6274 7642
rect 6326 7590 6338 7642
rect 6390 7590 6402 7642
rect 6454 7590 6466 7642
rect 6518 7590 9310 7642
rect 9362 7590 9374 7642
rect 9426 7590 9438 7642
rect 9490 7590 9502 7642
rect 9554 7590 9566 7642
rect 9618 7590 12410 7642
rect 12462 7590 12474 7642
rect 12526 7590 12538 7642
rect 12590 7590 12602 7642
rect 12654 7590 12666 7642
rect 12718 7590 15510 7642
rect 15562 7590 15574 7642
rect 15626 7590 15638 7642
rect 15690 7590 15702 7642
rect 15754 7590 15766 7642
rect 15818 7590 18610 7642
rect 18662 7590 18674 7642
rect 18726 7590 18738 7642
rect 18790 7590 18802 7642
rect 18854 7590 18866 7642
rect 18918 7590 18924 7642
rect 184 7568 18924 7590
rect 661 7531 719 7537
rect 661 7497 673 7531
rect 707 7528 719 7531
rect 750 7528 756 7540
rect 707 7500 756 7528
rect 707 7497 719 7500
rect 661 7491 719 7497
rect 750 7488 756 7500
rect 808 7488 814 7540
rect 1210 7488 1216 7540
rect 1268 7528 1274 7540
rect 3326 7528 3332 7540
rect 1268 7500 3332 7528
rect 1268 7488 1274 7500
rect 3326 7488 3332 7500
rect 3384 7488 3390 7540
rect 3602 7488 3608 7540
rect 3660 7528 3666 7540
rect 3660 7500 5304 7528
rect 3660 7488 3666 7500
rect 569 7463 627 7469
rect 569 7429 581 7463
rect 615 7460 627 7463
rect 934 7460 940 7472
rect 615 7432 940 7460
rect 615 7429 627 7432
rect 569 7423 627 7429
rect 934 7420 940 7432
rect 992 7420 998 7472
rect 2774 7420 2780 7472
rect 2832 7460 2838 7472
rect 3421 7463 3479 7469
rect 3421 7460 3433 7463
rect 2832 7432 3433 7460
rect 2832 7420 2838 7432
rect 3421 7429 3433 7432
rect 3467 7460 3479 7463
rect 3970 7460 3976 7472
rect 3467 7432 3976 7460
rect 3467 7429 3479 7432
rect 3421 7423 3479 7429
rect 3970 7420 3976 7432
rect 4028 7420 4034 7472
rect 4062 7420 4068 7472
rect 4120 7460 4126 7472
rect 4120 7432 4844 7460
rect 4120 7420 4126 7432
rect 753 7395 811 7401
rect 753 7361 765 7395
rect 799 7392 811 7395
rect 842 7392 848 7404
rect 799 7364 848 7392
rect 799 7361 811 7364
rect 753 7355 811 7361
rect 842 7352 848 7364
rect 900 7352 906 7404
rect 1302 7392 1308 7404
rect 1263 7364 1308 7392
rect 1302 7352 1308 7364
rect 1360 7392 1366 7404
rect 2130 7392 2136 7404
rect 1360 7364 2136 7392
rect 1360 7352 1366 7364
rect 2130 7352 2136 7364
rect 2188 7392 2194 7404
rect 2188 7364 3556 7392
rect 2188 7352 2194 7364
rect 474 7324 480 7336
rect 435 7296 480 7324
rect 474 7284 480 7296
rect 532 7284 538 7336
rect 1029 7327 1087 7333
rect 1029 7293 1041 7327
rect 1075 7324 1087 7327
rect 1118 7324 1124 7336
rect 1075 7296 1124 7324
rect 1075 7293 1087 7296
rect 1029 7287 1087 7293
rect 1118 7284 1124 7296
rect 1176 7284 1182 7336
rect 1210 7284 1216 7336
rect 1268 7324 1274 7336
rect 1268 7296 1313 7324
rect 1268 7284 1274 7296
rect 1394 7284 1400 7336
rect 1452 7324 1458 7336
rect 1489 7327 1547 7333
rect 1489 7324 1501 7327
rect 1452 7296 1501 7324
rect 1452 7284 1458 7296
rect 1489 7293 1501 7296
rect 1535 7293 1547 7327
rect 1489 7287 1547 7293
rect 2866 7284 2872 7336
rect 2924 7284 2930 7336
rect 3528 7333 3556 7364
rect 3786 7352 3792 7404
rect 3844 7392 3850 7404
rect 4816 7401 4844 7432
rect 4157 7395 4215 7401
rect 4157 7392 4169 7395
rect 3844 7364 4169 7392
rect 3844 7352 3850 7364
rect 4157 7361 4169 7364
rect 4203 7361 4215 7395
rect 4801 7395 4859 7401
rect 4157 7355 4215 7361
rect 4356 7364 4752 7392
rect 3513 7327 3571 7333
rect 3513 7293 3525 7327
rect 3559 7293 3571 7327
rect 3513 7287 3571 7293
rect 3697 7327 3755 7333
rect 3697 7293 3709 7327
rect 3743 7293 3755 7327
rect 4062 7324 4068 7336
rect 4023 7296 4068 7324
rect 3697 7287 3755 7293
rect 845 7191 903 7197
rect 845 7157 857 7191
rect 891 7188 903 7191
rect 1026 7188 1032 7200
rect 891 7160 1032 7188
rect 891 7157 903 7160
rect 845 7151 903 7157
rect 1026 7148 1032 7160
rect 1084 7148 1090 7200
rect 1146 7188 1174 7284
rect 1762 7216 1768 7268
rect 1820 7256 1826 7268
rect 3712 7256 3740 7287
rect 4062 7284 4068 7296
rect 4120 7284 4126 7336
rect 4246 7284 4252 7336
rect 4304 7324 4310 7336
rect 4356 7333 4384 7364
rect 4341 7327 4399 7333
rect 4341 7324 4353 7327
rect 4304 7296 4353 7324
rect 4304 7284 4310 7296
rect 4341 7293 4353 7296
rect 4387 7293 4399 7327
rect 4341 7287 4399 7293
rect 4430 7284 4436 7336
rect 4488 7324 4494 7336
rect 4617 7327 4675 7333
rect 4617 7324 4629 7327
rect 4488 7296 4629 7324
rect 4488 7284 4494 7296
rect 4617 7293 4629 7296
rect 4663 7293 4675 7327
rect 4724 7324 4752 7364
rect 4801 7361 4813 7395
rect 4847 7361 4859 7395
rect 4801 7355 4859 7361
rect 5276 7333 5304 7500
rect 5350 7488 5356 7540
rect 5408 7528 5414 7540
rect 7006 7528 7012 7540
rect 5408 7500 7012 7528
rect 5408 7488 5414 7500
rect 4985 7327 5043 7333
rect 4985 7324 4997 7327
rect 4724 7296 4997 7324
rect 4617 7287 4675 7293
rect 4985 7293 4997 7296
rect 5031 7293 5043 7327
rect 4985 7287 5043 7293
rect 5261 7327 5319 7333
rect 5261 7293 5273 7327
rect 5307 7293 5319 7327
rect 5534 7324 5540 7336
rect 5495 7296 5540 7324
rect 5261 7287 5319 7293
rect 5534 7284 5540 7296
rect 5592 7284 5598 7336
rect 6104 7333 6132 7500
rect 7006 7488 7012 7500
rect 7064 7488 7070 7540
rect 7650 7488 7656 7540
rect 7708 7528 7714 7540
rect 8297 7531 8355 7537
rect 8297 7528 8309 7531
rect 7708 7500 8309 7528
rect 7708 7488 7714 7500
rect 8297 7497 8309 7500
rect 8343 7497 8355 7531
rect 10134 7528 10140 7540
rect 8297 7491 8355 7497
rect 8404 7500 10140 7528
rect 8404 7460 8432 7500
rect 10134 7488 10140 7500
rect 10192 7488 10198 7540
rect 11330 7528 11336 7540
rect 11291 7500 11336 7528
rect 11330 7488 11336 7500
rect 11388 7488 11394 7540
rect 12986 7488 12992 7540
rect 13044 7528 13050 7540
rect 13081 7531 13139 7537
rect 13081 7528 13093 7531
rect 13044 7500 13093 7528
rect 13044 7488 13050 7500
rect 13081 7497 13093 7500
rect 13127 7497 13139 7531
rect 13081 7491 13139 7497
rect 16574 7488 16580 7540
rect 16632 7528 16638 7540
rect 18506 7528 18512 7540
rect 16632 7500 18512 7528
rect 16632 7488 16638 7500
rect 18506 7488 18512 7500
rect 18564 7488 18570 7540
rect 8220 7432 8432 7460
rect 6273 7395 6331 7401
rect 6273 7361 6285 7395
rect 6319 7392 6331 7395
rect 6546 7392 6552 7404
rect 6319 7364 6552 7392
rect 6319 7361 6331 7364
rect 6273 7355 6331 7361
rect 6546 7352 6552 7364
rect 6604 7352 6610 7404
rect 7650 7352 7656 7404
rect 7708 7392 7714 7404
rect 8220 7401 8248 7432
rect 8938 7420 8944 7472
rect 8996 7460 9002 7472
rect 8996 7432 9674 7460
rect 8996 7420 9002 7432
rect 8205 7395 8263 7401
rect 8205 7392 8217 7395
rect 7708 7364 8217 7392
rect 7708 7352 7714 7364
rect 8205 7361 8217 7364
rect 8251 7361 8263 7395
rect 8205 7355 8263 7361
rect 8389 7395 8447 7401
rect 8389 7361 8401 7395
rect 8435 7392 8447 7395
rect 9398 7392 9404 7404
rect 8435 7364 9076 7392
rect 9359 7364 9404 7392
rect 8435 7361 8447 7364
rect 8389 7355 8447 7361
rect 9048 7336 9076 7364
rect 9398 7352 9404 7364
rect 9456 7352 9462 7404
rect 9646 7392 9674 7432
rect 9766 7420 9772 7472
rect 9824 7460 9830 7472
rect 14366 7460 14372 7472
rect 9824 7432 14372 7460
rect 9824 7420 9830 7432
rect 14366 7420 14372 7432
rect 14424 7460 14430 7472
rect 14737 7463 14795 7469
rect 14737 7460 14749 7463
rect 14424 7432 14749 7460
rect 14424 7420 14430 7432
rect 14737 7429 14749 7432
rect 14783 7429 14795 7463
rect 14737 7423 14795 7429
rect 15010 7420 15016 7472
rect 15068 7460 15074 7472
rect 18322 7460 18328 7472
rect 15068 7432 16068 7460
rect 18283 7432 18328 7460
rect 15068 7420 15074 7432
rect 10321 7395 10379 7401
rect 10321 7392 10333 7395
rect 9646 7364 10333 7392
rect 10321 7361 10333 7364
rect 10367 7392 10379 7395
rect 11790 7392 11796 7404
rect 10367 7364 11796 7392
rect 10367 7361 10379 7364
rect 10321 7355 10379 7361
rect 11790 7352 11796 7364
rect 11848 7352 11854 7404
rect 15838 7392 15844 7404
rect 12820 7364 15844 7392
rect 6089 7327 6147 7333
rect 6089 7293 6101 7327
rect 6135 7293 6147 7327
rect 6638 7324 6644 7336
rect 6599 7296 6644 7324
rect 6089 7287 6147 7293
rect 6638 7284 6644 7296
rect 6696 7284 6702 7336
rect 8067 7327 8125 7333
rect 8067 7293 8079 7327
rect 8113 7324 8125 7327
rect 8481 7327 8539 7333
rect 8481 7324 8493 7327
rect 8113 7296 8493 7324
rect 8113 7293 8125 7296
rect 8067 7287 8125 7293
rect 8481 7293 8493 7296
rect 8527 7324 8539 7327
rect 8846 7324 8852 7336
rect 8527 7296 8852 7324
rect 8527 7293 8539 7296
rect 8481 7287 8539 7293
rect 8846 7284 8852 7296
rect 8904 7284 8910 7336
rect 9030 7324 9036 7336
rect 8991 7296 9036 7324
rect 9030 7284 9036 7296
rect 9088 7284 9094 7336
rect 9585 7327 9643 7333
rect 9585 7293 9597 7327
rect 9631 7324 9643 7327
rect 10410 7324 10416 7336
rect 9631 7296 10416 7324
rect 9631 7293 9643 7296
rect 9585 7287 9643 7293
rect 10410 7284 10416 7296
rect 10468 7284 10474 7336
rect 12820 7333 12848 7364
rect 15838 7352 15844 7364
rect 15896 7352 15902 7404
rect 16040 7392 16068 7432
rect 18322 7420 18328 7432
rect 18380 7420 18386 7472
rect 17218 7392 17224 7404
rect 16040 7364 17224 7392
rect 12805 7327 12863 7333
rect 12805 7293 12817 7327
rect 12851 7293 12863 7327
rect 13262 7324 13268 7336
rect 13223 7296 13268 7324
rect 12805 7287 12863 7293
rect 13262 7284 13268 7296
rect 13320 7284 13326 7336
rect 13372 7296 14504 7324
rect 5166 7256 5172 7268
rect 1820 7228 1865 7256
rect 3252 7228 3740 7256
rect 3804 7228 5172 7256
rect 1820 7216 1826 7228
rect 2774 7188 2780 7200
rect 1146 7160 2780 7188
rect 2774 7148 2780 7160
rect 2832 7188 2838 7200
rect 3252 7197 3280 7228
rect 3237 7191 3295 7197
rect 3237 7188 3249 7191
rect 2832 7160 3249 7188
rect 2832 7148 2838 7160
rect 3237 7157 3249 7160
rect 3283 7157 3295 7191
rect 3237 7151 3295 7157
rect 3418 7148 3424 7200
rect 3476 7188 3482 7200
rect 3605 7191 3663 7197
rect 3605 7188 3617 7191
rect 3476 7160 3617 7188
rect 3476 7148 3482 7160
rect 3605 7157 3617 7160
rect 3651 7188 3663 7191
rect 3804 7188 3832 7228
rect 5166 7216 5172 7228
rect 5224 7216 5230 7268
rect 5810 7256 5816 7268
rect 5771 7228 5816 7256
rect 5810 7216 5816 7228
rect 5868 7216 5874 7268
rect 6932 7228 7038 7256
rect 3970 7188 3976 7200
rect 3651 7160 3832 7188
rect 3883 7160 3976 7188
rect 3651 7157 3663 7160
rect 3605 7151 3663 7157
rect 3970 7148 3976 7160
rect 4028 7188 4034 7200
rect 4982 7188 4988 7200
rect 4028 7160 4988 7188
rect 4028 7148 4034 7160
rect 4982 7148 4988 7160
rect 5040 7148 5046 7200
rect 5258 7148 5264 7200
rect 5316 7188 5322 7200
rect 6932 7188 6960 7228
rect 8294 7216 8300 7268
rect 8352 7256 8358 7268
rect 8665 7259 8723 7265
rect 8665 7256 8677 7259
rect 8352 7228 8677 7256
rect 8352 7216 8358 7228
rect 8665 7225 8677 7228
rect 8711 7256 8723 7259
rect 9490 7256 9496 7268
rect 8711 7228 9496 7256
rect 8711 7225 8723 7228
rect 8665 7219 8723 7225
rect 9490 7216 9496 7228
rect 9548 7256 9554 7268
rect 9677 7259 9735 7265
rect 9677 7256 9689 7259
rect 9548 7228 9689 7256
rect 9548 7216 9554 7228
rect 9677 7225 9689 7228
rect 9723 7225 9735 7259
rect 10505 7259 10563 7265
rect 10505 7256 10517 7259
rect 9677 7219 9735 7225
rect 10060 7228 10517 7256
rect 10060 7197 10088 7228
rect 10505 7225 10517 7228
rect 10551 7225 10563 7259
rect 10505 7219 10563 7225
rect 12989 7259 13047 7265
rect 12989 7225 13001 7259
rect 13035 7225 13047 7259
rect 12989 7219 13047 7225
rect 13173 7259 13231 7265
rect 13173 7225 13185 7259
rect 13219 7256 13231 7259
rect 13372 7256 13400 7296
rect 13219 7228 13400 7256
rect 13219 7225 13231 7228
rect 13173 7219 13231 7225
rect 5316 7160 6960 7188
rect 10045 7191 10103 7197
rect 5316 7148 5322 7160
rect 10045 7157 10057 7191
rect 10091 7157 10103 7191
rect 10045 7151 10103 7157
rect 10873 7191 10931 7197
rect 10873 7157 10885 7191
rect 10919 7188 10931 7191
rect 11698 7188 11704 7200
rect 10919 7160 11704 7188
rect 10919 7157 10931 7160
rect 10873 7151 10931 7157
rect 11698 7148 11704 7160
rect 11756 7148 11762 7200
rect 13004 7188 13032 7219
rect 13446 7216 13452 7268
rect 13504 7256 13510 7268
rect 14476 7256 14504 7296
rect 15010 7284 15016 7336
rect 15068 7324 15074 7336
rect 15289 7327 15347 7333
rect 15289 7324 15301 7327
rect 15068 7296 15301 7324
rect 15068 7284 15074 7296
rect 15289 7293 15301 7296
rect 15335 7293 15347 7327
rect 15289 7287 15347 7293
rect 15443 7327 15501 7333
rect 15443 7293 15455 7327
rect 15489 7324 15501 7327
rect 15930 7324 15936 7336
rect 15489 7296 15936 7324
rect 15489 7293 15501 7296
rect 15443 7287 15501 7293
rect 15930 7284 15936 7296
rect 15988 7284 15994 7336
rect 16040 7333 16068 7364
rect 17218 7352 17224 7364
rect 17276 7352 17282 7404
rect 16040 7327 16113 7333
rect 16040 7296 16067 7327
rect 16055 7293 16067 7296
rect 16101 7293 16113 7327
rect 16206 7324 16212 7336
rect 16167 7296 16212 7324
rect 16055 7287 16113 7293
rect 16206 7284 16212 7296
rect 16264 7284 16270 7336
rect 16301 7327 16359 7333
rect 16301 7293 16313 7327
rect 16347 7293 16359 7327
rect 18506 7324 18512 7336
rect 18467 7296 18512 7324
rect 16301 7287 16359 7293
rect 15841 7259 15899 7265
rect 15841 7256 15853 7259
rect 13504 7228 13549 7256
rect 14476 7228 15853 7256
rect 13504 7216 13510 7228
rect 15841 7225 15853 7228
rect 15887 7225 15899 7259
rect 16316 7256 16344 7287
rect 18506 7284 18512 7296
rect 18564 7284 18570 7336
rect 15841 7219 15899 7225
rect 16224 7228 16344 7256
rect 16577 7259 16635 7265
rect 16224 7200 16252 7228
rect 16577 7225 16589 7259
rect 16623 7256 16635 7259
rect 16666 7256 16672 7268
rect 16623 7228 16672 7256
rect 16623 7225 16635 7228
rect 16577 7219 16635 7225
rect 16666 7216 16672 7228
rect 16724 7216 16730 7268
rect 16776 7228 17066 7256
rect 14734 7188 14740 7200
rect 13004 7160 14740 7188
rect 14734 7148 14740 7160
rect 14792 7148 14798 7200
rect 15657 7191 15715 7197
rect 15657 7157 15669 7191
rect 15703 7188 15715 7191
rect 15746 7188 15752 7200
rect 15703 7160 15752 7188
rect 15703 7157 15715 7160
rect 15657 7151 15715 7157
rect 15746 7148 15752 7160
rect 15804 7148 15810 7200
rect 16206 7148 16212 7200
rect 16264 7148 16270 7200
rect 16390 7148 16396 7200
rect 16448 7188 16454 7200
rect 16776 7188 16804 7228
rect 16448 7160 16804 7188
rect 18049 7191 18107 7197
rect 16448 7148 16454 7160
rect 18049 7157 18061 7191
rect 18095 7188 18107 7191
rect 18322 7188 18328 7200
rect 18095 7160 18328 7188
rect 18095 7157 18107 7160
rect 18049 7151 18107 7157
rect 18322 7148 18328 7160
rect 18380 7148 18386 7200
rect 184 7098 18860 7120
rect 184 7046 4660 7098
rect 4712 7046 4724 7098
rect 4776 7046 4788 7098
rect 4840 7046 4852 7098
rect 4904 7046 4916 7098
rect 4968 7046 7760 7098
rect 7812 7046 7824 7098
rect 7876 7046 7888 7098
rect 7940 7046 7952 7098
rect 8004 7046 8016 7098
rect 8068 7046 10860 7098
rect 10912 7046 10924 7098
rect 10976 7046 10988 7098
rect 11040 7046 11052 7098
rect 11104 7046 11116 7098
rect 11168 7046 13960 7098
rect 14012 7046 14024 7098
rect 14076 7046 14088 7098
rect 14140 7046 14152 7098
rect 14204 7046 14216 7098
rect 14268 7046 17060 7098
rect 17112 7046 17124 7098
rect 17176 7046 17188 7098
rect 17240 7046 17252 7098
rect 17304 7046 17316 7098
rect 17368 7046 18860 7098
rect 184 7024 18860 7046
rect 474 6944 480 6996
rect 532 6984 538 6996
rect 661 6987 719 6993
rect 661 6984 673 6987
rect 532 6956 673 6984
rect 532 6944 538 6956
rect 661 6953 673 6956
rect 707 6953 719 6987
rect 661 6947 719 6953
rect 1765 6987 1823 6993
rect 1765 6953 1777 6987
rect 1811 6984 1823 6987
rect 2130 6984 2136 6996
rect 1811 6956 2136 6984
rect 1811 6953 1823 6956
rect 1765 6947 1823 6953
rect 2130 6944 2136 6956
rect 2188 6944 2194 6996
rect 2406 6984 2412 6996
rect 2367 6956 2412 6984
rect 2406 6944 2412 6956
rect 2464 6984 2470 6996
rect 3234 6984 3240 6996
rect 2464 6956 3240 6984
rect 2464 6944 2470 6956
rect 3234 6944 3240 6956
rect 3292 6944 3298 6996
rect 3326 6944 3332 6996
rect 3384 6984 3390 6996
rect 3881 6987 3939 6993
rect 3881 6984 3893 6987
rect 3384 6956 3893 6984
rect 3384 6944 3390 6956
rect 3881 6953 3893 6956
rect 3927 6953 3939 6987
rect 3881 6947 3939 6953
rect 4246 6944 4252 6996
rect 4304 6984 4310 6996
rect 4801 6987 4859 6993
rect 4801 6984 4813 6987
rect 4304 6956 4813 6984
rect 4304 6944 4310 6956
rect 4801 6953 4813 6956
rect 4847 6953 4859 6987
rect 4801 6947 4859 6953
rect 1305 6919 1363 6925
rect 1305 6885 1317 6919
rect 1351 6916 1363 6919
rect 1351 6888 1900 6916
rect 1351 6885 1363 6888
rect 1305 6879 1363 6885
rect 750 6848 756 6860
rect 711 6820 756 6848
rect 750 6808 756 6820
rect 808 6808 814 6860
rect 842 6808 848 6860
rect 900 6848 906 6860
rect 1121 6851 1179 6857
rect 900 6820 945 6848
rect 900 6808 906 6820
rect 1121 6817 1133 6851
rect 1167 6848 1179 6851
rect 1872 6848 1900 6888
rect 3050 6876 3056 6928
rect 3108 6916 3114 6928
rect 3108 6888 3153 6916
rect 3108 6876 3114 6888
rect 4154 6876 4160 6928
rect 4212 6916 4218 6928
rect 4341 6919 4399 6925
rect 4341 6916 4353 6919
rect 4212 6888 4353 6916
rect 4212 6876 4218 6888
rect 4341 6885 4353 6888
rect 4387 6885 4399 6919
rect 4816 6916 4844 6947
rect 4982 6944 4988 6996
rect 5040 6984 5046 6996
rect 6822 6984 6828 6996
rect 5040 6956 6828 6984
rect 5040 6944 5046 6956
rect 6822 6944 6828 6956
rect 6880 6944 6886 6996
rect 8665 6987 8723 6993
rect 8665 6984 8677 6987
rect 7208 6956 8677 6984
rect 7208 6928 7236 6956
rect 8665 6953 8677 6956
rect 8711 6953 8723 6987
rect 8665 6947 8723 6953
rect 8754 6944 8760 6996
rect 8812 6984 8818 6996
rect 9125 6987 9183 6993
rect 9125 6984 9137 6987
rect 8812 6956 9137 6984
rect 8812 6944 8818 6956
rect 9125 6953 9137 6956
rect 9171 6984 9183 6987
rect 9398 6984 9404 6996
rect 9171 6956 9404 6984
rect 9171 6953 9183 6956
rect 9125 6947 9183 6953
rect 9398 6944 9404 6956
rect 9456 6944 9462 6996
rect 9674 6944 9680 6996
rect 9732 6984 9738 6996
rect 10318 6984 10324 6996
rect 9732 6956 10324 6984
rect 9732 6944 9738 6956
rect 10318 6944 10324 6956
rect 10376 6944 10382 6996
rect 12894 6944 12900 6996
rect 12952 6984 12958 6996
rect 13814 6984 13820 6996
rect 12952 6956 13820 6984
rect 12952 6944 12958 6956
rect 13814 6944 13820 6956
rect 13872 6984 13878 6996
rect 14826 6984 14832 6996
rect 13872 6956 14832 6984
rect 13872 6944 13878 6956
rect 4816 6888 7144 6916
rect 4341 6879 4399 6885
rect 2958 6848 2964 6860
rect 1167 6820 1808 6848
rect 1872 6820 2964 6848
rect 1167 6817 1179 6820
rect 1121 6811 1179 6817
rect 1486 6780 1492 6792
rect 1399 6752 1492 6780
rect 1486 6740 1492 6752
rect 1544 6740 1550 6792
rect 1670 6780 1676 6792
rect 1631 6752 1676 6780
rect 1670 6740 1676 6752
rect 1728 6740 1734 6792
rect 1780 6780 1808 6820
rect 2958 6808 2964 6820
rect 3016 6808 3022 6860
rect 3145 6851 3203 6857
rect 3145 6817 3157 6851
rect 3191 6848 3203 6851
rect 3694 6848 3700 6860
rect 3191 6820 3700 6848
rect 3191 6817 3203 6820
rect 3145 6811 3203 6817
rect 3694 6808 3700 6820
rect 3752 6808 3758 6860
rect 4246 6848 4252 6860
rect 4207 6820 4252 6848
rect 4246 6808 4252 6820
rect 4304 6808 4310 6860
rect 6914 6808 6920 6860
rect 6972 6848 6978 6860
rect 7009 6851 7067 6857
rect 7009 6848 7021 6851
rect 6972 6820 7021 6848
rect 6972 6808 6978 6820
rect 7009 6817 7021 6820
rect 7055 6817 7067 6851
rect 7116 6848 7144 6888
rect 7190 6876 7196 6928
rect 7248 6916 7254 6928
rect 8938 6916 8944 6928
rect 7248 6888 7293 6916
rect 7944 6888 8944 6916
rect 7248 6876 7254 6888
rect 7944 6860 7972 6888
rect 8938 6876 8944 6888
rect 8996 6876 9002 6928
rect 10134 6916 10140 6928
rect 9324 6888 10140 6916
rect 7116 6820 7420 6848
rect 7009 6811 7067 6817
rect 2317 6783 2375 6789
rect 2317 6780 2329 6783
rect 1780 6752 2329 6780
rect 2317 6749 2329 6752
rect 2363 6780 2375 6783
rect 2682 6780 2688 6792
rect 2363 6752 2688 6780
rect 2363 6749 2375 6752
rect 2317 6743 2375 6749
rect 2682 6740 2688 6752
rect 2740 6740 2746 6792
rect 3237 6783 3295 6789
rect 3237 6772 3249 6783
rect 3160 6749 3249 6772
rect 3283 6749 3295 6783
rect 3160 6744 3295 6749
rect 1504 6712 1532 6740
rect 3160 6712 3188 6744
rect 3237 6743 3295 6744
rect 4062 6740 4068 6792
rect 4120 6780 4126 6792
rect 4522 6780 4528 6792
rect 4120 6752 4528 6780
rect 4120 6740 4126 6752
rect 4522 6740 4528 6752
rect 4580 6740 4586 6792
rect 5534 6740 5540 6792
rect 5592 6780 5598 6792
rect 7282 6780 7288 6792
rect 5592 6752 7288 6780
rect 5592 6740 5598 6752
rect 7282 6740 7288 6752
rect 7340 6740 7346 6792
rect 7392 6780 7420 6820
rect 7558 6808 7564 6860
rect 7616 6848 7622 6860
rect 7653 6851 7711 6857
rect 7653 6848 7665 6851
rect 7616 6820 7665 6848
rect 7616 6808 7622 6820
rect 7653 6817 7665 6820
rect 7699 6817 7711 6851
rect 7834 6848 7840 6860
rect 7795 6820 7840 6848
rect 7653 6811 7711 6817
rect 7834 6808 7840 6820
rect 7892 6808 7898 6860
rect 7926 6808 7932 6860
rect 7984 6848 7990 6860
rect 8113 6851 8171 6857
rect 7984 6820 8029 6848
rect 7984 6808 7990 6820
rect 8113 6817 8125 6851
rect 8159 6848 8171 6851
rect 8386 6848 8392 6860
rect 8159 6820 8392 6848
rect 8159 6817 8171 6820
rect 8113 6811 8171 6817
rect 8386 6808 8392 6820
rect 8444 6808 8450 6860
rect 8570 6848 8576 6860
rect 8531 6820 8576 6848
rect 8570 6808 8576 6820
rect 8628 6808 8634 6860
rect 8846 6808 8852 6860
rect 8904 6848 8910 6860
rect 9125 6851 9183 6857
rect 9125 6848 9137 6851
rect 8904 6820 9137 6848
rect 8904 6808 8910 6820
rect 9125 6817 9137 6820
rect 9171 6848 9183 6851
rect 9214 6848 9220 6860
rect 9171 6820 9220 6848
rect 9171 6817 9183 6820
rect 9125 6811 9183 6817
rect 9214 6808 9220 6820
rect 9272 6808 9278 6860
rect 9324 6857 9352 6888
rect 10134 6876 10140 6888
rect 10192 6876 10198 6928
rect 12158 6876 12164 6928
rect 12216 6916 12222 6928
rect 12216 6888 12742 6916
rect 12216 6876 12222 6888
rect 9309 6851 9367 6857
rect 9309 6817 9321 6851
rect 9355 6817 9367 6851
rect 9490 6848 9496 6860
rect 9451 6820 9496 6848
rect 9309 6811 9367 6817
rect 9490 6808 9496 6820
rect 9548 6808 9554 6860
rect 9858 6848 9864 6860
rect 9819 6820 9864 6848
rect 9858 6808 9864 6820
rect 9916 6808 9922 6860
rect 11609 6851 11667 6857
rect 11609 6817 11621 6851
rect 11655 6848 11667 6851
rect 11882 6848 11888 6860
rect 11655 6820 11888 6848
rect 11655 6817 11667 6820
rect 11609 6811 11667 6817
rect 11882 6808 11888 6820
rect 11940 6808 11946 6860
rect 14200 6857 14228 6956
rect 14826 6944 14832 6956
rect 14884 6984 14890 6996
rect 16206 6984 16212 6996
rect 14884 6956 16212 6984
rect 14884 6944 14890 6956
rect 16206 6944 16212 6956
rect 16264 6984 16270 6996
rect 16853 6987 16911 6993
rect 16264 6956 16712 6984
rect 16264 6944 16270 6956
rect 15010 6916 15016 6928
rect 14844 6888 15016 6916
rect 14844 6860 14872 6888
rect 15010 6876 15016 6888
rect 15068 6876 15074 6928
rect 15102 6876 15108 6928
rect 15160 6876 15166 6928
rect 15286 6876 15292 6928
rect 15344 6916 15350 6928
rect 15381 6919 15439 6925
rect 15381 6916 15393 6919
rect 15344 6888 15393 6916
rect 15344 6876 15350 6888
rect 15381 6885 15393 6888
rect 15427 6885 15439 6919
rect 15381 6879 15439 6885
rect 16390 6876 16396 6928
rect 16448 6876 16454 6928
rect 11977 6851 12035 6857
rect 11977 6817 11989 6851
rect 12023 6848 12035 6851
rect 14185 6851 14243 6857
rect 12023 6820 12388 6848
rect 12023 6817 12035 6820
rect 11977 6811 12035 6817
rect 7745 6783 7803 6789
rect 7745 6780 7757 6783
rect 7392 6752 7757 6780
rect 7745 6749 7757 6752
rect 7791 6749 7803 6783
rect 7745 6743 7803 6749
rect 7852 6752 8708 6780
rect 1504 6684 3188 6712
rect 3789 6715 3847 6721
rect 3789 6681 3801 6715
rect 3835 6712 3847 6715
rect 3970 6712 3976 6724
rect 3835 6684 3976 6712
rect 3835 6681 3847 6684
rect 3789 6675 3847 6681
rect 3970 6672 3976 6684
rect 4028 6712 4034 6724
rect 4614 6712 4620 6724
rect 4028 6684 4620 6712
rect 4028 6672 4034 6684
rect 4614 6672 4620 6684
rect 4672 6712 4678 6724
rect 5721 6715 5779 6721
rect 4672 6684 5212 6712
rect 4672 6672 4678 6684
rect 937 6647 995 6653
rect 937 6613 949 6647
rect 983 6644 995 6647
rect 1118 6644 1124 6656
rect 983 6616 1124 6644
rect 983 6613 995 6616
rect 937 6607 995 6613
rect 1118 6604 1124 6616
rect 1176 6604 1182 6656
rect 1854 6604 1860 6656
rect 1912 6644 1918 6656
rect 2133 6647 2191 6653
rect 2133 6644 2145 6647
rect 1912 6616 2145 6644
rect 1912 6604 1918 6616
rect 2133 6613 2145 6616
rect 2179 6613 2191 6647
rect 2133 6607 2191 6613
rect 2685 6647 2743 6653
rect 2685 6613 2697 6647
rect 2731 6644 2743 6647
rect 2958 6644 2964 6656
rect 2731 6616 2964 6644
rect 2731 6613 2743 6616
rect 2685 6607 2743 6613
rect 2958 6604 2964 6616
rect 3016 6604 3022 6656
rect 3234 6604 3240 6656
rect 3292 6644 3298 6656
rect 3513 6647 3571 6653
rect 3513 6644 3525 6647
rect 3292 6616 3525 6644
rect 3292 6604 3298 6616
rect 3513 6613 3525 6616
rect 3559 6644 3571 6647
rect 4338 6644 4344 6656
rect 3559 6616 4344 6644
rect 3559 6613 3571 6616
rect 3513 6607 3571 6613
rect 4338 6604 4344 6616
rect 4396 6604 4402 6656
rect 5184 6653 5212 6684
rect 5721 6681 5733 6715
rect 5767 6712 5779 6715
rect 7006 6712 7012 6724
rect 5767 6684 7012 6712
rect 5767 6681 5779 6684
rect 5721 6675 5779 6681
rect 7006 6672 7012 6684
rect 7064 6672 7070 6724
rect 7374 6712 7380 6724
rect 7116 6684 7380 6712
rect 5169 6647 5227 6653
rect 5169 6613 5181 6647
rect 5215 6644 5227 6647
rect 5258 6644 5264 6656
rect 5215 6616 5264 6644
rect 5215 6613 5227 6616
rect 5169 6607 5227 6613
rect 5258 6604 5264 6616
rect 5316 6604 5322 6656
rect 6914 6604 6920 6656
rect 6972 6644 6978 6656
rect 7116 6644 7144 6684
rect 7374 6672 7380 6684
rect 7432 6712 7438 6724
rect 7650 6712 7656 6724
rect 7432 6684 7656 6712
rect 7432 6672 7438 6684
rect 7650 6672 7656 6684
rect 7708 6712 7714 6724
rect 7852 6712 7880 6752
rect 8205 6715 8263 6721
rect 8205 6712 8217 6715
rect 7708 6684 7880 6712
rect 7944 6684 8217 6712
rect 7708 6672 7714 6684
rect 6972 6616 7144 6644
rect 6972 6604 6978 6616
rect 7282 6604 7288 6656
rect 7340 6644 7346 6656
rect 7944 6644 7972 6684
rect 8205 6681 8217 6684
rect 8251 6681 8263 6715
rect 8680 6712 8708 6752
rect 8754 6740 8760 6792
rect 8812 6780 8818 6792
rect 9766 6780 9772 6792
rect 8812 6752 8857 6780
rect 9600 6752 9772 6780
rect 8812 6740 8818 6752
rect 9600 6712 9628 6752
rect 9766 6740 9772 6752
rect 9824 6740 9830 6792
rect 11698 6780 11704 6792
rect 11659 6752 11704 6780
rect 11698 6740 11704 6752
rect 11756 6740 11762 6792
rect 11790 6740 11796 6792
rect 11848 6780 11854 6792
rect 11992 6780 12020 6811
rect 11848 6752 12020 6780
rect 11848 6740 11854 6752
rect 12360 6721 12388 6820
rect 14185 6817 14197 6851
rect 14231 6817 14243 6851
rect 14185 6811 14243 6817
rect 14277 6851 14335 6857
rect 14277 6817 14289 6851
rect 14323 6817 14335 6851
rect 14277 6811 14335 6817
rect 14461 6851 14519 6857
rect 14461 6817 14473 6851
rect 14507 6848 14519 6851
rect 14642 6848 14648 6860
rect 14507 6820 14648 6848
rect 14507 6817 14519 6820
rect 14461 6811 14519 6817
rect 12437 6783 12495 6789
rect 12437 6749 12449 6783
rect 12483 6780 12495 6783
rect 12710 6780 12716 6792
rect 12483 6752 12716 6780
rect 12483 6749 12495 6752
rect 12437 6743 12495 6749
rect 12710 6740 12716 6752
rect 12768 6740 12774 6792
rect 13446 6780 13452 6792
rect 12912 6752 13452 6780
rect 8680 6684 9628 6712
rect 12345 6715 12403 6721
rect 8205 6675 8263 6681
rect 12345 6681 12357 6715
rect 12391 6712 12403 6715
rect 12912 6712 12940 6752
rect 13446 6740 13452 6752
rect 13504 6740 13510 6792
rect 13538 6740 13544 6792
rect 13596 6780 13602 6792
rect 13909 6783 13967 6789
rect 13909 6780 13921 6783
rect 13596 6752 13921 6780
rect 13596 6740 13602 6752
rect 13909 6749 13921 6752
rect 13955 6749 13967 6783
rect 14292 6780 14320 6811
rect 14642 6808 14648 6820
rect 14700 6808 14706 6860
rect 14826 6857 14832 6860
rect 14799 6851 14832 6857
rect 14799 6817 14811 6851
rect 14799 6811 14832 6817
rect 14826 6808 14832 6811
rect 14884 6808 14890 6860
rect 15120 6848 15148 6876
rect 14936 6820 15148 6848
rect 14936 6792 14964 6820
rect 14918 6780 14924 6792
rect 14292 6752 14924 6780
rect 13909 6743 13967 6749
rect 14918 6740 14924 6752
rect 14976 6740 14982 6792
rect 15105 6783 15163 6789
rect 15105 6749 15117 6783
rect 15151 6749 15163 6783
rect 15105 6743 15163 6749
rect 12391 6684 12940 6712
rect 14277 6715 14335 6721
rect 12391 6681 12403 6684
rect 12345 6675 12403 6681
rect 14277 6681 14289 6715
rect 14323 6712 14335 6715
rect 14458 6712 14464 6724
rect 14323 6684 14464 6712
rect 14323 6681 14335 6684
rect 14277 6675 14335 6681
rect 14458 6672 14464 6684
rect 14516 6672 14522 6724
rect 15010 6712 15016 6724
rect 14971 6684 15016 6712
rect 15010 6672 15016 6684
rect 15068 6672 15074 6724
rect 7340 6616 7972 6644
rect 7340 6604 7346 6616
rect 8386 6604 8392 6656
rect 8444 6644 8450 6656
rect 8846 6644 8852 6656
rect 8444 6616 8852 6644
rect 8444 6604 8450 6616
rect 8846 6604 8852 6616
rect 8904 6604 8910 6656
rect 8938 6604 8944 6656
rect 8996 6644 9002 6656
rect 11793 6647 11851 6653
rect 11793 6644 11805 6647
rect 8996 6616 11805 6644
rect 8996 6604 9002 6616
rect 11793 6613 11805 6616
rect 11839 6613 11851 6647
rect 11793 6607 11851 6613
rect 11885 6647 11943 6653
rect 11885 6613 11897 6647
rect 11931 6644 11943 6647
rect 11974 6644 11980 6656
rect 11931 6616 11980 6644
rect 11931 6613 11943 6616
rect 11885 6607 11943 6613
rect 11974 6604 11980 6616
rect 12032 6604 12038 6656
rect 12710 6604 12716 6656
rect 12768 6644 12774 6656
rect 13722 6644 13728 6656
rect 12768 6616 13728 6644
rect 12768 6604 12774 6616
rect 13722 6604 13728 6616
rect 13780 6604 13786 6656
rect 13906 6604 13912 6656
rect 13964 6644 13970 6656
rect 15120 6644 15148 6743
rect 16114 6740 16120 6792
rect 16172 6780 16178 6792
rect 16684 6780 16712 6956
rect 16853 6953 16865 6987
rect 16899 6953 16911 6987
rect 16853 6947 16911 6953
rect 16868 6848 16896 6947
rect 16942 6848 16948 6860
rect 16868 6820 16948 6848
rect 16942 6808 16948 6820
rect 17000 6808 17006 6860
rect 17126 6808 17132 6860
rect 17184 6848 17190 6860
rect 17293 6851 17351 6857
rect 17293 6848 17305 6851
rect 17184 6820 17305 6848
rect 17184 6808 17190 6820
rect 17293 6817 17305 6820
rect 17339 6817 17351 6851
rect 17293 6811 17351 6817
rect 17037 6783 17095 6789
rect 17037 6780 17049 6783
rect 16172 6752 16436 6780
rect 16684 6752 17049 6780
rect 16172 6740 16178 6752
rect 16408 6712 16436 6752
rect 17037 6749 17049 6752
rect 17083 6749 17095 6783
rect 17037 6743 17095 6749
rect 16408 6684 16988 6712
rect 16850 6644 16856 6656
rect 13964 6616 16856 6644
rect 13964 6604 13970 6616
rect 16850 6604 16856 6616
rect 16908 6604 16914 6656
rect 16960 6644 16988 6684
rect 18417 6647 18475 6653
rect 18417 6644 18429 6647
rect 16960 6616 18429 6644
rect 18417 6613 18429 6616
rect 18463 6613 18475 6647
rect 18417 6607 18475 6613
rect 184 6554 18924 6576
rect 184 6502 3110 6554
rect 3162 6502 3174 6554
rect 3226 6502 3238 6554
rect 3290 6502 3302 6554
rect 3354 6502 3366 6554
rect 3418 6502 6210 6554
rect 6262 6502 6274 6554
rect 6326 6502 6338 6554
rect 6390 6502 6402 6554
rect 6454 6502 6466 6554
rect 6518 6502 9310 6554
rect 9362 6502 9374 6554
rect 9426 6502 9438 6554
rect 9490 6502 9502 6554
rect 9554 6502 9566 6554
rect 9618 6502 12410 6554
rect 12462 6502 12474 6554
rect 12526 6502 12538 6554
rect 12590 6502 12602 6554
rect 12654 6502 12666 6554
rect 12718 6502 15510 6554
rect 15562 6502 15574 6554
rect 15626 6502 15638 6554
rect 15690 6502 15702 6554
rect 15754 6502 15766 6554
rect 15818 6502 18610 6554
rect 18662 6502 18674 6554
rect 18726 6502 18738 6554
rect 18790 6502 18802 6554
rect 18854 6502 18866 6554
rect 18918 6502 18924 6554
rect 184 6480 18924 6502
rect 566 6440 572 6452
rect 527 6412 572 6440
rect 566 6400 572 6412
rect 624 6400 630 6452
rect 1670 6400 1676 6452
rect 1728 6440 1734 6452
rect 4433 6443 4491 6449
rect 4433 6440 4445 6443
rect 1728 6412 4445 6440
rect 1728 6400 1734 6412
rect 4433 6409 4445 6412
rect 4479 6409 4491 6443
rect 4433 6403 4491 6409
rect 5994 6400 6000 6452
rect 6052 6440 6058 6452
rect 6270 6440 6276 6452
rect 6052 6412 6276 6440
rect 6052 6400 6058 6412
rect 6270 6400 6276 6412
rect 6328 6400 6334 6452
rect 6822 6400 6828 6452
rect 6880 6440 6886 6452
rect 9674 6440 9680 6452
rect 6880 6412 9680 6440
rect 6880 6400 6886 6412
rect 9674 6400 9680 6412
rect 9732 6400 9738 6452
rect 11314 6443 11372 6449
rect 11314 6440 11326 6443
rect 9876 6412 11326 6440
rect 753 6375 811 6381
rect 753 6341 765 6375
rect 799 6372 811 6375
rect 1118 6372 1124 6384
rect 799 6344 1124 6372
rect 799 6341 811 6344
rect 753 6335 811 6341
rect 1118 6332 1124 6344
rect 1176 6332 1182 6384
rect 2866 6332 2872 6384
rect 2924 6372 2930 6384
rect 3050 6372 3056 6384
rect 2924 6344 3056 6372
rect 2924 6332 2930 6344
rect 3050 6332 3056 6344
rect 3108 6332 3114 6384
rect 3234 6372 3240 6384
rect 3195 6344 3240 6372
rect 3234 6332 3240 6344
rect 3292 6332 3298 6384
rect 4249 6375 4307 6381
rect 4249 6341 4261 6375
rect 4295 6372 4307 6375
rect 4522 6372 4528 6384
rect 4295 6344 4528 6372
rect 4295 6341 4307 6344
rect 4249 6335 4307 6341
rect 4522 6332 4528 6344
rect 4580 6372 4586 6384
rect 4580 6344 5120 6372
rect 4580 6332 4586 6344
rect 1210 6264 1216 6316
rect 1268 6304 1274 6316
rect 1854 6304 1860 6316
rect 1268 6276 1716 6304
rect 1815 6276 1860 6304
rect 1268 6264 1274 6276
rect 842 6236 848 6248
rect 803 6208 848 6236
rect 842 6196 848 6208
rect 900 6196 906 6248
rect 1026 6236 1032 6248
rect 987 6208 1032 6236
rect 1026 6196 1032 6208
rect 1084 6196 1090 6248
rect 1302 6236 1308 6248
rect 1263 6208 1308 6236
rect 1302 6196 1308 6208
rect 1360 6196 1366 6248
rect 1486 6236 1492 6248
rect 1447 6208 1492 6236
rect 1486 6196 1492 6208
rect 1544 6196 1550 6248
rect 1688 6236 1716 6276
rect 1854 6264 1860 6276
rect 1912 6264 1918 6316
rect 2038 6304 2044 6316
rect 1964 6276 2044 6304
rect 1964 6236 1992 6276
rect 2038 6264 2044 6276
rect 2096 6304 2102 6316
rect 5092 6313 5120 6344
rect 8662 6332 8668 6384
rect 8720 6332 8726 6384
rect 8846 6332 8852 6384
rect 8904 6372 8910 6384
rect 9876 6372 9904 6412
rect 11314 6409 11326 6412
rect 11360 6409 11372 6443
rect 11314 6403 11372 6409
rect 11882 6400 11888 6452
rect 11940 6440 11946 6452
rect 11940 6412 12434 6440
rect 11940 6400 11946 6412
rect 8904 6344 9904 6372
rect 12406 6372 12434 6412
rect 12710 6400 12716 6452
rect 12768 6440 12774 6452
rect 15378 6440 15384 6452
rect 12768 6412 15384 6440
rect 12768 6400 12774 6412
rect 15378 6400 15384 6412
rect 15436 6400 15442 6452
rect 15657 6443 15715 6449
rect 15657 6409 15669 6443
rect 15703 6440 15715 6443
rect 15930 6440 15936 6452
rect 15703 6412 15936 6440
rect 15703 6409 15715 6412
rect 15657 6403 15715 6409
rect 15930 6400 15936 6412
rect 15988 6440 15994 6452
rect 16482 6440 16488 6452
rect 15988 6412 16488 6440
rect 15988 6400 15994 6412
rect 16482 6400 16488 6412
rect 16540 6400 16546 6452
rect 16666 6400 16672 6452
rect 16724 6440 16730 6452
rect 17681 6443 17739 6449
rect 17681 6440 17693 6443
rect 16724 6412 17693 6440
rect 16724 6400 16730 6412
rect 17681 6409 17693 6412
rect 17727 6409 17739 6443
rect 17681 6403 17739 6409
rect 18046 6400 18052 6452
rect 18104 6440 18110 6452
rect 18233 6443 18291 6449
rect 18233 6440 18245 6443
rect 18104 6412 18245 6440
rect 18104 6400 18110 6412
rect 18233 6409 18245 6412
rect 18279 6409 18291 6443
rect 18233 6403 18291 6409
rect 12406 6344 13400 6372
rect 8904 6332 8910 6344
rect 5077 6307 5135 6313
rect 2096 6276 3556 6304
rect 2096 6264 2102 6276
rect 3528 6245 3556 6276
rect 5077 6273 5089 6307
rect 5123 6304 5135 6307
rect 5534 6304 5540 6316
rect 5123 6276 5540 6304
rect 5123 6273 5135 6276
rect 5077 6267 5135 6273
rect 5534 6264 5540 6276
rect 5592 6264 5598 6316
rect 5902 6304 5908 6316
rect 5863 6276 5908 6304
rect 5902 6264 5908 6276
rect 5960 6264 5966 6316
rect 7190 6304 7196 6316
rect 6104 6276 7196 6304
rect 1688 6208 1992 6236
rect 3513 6239 3571 6245
rect 3513 6205 3525 6239
rect 3559 6205 3571 6239
rect 3513 6199 3571 6205
rect 3602 6196 3608 6248
rect 3660 6196 3666 6248
rect 3970 6236 3976 6248
rect 3931 6208 3976 6236
rect 3970 6196 3976 6208
rect 4028 6196 4034 6248
rect 5721 6239 5779 6245
rect 5721 6205 5733 6239
rect 5767 6236 5779 6239
rect 6104 6236 6132 6276
rect 7190 6264 7196 6276
rect 7248 6264 7254 6316
rect 8202 6264 8208 6316
rect 8260 6304 8266 6316
rect 8481 6307 8539 6313
rect 8481 6304 8493 6307
rect 8260 6276 8493 6304
rect 8260 6264 8266 6276
rect 8481 6273 8493 6276
rect 8527 6273 8539 6307
rect 8481 6267 8539 6273
rect 6270 6236 6276 6248
rect 5767 6208 6132 6236
rect 6231 6208 6276 6236
rect 5767 6205 5779 6208
rect 5721 6199 5779 6205
rect 6270 6196 6276 6208
rect 6328 6196 6334 6248
rect 6365 6239 6423 6245
rect 6365 6205 6377 6239
rect 6411 6205 6423 6239
rect 6365 6199 6423 6205
rect 3620 6168 3648 6196
rect 2898 6140 3648 6168
rect 3878 6128 3884 6180
rect 3936 6168 3942 6180
rect 4893 6171 4951 6177
rect 3936 6140 4200 6168
rect 3936 6128 3942 6140
rect 1213 6103 1271 6109
rect 1213 6069 1225 6103
rect 1259 6100 1271 6103
rect 3605 6103 3663 6109
rect 3605 6100 3617 6103
rect 1259 6072 3617 6100
rect 1259 6069 1271 6072
rect 1213 6063 1271 6069
rect 3605 6069 3617 6072
rect 3651 6100 3663 6103
rect 4062 6100 4068 6112
rect 3651 6072 4068 6100
rect 3651 6069 3663 6072
rect 3605 6063 3663 6069
rect 4062 6060 4068 6072
rect 4120 6060 4126 6112
rect 4172 6100 4200 6140
rect 4893 6137 4905 6171
rect 4939 6168 4951 6171
rect 5626 6168 5632 6180
rect 4939 6140 5632 6168
rect 4939 6137 4951 6140
rect 4893 6131 4951 6137
rect 5626 6128 5632 6140
rect 5684 6128 5690 6180
rect 6086 6128 6092 6180
rect 6144 6168 6150 6180
rect 6380 6168 6408 6199
rect 6546 6196 6552 6248
rect 6604 6236 6610 6248
rect 6822 6236 6828 6248
rect 6604 6208 6828 6236
rect 6604 6196 6610 6208
rect 6822 6196 6828 6208
rect 6880 6196 6886 6248
rect 8680 6245 8708 6332
rect 11057 6307 11115 6313
rect 11057 6273 11069 6307
rect 11103 6304 11115 6307
rect 12894 6304 12900 6316
rect 11103 6276 12900 6304
rect 11103 6273 11115 6276
rect 11057 6267 11115 6273
rect 12894 6264 12900 6276
rect 12952 6264 12958 6316
rect 8665 6239 8723 6245
rect 8665 6205 8677 6239
rect 8711 6205 8723 6239
rect 8846 6236 8852 6248
rect 8807 6208 8852 6236
rect 8665 6199 8723 6205
rect 8846 6196 8852 6208
rect 8904 6196 8910 6248
rect 8956 6208 11100 6236
rect 6144 6140 6408 6168
rect 6144 6128 6150 6140
rect 7650 6128 7656 6180
rect 7708 6128 7714 6180
rect 8205 6171 8263 6177
rect 8205 6137 8217 6171
rect 8251 6168 8263 6171
rect 8956 6168 8984 6208
rect 9122 6168 9128 6180
rect 8251 6140 8984 6168
rect 9083 6140 9128 6168
rect 8251 6137 8263 6140
rect 8205 6131 8263 6137
rect 9122 6128 9128 6140
rect 9180 6128 9186 6180
rect 10689 6171 10747 6177
rect 10689 6137 10701 6171
rect 10735 6137 10747 6171
rect 11072 6168 11100 6208
rect 11422 6168 11428 6180
rect 11072 6140 11428 6168
rect 10689 6131 10747 6137
rect 4801 6103 4859 6109
rect 4801 6100 4813 6103
rect 4172 6072 4813 6100
rect 4801 6069 4813 6072
rect 4847 6069 4859 6103
rect 4801 6063 4859 6069
rect 4982 6060 4988 6112
rect 5040 6100 5046 6112
rect 5353 6103 5411 6109
rect 5353 6100 5365 6103
rect 5040 6072 5365 6100
rect 5040 6060 5046 6072
rect 5353 6069 5365 6072
rect 5399 6069 5411 6103
rect 5810 6100 5816 6112
rect 5771 6072 5816 6100
rect 5353 6063 5411 6069
rect 5810 6060 5816 6072
rect 5868 6060 5874 6112
rect 5994 6060 6000 6112
rect 6052 6100 6058 6112
rect 6273 6103 6331 6109
rect 6273 6100 6285 6103
rect 6052 6072 6285 6100
rect 6052 6060 6058 6072
rect 6273 6069 6285 6072
rect 6319 6069 6331 6103
rect 6273 6063 6331 6069
rect 6733 6103 6791 6109
rect 6733 6069 6745 6103
rect 6779 6100 6791 6103
rect 7374 6100 7380 6112
rect 6779 6072 7380 6100
rect 6779 6069 6791 6072
rect 6733 6063 6791 6069
rect 7374 6060 7380 6072
rect 7432 6060 7438 6112
rect 8849 6103 8907 6109
rect 8849 6069 8861 6103
rect 8895 6100 8907 6103
rect 9214 6100 9220 6112
rect 8895 6072 9220 6100
rect 8895 6069 8907 6072
rect 8849 6063 8907 6069
rect 9214 6060 9220 6072
rect 9272 6060 9278 6112
rect 10704 6100 10732 6131
rect 11422 6128 11428 6140
rect 11480 6128 11486 6180
rect 12066 6128 12072 6180
rect 12124 6128 12130 6180
rect 13078 6168 13084 6180
rect 13039 6140 13084 6168
rect 13078 6128 13084 6140
rect 13136 6128 13142 6180
rect 13265 6171 13323 6177
rect 13265 6137 13277 6171
rect 13311 6168 13323 6171
rect 13372 6168 13400 6344
rect 13446 6332 13452 6384
rect 13504 6372 13510 6384
rect 13725 6375 13783 6381
rect 13725 6372 13737 6375
rect 13504 6344 13737 6372
rect 13504 6332 13510 6344
rect 13725 6341 13737 6344
rect 13771 6372 13783 6375
rect 13771 6344 14044 6372
rect 13771 6341 13783 6344
rect 13725 6335 13783 6341
rect 13906 6304 13912 6316
rect 13867 6276 13912 6304
rect 13906 6264 13912 6276
rect 13964 6264 13970 6316
rect 14016 6304 14044 6344
rect 17862 6332 17868 6384
rect 17920 6372 17926 6384
rect 18414 6372 18420 6384
rect 17920 6344 18420 6372
rect 17920 6332 17926 6344
rect 18414 6332 18420 6344
rect 18472 6332 18478 6384
rect 14550 6304 14556 6316
rect 14016 6276 14556 6304
rect 14550 6264 14556 6276
rect 14608 6264 14614 6316
rect 16574 6304 16580 6316
rect 15488 6276 16580 6304
rect 14185 6171 14243 6177
rect 13311 6140 14136 6168
rect 13311 6137 13323 6140
rect 13265 6131 13323 6137
rect 10873 6103 10931 6109
rect 10873 6100 10885 6103
rect 10704 6072 10885 6100
rect 10873 6069 10885 6072
rect 10919 6100 10931 6103
rect 12710 6100 12716 6112
rect 10919 6072 12716 6100
rect 10919 6069 10931 6072
rect 10873 6063 10931 6069
rect 12710 6060 12716 6072
rect 12768 6060 12774 6112
rect 13538 6100 13544 6112
rect 13499 6072 13544 6100
rect 13538 6060 13544 6072
rect 13596 6060 13602 6112
rect 14108 6100 14136 6140
rect 14185 6137 14197 6171
rect 14231 6168 14243 6171
rect 14458 6168 14464 6180
rect 14231 6140 14464 6168
rect 14231 6137 14243 6140
rect 14185 6131 14243 6137
rect 14458 6128 14464 6140
rect 14516 6128 14522 6180
rect 14918 6128 14924 6180
rect 14976 6128 14982 6180
rect 15488 6100 15516 6276
rect 16574 6264 16580 6276
rect 16632 6264 16638 6316
rect 15841 6239 15899 6245
rect 15841 6205 15853 6239
rect 15887 6205 15899 6239
rect 17770 6236 17776 6248
rect 17250 6208 17776 6236
rect 15841 6199 15899 6205
rect 15856 6168 15884 6199
rect 17770 6196 17776 6208
rect 17828 6196 17834 6248
rect 17865 6239 17923 6245
rect 17865 6205 17877 6239
rect 17911 6236 17923 6239
rect 17954 6236 17960 6248
rect 17911 6208 17960 6236
rect 17911 6205 17923 6208
rect 17865 6199 17923 6205
rect 17954 6196 17960 6208
rect 18012 6196 18018 6248
rect 18417 6239 18475 6245
rect 18417 6205 18429 6239
rect 18463 6236 18475 6239
rect 18966 6236 18972 6248
rect 18463 6208 18972 6236
rect 18463 6205 18475 6208
rect 18417 6199 18475 6205
rect 16114 6168 16120 6180
rect 15856 6140 15976 6168
rect 16075 6140 16120 6168
rect 14108 6072 15516 6100
rect 15948 6100 15976 6140
rect 16114 6128 16120 6140
rect 16172 6128 16178 6180
rect 18046 6168 18052 6180
rect 17512 6140 17908 6168
rect 18007 6140 18052 6168
rect 16206 6100 16212 6112
rect 15948 6072 16212 6100
rect 16206 6060 16212 6072
rect 16264 6060 16270 6112
rect 16298 6060 16304 6112
rect 16356 6100 16362 6112
rect 17512 6100 17540 6140
rect 16356 6072 17540 6100
rect 17589 6103 17647 6109
rect 16356 6060 16362 6072
rect 17589 6069 17601 6103
rect 17635 6100 17647 6103
rect 17678 6100 17684 6112
rect 17635 6072 17684 6100
rect 17635 6069 17647 6072
rect 17589 6063 17647 6069
rect 17678 6060 17684 6072
rect 17736 6060 17742 6112
rect 17880 6100 17908 6140
rect 18046 6128 18052 6140
rect 18104 6128 18110 6180
rect 18432 6100 18460 6199
rect 18966 6196 18972 6208
rect 19024 6196 19030 6248
rect 17880 6072 18460 6100
rect 184 6010 18860 6032
rect 184 5958 4660 6010
rect 4712 5958 4724 6010
rect 4776 5958 4788 6010
rect 4840 5958 4852 6010
rect 4904 5958 4916 6010
rect 4968 5958 7760 6010
rect 7812 5958 7824 6010
rect 7876 5958 7888 6010
rect 7940 5958 7952 6010
rect 8004 5958 8016 6010
rect 8068 5958 10860 6010
rect 10912 5958 10924 6010
rect 10976 5958 10988 6010
rect 11040 5958 11052 6010
rect 11104 5958 11116 6010
rect 11168 5958 13960 6010
rect 14012 5958 14024 6010
rect 14076 5958 14088 6010
rect 14140 5958 14152 6010
rect 14204 5958 14216 6010
rect 14268 5958 17060 6010
rect 17112 5958 17124 6010
rect 17176 5958 17188 6010
rect 17240 5958 17252 6010
rect 17304 5958 17316 6010
rect 17368 5958 18860 6010
rect 184 5936 18860 5958
rect 1213 5899 1271 5905
rect 1213 5865 1225 5899
rect 1259 5896 1271 5899
rect 1486 5896 1492 5908
rect 1259 5868 1492 5896
rect 1259 5865 1271 5868
rect 1213 5859 1271 5865
rect 1486 5856 1492 5868
rect 1544 5856 1550 5908
rect 1578 5856 1584 5908
rect 1636 5856 1642 5908
rect 2501 5899 2559 5905
rect 2501 5865 2513 5899
rect 2547 5865 2559 5899
rect 2501 5859 2559 5865
rect 2777 5899 2835 5905
rect 2777 5865 2789 5899
rect 2823 5896 2835 5899
rect 3050 5896 3056 5908
rect 2823 5868 3056 5896
rect 2823 5865 2835 5868
rect 2777 5859 2835 5865
rect 1397 5831 1455 5837
rect 1397 5797 1409 5831
rect 1443 5828 1455 5831
rect 1596 5828 1624 5856
rect 2516 5828 2544 5859
rect 3050 5856 3056 5868
rect 3108 5856 3114 5908
rect 3510 5856 3516 5908
rect 3568 5896 3574 5908
rect 3878 5896 3884 5908
rect 3568 5868 3884 5896
rect 3568 5856 3574 5868
rect 3878 5856 3884 5868
rect 3936 5896 3942 5908
rect 5721 5899 5779 5905
rect 5721 5896 5733 5899
rect 3936 5868 5733 5896
rect 3936 5856 3942 5868
rect 5721 5865 5733 5868
rect 5767 5896 5779 5899
rect 6914 5896 6920 5908
rect 5767 5868 6920 5896
rect 5767 5865 5779 5868
rect 5721 5859 5779 5865
rect 6914 5856 6920 5868
rect 6972 5896 6978 5908
rect 8202 5896 8208 5908
rect 6972 5868 8208 5896
rect 6972 5856 6978 5868
rect 8202 5856 8208 5868
rect 8260 5856 8266 5908
rect 8570 5856 8576 5908
rect 8628 5896 8634 5908
rect 9033 5899 9091 5905
rect 9033 5896 9045 5899
rect 8628 5868 9045 5896
rect 8628 5856 8634 5868
rect 9033 5865 9045 5868
rect 9079 5865 9091 5899
rect 9033 5859 9091 5865
rect 9861 5899 9919 5905
rect 9861 5865 9873 5899
rect 9907 5896 9919 5899
rect 9950 5896 9956 5908
rect 9907 5868 9956 5896
rect 9907 5865 9919 5868
rect 9861 5859 9919 5865
rect 9950 5856 9956 5868
rect 10008 5856 10014 5908
rect 11348 5868 14412 5896
rect 3786 5828 3792 5840
rect 1443 5800 1624 5828
rect 1688 5800 2452 5828
rect 2516 5800 3792 5828
rect 1443 5797 1455 5800
rect 1397 5791 1455 5797
rect 1213 5763 1271 5769
rect 1213 5729 1225 5763
rect 1259 5760 1271 5763
rect 1486 5760 1492 5772
rect 1259 5732 1492 5760
rect 1259 5729 1271 5732
rect 1213 5723 1271 5729
rect 1486 5720 1492 5732
rect 1544 5720 1550 5772
rect 1688 5769 1716 5800
rect 1581 5763 1639 5769
rect 1581 5729 1593 5763
rect 1627 5729 1639 5763
rect 1581 5723 1639 5729
rect 1673 5763 1731 5769
rect 1673 5729 1685 5763
rect 1719 5729 1731 5763
rect 1673 5723 1731 5729
rect 1765 5763 1823 5769
rect 1765 5729 1777 5763
rect 1811 5729 1823 5763
rect 2130 5760 2136 5772
rect 2091 5732 2136 5760
rect 1765 5723 1823 5729
rect 934 5652 940 5704
rect 992 5692 998 5704
rect 1596 5692 1624 5723
rect 992 5664 1624 5692
rect 992 5652 998 5664
rect 1780 5624 1808 5723
rect 2130 5720 2136 5732
rect 2188 5720 2194 5772
rect 2424 5760 2452 5800
rect 3786 5788 3792 5800
rect 3844 5788 3850 5840
rect 4062 5828 4068 5840
rect 4023 5800 4068 5828
rect 4062 5788 4068 5800
rect 4120 5788 4126 5840
rect 4157 5831 4215 5837
rect 4157 5797 4169 5831
rect 4203 5797 4215 5831
rect 4157 5791 4215 5797
rect 2590 5760 2596 5772
rect 2424 5732 2596 5760
rect 2590 5720 2596 5732
rect 2648 5720 2654 5772
rect 2774 5720 2780 5772
rect 2832 5760 2838 5772
rect 3145 5763 3203 5769
rect 3145 5760 3157 5763
rect 2832 5732 3157 5760
rect 2832 5720 2838 5732
rect 3145 5729 3157 5732
rect 3191 5729 3203 5763
rect 4172 5760 4200 5791
rect 4338 5788 4344 5840
rect 4396 5828 4402 5840
rect 4617 5831 4675 5837
rect 4617 5828 4629 5831
rect 4396 5800 4629 5828
rect 4396 5788 4402 5800
rect 4617 5797 4629 5800
rect 4663 5797 4675 5831
rect 4617 5791 4675 5797
rect 7009 5831 7067 5837
rect 7009 5797 7021 5831
rect 7055 5828 7067 5831
rect 9122 5828 9128 5840
rect 7055 5800 9128 5828
rect 7055 5797 7067 5800
rect 7009 5791 7067 5797
rect 9122 5788 9128 5800
rect 9180 5788 9186 5840
rect 9674 5828 9680 5840
rect 9232 5800 9680 5828
rect 4172 5732 4844 5760
rect 3145 5723 3203 5729
rect 2038 5692 2044 5704
rect 1999 5664 2044 5692
rect 2038 5652 2044 5664
rect 2096 5652 2102 5704
rect 2222 5692 2228 5704
rect 2148 5664 2228 5692
rect 2148 5624 2176 5664
rect 2222 5652 2228 5664
rect 2280 5692 2286 5704
rect 4341 5695 4399 5701
rect 4341 5692 4353 5695
rect 2280 5664 4353 5692
rect 2280 5652 2286 5664
rect 4341 5661 4353 5664
rect 4387 5692 4399 5695
rect 4522 5692 4528 5704
rect 4387 5664 4528 5692
rect 4387 5661 4399 5664
rect 4341 5655 4399 5661
rect 4522 5652 4528 5664
rect 4580 5652 4586 5704
rect 3694 5624 3700 5636
rect 1780 5596 2176 5624
rect 3655 5596 3700 5624
rect 3694 5584 3700 5596
rect 3752 5584 3758 5636
rect 4816 5624 4844 5732
rect 5810 5720 5816 5772
rect 5868 5760 5874 5772
rect 7101 5763 7159 5769
rect 7101 5760 7113 5763
rect 5868 5732 7113 5760
rect 5868 5720 5874 5732
rect 7101 5729 7113 5732
rect 7147 5729 7159 5763
rect 7101 5723 7159 5729
rect 7285 5763 7343 5769
rect 7285 5729 7297 5763
rect 7331 5760 7343 5763
rect 7374 5760 7380 5772
rect 7331 5732 7380 5760
rect 7331 5729 7343 5732
rect 7285 5723 7343 5729
rect 5169 5695 5227 5701
rect 5169 5661 5181 5695
rect 5215 5692 5227 5695
rect 5902 5692 5908 5704
rect 5215 5664 5908 5692
rect 5215 5661 5227 5664
rect 5169 5655 5227 5661
rect 5902 5652 5908 5664
rect 5960 5692 5966 5704
rect 6270 5692 6276 5704
rect 5960 5664 6276 5692
rect 5960 5652 5966 5664
rect 6270 5652 6276 5664
rect 6328 5652 6334 5704
rect 7116 5692 7144 5723
rect 7374 5720 7380 5732
rect 7432 5760 7438 5772
rect 7653 5763 7711 5769
rect 7653 5760 7665 5763
rect 7432 5732 7665 5760
rect 7432 5720 7438 5732
rect 7653 5729 7665 5732
rect 7699 5760 7711 5763
rect 7742 5760 7748 5772
rect 7699 5732 7748 5760
rect 7699 5729 7711 5732
rect 7653 5723 7711 5729
rect 7742 5720 7748 5732
rect 7800 5720 7806 5772
rect 7926 5760 7932 5772
rect 7887 5732 7932 5760
rect 7926 5720 7932 5732
rect 7984 5720 7990 5772
rect 8478 5720 8484 5772
rect 8536 5760 8542 5772
rect 8573 5763 8631 5769
rect 8573 5760 8585 5763
rect 8536 5732 8585 5760
rect 8536 5720 8542 5732
rect 8573 5729 8585 5732
rect 8619 5729 8631 5763
rect 8573 5723 8631 5729
rect 8665 5763 8723 5769
rect 8665 5729 8677 5763
rect 8711 5760 8723 5763
rect 9232 5760 9260 5800
rect 9674 5788 9680 5800
rect 9732 5828 9738 5840
rect 10042 5828 10048 5840
rect 9732 5800 10048 5828
rect 9732 5788 9738 5800
rect 10042 5788 10048 5800
rect 10100 5788 10106 5840
rect 10686 5788 10692 5840
rect 10744 5788 10750 5840
rect 11348 5837 11376 5868
rect 11333 5831 11391 5837
rect 11333 5797 11345 5831
rect 11379 5797 11391 5831
rect 11333 5791 11391 5797
rect 11422 5788 11428 5840
rect 11480 5828 11486 5840
rect 12069 5831 12127 5837
rect 12069 5828 12081 5831
rect 11480 5800 12081 5828
rect 11480 5788 11486 5800
rect 12069 5797 12081 5800
rect 12115 5797 12127 5831
rect 12618 5828 12624 5840
rect 12069 5791 12127 5797
rect 12406 5800 12624 5828
rect 9398 5760 9404 5772
rect 8711 5732 9260 5760
rect 9359 5732 9404 5760
rect 8711 5729 8723 5732
rect 8665 5723 8723 5729
rect 9398 5720 9404 5732
rect 9456 5720 9462 5772
rect 11698 5760 11704 5772
rect 11659 5732 11704 5760
rect 11698 5720 11704 5732
rect 11756 5720 11762 5772
rect 11882 5760 11888 5772
rect 11843 5732 11888 5760
rect 11882 5720 11888 5732
rect 11940 5720 11946 5772
rect 12406 5760 12434 5800
rect 12618 5788 12624 5800
rect 12676 5788 12682 5840
rect 12713 5831 12771 5837
rect 12713 5797 12725 5831
rect 12759 5828 12771 5831
rect 12986 5828 12992 5840
rect 12759 5800 12992 5828
rect 12759 5797 12771 5800
rect 12713 5791 12771 5797
rect 12986 5788 12992 5800
rect 13044 5788 13050 5840
rect 14384 5828 14412 5868
rect 14458 5856 14464 5908
rect 14516 5896 14522 5908
rect 14645 5899 14703 5905
rect 14645 5896 14657 5899
rect 14516 5868 14657 5896
rect 14516 5856 14522 5868
rect 14645 5865 14657 5868
rect 14691 5865 14703 5899
rect 17126 5896 17132 5908
rect 14645 5859 14703 5865
rect 14844 5868 17132 5896
rect 14844 5828 14872 5868
rect 17126 5856 17132 5868
rect 17184 5856 17190 5908
rect 17310 5856 17316 5908
rect 17368 5896 17374 5908
rect 17494 5896 17500 5908
rect 17368 5868 17500 5896
rect 17368 5856 17374 5868
rect 17494 5856 17500 5868
rect 17552 5856 17558 5908
rect 17865 5899 17923 5905
rect 17865 5865 17877 5899
rect 17911 5896 17923 5899
rect 18046 5896 18052 5908
rect 17911 5868 18052 5896
rect 17911 5865 17923 5868
rect 17865 5859 17923 5865
rect 18046 5856 18052 5868
rect 18104 5856 18110 5908
rect 14384 5800 14872 5828
rect 15102 5788 15108 5840
rect 15160 5788 15166 5840
rect 16022 5788 16028 5840
rect 16080 5828 16086 5840
rect 16117 5831 16175 5837
rect 16117 5828 16129 5831
rect 16080 5800 16129 5828
rect 16080 5788 16086 5800
rect 16117 5797 16129 5800
rect 16163 5797 16175 5831
rect 16117 5791 16175 5797
rect 16390 5788 16396 5840
rect 16448 5828 16454 5840
rect 16853 5831 16911 5837
rect 16448 5800 16528 5828
rect 16448 5788 16454 5800
rect 14458 5760 14464 5772
rect 11992 5732 12434 5760
rect 13846 5732 14464 5760
rect 7116 5664 7880 5692
rect 7852 5636 7880 5664
rect 8754 5652 8760 5704
rect 8812 5692 8818 5704
rect 8812 5664 8857 5692
rect 8812 5652 8818 5664
rect 9030 5652 9036 5704
rect 9088 5692 9094 5704
rect 9493 5695 9551 5701
rect 9493 5692 9505 5695
rect 9088 5664 9505 5692
rect 9088 5652 9094 5664
rect 9493 5661 9505 5664
rect 9539 5692 9551 5695
rect 9539 5664 11560 5692
rect 9539 5661 9551 5664
rect 9493 5655 9551 5661
rect 5718 5624 5724 5636
rect 4816 5596 5724 5624
rect 5718 5584 5724 5596
rect 5776 5584 5782 5636
rect 7006 5584 7012 5636
rect 7064 5624 7070 5636
rect 7745 5627 7803 5633
rect 7745 5624 7757 5627
rect 7064 5596 7757 5624
rect 7064 5584 7070 5596
rect 7745 5593 7757 5596
rect 7791 5593 7803 5627
rect 7745 5587 7803 5593
rect 7834 5584 7840 5636
rect 7892 5624 7898 5636
rect 8113 5627 8171 5633
rect 7892 5596 7937 5624
rect 7892 5584 7898 5596
rect 8113 5593 8125 5627
rect 8159 5624 8171 5627
rect 11532 5624 11560 5664
rect 11606 5652 11612 5704
rect 11664 5692 11670 5704
rect 11664 5664 11709 5692
rect 11664 5652 11670 5664
rect 11992 5624 12020 5732
rect 14458 5720 14464 5732
rect 14516 5720 14522 5772
rect 16500 5769 16528 5800
rect 16853 5797 16865 5831
rect 16899 5828 16911 5831
rect 18138 5828 18144 5840
rect 16899 5800 18144 5828
rect 16899 5797 16911 5800
rect 16853 5791 16911 5797
rect 18138 5788 18144 5800
rect 18196 5788 18202 5840
rect 18414 5828 18420 5840
rect 18248 5800 18420 5828
rect 16485 5763 16543 5769
rect 16485 5729 16497 5763
rect 16531 5729 16543 5763
rect 16485 5723 16543 5729
rect 16639 5763 16697 5769
rect 16639 5729 16651 5763
rect 16685 5760 16697 5763
rect 16758 5760 16764 5772
rect 16685 5732 16764 5760
rect 16685 5729 16697 5732
rect 16639 5723 16697 5729
rect 16758 5720 16764 5732
rect 16816 5720 16822 5772
rect 17218 5720 17224 5772
rect 17276 5760 17282 5772
rect 17405 5763 17463 5769
rect 17405 5760 17417 5763
rect 17276 5732 17417 5760
rect 17276 5720 17282 5732
rect 17405 5729 17417 5732
rect 17451 5729 17463 5763
rect 18046 5760 18052 5772
rect 17959 5732 18052 5760
rect 17405 5723 17463 5729
rect 18046 5720 18052 5732
rect 18104 5760 18110 5772
rect 18248 5760 18276 5800
rect 18414 5788 18420 5800
rect 18472 5788 18478 5840
rect 18104 5732 18276 5760
rect 18325 5763 18383 5769
rect 18104 5720 18110 5732
rect 18325 5729 18337 5763
rect 18371 5729 18383 5763
rect 18325 5723 18383 5729
rect 12426 5695 12484 5701
rect 12426 5692 12438 5695
rect 8159 5596 10364 5624
rect 11532 5596 12020 5624
rect 12360 5664 12438 5692
rect 12360 5624 12388 5664
rect 12426 5661 12438 5664
rect 12472 5661 12484 5695
rect 12426 5655 12484 5661
rect 12710 5652 12716 5704
rect 12768 5692 12774 5704
rect 13078 5692 13084 5704
rect 12768 5664 13084 5692
rect 12768 5652 12774 5664
rect 13078 5652 13084 5664
rect 13136 5692 13142 5704
rect 16393 5695 16451 5701
rect 13136 5664 16344 5692
rect 13136 5652 13142 5664
rect 12360 5596 12434 5624
rect 8159 5593 8171 5596
rect 8113 5587 8171 5593
rect 753 5559 811 5565
rect 753 5525 765 5559
rect 799 5556 811 5559
rect 1394 5556 1400 5568
rect 799 5528 1400 5556
rect 799 5525 811 5528
rect 753 5519 811 5525
rect 1394 5516 1400 5528
rect 1452 5516 1458 5568
rect 3513 5559 3571 5565
rect 3513 5525 3525 5559
rect 3559 5556 3571 5559
rect 4430 5556 4436 5568
rect 3559 5528 4436 5556
rect 3559 5525 3571 5528
rect 3513 5519 3571 5525
rect 4430 5516 4436 5528
rect 4488 5516 4494 5568
rect 4893 5559 4951 5565
rect 4893 5525 4905 5559
rect 4939 5556 4951 5559
rect 5258 5556 5264 5568
rect 4939 5528 5264 5556
rect 4939 5525 4951 5528
rect 4893 5519 4951 5525
rect 5258 5516 5264 5528
rect 5316 5516 5322 5568
rect 7285 5559 7343 5565
rect 7285 5525 7297 5559
rect 7331 5556 7343 5559
rect 7650 5556 7656 5568
rect 7331 5528 7656 5556
rect 7331 5525 7343 5528
rect 7285 5519 7343 5525
rect 7650 5516 7656 5528
rect 7708 5516 7714 5568
rect 8202 5556 8208 5568
rect 8163 5528 8208 5556
rect 8202 5516 8208 5528
rect 8260 5516 8266 5568
rect 10336 5556 10364 5596
rect 11698 5556 11704 5568
rect 10336 5528 11704 5556
rect 11698 5516 11704 5528
rect 11756 5516 11762 5568
rect 12158 5516 12164 5568
rect 12216 5556 12222 5568
rect 12253 5559 12311 5565
rect 12253 5556 12265 5559
rect 12216 5528 12265 5556
rect 12216 5516 12222 5528
rect 12253 5525 12265 5528
rect 12299 5525 12311 5559
rect 12406 5556 12434 5596
rect 13446 5556 13452 5568
rect 12406 5528 13452 5556
rect 12253 5519 12311 5525
rect 13446 5516 13452 5528
rect 13504 5516 13510 5568
rect 13814 5516 13820 5568
rect 13872 5556 13878 5568
rect 14185 5559 14243 5565
rect 14185 5556 14197 5559
rect 13872 5528 14197 5556
rect 13872 5516 13878 5528
rect 14185 5525 14197 5528
rect 14231 5525 14243 5559
rect 14185 5519 14243 5525
rect 14369 5559 14427 5565
rect 14369 5525 14381 5559
rect 14415 5556 14427 5559
rect 15102 5556 15108 5568
rect 14415 5528 15108 5556
rect 14415 5525 14427 5528
rect 14369 5519 14427 5525
rect 15102 5516 15108 5528
rect 15160 5516 15166 5568
rect 16316 5556 16344 5664
rect 16393 5661 16405 5695
rect 16439 5692 16451 5695
rect 16850 5692 16856 5704
rect 16439 5664 16856 5692
rect 16439 5661 16451 5664
rect 16393 5655 16451 5661
rect 16850 5652 16856 5664
rect 16908 5652 16914 5704
rect 17494 5692 17500 5704
rect 17455 5664 17500 5692
rect 17494 5652 17500 5664
rect 17552 5652 17558 5704
rect 17589 5695 17647 5701
rect 17589 5661 17601 5695
rect 17635 5661 17647 5695
rect 17589 5655 17647 5661
rect 16666 5584 16672 5636
rect 16724 5624 16730 5636
rect 17218 5624 17224 5636
rect 16724 5596 17224 5624
rect 16724 5584 16730 5596
rect 17218 5584 17224 5596
rect 17276 5584 17282 5636
rect 16850 5556 16856 5568
rect 16316 5528 16856 5556
rect 16850 5516 16856 5528
rect 16908 5516 16914 5568
rect 17034 5556 17040 5568
rect 16995 5528 17040 5556
rect 17034 5516 17040 5528
rect 17092 5516 17098 5568
rect 17604 5556 17632 5655
rect 17770 5652 17776 5704
rect 17828 5692 17834 5704
rect 18233 5695 18291 5701
rect 18233 5692 18245 5695
rect 17828 5664 18245 5692
rect 17828 5652 17834 5664
rect 18233 5661 18245 5664
rect 18279 5661 18291 5695
rect 18233 5655 18291 5661
rect 18340 5636 18368 5723
rect 17678 5584 17684 5636
rect 17736 5624 17742 5636
rect 18141 5627 18199 5633
rect 18141 5624 18153 5627
rect 17736 5596 18153 5624
rect 17736 5584 17742 5596
rect 18141 5593 18153 5596
rect 18187 5593 18199 5627
rect 18141 5587 18199 5593
rect 18322 5584 18328 5636
rect 18380 5584 18386 5636
rect 18230 5556 18236 5568
rect 17604 5528 18236 5556
rect 18230 5516 18236 5528
rect 18288 5516 18294 5568
rect 184 5466 18924 5488
rect 184 5414 3110 5466
rect 3162 5414 3174 5466
rect 3226 5414 3238 5466
rect 3290 5414 3302 5466
rect 3354 5414 3366 5466
rect 3418 5414 6210 5466
rect 6262 5414 6274 5466
rect 6326 5414 6338 5466
rect 6390 5414 6402 5466
rect 6454 5414 6466 5466
rect 6518 5414 9310 5466
rect 9362 5414 9374 5466
rect 9426 5414 9438 5466
rect 9490 5414 9502 5466
rect 9554 5414 9566 5466
rect 9618 5414 12410 5466
rect 12462 5414 12474 5466
rect 12526 5414 12538 5466
rect 12590 5414 12602 5466
rect 12654 5414 12666 5466
rect 12718 5414 15510 5466
rect 15562 5414 15574 5466
rect 15626 5414 15638 5466
rect 15690 5414 15702 5466
rect 15754 5414 15766 5466
rect 15818 5414 18610 5466
rect 18662 5414 18674 5466
rect 18726 5414 18738 5466
rect 18790 5414 18802 5466
rect 18854 5414 18866 5466
rect 18918 5414 18924 5466
rect 184 5392 18924 5414
rect 1489 5355 1547 5361
rect 1489 5321 1501 5355
rect 1535 5352 1547 5355
rect 1946 5352 1952 5364
rect 1535 5324 1952 5352
rect 1535 5321 1547 5324
rect 1489 5315 1547 5321
rect 1946 5312 1952 5324
rect 2004 5312 2010 5364
rect 5626 5312 5632 5364
rect 5684 5352 5690 5364
rect 5813 5355 5871 5361
rect 5813 5352 5825 5355
rect 5684 5324 5825 5352
rect 5684 5312 5690 5324
rect 5813 5321 5825 5324
rect 5859 5321 5871 5355
rect 5813 5315 5871 5321
rect 6457 5355 6515 5361
rect 6457 5321 6469 5355
rect 6503 5352 6515 5355
rect 6546 5352 6552 5364
rect 6503 5324 6552 5352
rect 6503 5321 6515 5324
rect 6457 5315 6515 5321
rect 6546 5312 6552 5324
rect 6604 5312 6610 5364
rect 7190 5312 7196 5364
rect 7248 5352 7254 5364
rect 7377 5355 7435 5361
rect 7377 5352 7389 5355
rect 7248 5324 7389 5352
rect 7248 5312 7254 5324
rect 7377 5321 7389 5324
rect 7423 5321 7435 5355
rect 7377 5315 7435 5321
rect 7834 5312 7840 5364
rect 7892 5352 7898 5364
rect 8478 5352 8484 5364
rect 7892 5324 8484 5352
rect 7892 5312 7898 5324
rect 8478 5312 8484 5324
rect 8536 5312 8542 5364
rect 8846 5352 8852 5364
rect 8807 5324 8852 5352
rect 8846 5312 8852 5324
rect 8904 5312 8910 5364
rect 10226 5352 10232 5364
rect 8956 5324 10232 5352
rect 7742 5244 7748 5296
rect 7800 5284 7806 5296
rect 8956 5284 8984 5324
rect 10226 5312 10232 5324
rect 10284 5312 10290 5364
rect 13170 5312 13176 5364
rect 13228 5352 13234 5364
rect 15841 5355 15899 5361
rect 13228 5324 15516 5352
rect 13228 5312 13234 5324
rect 13081 5287 13139 5293
rect 13081 5284 13093 5287
rect 7800 5256 8984 5284
rect 12406 5256 13093 5284
rect 7800 5244 7806 5256
rect 1486 5176 1492 5228
rect 1544 5216 1550 5228
rect 3237 5219 3295 5225
rect 3237 5216 3249 5219
rect 1544 5188 3249 5216
rect 1544 5176 1550 5188
rect 3237 5185 3249 5188
rect 3283 5185 3295 5219
rect 3878 5216 3884 5228
rect 3839 5188 3884 5216
rect 3237 5179 3295 5185
rect 3878 5176 3884 5188
rect 3936 5176 3942 5228
rect 4154 5176 4160 5228
rect 4212 5216 4218 5228
rect 6730 5216 6736 5228
rect 4212 5188 5028 5216
rect 6691 5188 6736 5216
rect 4212 5176 4218 5188
rect 4246 5148 4252 5160
rect 4207 5120 4252 5148
rect 4246 5108 4252 5120
rect 4304 5108 4310 5160
rect 5000 5148 5028 5188
rect 6730 5176 6736 5188
rect 6788 5176 6794 5228
rect 7006 5176 7012 5228
rect 7064 5216 7070 5228
rect 8021 5219 8079 5225
rect 7064 5188 7512 5216
rect 7064 5176 7070 5188
rect 5813 5151 5871 5157
rect 5813 5148 5825 5151
rect 5000 5120 5825 5148
rect 5813 5117 5825 5120
rect 5859 5117 5871 5151
rect 5994 5148 6000 5160
rect 5955 5120 6000 5148
rect 5813 5111 5871 5117
rect 5994 5108 6000 5120
rect 6052 5108 6058 5160
rect 6086 5108 6092 5160
rect 6144 5148 6150 5160
rect 6825 5151 6883 5157
rect 6825 5148 6837 5151
rect 6144 5120 6837 5148
rect 6144 5108 6150 5120
rect 6825 5117 6837 5120
rect 6871 5117 6883 5151
rect 6825 5111 6883 5117
rect 6917 5151 6975 5157
rect 6917 5117 6929 5151
rect 6963 5148 6975 5151
rect 7282 5148 7288 5160
rect 6963 5120 7288 5148
rect 6963 5117 6975 5120
rect 6917 5111 6975 5117
rect 7282 5108 7288 5120
rect 7340 5108 7346 5160
rect 7484 5148 7512 5188
rect 8021 5185 8033 5219
rect 8067 5216 8079 5219
rect 8110 5216 8116 5228
rect 8067 5188 8116 5216
rect 8067 5185 8079 5188
rect 8021 5179 8079 5185
rect 8110 5176 8116 5188
rect 8168 5216 8174 5228
rect 8757 5219 8815 5225
rect 8757 5216 8769 5219
rect 8168 5188 8769 5216
rect 8168 5176 8174 5188
rect 8757 5185 8769 5188
rect 8803 5185 8815 5219
rect 8757 5179 8815 5185
rect 8846 5176 8852 5228
rect 8904 5216 8910 5228
rect 8941 5219 8999 5225
rect 8941 5216 8953 5219
rect 8904 5188 8953 5216
rect 8904 5176 8910 5188
rect 8941 5185 8953 5188
rect 8987 5185 8999 5219
rect 8941 5179 8999 5185
rect 9214 5176 9220 5228
rect 9272 5216 9278 5228
rect 9401 5219 9459 5225
rect 9401 5216 9413 5219
rect 9272 5188 9413 5216
rect 9272 5176 9278 5188
rect 9401 5185 9413 5188
rect 9447 5185 9459 5219
rect 9401 5179 9459 5185
rect 9582 5176 9588 5228
rect 9640 5216 9646 5228
rect 12406 5216 12434 5256
rect 13081 5253 13093 5256
rect 13127 5253 13139 5287
rect 13081 5247 13139 5253
rect 14734 5244 14740 5296
rect 14792 5284 14798 5296
rect 15381 5287 15439 5293
rect 15381 5284 15393 5287
rect 14792 5256 15393 5284
rect 14792 5244 14798 5256
rect 15381 5253 15393 5256
rect 15427 5253 15439 5287
rect 15381 5247 15439 5253
rect 14366 5216 14372 5228
rect 9640 5188 12434 5216
rect 12820 5188 14372 5216
rect 9640 5176 9646 5188
rect 8297 5151 8355 5157
rect 8297 5148 8309 5151
rect 7484 5120 8309 5148
rect 8297 5117 8309 5120
rect 8343 5117 8355 5151
rect 8297 5111 8355 5117
rect 8665 5151 8723 5157
rect 8665 5117 8677 5151
rect 8711 5117 8723 5151
rect 9030 5148 9036 5160
rect 8991 5120 9036 5148
rect 8665 5111 8723 5117
rect 2958 5080 2964 5092
rect 2530 5052 2774 5080
rect 2919 5052 2964 5080
rect 2746 5012 2774 5052
rect 2958 5040 2964 5052
rect 3016 5040 3022 5092
rect 5350 5080 5356 5092
rect 5263 5052 5356 5080
rect 5350 5040 5356 5052
rect 5408 5080 5414 5092
rect 5408 5052 5488 5080
rect 5408 5040 5414 5052
rect 3602 5012 3608 5024
rect 2746 4984 3608 5012
rect 3602 4972 3608 4984
rect 3660 4972 3666 5024
rect 3697 5015 3755 5021
rect 3697 4981 3709 5015
rect 3743 5012 3755 5015
rect 5166 5012 5172 5024
rect 3743 4984 5172 5012
rect 3743 4981 3755 4984
rect 3697 4975 3755 4981
rect 5166 4972 5172 4984
rect 5224 4972 5230 5024
rect 5460 5012 5488 5052
rect 5534 5040 5540 5092
rect 5592 5080 5598 5092
rect 5721 5083 5779 5089
rect 5721 5080 5733 5083
rect 5592 5052 5733 5080
rect 5592 5040 5598 5052
rect 5721 5049 5733 5052
rect 5767 5080 5779 5083
rect 7006 5080 7012 5092
rect 5767 5052 7012 5080
rect 5767 5049 5779 5052
rect 5721 5043 5779 5049
rect 7006 5040 7012 5052
rect 7064 5040 7070 5092
rect 7098 5040 7104 5092
rect 7156 5080 7162 5092
rect 7745 5083 7803 5089
rect 7745 5080 7757 5083
rect 7156 5052 7757 5080
rect 7156 5040 7162 5052
rect 7745 5049 7757 5052
rect 7791 5049 7803 5083
rect 8202 5080 8208 5092
rect 8163 5052 8208 5080
rect 7745 5043 7803 5049
rect 8202 5040 8208 5052
rect 8260 5040 8266 5092
rect 6822 5012 6828 5024
rect 5460 4984 6828 5012
rect 6822 4972 6828 4984
rect 6880 4972 6886 5024
rect 7282 5012 7288 5024
rect 7243 4984 7288 5012
rect 7282 4972 7288 4984
rect 7340 4972 7346 5024
rect 7374 4972 7380 5024
rect 7432 5012 7438 5024
rect 7837 5015 7895 5021
rect 7837 5012 7849 5015
rect 7432 4984 7849 5012
rect 7432 4972 7438 4984
rect 7837 4981 7849 4984
rect 7883 4981 7895 5015
rect 7837 4975 7895 4981
rect 7926 4972 7932 5024
rect 7984 5012 7990 5024
rect 8680 5012 8708 5111
rect 9030 5108 9036 5120
rect 9088 5108 9094 5160
rect 12820 5157 12848 5188
rect 14366 5176 14372 5188
rect 14424 5176 14430 5228
rect 14458 5176 14464 5228
rect 14516 5216 14522 5228
rect 15488 5216 15516 5324
rect 15841 5321 15853 5355
rect 15887 5352 15899 5355
rect 16114 5352 16120 5364
rect 15887 5324 16120 5352
rect 15887 5321 15899 5324
rect 15841 5315 15899 5321
rect 16114 5312 16120 5324
rect 16172 5312 16178 5364
rect 17405 5355 17463 5361
rect 16316 5324 17356 5352
rect 16316 5225 16344 5324
rect 16482 5244 16488 5296
rect 16540 5284 16546 5296
rect 17126 5284 17132 5296
rect 16540 5256 17132 5284
rect 16540 5244 16546 5256
rect 17126 5244 17132 5256
rect 17184 5244 17190 5296
rect 17328 5284 17356 5324
rect 17405 5321 17417 5355
rect 17451 5352 17463 5355
rect 17494 5352 17500 5364
rect 17451 5324 17500 5352
rect 17451 5321 17463 5324
rect 17405 5315 17463 5321
rect 17494 5312 17500 5324
rect 17552 5312 17558 5364
rect 17862 5312 17868 5364
rect 17920 5352 17926 5364
rect 17957 5355 18015 5361
rect 17957 5352 17969 5355
rect 17920 5324 17969 5352
rect 17920 5312 17926 5324
rect 17957 5321 17969 5324
rect 18003 5321 18015 5355
rect 17957 5315 18015 5321
rect 17328 5256 17448 5284
rect 16301 5219 16359 5225
rect 14516 5188 14964 5216
rect 15488 5188 15700 5216
rect 14516 5176 14522 5188
rect 12805 5151 12863 5157
rect 12805 5117 12817 5151
rect 12851 5117 12863 5151
rect 12805 5111 12863 5117
rect 12894 5108 12900 5160
rect 12952 5148 12958 5160
rect 12952 5120 12997 5148
rect 12952 5108 12958 5120
rect 13078 5108 13084 5160
rect 13136 5148 13142 5160
rect 13446 5148 13452 5160
rect 13136 5120 13181 5148
rect 13407 5120 13452 5148
rect 13136 5108 13142 5120
rect 13446 5108 13452 5120
rect 13504 5108 13510 5160
rect 10686 5080 10692 5092
rect 10442 5052 10692 5080
rect 10686 5040 10692 5052
rect 10744 5080 10750 5092
rect 12250 5080 12256 5092
rect 10744 5052 12256 5080
rect 10744 5040 10750 5052
rect 12250 5040 12256 5052
rect 12308 5040 12314 5092
rect 12434 5040 12440 5092
rect 12492 5080 12498 5092
rect 13464 5080 13492 5108
rect 12492 5052 13492 5080
rect 13725 5083 13783 5089
rect 12492 5040 12498 5052
rect 13725 5049 13737 5083
rect 13771 5080 13783 5083
rect 13814 5080 13820 5092
rect 13771 5052 13820 5080
rect 13771 5049 13783 5052
rect 13725 5043 13783 5049
rect 13814 5040 13820 5052
rect 13872 5040 13878 5092
rect 14936 5080 14964 5188
rect 15194 5108 15200 5160
rect 15252 5148 15258 5160
rect 15289 5151 15347 5157
rect 15289 5148 15301 5151
rect 15252 5120 15301 5148
rect 15252 5108 15258 5120
rect 15289 5117 15301 5120
rect 15335 5117 15347 5151
rect 15562 5148 15568 5160
rect 15523 5120 15568 5148
rect 15289 5111 15347 5117
rect 15562 5108 15568 5120
rect 15620 5108 15626 5160
rect 15672 5148 15700 5188
rect 16301 5185 16313 5219
rect 16347 5185 16359 5219
rect 16301 5179 16359 5185
rect 16393 5219 16451 5225
rect 16393 5185 16405 5219
rect 16439 5216 16451 5219
rect 16666 5216 16672 5228
rect 16439 5188 16672 5216
rect 16439 5185 16451 5188
rect 16393 5179 16451 5185
rect 16666 5176 16672 5188
rect 16724 5216 16730 5228
rect 16945 5219 17003 5225
rect 16945 5216 16957 5219
rect 16724 5188 16957 5216
rect 16724 5176 16730 5188
rect 16945 5185 16957 5188
rect 16991 5185 17003 5219
rect 16945 5179 17003 5185
rect 16761 5151 16819 5157
rect 16761 5148 16773 5151
rect 15672 5120 16773 5148
rect 16761 5117 16773 5120
rect 16807 5117 16819 5151
rect 16761 5111 16819 5117
rect 16850 5108 16856 5160
rect 16908 5148 16914 5160
rect 17129 5151 17187 5157
rect 16908 5120 16953 5148
rect 16908 5108 16914 5120
rect 17129 5117 17141 5151
rect 17175 5117 17187 5151
rect 17129 5111 17187 5117
rect 15010 5080 15016 5092
rect 14936 5066 15016 5080
rect 14950 5052 15016 5066
rect 15010 5040 15016 5052
rect 15068 5040 15074 5092
rect 15473 5083 15531 5089
rect 15473 5049 15485 5083
rect 15519 5080 15531 5083
rect 15838 5080 15844 5092
rect 15519 5052 15844 5080
rect 15519 5049 15531 5052
rect 15473 5043 15531 5049
rect 15838 5040 15844 5052
rect 15896 5040 15902 5092
rect 16209 5083 16267 5089
rect 16209 5049 16221 5083
rect 16255 5080 16267 5083
rect 17034 5080 17040 5092
rect 16255 5052 17040 5080
rect 16255 5049 16267 5052
rect 16209 5043 16267 5049
rect 17034 5040 17040 5052
rect 17092 5040 17098 5092
rect 17144 5080 17172 5111
rect 17218 5108 17224 5160
rect 17276 5148 17282 5160
rect 17420 5148 17448 5256
rect 17586 5176 17592 5228
rect 17644 5216 17650 5228
rect 17770 5216 17776 5228
rect 17644 5188 17776 5216
rect 17644 5176 17650 5188
rect 17770 5176 17776 5188
rect 17828 5176 17834 5228
rect 17678 5148 17684 5160
rect 17276 5120 17321 5148
rect 17420 5120 17684 5148
rect 17276 5108 17282 5120
rect 17678 5108 17684 5120
rect 17736 5108 17742 5160
rect 18046 5108 18052 5160
rect 18104 5148 18110 5160
rect 18233 5151 18291 5157
rect 18233 5148 18245 5151
rect 18104 5120 18245 5148
rect 18104 5108 18110 5120
rect 18233 5117 18245 5120
rect 18279 5117 18291 5151
rect 18233 5111 18291 5117
rect 17310 5080 17316 5092
rect 17144 5052 17316 5080
rect 17310 5040 17316 5052
rect 17368 5080 17374 5092
rect 17586 5080 17592 5092
rect 17368 5052 17592 5080
rect 17368 5040 17374 5052
rect 17586 5040 17592 5052
rect 17644 5040 17650 5092
rect 18138 5040 18144 5092
rect 18196 5080 18202 5092
rect 18325 5083 18383 5089
rect 18325 5080 18337 5083
rect 18196 5052 18337 5080
rect 18196 5040 18202 5052
rect 18325 5049 18337 5052
rect 18371 5049 18383 5083
rect 18325 5043 18383 5049
rect 18509 5083 18567 5089
rect 18509 5049 18521 5083
rect 18555 5080 18567 5083
rect 19150 5080 19156 5092
rect 18555 5052 19156 5080
rect 18555 5049 18567 5052
rect 18509 5043 18567 5049
rect 19150 5040 19156 5052
rect 19208 5040 19214 5092
rect 9858 5012 9864 5024
rect 7984 4984 9864 5012
rect 7984 4972 7990 4984
rect 9858 4972 9864 4984
rect 9916 4972 9922 5024
rect 10778 4972 10784 5024
rect 10836 5021 10842 5024
rect 10836 5015 10885 5021
rect 10836 4981 10839 5015
rect 10873 4981 10885 5015
rect 10836 4975 10885 4981
rect 10836 4972 10842 4975
rect 11422 4972 11428 5024
rect 11480 5012 11486 5024
rect 11517 5015 11575 5021
rect 11517 5012 11529 5015
rect 11480 4984 11529 5012
rect 11480 4972 11486 4984
rect 11517 4981 11529 4984
rect 11563 4981 11575 5015
rect 11517 4975 11575 4981
rect 12158 4972 12164 5024
rect 12216 5012 12222 5024
rect 13265 5015 13323 5021
rect 13265 5012 13277 5015
rect 12216 4984 13277 5012
rect 12216 4972 12222 4984
rect 13265 4981 13277 4984
rect 13311 5012 13323 5015
rect 13354 5012 13360 5024
rect 13311 4984 13360 5012
rect 13311 4981 13323 4984
rect 13265 4975 13323 4981
rect 13354 4972 13360 4984
rect 13412 4972 13418 5024
rect 15194 5012 15200 5024
rect 15155 4984 15200 5012
rect 15194 4972 15200 4984
rect 15252 4972 15258 5024
rect 16761 5015 16819 5021
rect 16761 4981 16773 5015
rect 16807 5012 16819 5015
rect 17402 5012 17408 5024
rect 16807 4984 17408 5012
rect 16807 4981 16819 4984
rect 16761 4975 16819 4981
rect 17402 4972 17408 4984
rect 17460 4972 17466 5024
rect 18414 5012 18420 5024
rect 18375 4984 18420 5012
rect 18414 4972 18420 4984
rect 18472 4972 18478 5024
rect 184 4922 18860 4944
rect 184 4870 4660 4922
rect 4712 4870 4724 4922
rect 4776 4870 4788 4922
rect 4840 4870 4852 4922
rect 4904 4870 4916 4922
rect 4968 4870 7760 4922
rect 7812 4870 7824 4922
rect 7876 4870 7888 4922
rect 7940 4870 7952 4922
rect 8004 4870 8016 4922
rect 8068 4870 10860 4922
rect 10912 4870 10924 4922
rect 10976 4870 10988 4922
rect 11040 4870 11052 4922
rect 11104 4870 11116 4922
rect 11168 4870 13960 4922
rect 14012 4870 14024 4922
rect 14076 4870 14088 4922
rect 14140 4870 14152 4922
rect 14204 4870 14216 4922
rect 14268 4870 17060 4922
rect 17112 4870 17124 4922
rect 17176 4870 17188 4922
rect 17240 4870 17252 4922
rect 17304 4870 17316 4922
rect 17368 4870 18860 4922
rect 184 4848 18860 4870
rect 2498 4768 2504 4820
rect 2556 4808 2562 4820
rect 2958 4808 2964 4820
rect 2556 4780 2964 4808
rect 2556 4768 2562 4780
rect 2958 4768 2964 4780
rect 3016 4768 3022 4820
rect 4246 4768 4252 4820
rect 4304 4808 4310 4820
rect 6365 4811 6423 4817
rect 6365 4808 6377 4811
rect 4304 4780 6377 4808
rect 4304 4768 4310 4780
rect 6365 4777 6377 4780
rect 6411 4777 6423 4811
rect 6365 4771 6423 4777
rect 6546 4768 6552 4820
rect 6604 4808 6610 4820
rect 6825 4811 6883 4817
rect 6604 4780 6776 4808
rect 6604 4768 6610 4780
rect 3510 4740 3516 4752
rect 3160 4712 3516 4740
rect 2498 4632 2504 4684
rect 2556 4672 2562 4684
rect 3160 4681 3188 4712
rect 3510 4700 3516 4712
rect 3568 4700 3574 4752
rect 4706 4740 4712 4752
rect 4619 4712 4712 4740
rect 4706 4700 4712 4712
rect 4764 4740 4770 4752
rect 5350 4740 5356 4752
rect 4764 4712 5356 4740
rect 4764 4700 4770 4712
rect 5350 4700 5356 4712
rect 5408 4700 5414 4752
rect 5629 4743 5687 4749
rect 5629 4709 5641 4743
rect 5675 4740 5687 4743
rect 6638 4740 6644 4752
rect 5675 4712 6644 4740
rect 5675 4709 5687 4712
rect 5629 4703 5687 4709
rect 6638 4700 6644 4712
rect 6696 4700 6702 4752
rect 6748 4740 6776 4780
rect 6825 4777 6837 4811
rect 6871 4808 6883 4811
rect 7006 4808 7012 4820
rect 6871 4780 7012 4808
rect 6871 4777 6883 4780
rect 6825 4771 6883 4777
rect 7006 4768 7012 4780
rect 7064 4808 7070 4820
rect 7742 4808 7748 4820
rect 7064 4780 7748 4808
rect 7064 4768 7070 4780
rect 7742 4768 7748 4780
rect 7800 4808 7806 4820
rect 8205 4811 8263 4817
rect 7800 4780 8064 4808
rect 7800 4768 7806 4780
rect 7469 4743 7527 4749
rect 7469 4740 7481 4743
rect 6748 4712 7481 4740
rect 7469 4709 7481 4712
rect 7515 4709 7527 4743
rect 7469 4703 7527 4709
rect 7650 4700 7656 4752
rect 7708 4740 7714 4752
rect 7926 4740 7932 4752
rect 7708 4712 7932 4740
rect 7708 4700 7714 4712
rect 7926 4700 7932 4712
rect 7984 4700 7990 4752
rect 8036 4749 8064 4780
rect 8205 4777 8217 4811
rect 8251 4808 8263 4811
rect 8662 4808 8668 4820
rect 8251 4780 8668 4808
rect 8251 4777 8263 4780
rect 8205 4771 8263 4777
rect 8662 4768 8668 4780
rect 8720 4768 8726 4820
rect 9030 4768 9036 4820
rect 9088 4808 9094 4820
rect 9401 4811 9459 4817
rect 9401 4808 9413 4811
rect 9088 4780 9413 4808
rect 9088 4768 9094 4780
rect 9401 4777 9413 4780
rect 9447 4808 9459 4811
rect 9950 4808 9956 4820
rect 9447 4780 9956 4808
rect 9447 4777 9459 4780
rect 9401 4771 9459 4777
rect 9950 4768 9956 4780
rect 10008 4768 10014 4820
rect 11422 4768 11428 4820
rect 11480 4808 11486 4820
rect 12434 4808 12440 4820
rect 11480 4780 12440 4808
rect 11480 4768 11486 4780
rect 12434 4768 12440 4780
rect 12492 4768 12498 4820
rect 12986 4768 12992 4820
rect 13044 4808 13050 4820
rect 14642 4808 14648 4820
rect 13044 4780 14136 4808
rect 14603 4780 14648 4808
rect 13044 4768 13050 4780
rect 8021 4743 8079 4749
rect 8021 4709 8033 4743
rect 8067 4709 8079 4743
rect 8021 4703 8079 4709
rect 3145 4675 3203 4681
rect 3145 4672 3157 4675
rect 2556 4644 3157 4672
rect 2556 4632 2562 4644
rect 3145 4641 3157 4644
rect 3191 4641 3203 4675
rect 3145 4635 3203 4641
rect 5169 4675 5227 4681
rect 5169 4641 5181 4675
rect 5215 4641 5227 4675
rect 5169 4635 5227 4641
rect 3421 4607 3479 4613
rect 3421 4573 3433 4607
rect 3467 4604 3479 4607
rect 4982 4604 4988 4616
rect 3467 4576 4988 4604
rect 3467 4573 3479 4576
rect 3421 4567 3479 4573
rect 4982 4564 4988 4576
rect 5040 4564 5046 4616
rect 5184 4604 5212 4635
rect 5258 4632 5264 4684
rect 5316 4672 5322 4684
rect 5445 4675 5503 4681
rect 5445 4672 5457 4675
rect 5316 4644 5457 4672
rect 5316 4632 5322 4644
rect 5445 4641 5457 4644
rect 5491 4672 5503 4675
rect 5902 4672 5908 4684
rect 5491 4644 5908 4672
rect 5491 4641 5503 4644
rect 5445 4635 5503 4641
rect 5902 4632 5908 4644
rect 5960 4632 5966 4684
rect 6086 4672 6092 4684
rect 6047 4644 6092 4672
rect 6086 4632 6092 4644
rect 6144 4632 6150 4684
rect 6546 4632 6552 4684
rect 6604 4672 6610 4684
rect 6733 4675 6791 4681
rect 6733 4672 6745 4675
rect 6604 4644 6745 4672
rect 6604 4632 6610 4644
rect 6733 4641 6745 4644
rect 6779 4641 6791 4675
rect 7190 4672 7196 4684
rect 6733 4635 6791 4641
rect 7024 4644 7196 4672
rect 5184 4576 5948 4604
rect 5258 4536 5264 4548
rect 4816 4508 5264 4536
rect 2958 4428 2964 4480
rect 3016 4468 3022 4480
rect 4816 4468 4844 4508
rect 5258 4496 5264 4508
rect 5316 4496 5322 4548
rect 5353 4539 5411 4545
rect 5353 4505 5365 4539
rect 5399 4536 5411 4539
rect 5442 4536 5448 4548
rect 5399 4508 5448 4536
rect 5399 4505 5411 4508
rect 5353 4499 5411 4505
rect 5442 4496 5448 4508
rect 5500 4496 5506 4548
rect 5718 4536 5724 4548
rect 5679 4508 5724 4536
rect 5718 4496 5724 4508
rect 5776 4496 5782 4548
rect 5920 4536 5948 4576
rect 5994 4564 6000 4616
rect 6052 4604 6058 4616
rect 7024 4613 7052 4644
rect 7190 4632 7196 4644
rect 7248 4672 7254 4684
rect 7745 4675 7803 4681
rect 7745 4672 7757 4675
rect 7248 4644 7757 4672
rect 7248 4632 7254 4644
rect 7745 4641 7757 4644
rect 7791 4641 7803 4675
rect 7745 4635 7803 4641
rect 7837 4675 7895 4681
rect 7837 4641 7849 4675
rect 7883 4641 7895 4675
rect 8036 4672 8064 4703
rect 8478 4700 8484 4752
rect 8536 4740 8542 4752
rect 12250 4740 12256 4752
rect 8536 4712 9996 4740
rect 11822 4712 12256 4740
rect 8536 4700 8542 4712
rect 8036 4644 8616 4672
rect 7837 4635 7895 4641
rect 7009 4607 7067 4613
rect 6052 4576 6097 4604
rect 6052 4564 6058 4576
rect 7009 4573 7021 4607
rect 7055 4573 7067 4607
rect 7009 4567 7067 4573
rect 7650 4536 7656 4548
rect 5920 4508 7656 4536
rect 7650 4496 7656 4508
rect 7708 4496 7714 4548
rect 7852 4536 7880 4635
rect 8297 4607 8355 4613
rect 8297 4573 8309 4607
rect 8343 4604 8355 4607
rect 8478 4604 8484 4616
rect 8343 4576 8484 4604
rect 8343 4573 8355 4576
rect 8297 4567 8355 4573
rect 8478 4564 8484 4576
rect 8536 4564 8542 4616
rect 8588 4604 8616 4644
rect 8846 4632 8852 4684
rect 8904 4672 8910 4684
rect 9214 4672 9220 4684
rect 8904 4644 9220 4672
rect 8904 4632 8910 4644
rect 9214 4632 9220 4644
rect 9272 4672 9278 4684
rect 9309 4675 9367 4681
rect 9309 4672 9321 4675
rect 9272 4644 9321 4672
rect 9272 4632 9278 4644
rect 9309 4641 9321 4644
rect 9355 4641 9367 4675
rect 9582 4672 9588 4684
rect 9309 4635 9367 4641
rect 9508 4644 9588 4672
rect 9508 4613 9536 4644
rect 9582 4632 9588 4644
rect 9640 4632 9646 4684
rect 9968 4681 9996 4712
rect 12250 4700 12256 4712
rect 12308 4700 12314 4752
rect 12452 4740 12480 4768
rect 12452 4712 12756 4740
rect 9953 4675 10011 4681
rect 9953 4641 9965 4675
rect 9999 4641 10011 4675
rect 10226 4672 10232 4684
rect 10187 4644 10232 4672
rect 9953 4635 10011 4641
rect 10226 4632 10232 4644
rect 10284 4632 10290 4684
rect 12437 4675 12495 4681
rect 12437 4672 12449 4675
rect 11808 4644 12449 4672
rect 9493 4607 9551 4613
rect 8588 4576 9076 4604
rect 8570 4536 8576 4548
rect 7852 4508 8576 4536
rect 8570 4496 8576 4508
rect 8628 4496 8634 4548
rect 8665 4539 8723 4545
rect 8665 4505 8677 4539
rect 8711 4536 8723 4539
rect 8941 4539 8999 4545
rect 8941 4536 8953 4539
rect 8711 4508 8953 4536
rect 8711 4505 8723 4508
rect 8665 4499 8723 4505
rect 8941 4505 8953 4508
rect 8987 4505 8999 4539
rect 9048 4536 9076 4576
rect 9493 4573 9505 4607
rect 9539 4573 9551 4607
rect 9858 4604 9864 4616
rect 9819 4576 9864 4604
rect 9493 4567 9551 4573
rect 9858 4564 9864 4576
rect 9916 4564 9922 4616
rect 10318 4604 10324 4616
rect 10279 4576 10324 4604
rect 10318 4564 10324 4576
rect 10376 4564 10382 4616
rect 10594 4604 10600 4616
rect 10555 4576 10600 4604
rect 10594 4564 10600 4576
rect 10652 4564 10658 4616
rect 11054 4564 11060 4616
rect 11112 4604 11118 4616
rect 11808 4604 11836 4644
rect 12437 4641 12449 4644
rect 12483 4641 12495 4675
rect 12618 4672 12624 4684
rect 12579 4644 12624 4672
rect 12437 4635 12495 4641
rect 12618 4632 12624 4644
rect 12676 4632 12682 4684
rect 12728 4681 12756 4712
rect 12713 4675 12771 4681
rect 12713 4641 12725 4675
rect 12759 4641 12771 4675
rect 14108 4672 14136 4780
rect 14642 4768 14648 4780
rect 14700 4768 14706 4820
rect 16485 4811 16543 4817
rect 16485 4808 16497 4811
rect 14752 4780 16497 4808
rect 14550 4700 14556 4752
rect 14608 4740 14614 4752
rect 14752 4740 14780 4780
rect 16485 4777 16497 4780
rect 16531 4777 16543 4811
rect 16485 4771 16543 4777
rect 16850 4768 16856 4820
rect 16908 4808 16914 4820
rect 17586 4808 17592 4820
rect 16908 4780 17592 4808
rect 16908 4768 16914 4780
rect 17586 4768 17592 4780
rect 17644 4768 17650 4820
rect 17954 4768 17960 4820
rect 18012 4808 18018 4820
rect 18417 4811 18475 4817
rect 18417 4808 18429 4811
rect 18012 4780 18429 4808
rect 18012 4768 18018 4780
rect 18417 4777 18429 4780
rect 18463 4777 18475 4811
rect 18417 4771 18475 4777
rect 14608 4712 14780 4740
rect 14608 4700 14614 4712
rect 15746 4700 15752 4752
rect 15804 4749 15810 4752
rect 15804 4740 15816 4749
rect 16114 4740 16120 4752
rect 15804 4712 15849 4740
rect 16075 4712 16120 4740
rect 15804 4703 15816 4712
rect 15804 4700 15810 4703
rect 16114 4700 16120 4712
rect 16172 4700 16178 4752
rect 14458 4672 14464 4684
rect 14108 4658 14464 4672
rect 14122 4644 14464 4658
rect 12713 4635 12771 4641
rect 14458 4632 14464 4644
rect 14516 4632 14522 4684
rect 16393 4675 16451 4681
rect 16393 4672 16405 4675
rect 14568 4644 16405 4672
rect 11112 4576 11836 4604
rect 12069 4607 12127 4613
rect 11112 4564 11118 4576
rect 12069 4573 12081 4607
rect 12115 4604 12127 4607
rect 12989 4607 13047 4613
rect 12989 4604 13001 4607
rect 12115 4576 13001 4604
rect 12115 4573 12127 4576
rect 12069 4567 12127 4573
rect 12989 4573 13001 4576
rect 13035 4573 13047 4607
rect 12989 4567 13047 4573
rect 13722 4564 13728 4616
rect 13780 4604 13786 4616
rect 14568 4604 14596 4644
rect 16393 4641 16405 4644
rect 16439 4641 16451 4675
rect 16393 4635 16451 4641
rect 16574 4632 16580 4684
rect 16632 4672 16638 4684
rect 17218 4672 17224 4684
rect 16632 4644 17224 4672
rect 16632 4632 16638 4644
rect 17218 4632 17224 4644
rect 17276 4632 17282 4684
rect 17865 4675 17923 4681
rect 17865 4672 17877 4675
rect 17328 4644 17877 4672
rect 13780 4576 14596 4604
rect 16025 4607 16083 4613
rect 13780 4564 13786 4576
rect 16025 4573 16037 4607
rect 16071 4604 16083 4607
rect 16206 4604 16212 4616
rect 16071 4576 16212 4604
rect 16071 4573 16083 4576
rect 16025 4567 16083 4573
rect 16206 4564 16212 4576
rect 16264 4564 16270 4616
rect 16666 4564 16672 4616
rect 16724 4604 16730 4616
rect 17328 4604 17356 4644
rect 17865 4641 17877 4644
rect 17911 4641 17923 4675
rect 18138 4672 18144 4684
rect 18099 4644 18144 4672
rect 17865 4635 17923 4641
rect 18138 4632 18144 4644
rect 18196 4632 18202 4684
rect 18322 4672 18328 4684
rect 18283 4644 18328 4672
rect 18322 4632 18328 4644
rect 18380 4632 18386 4684
rect 19058 4604 19064 4616
rect 16724 4576 17356 4604
rect 17420 4576 19064 4604
rect 16724 4564 16730 4576
rect 10045 4539 10103 4545
rect 10045 4536 10057 4539
rect 9048 4508 10057 4536
rect 8941 4499 8999 4505
rect 10045 4505 10057 4508
rect 10091 4505 10103 4539
rect 17420 4536 17448 4576
rect 19058 4564 19064 4576
rect 19116 4564 19122 4616
rect 10045 4499 10103 4505
rect 16040 4508 17448 4536
rect 3016 4440 4844 4468
rect 4893 4471 4951 4477
rect 3016 4428 3022 4440
rect 4893 4437 4905 4471
rect 4939 4468 4951 4471
rect 5810 4468 5816 4480
rect 4939 4440 5816 4468
rect 4939 4437 4951 4440
rect 4893 4431 4951 4437
rect 5810 4428 5816 4440
rect 5868 4428 5874 4480
rect 6086 4428 6092 4480
rect 6144 4468 6150 4480
rect 7193 4471 7251 4477
rect 7193 4468 7205 4471
rect 6144 4440 7205 4468
rect 6144 4428 6150 4440
rect 7193 4437 7205 4440
rect 7239 4437 7251 4471
rect 7193 4431 7251 4437
rect 8757 4471 8815 4477
rect 8757 4437 8769 4471
rect 8803 4468 8815 4471
rect 10134 4468 10140 4480
rect 8803 4440 10140 4468
rect 8803 4437 8815 4440
rect 8757 4431 8815 4437
rect 10134 4428 10140 4440
rect 10192 4428 10198 4480
rect 10229 4471 10287 4477
rect 10229 4437 10241 4471
rect 10275 4468 10287 4471
rect 11882 4468 11888 4480
rect 10275 4440 11888 4468
rect 10275 4437 10287 4440
rect 10229 4431 10287 4437
rect 11882 4428 11888 4440
rect 11940 4428 11946 4480
rect 11974 4428 11980 4480
rect 12032 4468 12038 4480
rect 12253 4471 12311 4477
rect 12253 4468 12265 4471
rect 12032 4440 12265 4468
rect 12032 4428 12038 4440
rect 12253 4437 12265 4440
rect 12299 4437 12311 4471
rect 12253 4431 12311 4437
rect 13078 4428 13084 4480
rect 13136 4468 13142 4480
rect 13722 4468 13728 4480
rect 13136 4440 13728 4468
rect 13136 4428 13142 4440
rect 13722 4428 13728 4440
rect 13780 4428 13786 4480
rect 14458 4468 14464 4480
rect 14419 4440 14464 4468
rect 14458 4428 14464 4440
rect 14516 4428 14522 4480
rect 14642 4428 14648 4480
rect 14700 4468 14706 4480
rect 14918 4468 14924 4480
rect 14700 4440 14924 4468
rect 14700 4428 14706 4440
rect 14918 4428 14924 4440
rect 14976 4428 14982 4480
rect 15838 4428 15844 4480
rect 15896 4468 15902 4480
rect 16040 4468 16068 4508
rect 17586 4496 17592 4548
rect 17644 4536 17650 4548
rect 17957 4539 18015 4545
rect 17957 4536 17969 4539
rect 17644 4508 17969 4536
rect 17644 4496 17650 4508
rect 17957 4505 17969 4508
rect 18003 4505 18015 4539
rect 17957 4499 18015 4505
rect 18049 4539 18107 4545
rect 18049 4505 18061 4539
rect 18095 4536 18107 4539
rect 18230 4536 18236 4548
rect 18095 4508 18236 4536
rect 18095 4505 18107 4508
rect 18049 4499 18107 4505
rect 18230 4496 18236 4508
rect 18288 4496 18294 4548
rect 17310 4468 17316 4480
rect 15896 4440 16068 4468
rect 17271 4440 17316 4468
rect 15896 4428 15902 4440
rect 17310 4428 17316 4440
rect 17368 4428 17374 4480
rect 17402 4428 17408 4480
rect 17460 4468 17466 4480
rect 17681 4471 17739 4477
rect 17681 4468 17693 4471
rect 17460 4440 17693 4468
rect 17460 4428 17466 4440
rect 17681 4437 17693 4440
rect 17727 4437 17739 4471
rect 17681 4431 17739 4437
rect 184 4378 18924 4400
rect 184 4326 3110 4378
rect 3162 4326 3174 4378
rect 3226 4326 3238 4378
rect 3290 4326 3302 4378
rect 3354 4326 3366 4378
rect 3418 4326 6210 4378
rect 6262 4326 6274 4378
rect 6326 4326 6338 4378
rect 6390 4326 6402 4378
rect 6454 4326 6466 4378
rect 6518 4326 9310 4378
rect 9362 4326 9374 4378
rect 9426 4326 9438 4378
rect 9490 4326 9502 4378
rect 9554 4326 9566 4378
rect 9618 4326 12410 4378
rect 12462 4326 12474 4378
rect 12526 4326 12538 4378
rect 12590 4326 12602 4378
rect 12654 4326 12666 4378
rect 12718 4326 15510 4378
rect 15562 4326 15574 4378
rect 15626 4326 15638 4378
rect 15690 4326 15702 4378
rect 15754 4326 15766 4378
rect 15818 4326 18610 4378
rect 18662 4326 18674 4378
rect 18726 4326 18738 4378
rect 18790 4326 18802 4378
rect 18854 4326 18866 4378
rect 18918 4326 18924 4378
rect 184 4304 18924 4326
rect 1118 4224 1124 4276
rect 1176 4264 1182 4276
rect 4065 4267 4123 4273
rect 4065 4264 4077 4267
rect 1176 4236 4077 4264
rect 1176 4224 1182 4236
rect 4065 4233 4077 4236
rect 4111 4264 4123 4267
rect 5994 4264 6000 4276
rect 4111 4236 6000 4264
rect 4111 4233 4123 4236
rect 4065 4227 4123 4233
rect 5994 4224 6000 4236
rect 6052 4224 6058 4276
rect 6730 4224 6736 4276
rect 6788 4264 6794 4276
rect 6788 4236 7512 4264
rect 6788 4224 6794 4236
rect 4706 4196 4712 4208
rect 3620 4168 4712 4196
rect 3620 4072 3648 4168
rect 4706 4156 4712 4168
rect 4764 4156 4770 4208
rect 7101 4199 7159 4205
rect 7101 4196 7113 4199
rect 6380 4168 7113 4196
rect 3697 4131 3755 4137
rect 3697 4097 3709 4131
rect 3743 4097 3755 4131
rect 3697 4091 3755 4097
rect 4249 4131 4307 4137
rect 4249 4097 4261 4131
rect 4295 4128 4307 4131
rect 4338 4128 4344 4140
rect 4295 4100 4344 4128
rect 4295 4097 4307 4100
rect 4249 4091 4307 4097
rect 1949 4063 2007 4069
rect 1949 4029 1961 4063
rect 1995 4029 2007 4063
rect 3602 4060 3608 4072
rect 3358 4032 3608 4060
rect 1949 4023 2007 4029
rect 1964 3924 1992 4023
rect 3602 4020 3608 4032
rect 3660 4020 3666 4072
rect 3712 4060 3740 4091
rect 4338 4088 4344 4100
rect 4396 4088 4402 4140
rect 4982 4128 4988 4140
rect 4895 4100 4988 4128
rect 4982 4088 4988 4100
rect 5040 4128 5046 4140
rect 5813 4131 5871 4137
rect 5813 4128 5825 4131
rect 5040 4100 5825 4128
rect 5040 4088 5046 4100
rect 5813 4097 5825 4100
rect 5859 4097 5871 4131
rect 5813 4091 5871 4097
rect 4154 4060 4160 4072
rect 3712 4032 4160 4060
rect 4154 4020 4160 4032
rect 4212 4060 4218 4072
rect 5166 4060 5172 4072
rect 4212 4032 5172 4060
rect 4212 4020 4218 4032
rect 5166 4020 5172 4032
rect 5224 4020 5230 4072
rect 2222 3992 2228 4004
rect 2183 3964 2228 3992
rect 2222 3952 2228 3964
rect 2280 3952 2286 4004
rect 5828 3992 5856 4091
rect 5902 4088 5908 4140
rect 5960 4128 5966 4140
rect 6089 4131 6147 4137
rect 6089 4128 6101 4131
rect 5960 4100 6101 4128
rect 5960 4088 5966 4100
rect 6089 4097 6101 4100
rect 6135 4128 6147 4131
rect 6178 4128 6184 4140
rect 6135 4100 6184 4128
rect 6135 4097 6147 4100
rect 6089 4091 6147 4097
rect 6178 4088 6184 4100
rect 6236 4088 6242 4140
rect 6086 3992 6092 4004
rect 3620 3964 5212 3992
rect 5828 3964 6092 3992
rect 2498 3924 2504 3936
rect 1964 3896 2504 3924
rect 2498 3884 2504 3896
rect 2556 3884 2562 3936
rect 2590 3884 2596 3936
rect 2648 3924 2654 3936
rect 3620 3924 3648 3964
rect 4338 3924 4344 3936
rect 2648 3896 3648 3924
rect 4299 3896 4344 3924
rect 2648 3884 2654 3896
rect 4338 3884 4344 3896
rect 4396 3884 4402 3936
rect 4522 3884 4528 3936
rect 4580 3924 4586 3936
rect 4709 3927 4767 3933
rect 4709 3924 4721 3927
rect 4580 3896 4721 3924
rect 4580 3884 4586 3896
rect 4709 3893 4721 3896
rect 4755 3893 4767 3927
rect 4709 3887 4767 3893
rect 4801 3927 4859 3933
rect 4801 3893 4813 3927
rect 4847 3924 4859 3927
rect 5074 3924 5080 3936
rect 4847 3896 5080 3924
rect 4847 3893 4859 3896
rect 4801 3887 4859 3893
rect 5074 3884 5080 3896
rect 5132 3884 5138 3936
rect 5184 3933 5212 3964
rect 6086 3952 6092 3964
rect 6144 3952 6150 4004
rect 5169 3927 5227 3933
rect 5169 3893 5181 3927
rect 5215 3893 5227 3927
rect 5169 3887 5227 3893
rect 5258 3884 5264 3936
rect 5316 3924 5322 3936
rect 5537 3927 5595 3933
rect 5537 3924 5549 3927
rect 5316 3896 5549 3924
rect 5316 3884 5322 3896
rect 5537 3893 5549 3896
rect 5583 3893 5595 3927
rect 5537 3887 5595 3893
rect 5629 3927 5687 3933
rect 5629 3893 5641 3927
rect 5675 3924 5687 3927
rect 6380 3924 6408 4168
rect 7101 4165 7113 4168
rect 7147 4165 7159 4199
rect 7101 4159 7159 4165
rect 6457 4131 6515 4137
rect 6457 4097 6469 4131
rect 6503 4097 6515 4131
rect 6457 4091 6515 4097
rect 6549 4131 6607 4137
rect 6549 4097 6561 4131
rect 6595 4128 6607 4131
rect 6638 4128 6644 4140
rect 6595 4100 6644 4128
rect 6595 4097 6607 4100
rect 6549 4091 6607 4097
rect 6472 4060 6500 4091
rect 6638 4088 6644 4100
rect 6696 4088 6702 4140
rect 6822 4088 6828 4140
rect 6880 4128 6886 4140
rect 7190 4128 7196 4140
rect 6880 4100 7196 4128
rect 6880 4088 6886 4100
rect 7190 4088 7196 4100
rect 7248 4128 7254 4140
rect 7377 4131 7435 4137
rect 7377 4128 7389 4131
rect 7248 4100 7389 4128
rect 7248 4088 7254 4100
rect 7377 4097 7389 4100
rect 7423 4097 7435 4131
rect 7377 4091 7435 4097
rect 6472 4032 7144 4060
rect 6546 3952 6552 4004
rect 6604 3992 6610 4004
rect 7116 3992 7144 4032
rect 7392 3992 7420 4091
rect 7484 4069 7512 4236
rect 9214 4224 9220 4276
rect 9272 4264 9278 4276
rect 9272 4236 9904 4264
rect 9272 4224 9278 4236
rect 8294 4156 8300 4208
rect 8352 4156 8358 4208
rect 8312 4128 8340 4156
rect 8938 4128 8944 4140
rect 8174 4100 8340 4128
rect 8496 4100 8944 4128
rect 7469 4063 7527 4069
rect 7469 4029 7481 4063
rect 7515 4029 7527 4063
rect 7742 4060 7748 4072
rect 7703 4032 7748 4060
rect 7469 4023 7527 4029
rect 7742 4020 7748 4032
rect 7800 4020 7806 4072
rect 7926 4060 7932 4072
rect 7887 4032 7932 4060
rect 7926 4020 7932 4032
rect 7984 4020 7990 4072
rect 8018 4020 8024 4072
rect 8076 4060 8082 4072
rect 8174 4069 8202 4100
rect 8159 4063 8217 4069
rect 8076 4032 8121 4060
rect 8076 4020 8082 4032
rect 8159 4029 8171 4063
rect 8205 4029 8217 4063
rect 8159 4023 8217 4029
rect 8294 4020 8300 4072
rect 8352 4060 8358 4072
rect 8496 4069 8524 4100
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 8481 4063 8539 4069
rect 8352 4032 8397 4060
rect 8352 4020 8358 4032
rect 8481 4029 8493 4063
rect 8527 4029 8539 4063
rect 8662 4060 8668 4072
rect 8623 4032 8668 4060
rect 8481 4023 8539 4029
rect 8662 4020 8668 4032
rect 8720 4020 8726 4072
rect 9030 4060 9036 4072
rect 8991 4032 9036 4060
rect 9030 4020 9036 4032
rect 9088 4020 9094 4072
rect 9876 4060 9904 4236
rect 10594 4224 10600 4276
rect 10652 4264 10658 4276
rect 15838 4264 15844 4276
rect 10652 4236 15844 4264
rect 10652 4224 10658 4236
rect 15838 4224 15844 4236
rect 15896 4224 15902 4276
rect 16104 4267 16162 4273
rect 16104 4233 16116 4267
rect 16150 4264 16162 4267
rect 17954 4264 17960 4276
rect 16150 4236 17960 4264
rect 16150 4233 16162 4236
rect 16104 4227 16162 4233
rect 17954 4224 17960 4236
rect 18012 4224 18018 4276
rect 15243 4199 15301 4205
rect 15243 4196 15255 4199
rect 14844 4168 15255 4196
rect 10459 4131 10517 4137
rect 10459 4097 10471 4131
rect 10505 4128 10517 4131
rect 11422 4128 11428 4140
rect 10505 4100 11100 4128
rect 11383 4100 11428 4128
rect 10505 4097 10517 4100
rect 10459 4091 10517 4097
rect 11072 4072 11100 4100
rect 11422 4088 11428 4100
rect 11480 4088 11486 4140
rect 13446 4088 13452 4140
rect 13504 4128 13510 4140
rect 13504 4100 13549 4128
rect 13504 4088 13510 4100
rect 13722 4088 13728 4140
rect 13780 4128 13786 4140
rect 14844 4128 14872 4168
rect 15243 4165 15255 4168
rect 15289 4165 15301 4199
rect 15243 4159 15301 4165
rect 17218 4156 17224 4208
rect 17276 4196 17282 4208
rect 17770 4196 17776 4208
rect 17276 4168 17776 4196
rect 17276 4156 17282 4168
rect 17770 4156 17776 4168
rect 17828 4156 17834 4208
rect 18046 4196 18052 4208
rect 18007 4168 18052 4196
rect 18046 4156 18052 4168
rect 18104 4156 18110 4208
rect 13780 4100 14872 4128
rect 13780 4088 13786 4100
rect 10778 4060 10784 4072
rect 9876 4032 10784 4060
rect 10778 4020 10784 4032
rect 10836 4020 10842 4072
rect 11054 4060 11060 4072
rect 11015 4032 11060 4060
rect 11054 4020 11060 4032
rect 11112 4020 11118 4072
rect 11241 4063 11299 4069
rect 11241 4029 11253 4063
rect 11287 4060 11299 4063
rect 11330 4060 11336 4072
rect 11287 4032 11336 4060
rect 11287 4029 11299 4032
rect 11241 4023 11299 4029
rect 11330 4020 11336 4032
rect 11388 4020 11394 4072
rect 11793 4063 11851 4069
rect 11793 4029 11805 4063
rect 11839 4060 11851 4063
rect 11882 4060 11888 4072
rect 11839 4032 11888 4060
rect 11839 4029 11851 4032
rect 11793 4023 11851 4029
rect 11882 4020 11888 4032
rect 11940 4020 11946 4072
rect 13219 4063 13277 4069
rect 13219 4029 13231 4063
rect 13265 4060 13277 4063
rect 13817 4063 13875 4069
rect 13817 4060 13829 4063
rect 13265 4054 13492 4060
rect 13556 4054 13829 4060
rect 13265 4032 13829 4054
rect 13265 4029 13277 4032
rect 13219 4023 13277 4029
rect 13464 4026 13584 4032
rect 13817 4029 13829 4032
rect 13863 4029 13875 4063
rect 14844 4060 14872 4100
rect 14918 4088 14924 4140
rect 14976 4128 14982 4140
rect 15841 4131 15899 4137
rect 15841 4128 15853 4131
rect 14976 4100 15853 4128
rect 14976 4088 14982 4100
rect 15841 4097 15853 4100
rect 15887 4097 15899 4131
rect 15841 4091 15899 4097
rect 16114 4088 16120 4140
rect 16172 4128 16178 4140
rect 16574 4128 16580 4140
rect 16172 4100 16580 4128
rect 16172 4088 16178 4100
rect 16574 4088 16580 4100
rect 16632 4088 16638 4140
rect 16758 4088 16764 4140
rect 16816 4128 16822 4140
rect 18230 4128 18236 4140
rect 16816 4100 17724 4128
rect 18191 4100 18236 4128
rect 16816 4088 16822 4100
rect 14844 4032 15148 4060
rect 13817 4023 13875 4029
rect 6604 3964 7052 3992
rect 7116 3964 7236 3992
rect 7392 3964 8248 3992
rect 6604 3952 6610 3964
rect 5675 3896 6408 3924
rect 6641 3927 6699 3933
rect 5675 3893 5687 3896
rect 5629 3887 5687 3893
rect 6641 3893 6653 3927
rect 6687 3924 6699 3927
rect 6730 3924 6736 3936
rect 6687 3896 6736 3924
rect 6687 3893 6699 3896
rect 6641 3887 6699 3893
rect 6730 3884 6736 3896
rect 6788 3884 6794 3936
rect 7024 3933 7052 3964
rect 7009 3927 7067 3933
rect 7009 3893 7021 3927
rect 7055 3893 7067 3927
rect 7208 3924 7236 3964
rect 8220 3936 8248 3964
rect 9766 3952 9772 4004
rect 9824 3952 9830 4004
rect 10689 3995 10747 4001
rect 10689 3992 10701 3995
rect 10152 3964 10701 3992
rect 7745 3927 7803 3933
rect 7745 3924 7757 3927
rect 7208 3896 7757 3924
rect 7009 3887 7067 3893
rect 7745 3893 7757 3896
rect 7791 3924 7803 3927
rect 8110 3924 8116 3936
rect 7791 3896 8116 3924
rect 7791 3893 7803 3896
rect 7745 3887 7803 3893
rect 8110 3884 8116 3896
rect 8168 3884 8174 3936
rect 8202 3884 8208 3936
rect 8260 3884 8266 3936
rect 8386 3924 8392 3936
rect 8347 3896 8392 3924
rect 8386 3884 8392 3896
rect 8444 3884 8450 3936
rect 8570 3884 8576 3936
rect 8628 3924 8634 3936
rect 10152 3924 10180 3964
rect 10689 3961 10701 3964
rect 10735 3961 10747 3995
rect 12986 3992 12992 4004
rect 12834 3964 12992 3992
rect 10689 3955 10747 3961
rect 12986 3952 12992 3964
rect 13044 3952 13050 4004
rect 15010 3992 15016 4004
rect 14858 3964 15016 3992
rect 15010 3952 15016 3964
rect 15068 3952 15074 4004
rect 15120 3992 15148 4032
rect 15194 4020 15200 4072
rect 15252 4060 15258 4072
rect 17696 4069 17724 4100
rect 18230 4088 18236 4100
rect 18288 4128 18294 4140
rect 18598 4128 18604 4140
rect 18288 4100 18604 4128
rect 18288 4088 18294 4100
rect 18598 4088 18604 4100
rect 18656 4088 18662 4140
rect 15473 4063 15531 4069
rect 15473 4060 15485 4063
rect 15252 4032 15485 4060
rect 15252 4020 15258 4032
rect 15473 4029 15485 4032
rect 15519 4029 15531 4063
rect 15473 4023 15531 4029
rect 17681 4063 17739 4069
rect 17681 4029 17693 4063
rect 17727 4029 17739 4063
rect 17681 4023 17739 4029
rect 17774 4063 17832 4069
rect 17774 4029 17786 4063
rect 17820 4029 17832 4063
rect 17774 4023 17832 4029
rect 16114 3992 16120 4004
rect 15120 3964 16120 3992
rect 16114 3952 16120 3964
rect 16172 3952 16178 4004
rect 16574 3952 16580 4004
rect 16632 3952 16638 4004
rect 17789 3992 17817 4023
rect 18046 4020 18052 4072
rect 18104 4060 18110 4072
rect 18417 4063 18475 4069
rect 18417 4060 18429 4063
rect 18104 4032 18429 4060
rect 18104 4020 18110 4032
rect 18417 4029 18429 4032
rect 18463 4029 18475 4063
rect 18417 4023 18475 4029
rect 18506 4020 18512 4072
rect 18564 4060 18570 4072
rect 18564 4032 18609 4060
rect 18564 4020 18570 4032
rect 17512 3964 17817 3992
rect 8628 3896 10180 3924
rect 8628 3884 8634 3896
rect 10778 3884 10784 3936
rect 10836 3924 10842 3936
rect 11057 3927 11115 3933
rect 11057 3924 11069 3927
rect 10836 3896 11069 3924
rect 10836 3884 10842 3896
rect 11057 3893 11069 3896
rect 11103 3893 11115 3927
rect 11057 3887 11115 3893
rect 15194 3884 15200 3936
rect 15252 3924 15258 3936
rect 15565 3927 15623 3933
rect 15565 3924 15577 3927
rect 15252 3896 15577 3924
rect 15252 3884 15258 3896
rect 15565 3893 15577 3896
rect 15611 3893 15623 3927
rect 15565 3887 15623 3893
rect 15930 3884 15936 3936
rect 15988 3924 15994 3936
rect 16482 3924 16488 3936
rect 15988 3896 16488 3924
rect 15988 3884 15994 3896
rect 16482 3884 16488 3896
rect 16540 3884 16546 3936
rect 17126 3884 17132 3936
rect 17184 3924 17190 3936
rect 17512 3924 17540 3964
rect 17184 3896 17540 3924
rect 17589 3927 17647 3933
rect 17184 3884 17190 3896
rect 17589 3893 17601 3927
rect 17635 3924 17647 3927
rect 17678 3924 17684 3936
rect 17635 3896 17684 3924
rect 17635 3893 17647 3896
rect 17589 3887 17647 3893
rect 17678 3884 17684 3896
rect 17736 3884 17742 3936
rect 18230 3924 18236 3936
rect 18191 3896 18236 3924
rect 18230 3884 18236 3896
rect 18288 3884 18294 3936
rect 184 3834 18860 3856
rect 184 3782 4660 3834
rect 4712 3782 4724 3834
rect 4776 3782 4788 3834
rect 4840 3782 4852 3834
rect 4904 3782 4916 3834
rect 4968 3782 7760 3834
rect 7812 3782 7824 3834
rect 7876 3782 7888 3834
rect 7940 3782 7952 3834
rect 8004 3782 8016 3834
rect 8068 3782 10860 3834
rect 10912 3782 10924 3834
rect 10976 3782 10988 3834
rect 11040 3782 11052 3834
rect 11104 3782 11116 3834
rect 11168 3782 13960 3834
rect 14012 3782 14024 3834
rect 14076 3782 14088 3834
rect 14140 3782 14152 3834
rect 14204 3782 14216 3834
rect 14268 3782 17060 3834
rect 17112 3782 17124 3834
rect 17176 3782 17188 3834
rect 17240 3782 17252 3834
rect 17304 3782 17316 3834
rect 17368 3782 18860 3834
rect 184 3760 18860 3782
rect 2222 3680 2228 3732
rect 2280 3720 2286 3732
rect 2501 3723 2559 3729
rect 2501 3720 2513 3723
rect 2280 3692 2513 3720
rect 2280 3680 2286 3692
rect 2501 3689 2513 3692
rect 2547 3689 2559 3723
rect 4246 3720 4252 3732
rect 2501 3683 2559 3689
rect 2746 3692 4252 3720
rect 2133 3655 2191 3661
rect 2133 3621 2145 3655
rect 2179 3652 2191 3655
rect 2746 3652 2774 3692
rect 4246 3680 4252 3692
rect 4304 3680 4310 3732
rect 5074 3680 5080 3732
rect 5132 3720 5138 3732
rect 7285 3723 7343 3729
rect 7285 3720 7297 3723
rect 5132 3692 7297 3720
rect 5132 3680 5138 3692
rect 7285 3689 7297 3692
rect 7331 3720 7343 3723
rect 7331 3692 8064 3720
rect 7331 3689 7343 3692
rect 7285 3683 7343 3689
rect 2179 3624 2774 3652
rect 2179 3621 2191 3624
rect 2133 3615 2191 3621
rect 3602 3612 3608 3664
rect 3660 3612 3666 3664
rect 4430 3612 4436 3664
rect 4488 3652 4494 3664
rect 4709 3655 4767 3661
rect 4709 3652 4721 3655
rect 4488 3624 4721 3652
rect 4488 3612 4494 3624
rect 4709 3621 4721 3624
rect 4755 3652 4767 3655
rect 4982 3652 4988 3664
rect 4755 3624 4988 3652
rect 4755 3621 4767 3624
rect 4709 3615 4767 3621
rect 4982 3612 4988 3624
rect 5040 3612 5046 3664
rect 5350 3612 5356 3664
rect 5408 3652 5414 3664
rect 6089 3655 6147 3661
rect 6089 3652 6101 3655
rect 5408 3624 6101 3652
rect 5408 3612 5414 3624
rect 6089 3621 6101 3624
rect 6135 3652 6147 3655
rect 6135 3624 7788 3652
rect 6135 3621 6147 3624
rect 6089 3615 6147 3621
rect 7760 3596 7788 3624
rect 2041 3587 2099 3593
rect 2041 3553 2053 3587
rect 2087 3584 2099 3587
rect 2590 3584 2596 3596
rect 2087 3556 2596 3584
rect 2087 3553 2099 3556
rect 2041 3547 2099 3553
rect 2590 3544 2596 3556
rect 2648 3544 2654 3596
rect 4890 3584 4896 3596
rect 4851 3556 4896 3584
rect 4890 3544 4896 3556
rect 4948 3544 4954 3596
rect 5166 3584 5172 3596
rect 5127 3556 5172 3584
rect 5166 3544 5172 3556
rect 5224 3544 5230 3596
rect 5707 3587 5765 3593
rect 5707 3553 5719 3587
rect 5753 3584 5765 3587
rect 5810 3584 5816 3596
rect 5753 3556 5816 3584
rect 5753 3553 5765 3556
rect 5707 3547 5765 3553
rect 5810 3544 5816 3556
rect 5868 3544 5874 3596
rect 6365 3587 6423 3593
rect 6365 3553 6377 3587
rect 6411 3553 6423 3587
rect 6365 3547 6423 3553
rect 6457 3587 6515 3593
rect 6457 3553 6469 3587
rect 6503 3553 6515 3587
rect 6457 3547 6515 3553
rect 1949 3519 2007 3525
rect 1949 3485 1961 3519
rect 1995 3485 2007 3519
rect 1949 3479 2007 3485
rect 1964 3448 1992 3479
rect 2498 3476 2504 3528
rect 2556 3516 2562 3528
rect 2685 3519 2743 3525
rect 2685 3516 2697 3519
rect 2556 3488 2697 3516
rect 2556 3476 2562 3488
rect 2685 3485 2697 3488
rect 2731 3485 2743 3519
rect 2958 3516 2964 3528
rect 2919 3488 2964 3516
rect 2685 3479 2743 3485
rect 2958 3476 2964 3488
rect 3016 3476 3022 3528
rect 5534 3516 5540 3528
rect 5495 3488 5540 3516
rect 5534 3476 5540 3488
rect 5592 3476 5598 3528
rect 6086 3476 6092 3528
rect 6144 3516 6150 3528
rect 6380 3516 6408 3547
rect 6144 3488 6408 3516
rect 6472 3516 6500 3547
rect 6546 3544 6552 3596
rect 6604 3584 6610 3596
rect 6604 3556 6649 3584
rect 6604 3544 6610 3556
rect 6730 3544 6736 3596
rect 6788 3584 6794 3596
rect 6825 3587 6883 3593
rect 6825 3584 6837 3587
rect 6788 3556 6837 3584
rect 6788 3544 6794 3556
rect 6825 3553 6837 3556
rect 6871 3553 6883 3587
rect 6825 3547 6883 3553
rect 7101 3587 7159 3593
rect 7101 3553 7113 3587
rect 7147 3584 7159 3587
rect 7190 3584 7196 3596
rect 7147 3556 7196 3584
rect 7147 3553 7159 3556
rect 7101 3547 7159 3553
rect 7190 3544 7196 3556
rect 7248 3544 7254 3596
rect 7742 3584 7748 3596
rect 7655 3556 7748 3584
rect 7742 3544 7748 3556
rect 7800 3544 7806 3596
rect 7926 3593 7932 3596
rect 7910 3587 7932 3593
rect 7910 3553 7922 3587
rect 7910 3547 7932 3553
rect 7926 3544 7932 3547
rect 7984 3544 7990 3596
rect 8036 3593 8064 3692
rect 8110 3680 8116 3732
rect 8168 3680 8174 3732
rect 8202 3680 8208 3732
rect 8260 3720 8266 3732
rect 8260 3692 8432 3720
rect 8260 3680 8266 3692
rect 8128 3652 8156 3680
rect 8294 3652 8300 3664
rect 8128 3624 8300 3652
rect 8294 3612 8300 3624
rect 8352 3612 8358 3664
rect 8404 3652 8432 3692
rect 8662 3680 8668 3732
rect 8720 3720 8726 3732
rect 9953 3723 10011 3729
rect 9953 3720 9965 3723
rect 8720 3692 9965 3720
rect 8720 3680 8726 3692
rect 9953 3689 9965 3692
rect 9999 3689 10011 3723
rect 9953 3683 10011 3689
rect 10042 3680 10048 3732
rect 10100 3720 10106 3732
rect 13357 3723 13415 3729
rect 13357 3720 13369 3723
rect 10100 3692 13369 3720
rect 10100 3680 10106 3692
rect 13357 3689 13369 3692
rect 13403 3720 13415 3723
rect 13446 3720 13452 3732
rect 13403 3692 13452 3720
rect 13403 3689 13415 3692
rect 13357 3683 13415 3689
rect 13446 3680 13452 3692
rect 13504 3680 13510 3732
rect 13541 3723 13599 3729
rect 13541 3689 13553 3723
rect 13587 3720 13599 3723
rect 13814 3720 13820 3732
rect 13587 3692 13820 3720
rect 13587 3689 13599 3692
rect 13541 3683 13599 3689
rect 13814 3680 13820 3692
rect 13872 3680 13878 3732
rect 13998 3680 14004 3732
rect 14056 3720 14062 3732
rect 14277 3723 14335 3729
rect 14277 3720 14289 3723
rect 14056 3692 14289 3720
rect 14056 3680 14062 3692
rect 14277 3689 14289 3692
rect 14323 3720 14335 3723
rect 14323 3692 14596 3720
rect 14323 3689 14335 3692
rect 14277 3683 14335 3689
rect 8754 3652 8760 3664
rect 8404 3624 8616 3652
rect 8715 3624 8760 3652
rect 8021 3587 8079 3593
rect 8021 3553 8033 3587
rect 8067 3553 8079 3587
rect 8021 3547 8079 3553
rect 8205 3587 8263 3593
rect 8205 3553 8217 3587
rect 8251 3553 8263 3587
rect 8588 3584 8616 3624
rect 8754 3612 8760 3624
rect 8812 3612 8818 3664
rect 9122 3612 9128 3664
rect 9180 3652 9186 3664
rect 10321 3655 10379 3661
rect 10321 3652 10333 3655
rect 9180 3624 10333 3652
rect 9180 3612 9186 3624
rect 10321 3621 10333 3624
rect 10367 3621 10379 3655
rect 10321 3615 10379 3621
rect 12894 3612 12900 3664
rect 12952 3652 12958 3664
rect 14568 3652 14596 3692
rect 14826 3680 14832 3732
rect 14884 3720 14890 3732
rect 14884 3692 14929 3720
rect 14884 3680 14890 3692
rect 15194 3680 15200 3732
rect 15252 3720 15258 3732
rect 18325 3723 18383 3729
rect 15252 3692 17264 3720
rect 15252 3680 15258 3692
rect 17037 3655 17095 3661
rect 17037 3652 17049 3655
rect 12952 3624 13308 3652
rect 14568 3624 17049 3652
rect 12952 3612 12958 3624
rect 8665 3587 8723 3593
rect 8665 3584 8677 3587
rect 8588 3556 8677 3584
rect 8205 3547 8263 3553
rect 8665 3553 8677 3556
rect 8711 3553 8723 3587
rect 8846 3584 8852 3596
rect 8807 3556 8852 3584
rect 8665 3547 8723 3553
rect 6638 3516 6644 3528
rect 6472 3488 6644 3516
rect 6144 3476 6150 3488
rect 6638 3476 6644 3488
rect 6696 3476 6702 3528
rect 7282 3476 7288 3528
rect 7340 3516 7346 3528
rect 7469 3519 7527 3525
rect 7469 3516 7481 3519
rect 7340 3488 7481 3516
rect 7340 3476 7346 3488
rect 7469 3485 7481 3488
rect 7515 3485 7527 3519
rect 7469 3479 7527 3485
rect 4525 3451 4583 3457
rect 1964 3420 2084 3448
rect 2056 3380 2084 3420
rect 4525 3417 4537 3451
rect 4571 3448 4583 3451
rect 5994 3448 6000 3460
rect 4571 3420 6000 3448
rect 4571 3417 4583 3420
rect 4525 3411 4583 3417
rect 5994 3408 6000 3420
rect 6052 3408 6058 3460
rect 6733 3451 6791 3457
rect 6733 3417 6745 3451
rect 6779 3448 6791 3451
rect 7098 3448 7104 3460
rect 6779 3420 7104 3448
rect 6779 3417 6791 3420
rect 6733 3411 6791 3417
rect 7098 3408 7104 3420
rect 7156 3408 7162 3460
rect 2866 3380 2872 3392
rect 2056 3352 2872 3380
rect 2866 3340 2872 3352
rect 2924 3380 2930 3392
rect 4062 3380 4068 3392
rect 2924 3352 4068 3380
rect 2924 3340 2930 3352
rect 4062 3340 4068 3352
rect 4120 3340 4126 3392
rect 4433 3383 4491 3389
rect 4433 3349 4445 3383
rect 4479 3380 4491 3383
rect 4614 3380 4620 3392
rect 4479 3352 4620 3380
rect 4479 3349 4491 3352
rect 4433 3343 4491 3349
rect 4614 3340 4620 3352
rect 4672 3340 4678 3392
rect 4982 3340 4988 3392
rect 5040 3380 5046 3392
rect 5258 3380 5264 3392
rect 5040 3352 5264 3380
rect 5040 3340 5046 3352
rect 5258 3340 5264 3352
rect 5316 3340 5322 3392
rect 5902 3380 5908 3392
rect 5863 3352 5908 3380
rect 5902 3340 5908 3352
rect 5960 3340 5966 3392
rect 6822 3340 6828 3392
rect 6880 3380 6886 3392
rect 6917 3383 6975 3389
rect 6917 3380 6929 3383
rect 6880 3352 6929 3380
rect 6880 3340 6886 3352
rect 6917 3349 6929 3352
rect 6963 3349 6975 3383
rect 6917 3343 6975 3349
rect 7650 3340 7656 3392
rect 7708 3380 7714 3392
rect 7745 3383 7803 3389
rect 7745 3380 7757 3383
rect 7708 3352 7757 3380
rect 7708 3340 7714 3352
rect 7745 3349 7757 3352
rect 7791 3349 7803 3383
rect 8018 3380 8024 3392
rect 7979 3352 8024 3380
rect 7745 3343 7803 3349
rect 8018 3340 8024 3352
rect 8076 3340 8082 3392
rect 8110 3340 8116 3392
rect 8168 3380 8174 3392
rect 8220 3380 8248 3547
rect 8846 3544 8852 3556
rect 8904 3544 8910 3596
rect 8938 3544 8944 3596
rect 8996 3584 9002 3596
rect 9217 3587 9275 3593
rect 9217 3584 9229 3587
rect 8996 3556 9229 3584
rect 8996 3544 9002 3556
rect 9217 3553 9229 3556
rect 9263 3584 9275 3587
rect 9766 3584 9772 3596
rect 9263 3556 9772 3584
rect 9263 3553 9275 3556
rect 9217 3547 9275 3553
rect 9766 3544 9772 3556
rect 9824 3544 9830 3596
rect 9950 3584 9956 3596
rect 9911 3556 9956 3584
rect 9950 3544 9956 3556
rect 10008 3584 10014 3596
rect 11606 3584 11612 3596
rect 10008 3556 11612 3584
rect 10008 3544 10014 3556
rect 11606 3544 11612 3556
rect 11664 3584 11670 3596
rect 11885 3587 11943 3593
rect 11885 3584 11897 3587
rect 11664 3556 11897 3584
rect 11664 3544 11670 3556
rect 11885 3553 11897 3556
rect 11931 3553 11943 3587
rect 13078 3584 13084 3596
rect 13039 3556 13084 3584
rect 11885 3547 11943 3553
rect 13078 3544 13084 3556
rect 13136 3544 13142 3596
rect 13280 3593 13308 3624
rect 17037 3621 17049 3624
rect 17083 3621 17095 3655
rect 17037 3615 17095 3621
rect 17126 3612 17132 3664
rect 17184 3612 17190 3664
rect 13265 3587 13323 3593
rect 13265 3553 13277 3587
rect 13311 3553 13323 3587
rect 13265 3547 13323 3553
rect 13708 3587 13766 3593
rect 13708 3553 13720 3587
rect 13754 3584 13766 3587
rect 13754 3553 13768 3584
rect 13708 3547 13768 3553
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3516 8447 3519
rect 8754 3516 8760 3528
rect 8435 3488 8760 3516
rect 8435 3485 8447 3488
rect 8389 3479 8447 3485
rect 8754 3476 8760 3488
rect 8812 3476 8818 3528
rect 9493 3519 9551 3525
rect 9493 3485 9505 3519
rect 9539 3516 9551 3519
rect 10686 3516 10692 3528
rect 9539 3488 10692 3516
rect 9539 3485 9551 3488
rect 9493 3479 9551 3485
rect 10686 3476 10692 3488
rect 10744 3476 10750 3528
rect 12158 3476 12164 3528
rect 12216 3516 12222 3528
rect 12253 3519 12311 3525
rect 12253 3516 12265 3519
rect 12216 3488 12265 3516
rect 12216 3476 12222 3488
rect 12253 3485 12265 3488
rect 12299 3485 12311 3519
rect 12253 3479 12311 3485
rect 12805 3519 12863 3525
rect 12805 3485 12817 3519
rect 12851 3485 12863 3519
rect 12805 3479 12863 3485
rect 12820 3448 12848 3479
rect 12986 3476 12992 3528
rect 13044 3516 13050 3528
rect 13538 3516 13544 3528
rect 13044 3488 13544 3516
rect 13044 3476 13050 3488
rect 13538 3476 13544 3488
rect 13596 3476 13602 3528
rect 13740 3516 13768 3547
rect 13814 3544 13820 3596
rect 13872 3584 13878 3596
rect 14093 3587 14151 3593
rect 13872 3556 13917 3584
rect 13872 3544 13878 3556
rect 14093 3553 14105 3587
rect 14139 3553 14151 3587
rect 14093 3547 14151 3553
rect 14108 3516 14136 3547
rect 14182 3544 14188 3596
rect 14240 3584 14246 3596
rect 14471 3587 14529 3593
rect 14240 3556 14285 3584
rect 14240 3544 14246 3556
rect 14471 3553 14483 3587
rect 14517 3584 14529 3587
rect 14517 3556 14842 3584
rect 14517 3553 14529 3556
rect 14471 3547 14529 3553
rect 14366 3516 14372 3528
rect 13740 3488 13860 3516
rect 14108 3488 14372 3516
rect 13832 3460 13860 3488
rect 14366 3476 14372 3488
rect 14424 3476 14430 3528
rect 14642 3476 14648 3528
rect 14700 3516 14706 3528
rect 14700 3488 14745 3516
rect 14700 3476 14706 3488
rect 13722 3448 13728 3460
rect 8864 3420 13728 3448
rect 8478 3380 8484 3392
rect 8168 3352 8248 3380
rect 8439 3352 8484 3380
rect 8168 3340 8174 3352
rect 8478 3340 8484 3352
rect 8536 3340 8542 3392
rect 8570 3340 8576 3392
rect 8628 3380 8634 3392
rect 8864 3380 8892 3420
rect 13722 3408 13728 3420
rect 13780 3408 13786 3460
rect 13814 3408 13820 3460
rect 13872 3408 13878 3460
rect 14001 3451 14059 3457
rect 14001 3417 14013 3451
rect 14047 3448 14059 3451
rect 14660 3448 14688 3476
rect 14047 3420 14688 3448
rect 14047 3417 14059 3420
rect 14001 3411 14059 3417
rect 14814 3392 14842 3556
rect 15930 3544 15936 3596
rect 15988 3593 15994 3596
rect 15988 3584 16000 3593
rect 16206 3584 16212 3596
rect 15988 3556 16033 3584
rect 16167 3556 16212 3584
rect 15988 3547 16000 3556
rect 15988 3544 15994 3547
rect 16206 3544 16212 3556
rect 16264 3544 16270 3596
rect 16482 3584 16488 3596
rect 16443 3556 16488 3584
rect 16482 3544 16488 3556
rect 16540 3544 16546 3596
rect 16853 3587 16911 3593
rect 16853 3553 16865 3587
rect 16899 3584 16911 3587
rect 17144 3584 17172 3612
rect 16899 3556 17172 3584
rect 17236 3584 17264 3692
rect 18325 3689 18337 3723
rect 18371 3720 18383 3723
rect 19058 3720 19064 3732
rect 18371 3692 19064 3720
rect 18371 3689 18383 3692
rect 18325 3683 18383 3689
rect 19058 3680 19064 3692
rect 19116 3680 19122 3732
rect 18230 3652 18236 3664
rect 17972 3624 18236 3652
rect 17313 3587 17371 3593
rect 17313 3584 17325 3587
rect 17236 3556 17325 3584
rect 16899 3553 16911 3556
rect 16853 3547 16911 3553
rect 17313 3553 17325 3556
rect 17359 3553 17371 3587
rect 17678 3584 17684 3596
rect 17639 3556 17684 3584
rect 17313 3547 17371 3553
rect 17678 3544 17684 3556
rect 17736 3544 17742 3596
rect 17972 3593 18000 3624
rect 18230 3612 18236 3624
rect 18288 3612 18294 3664
rect 17957 3587 18015 3593
rect 17957 3553 17969 3587
rect 18003 3553 18015 3587
rect 17957 3547 18015 3553
rect 18049 3587 18107 3593
rect 18049 3553 18061 3587
rect 18095 3584 18107 3587
rect 18414 3584 18420 3596
rect 18095 3556 18420 3584
rect 18095 3553 18107 3556
rect 18049 3547 18107 3553
rect 18414 3544 18420 3556
rect 18472 3544 18478 3596
rect 18509 3587 18567 3593
rect 18509 3553 18521 3587
rect 18555 3584 18567 3587
rect 18874 3584 18880 3596
rect 18555 3556 18880 3584
rect 18555 3553 18567 3556
rect 18509 3547 18567 3553
rect 18874 3544 18880 3556
rect 18932 3544 18938 3596
rect 17129 3519 17187 3525
rect 17129 3516 17141 3519
rect 16224 3488 17141 3516
rect 16224 3460 16252 3488
rect 17129 3485 17141 3488
rect 17175 3485 17187 3519
rect 17129 3479 17187 3485
rect 17218 3476 17224 3528
rect 17276 3516 17282 3528
rect 17276 3488 17321 3516
rect 17276 3476 17282 3488
rect 17494 3476 17500 3528
rect 17552 3516 17558 3528
rect 17589 3519 17647 3525
rect 17589 3516 17601 3519
rect 17552 3488 17601 3516
rect 17552 3476 17558 3488
rect 17589 3485 17601 3488
rect 17635 3485 17647 3519
rect 17589 3479 17647 3485
rect 17773 3519 17831 3525
rect 17773 3485 17785 3519
rect 17819 3516 17831 3519
rect 18598 3516 18604 3528
rect 17819 3488 18604 3516
rect 17819 3485 17831 3488
rect 17773 3479 17831 3485
rect 18432 3460 18460 3488
rect 18598 3476 18604 3488
rect 18656 3476 18662 3528
rect 16206 3408 16212 3460
rect 16264 3408 16270 3460
rect 16298 3408 16304 3460
rect 16356 3448 16362 3460
rect 16482 3448 16488 3460
rect 16356 3420 16488 3448
rect 16356 3408 16362 3420
rect 16482 3408 16488 3420
rect 16540 3408 16546 3460
rect 17954 3408 17960 3460
rect 18012 3448 18018 3460
rect 18233 3451 18291 3457
rect 18233 3448 18245 3451
rect 18012 3420 18245 3448
rect 18012 3408 18018 3420
rect 18233 3417 18245 3420
rect 18279 3417 18291 3451
rect 18233 3411 18291 3417
rect 18414 3408 18420 3460
rect 18472 3408 18478 3460
rect 9122 3380 9128 3392
rect 8628 3352 8892 3380
rect 9083 3352 9128 3380
rect 8628 3340 8634 3352
rect 9122 3340 9128 3352
rect 9180 3340 9186 3392
rect 9214 3340 9220 3392
rect 9272 3380 9278 3392
rect 12066 3380 12072 3392
rect 9272 3352 12072 3380
rect 9272 3340 9278 3352
rect 12066 3340 12072 3352
rect 12124 3340 12130 3392
rect 12250 3340 12256 3392
rect 12308 3380 12314 3392
rect 12986 3380 12992 3392
rect 12308 3352 12992 3380
rect 12308 3340 12314 3352
rect 12986 3340 12992 3352
rect 13044 3340 13050 3392
rect 13446 3340 13452 3392
rect 13504 3380 13510 3392
rect 13906 3380 13912 3392
rect 13504 3352 13912 3380
rect 13504 3340 13510 3352
rect 13906 3340 13912 3352
rect 13964 3340 13970 3392
rect 14090 3340 14096 3392
rect 14148 3380 14154 3392
rect 14461 3383 14519 3389
rect 14461 3380 14473 3383
rect 14148 3352 14473 3380
rect 14148 3340 14154 3352
rect 14461 3349 14473 3352
rect 14507 3349 14519 3383
rect 14814 3380 14832 3392
rect 14739 3352 14832 3380
rect 14461 3343 14519 3349
rect 14826 3340 14832 3352
rect 14884 3380 14890 3392
rect 16666 3380 16672 3392
rect 14884 3352 16672 3380
rect 14884 3340 14890 3352
rect 16666 3340 16672 3352
rect 16724 3340 16730 3392
rect 17497 3383 17555 3389
rect 17497 3349 17509 3383
rect 17543 3380 17555 3383
rect 17770 3380 17776 3392
rect 17543 3352 17776 3380
rect 17543 3349 17555 3352
rect 17497 3343 17555 3349
rect 17770 3340 17776 3352
rect 17828 3340 17834 3392
rect 184 3290 18924 3312
rect 184 3238 3110 3290
rect 3162 3238 3174 3290
rect 3226 3238 3238 3290
rect 3290 3238 3302 3290
rect 3354 3238 3366 3290
rect 3418 3238 6210 3290
rect 6262 3238 6274 3290
rect 6326 3238 6338 3290
rect 6390 3238 6402 3290
rect 6454 3238 6466 3290
rect 6518 3238 9310 3290
rect 9362 3238 9374 3290
rect 9426 3238 9438 3290
rect 9490 3238 9502 3290
rect 9554 3238 9566 3290
rect 9618 3238 12410 3290
rect 12462 3238 12474 3290
rect 12526 3238 12538 3290
rect 12590 3238 12602 3290
rect 12654 3238 12666 3290
rect 12718 3238 15510 3290
rect 15562 3238 15574 3290
rect 15626 3238 15638 3290
rect 15690 3238 15702 3290
rect 15754 3238 15766 3290
rect 15818 3238 18610 3290
rect 18662 3238 18674 3290
rect 18726 3238 18738 3290
rect 18790 3238 18802 3290
rect 18854 3238 18866 3290
rect 18918 3238 18924 3290
rect 184 3216 18924 3238
rect 2958 3136 2964 3188
rect 3016 3176 3022 3188
rect 3881 3179 3939 3185
rect 3881 3176 3893 3179
rect 3016 3148 3893 3176
rect 3016 3136 3022 3148
rect 3881 3145 3893 3148
rect 3927 3145 3939 3179
rect 3881 3139 3939 3145
rect 4062 3136 4068 3188
rect 4120 3176 4126 3188
rect 6273 3179 6331 3185
rect 6273 3176 6285 3179
rect 4120 3148 6285 3176
rect 4120 3136 4126 3148
rect 2225 3043 2283 3049
rect 2225 3009 2237 3043
rect 2271 3040 2283 3043
rect 2774 3040 2780 3052
rect 2271 3012 2780 3040
rect 2271 3009 2283 3012
rect 2225 3003 2283 3009
rect 2774 3000 2780 3012
rect 2832 3000 2838 3052
rect 4338 3040 4344 3052
rect 4299 3012 4344 3040
rect 4338 3000 4344 3012
rect 4396 3000 4402 3052
rect 4540 3049 4568 3148
rect 6273 3145 6285 3148
rect 6319 3145 6331 3179
rect 7466 3176 7472 3188
rect 7427 3148 7472 3176
rect 6273 3139 6331 3145
rect 7466 3136 7472 3148
rect 7524 3136 7530 3188
rect 7558 3136 7564 3188
rect 7616 3176 7622 3188
rect 7745 3179 7803 3185
rect 7745 3176 7757 3179
rect 7616 3148 7757 3176
rect 7616 3136 7622 3148
rect 7745 3145 7757 3148
rect 7791 3145 7803 3179
rect 8478 3176 8484 3188
rect 7745 3139 7803 3145
rect 7852 3148 8484 3176
rect 6454 3068 6460 3120
rect 6512 3108 6518 3120
rect 6730 3108 6736 3120
rect 6512 3080 6736 3108
rect 6512 3068 6518 3080
rect 6730 3068 6736 3080
rect 6788 3108 6794 3120
rect 6788 3080 7328 3108
rect 6788 3068 6794 3080
rect 4525 3043 4583 3049
rect 4525 3009 4537 3043
rect 4571 3009 4583 3043
rect 4525 3003 4583 3009
rect 5353 3043 5411 3049
rect 5353 3009 5365 3043
rect 5399 3040 5411 3043
rect 6086 3040 6092 3052
rect 5399 3012 6092 3040
rect 5399 3009 5411 3012
rect 5353 3003 5411 3009
rect 6086 3000 6092 3012
rect 6144 3040 6150 3052
rect 7300 3049 7328 3080
rect 7374 3068 7380 3120
rect 7432 3108 7438 3120
rect 7432 3080 7477 3108
rect 7432 3068 7438 3080
rect 6825 3043 6883 3049
rect 6144 3012 6776 3040
rect 6144 3000 6150 3012
rect 1854 2972 1860 2984
rect 1815 2944 1860 2972
rect 1854 2932 1860 2944
rect 1912 2932 1918 2984
rect 3602 2972 3608 2984
rect 3252 2944 3608 2972
rect 3252 2890 3280 2944
rect 3602 2932 3608 2944
rect 3660 2932 3666 2984
rect 4246 2972 4252 2984
rect 4159 2944 4252 2972
rect 4246 2932 4252 2944
rect 4304 2972 4310 2984
rect 4614 2972 4620 2984
rect 4304 2944 4620 2972
rect 4304 2932 4310 2944
rect 4614 2932 4620 2944
rect 4672 2972 4678 2984
rect 5629 2975 5687 2981
rect 5629 2972 5641 2975
rect 4672 2944 5641 2972
rect 4672 2932 4678 2944
rect 5629 2941 5641 2944
rect 5675 2941 5687 2975
rect 5629 2935 5687 2941
rect 5994 2932 6000 2984
rect 6052 2972 6058 2984
rect 6748 2981 6776 3012
rect 6825 3009 6837 3043
rect 6871 3009 6883 3043
rect 6825 3003 6883 3009
rect 7285 3043 7343 3049
rect 7285 3009 7297 3043
rect 7331 3040 7343 3043
rect 7852 3040 7880 3148
rect 8478 3136 8484 3148
rect 8536 3176 8542 3188
rect 9214 3176 9220 3188
rect 8536 3148 9220 3176
rect 8536 3136 8542 3148
rect 9214 3136 9220 3148
rect 9272 3136 9278 3188
rect 11238 3176 11244 3188
rect 9784 3148 11244 3176
rect 7926 3068 7932 3120
rect 7984 3108 7990 3120
rect 8205 3111 8263 3117
rect 8205 3108 8217 3111
rect 7984 3080 8217 3108
rect 7984 3068 7990 3080
rect 8205 3077 8217 3080
rect 8251 3077 8263 3111
rect 8205 3071 8263 3077
rect 8294 3068 8300 3120
rect 8352 3108 8358 3120
rect 9493 3111 9551 3117
rect 9493 3108 9505 3111
rect 8352 3080 9505 3108
rect 8352 3068 8358 3080
rect 9493 3077 9505 3080
rect 9539 3077 9551 3111
rect 9493 3071 9551 3077
rect 7331 3012 7880 3040
rect 7331 3009 7343 3012
rect 7285 3003 7343 3009
rect 6641 2975 6699 2981
rect 6641 2972 6653 2975
rect 6052 2944 6653 2972
rect 6052 2932 6058 2944
rect 6641 2941 6653 2944
rect 6687 2941 6699 2975
rect 6641 2935 6699 2941
rect 6733 2975 6791 2981
rect 6733 2941 6745 2975
rect 6779 2941 6791 2975
rect 6840 2972 6868 3003
rect 8110 3000 8116 3052
rect 8168 3040 8174 3052
rect 8662 3040 8668 3052
rect 8168 3012 8668 3040
rect 8168 3000 8174 3012
rect 8662 3000 8668 3012
rect 8720 3040 8726 3052
rect 8757 3043 8815 3049
rect 8757 3040 8769 3043
rect 8720 3012 8769 3040
rect 8720 3000 8726 3012
rect 8757 3009 8769 3012
rect 8803 3009 8815 3043
rect 8757 3003 8815 3009
rect 8938 3000 8944 3052
rect 8996 3040 9002 3052
rect 9033 3043 9091 3049
rect 9033 3040 9045 3043
rect 8996 3012 9045 3040
rect 8996 3000 9002 3012
rect 9033 3009 9045 3012
rect 9079 3009 9091 3043
rect 9033 3003 9091 3009
rect 9125 3043 9183 3049
rect 9125 3009 9137 3043
rect 9171 3040 9183 3043
rect 9582 3040 9588 3052
rect 9171 3012 9588 3040
rect 9171 3009 9183 3012
rect 9125 3003 9183 3009
rect 9582 3000 9588 3012
rect 9640 3040 9646 3052
rect 9677 3043 9735 3049
rect 9677 3040 9689 3043
rect 9640 3012 9689 3040
rect 9640 3000 9646 3012
rect 9677 3009 9689 3012
rect 9723 3009 9735 3043
rect 9677 3003 9735 3009
rect 7377 2975 7435 2981
rect 6840 2944 7328 2972
rect 6733 2935 6791 2941
rect 3694 2904 3700 2916
rect 3655 2876 3700 2904
rect 3694 2864 3700 2876
rect 3752 2864 3758 2916
rect 4798 2904 4804 2916
rect 4264 2876 4804 2904
rect 1394 2796 1400 2848
rect 1452 2836 1458 2848
rect 4264 2836 4292 2876
rect 4798 2864 4804 2876
rect 4856 2864 4862 2916
rect 4890 2864 4896 2916
rect 4948 2904 4954 2916
rect 6086 2904 6092 2916
rect 4948 2876 5948 2904
rect 6047 2876 6092 2904
rect 4948 2864 4954 2876
rect 1452 2808 4292 2836
rect 1452 2796 1458 2808
rect 4338 2796 4344 2848
rect 4396 2836 4402 2848
rect 4709 2839 4767 2845
rect 4709 2836 4721 2839
rect 4396 2808 4721 2836
rect 4396 2796 4402 2808
rect 4709 2805 4721 2808
rect 4755 2805 4767 2839
rect 5074 2836 5080 2848
rect 5035 2808 5080 2836
rect 4709 2799 4767 2805
rect 5074 2796 5080 2808
rect 5132 2796 5138 2848
rect 5169 2839 5227 2845
rect 5169 2805 5181 2839
rect 5215 2836 5227 2839
rect 5350 2836 5356 2848
rect 5215 2808 5356 2836
rect 5215 2805 5227 2808
rect 5169 2799 5227 2805
rect 5350 2796 5356 2808
rect 5408 2796 5414 2848
rect 5920 2836 5948 2876
rect 6086 2864 6092 2876
rect 6144 2864 6150 2916
rect 6748 2904 6776 2935
rect 7006 2904 7012 2916
rect 6748 2876 7012 2904
rect 7006 2864 7012 2876
rect 7064 2864 7070 2916
rect 7101 2907 7159 2913
rect 7101 2873 7113 2907
rect 7147 2904 7159 2907
rect 7190 2904 7196 2916
rect 7147 2876 7196 2904
rect 7147 2873 7159 2876
rect 7101 2867 7159 2873
rect 7190 2864 7196 2876
rect 7248 2864 7254 2916
rect 7300 2904 7328 2944
rect 7377 2941 7389 2975
rect 7423 2972 7435 2975
rect 7466 2972 7472 2984
rect 7423 2944 7472 2972
rect 7423 2941 7435 2944
rect 7377 2935 7435 2941
rect 7466 2932 7472 2944
rect 7524 2932 7530 2984
rect 7742 2972 7748 2984
rect 7703 2944 7748 2972
rect 7742 2932 7748 2944
rect 7800 2932 7806 2984
rect 7834 2932 7840 2984
rect 7892 2972 7898 2984
rect 7929 2975 7987 2981
rect 7929 2972 7941 2975
rect 7892 2944 7941 2972
rect 7892 2932 7898 2944
rect 7929 2941 7941 2944
rect 7975 2941 7987 2975
rect 8386 2972 8392 2984
rect 8299 2944 8392 2972
rect 7929 2935 7987 2941
rect 8386 2932 8392 2944
rect 8444 2972 8450 2984
rect 8570 2972 8576 2984
rect 8444 2944 8576 2972
rect 8444 2932 8450 2944
rect 8570 2932 8576 2944
rect 8628 2932 8634 2984
rect 9217 2975 9275 2981
rect 9217 2941 9229 2975
rect 9263 2941 9275 2975
rect 9217 2935 9275 2941
rect 8294 2904 8300 2916
rect 7300 2876 8300 2904
rect 8294 2864 8300 2876
rect 8352 2864 8358 2916
rect 8846 2864 8852 2916
rect 8904 2904 8910 2916
rect 8941 2907 8999 2913
rect 8941 2904 8953 2907
rect 8904 2876 8953 2904
rect 8904 2864 8910 2876
rect 8941 2873 8953 2876
rect 8987 2873 8999 2907
rect 9232 2904 9260 2935
rect 9306 2932 9312 2984
rect 9364 2972 9370 2984
rect 9784 2981 9812 3148
rect 11238 3136 11244 3148
rect 11296 3136 11302 3188
rect 11330 3136 11336 3188
rect 11388 3185 11394 3188
rect 11388 3179 11437 3185
rect 11388 3145 11391 3179
rect 11425 3176 11437 3179
rect 13446 3176 13452 3188
rect 11425 3148 13452 3176
rect 11425 3145 11437 3148
rect 11388 3139 11437 3145
rect 11388 3136 11394 3139
rect 13446 3136 13452 3148
rect 13504 3136 13510 3188
rect 13541 3179 13599 3185
rect 13541 3145 13553 3179
rect 13587 3176 13599 3179
rect 13998 3176 14004 3188
rect 13587 3148 14004 3176
rect 13587 3145 13599 3148
rect 13541 3139 13599 3145
rect 13998 3136 14004 3148
rect 14056 3136 14062 3188
rect 17126 3136 17132 3188
rect 17184 3176 17190 3188
rect 17494 3176 17500 3188
rect 17184 3148 17500 3176
rect 17184 3136 17190 3148
rect 17494 3136 17500 3148
rect 17552 3176 17558 3188
rect 17862 3176 17868 3188
rect 17552 3148 17868 3176
rect 17552 3136 17558 3148
rect 17862 3136 17868 3148
rect 17920 3136 17926 3188
rect 18046 3176 18052 3188
rect 18007 3148 18052 3176
rect 18046 3136 18052 3148
rect 18104 3136 18110 3188
rect 15286 3068 15292 3120
rect 15344 3108 15350 3120
rect 15746 3108 15752 3120
rect 15344 3080 15752 3108
rect 15344 3068 15350 3080
rect 15746 3068 15752 3080
rect 15804 3068 15810 3120
rect 17310 3068 17316 3120
rect 17368 3108 17374 3120
rect 18325 3111 18383 3117
rect 18325 3108 18337 3111
rect 17368 3080 18337 3108
rect 17368 3068 17374 3080
rect 18325 3077 18337 3080
rect 18371 3077 18383 3111
rect 18325 3071 18383 3077
rect 10502 3040 10508 3052
rect 10428 3012 10508 3040
rect 9401 2975 9459 2981
rect 9401 2972 9413 2975
rect 9364 2944 9413 2972
rect 9364 2932 9370 2944
rect 9401 2941 9413 2944
rect 9447 2941 9459 2975
rect 9401 2935 9459 2941
rect 9769 2975 9827 2981
rect 9769 2941 9781 2975
rect 9815 2941 9827 2975
rect 9769 2935 9827 2941
rect 10134 2932 10140 2984
rect 10192 2972 10198 2984
rect 10321 2975 10379 2981
rect 10321 2972 10333 2975
rect 10192 2944 10333 2972
rect 10192 2932 10198 2944
rect 10321 2941 10333 2944
rect 10367 2941 10379 2975
rect 10321 2935 10379 2941
rect 10428 2904 10456 3012
rect 10502 3000 10508 3012
rect 10560 3000 10566 3052
rect 10873 3043 10931 3049
rect 10873 3009 10885 3043
rect 10919 3040 10931 3043
rect 12986 3040 12992 3052
rect 10919 3012 12992 3040
rect 10919 3009 10931 3012
rect 10873 3003 10931 3009
rect 12986 3000 12992 3012
rect 13044 3000 13050 3052
rect 13173 3043 13231 3049
rect 13173 3009 13185 3043
rect 13219 3040 13231 3043
rect 13725 3043 13783 3049
rect 13219 3012 13584 3040
rect 13219 3009 13231 3012
rect 13173 3003 13231 3009
rect 10689 2975 10747 2981
rect 10689 2941 10701 2975
rect 10735 2972 10747 2975
rect 10778 2972 10784 2984
rect 10735 2944 10784 2972
rect 10735 2941 10747 2944
rect 10689 2935 10747 2941
rect 10778 2932 10784 2944
rect 10836 2932 10842 2984
rect 11974 2972 11980 2984
rect 11348 2944 11980 2972
rect 9232 2876 10456 2904
rect 10487 2907 10545 2913
rect 8941 2867 8999 2873
rect 10487 2873 10499 2907
rect 10533 2904 10545 2907
rect 11348 2904 11376 2944
rect 11974 2932 11980 2944
rect 12032 2932 12038 2984
rect 12710 2932 12716 2984
rect 12768 2972 12774 2984
rect 12805 2975 12863 2981
rect 12805 2972 12817 2975
rect 12768 2944 12817 2972
rect 12768 2932 12774 2944
rect 12805 2941 12817 2944
rect 12851 2941 12863 2975
rect 12805 2935 12863 2941
rect 10533 2876 11376 2904
rect 10533 2873 10545 2876
rect 10487 2867 10545 2873
rect 6730 2836 6736 2848
rect 5920 2808 6736 2836
rect 6730 2796 6736 2808
rect 6788 2796 6794 2848
rect 7466 2796 7472 2848
rect 7524 2836 7530 2848
rect 7926 2836 7932 2848
rect 7524 2808 7932 2836
rect 7524 2796 7530 2808
rect 7926 2796 7932 2808
rect 7984 2796 7990 2848
rect 8662 2796 8668 2848
rect 8720 2836 8726 2848
rect 8757 2839 8815 2845
rect 8757 2836 8769 2839
rect 8720 2808 8769 2836
rect 8720 2796 8726 2808
rect 8757 2805 8769 2808
rect 8803 2805 8815 2839
rect 8956 2836 8984 2867
rect 12250 2864 12256 2916
rect 12308 2864 12314 2916
rect 13188 2904 13216 3003
rect 13446 2972 13452 2984
rect 13407 2944 13452 2972
rect 13446 2932 13452 2944
rect 13504 2932 13510 2984
rect 13556 2972 13584 3012
rect 13725 3009 13737 3043
rect 13771 3040 13783 3043
rect 14090 3040 14096 3052
rect 13771 3012 14096 3040
rect 13771 3009 13783 3012
rect 13725 3003 13783 3009
rect 14090 3000 14096 3012
rect 14148 3000 14154 3052
rect 14918 3000 14924 3052
rect 14976 3040 14982 3052
rect 15841 3043 15899 3049
rect 15841 3040 15853 3043
rect 14976 3012 15853 3040
rect 14976 3000 14982 3012
rect 15841 3009 15853 3012
rect 15887 3009 15899 3043
rect 15841 3003 15899 3009
rect 16117 3043 16175 3049
rect 16117 3009 16129 3043
rect 16163 3040 16175 3043
rect 17402 3040 17408 3052
rect 16163 3012 17408 3040
rect 16163 3009 16175 3012
rect 16117 3003 16175 3009
rect 17402 3000 17408 3012
rect 17460 3000 17466 3052
rect 13814 2972 13820 2984
rect 13556 2944 13820 2972
rect 13814 2932 13820 2944
rect 13872 2932 13878 2984
rect 14182 2972 14188 2984
rect 14143 2944 14188 2972
rect 14182 2932 14188 2944
rect 14240 2932 14246 2984
rect 17586 2932 17592 2984
rect 17644 2972 17650 2984
rect 17681 2975 17739 2981
rect 17681 2972 17693 2975
rect 17644 2944 17693 2972
rect 17644 2932 17650 2944
rect 17681 2941 17693 2944
rect 17727 2941 17739 2975
rect 17862 2972 17868 2984
rect 17823 2944 17868 2972
rect 17681 2935 17739 2941
rect 17862 2932 17868 2944
rect 17920 2932 17926 2984
rect 18509 2975 18567 2981
rect 18509 2941 18521 2975
rect 18555 2972 18567 2975
rect 18966 2972 18972 2984
rect 18555 2944 18972 2972
rect 18555 2941 18567 2944
rect 18509 2935 18567 2941
rect 13142 2876 13216 2904
rect 10594 2836 10600 2848
rect 8956 2808 10600 2836
rect 8757 2799 8815 2805
rect 10594 2796 10600 2808
rect 10652 2796 10658 2848
rect 11149 2839 11207 2845
rect 11149 2805 11161 2839
rect 11195 2836 11207 2839
rect 11238 2836 11244 2848
rect 11195 2808 11244 2836
rect 11195 2805 11207 2808
rect 11149 2799 11207 2805
rect 11238 2796 11244 2808
rect 11296 2796 11302 2848
rect 11606 2796 11612 2848
rect 11664 2836 11670 2848
rect 13142 2836 13170 2876
rect 13262 2864 13268 2916
rect 13320 2904 13326 2916
rect 13725 2907 13783 2913
rect 13725 2904 13737 2907
rect 13320 2876 13737 2904
rect 13320 2864 13326 2876
rect 13725 2873 13737 2876
rect 13771 2873 13783 2907
rect 13725 2867 13783 2873
rect 14550 2864 14556 2916
rect 14608 2864 14614 2916
rect 18524 2904 18552 2935
rect 18966 2932 18972 2944
rect 19024 2932 19030 2984
rect 15258 2876 16606 2904
rect 17420 2876 18552 2904
rect 11664 2808 13170 2836
rect 11664 2796 11670 2808
rect 13906 2796 13912 2848
rect 13964 2836 13970 2848
rect 14559 2836 14587 2864
rect 15102 2836 15108 2848
rect 13964 2808 15108 2836
rect 13964 2796 13970 2808
rect 15102 2796 15108 2808
rect 15160 2836 15166 2848
rect 15258 2836 15286 2876
rect 15160 2808 15286 2836
rect 15611 2839 15669 2845
rect 15160 2796 15166 2808
rect 15611 2805 15623 2839
rect 15657 2836 15669 2839
rect 15838 2836 15844 2848
rect 15657 2808 15844 2836
rect 15657 2805 15669 2808
rect 15611 2799 15669 2805
rect 15838 2796 15844 2808
rect 15896 2796 15902 2848
rect 15930 2796 15936 2848
rect 15988 2836 15994 2848
rect 17420 2836 17448 2876
rect 15988 2808 17448 2836
rect 17589 2839 17647 2845
rect 15988 2796 15994 2808
rect 17589 2805 17601 2839
rect 17635 2836 17647 2839
rect 17770 2836 17776 2848
rect 17635 2808 17776 2836
rect 17635 2805 17647 2808
rect 17589 2799 17647 2805
rect 17770 2796 17776 2808
rect 17828 2796 17834 2848
rect 184 2746 18860 2768
rect 184 2694 4660 2746
rect 4712 2694 4724 2746
rect 4776 2694 4788 2746
rect 4840 2694 4852 2746
rect 4904 2694 4916 2746
rect 4968 2694 7760 2746
rect 7812 2694 7824 2746
rect 7876 2694 7888 2746
rect 7940 2694 7952 2746
rect 8004 2694 8016 2746
rect 8068 2694 10860 2746
rect 10912 2694 10924 2746
rect 10976 2694 10988 2746
rect 11040 2694 11052 2746
rect 11104 2694 11116 2746
rect 11168 2694 13960 2746
rect 14012 2694 14024 2746
rect 14076 2694 14088 2746
rect 14140 2694 14152 2746
rect 14204 2694 14216 2746
rect 14268 2694 17060 2746
rect 17112 2694 17124 2746
rect 17176 2694 17188 2746
rect 17240 2694 17252 2746
rect 17304 2694 17316 2746
rect 17368 2694 18860 2746
rect 184 2672 18860 2694
rect 2774 2592 2780 2644
rect 2832 2632 2838 2644
rect 2869 2635 2927 2641
rect 2869 2632 2881 2635
rect 2832 2604 2881 2632
rect 2832 2592 2838 2604
rect 2869 2601 2881 2604
rect 2915 2601 2927 2635
rect 2869 2595 2927 2601
rect 3329 2635 3387 2641
rect 3329 2601 3341 2635
rect 3375 2632 3387 2635
rect 4338 2632 4344 2644
rect 3375 2604 4344 2632
rect 3375 2601 3387 2604
rect 3329 2595 3387 2601
rect 4338 2592 4344 2604
rect 4396 2592 4402 2644
rect 5169 2635 5227 2641
rect 5169 2601 5181 2635
rect 5215 2632 5227 2635
rect 5534 2632 5540 2644
rect 5215 2604 5540 2632
rect 5215 2601 5227 2604
rect 5169 2595 5227 2601
rect 5534 2592 5540 2604
rect 5592 2632 5598 2644
rect 6178 2632 6184 2644
rect 5592 2604 6184 2632
rect 5592 2592 5598 2604
rect 6178 2592 6184 2604
rect 6236 2592 6242 2644
rect 6454 2592 6460 2644
rect 6512 2592 6518 2644
rect 7190 2592 7196 2644
rect 7248 2632 7254 2644
rect 8754 2632 8760 2644
rect 7248 2604 8760 2632
rect 7248 2592 7254 2604
rect 1854 2524 1860 2576
rect 1912 2564 1918 2576
rect 1949 2567 2007 2573
rect 1949 2564 1961 2567
rect 1912 2536 1961 2564
rect 1912 2524 1918 2536
rect 1949 2533 1961 2536
rect 1995 2533 2007 2567
rect 1949 2527 2007 2533
rect 4172 2536 5120 2564
rect 2317 2499 2375 2505
rect 2317 2465 2329 2499
rect 2363 2496 2375 2499
rect 2498 2496 2504 2508
rect 2363 2468 2504 2496
rect 2363 2465 2375 2468
rect 2317 2459 2375 2465
rect 2498 2456 2504 2468
rect 2556 2456 2562 2508
rect 3237 2499 3295 2505
rect 3237 2465 3249 2499
rect 3283 2496 3295 2499
rect 3694 2496 3700 2508
rect 3283 2468 3700 2496
rect 3283 2465 3295 2468
rect 3237 2459 3295 2465
rect 3694 2456 3700 2468
rect 3752 2496 3758 2508
rect 3881 2499 3939 2505
rect 3881 2496 3893 2499
rect 3752 2468 3893 2496
rect 3752 2456 3758 2468
rect 3881 2465 3893 2468
rect 3927 2496 3939 2499
rect 4172 2496 4200 2536
rect 3927 2468 4200 2496
rect 3927 2465 3939 2468
rect 3881 2459 3939 2465
rect 3421 2431 3479 2437
rect 3421 2397 3433 2431
rect 3467 2397 3479 2431
rect 3786 2428 3792 2440
rect 3747 2400 3792 2428
rect 3421 2391 3479 2397
rect 2866 2320 2872 2372
rect 2924 2360 2930 2372
rect 3436 2360 3464 2391
rect 3786 2388 3792 2400
rect 3844 2388 3850 2440
rect 4172 2428 4200 2468
rect 4246 2456 4252 2508
rect 4304 2496 4310 2508
rect 5092 2505 5120 2536
rect 5994 2524 6000 2576
rect 6052 2564 6058 2576
rect 6472 2564 6500 2592
rect 6052 2536 6776 2564
rect 6052 2524 6058 2536
rect 4709 2499 4767 2505
rect 4709 2496 4721 2499
rect 4304 2468 4721 2496
rect 4304 2456 4310 2468
rect 4709 2465 4721 2468
rect 4755 2465 4767 2499
rect 4709 2459 4767 2465
rect 5077 2499 5135 2505
rect 5077 2465 5089 2499
rect 5123 2496 5135 2499
rect 5166 2496 5172 2508
rect 5123 2468 5172 2496
rect 5123 2465 5135 2468
rect 5077 2459 5135 2465
rect 4433 2431 4491 2437
rect 4433 2428 4445 2431
rect 4172 2400 4445 2428
rect 4433 2397 4445 2400
rect 4479 2397 4491 2431
rect 4724 2428 4752 2459
rect 5166 2456 5172 2468
rect 5224 2456 5230 2508
rect 5261 2499 5319 2505
rect 5261 2465 5273 2499
rect 5307 2465 5319 2499
rect 5718 2496 5724 2508
rect 5679 2468 5724 2496
rect 5261 2459 5319 2465
rect 5276 2428 5304 2459
rect 5718 2456 5724 2468
rect 5776 2456 5782 2508
rect 6086 2496 6092 2508
rect 6047 2468 6092 2496
rect 6086 2456 6092 2468
rect 6144 2456 6150 2508
rect 6748 2505 6776 2536
rect 7300 2505 7328 2604
rect 8754 2592 8760 2604
rect 8812 2592 8818 2644
rect 9030 2592 9036 2644
rect 9088 2632 9094 2644
rect 9309 2635 9367 2641
rect 9309 2632 9321 2635
rect 9088 2604 9321 2632
rect 9088 2592 9094 2604
rect 9309 2601 9321 2604
rect 9355 2601 9367 2635
rect 9309 2595 9367 2601
rect 10594 2592 10600 2644
rect 10652 2632 10658 2644
rect 12158 2632 12164 2644
rect 10652 2604 12164 2632
rect 10652 2592 10658 2604
rect 12158 2592 12164 2604
rect 12216 2592 12222 2644
rect 12250 2592 12256 2644
rect 12308 2592 12314 2644
rect 14274 2592 14280 2644
rect 14332 2632 14338 2644
rect 16301 2635 16359 2641
rect 14332 2604 14964 2632
rect 14332 2592 14338 2604
rect 9766 2564 9772 2576
rect 8970 2536 9772 2564
rect 9766 2524 9772 2536
rect 9824 2524 9830 2576
rect 12268 2564 12296 2592
rect 10902 2536 12296 2564
rect 13538 2524 13544 2576
rect 13596 2524 13602 2576
rect 13906 2524 13912 2576
rect 13964 2564 13970 2576
rect 14642 2564 14648 2576
rect 13964 2536 14648 2564
rect 13964 2524 13970 2536
rect 14642 2524 14648 2536
rect 14700 2524 14706 2576
rect 14936 2508 14964 2604
rect 16301 2601 16313 2635
rect 16347 2632 16359 2635
rect 19150 2632 19156 2644
rect 16347 2604 19156 2632
rect 16347 2601 16359 2604
rect 16301 2595 16359 2601
rect 19150 2592 19156 2604
rect 19208 2592 19214 2644
rect 16761 2567 16819 2573
rect 16761 2533 16773 2567
rect 16807 2564 16819 2567
rect 16850 2564 16856 2576
rect 16807 2536 16856 2564
rect 16807 2533 16819 2536
rect 16761 2527 16819 2533
rect 16850 2524 16856 2536
rect 16908 2524 16914 2576
rect 17126 2524 17132 2576
rect 17184 2564 17190 2576
rect 17184 2536 18092 2564
rect 17184 2524 17190 2536
rect 18064 2508 18092 2536
rect 6457 2499 6515 2505
rect 6457 2465 6469 2499
rect 6503 2465 6515 2499
rect 6457 2459 6515 2465
rect 6733 2499 6791 2505
rect 6733 2465 6745 2499
rect 6779 2465 6791 2499
rect 6733 2459 6791 2465
rect 7285 2499 7343 2505
rect 7285 2465 7297 2499
rect 7331 2465 7343 2499
rect 7285 2459 7343 2465
rect 4724 2400 5304 2428
rect 6472 2428 6500 2459
rect 9122 2456 9128 2508
rect 9180 2496 9186 2508
rect 9582 2496 9588 2508
rect 9180 2468 9444 2496
rect 9543 2468 9588 2496
rect 9180 2456 9186 2468
rect 7374 2428 7380 2440
rect 6472 2400 7380 2428
rect 4433 2391 4491 2397
rect 7374 2388 7380 2400
rect 7432 2388 7438 2440
rect 7469 2431 7527 2437
rect 7469 2397 7481 2431
rect 7515 2397 7527 2431
rect 7742 2428 7748 2440
rect 7703 2400 7748 2428
rect 7469 2391 7527 2397
rect 2924 2332 3464 2360
rect 3804 2360 3832 2388
rect 4525 2363 4583 2369
rect 4525 2360 4537 2363
rect 3804 2332 4537 2360
rect 2924 2320 2930 2332
rect 4525 2329 4537 2332
rect 4571 2329 4583 2363
rect 5074 2360 5080 2372
rect 4525 2323 4583 2329
rect 4632 2332 5080 2360
rect 4157 2295 4215 2301
rect 4157 2261 4169 2295
rect 4203 2292 4215 2295
rect 4632 2292 4660 2332
rect 5074 2320 5080 2332
rect 5132 2320 5138 2372
rect 7282 2320 7288 2372
rect 7340 2360 7346 2372
rect 7484 2360 7512 2391
rect 7742 2388 7748 2400
rect 7800 2388 7806 2440
rect 9309 2431 9367 2437
rect 9309 2428 9321 2431
rect 8864 2400 9321 2428
rect 8864 2372 8892 2400
rect 9309 2397 9321 2400
rect 9355 2397 9367 2431
rect 9309 2391 9367 2397
rect 7340 2332 7512 2360
rect 7340 2320 7346 2332
rect 8846 2320 8852 2372
rect 8904 2320 8910 2372
rect 8938 2320 8944 2372
rect 8996 2360 9002 2372
rect 9416 2360 9444 2468
rect 9582 2456 9588 2468
rect 9640 2456 9646 2508
rect 11606 2496 11612 2508
rect 11567 2468 11612 2496
rect 11606 2456 11612 2468
rect 11664 2496 11670 2508
rect 12253 2499 12311 2505
rect 12253 2496 12265 2499
rect 11664 2468 12265 2496
rect 11664 2456 11670 2468
rect 12253 2465 12265 2468
rect 12299 2465 12311 2499
rect 14182 2496 14188 2508
rect 14143 2468 14188 2496
rect 12253 2459 12311 2465
rect 14182 2456 14188 2468
rect 14240 2456 14246 2508
rect 14369 2499 14427 2505
rect 14369 2465 14381 2499
rect 14415 2496 14427 2499
rect 14734 2496 14740 2508
rect 14415 2468 14740 2496
rect 14415 2465 14427 2468
rect 14369 2459 14427 2465
rect 14734 2456 14740 2468
rect 14792 2456 14798 2508
rect 14918 2496 14924 2508
rect 14831 2468 14924 2496
rect 14918 2456 14924 2468
rect 14976 2456 14982 2508
rect 15194 2505 15200 2508
rect 15177 2499 15200 2505
rect 15177 2496 15189 2499
rect 15028 2468 15189 2496
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 11333 2431 11391 2437
rect 11333 2428 11345 2431
rect 9732 2400 11345 2428
rect 9732 2388 9738 2400
rect 11333 2397 11345 2400
rect 11379 2397 11391 2431
rect 12529 2431 12587 2437
rect 12529 2428 12541 2431
rect 11333 2391 11391 2397
rect 12268 2400 12541 2428
rect 12268 2372 12296 2400
rect 12529 2397 12541 2400
rect 12575 2397 12587 2431
rect 12529 2391 12587 2397
rect 13722 2388 13728 2440
rect 13780 2428 13786 2440
rect 15028 2428 15056 2468
rect 15177 2465 15189 2468
rect 15252 2496 15258 2508
rect 15252 2468 15325 2496
rect 15177 2459 15200 2465
rect 15194 2456 15200 2459
rect 15252 2456 15258 2468
rect 16666 2456 16672 2508
rect 16724 2456 16730 2508
rect 17034 2456 17040 2508
rect 17092 2496 17098 2508
rect 17405 2499 17463 2505
rect 17405 2496 17417 2499
rect 17092 2468 17417 2496
rect 17092 2456 17098 2468
rect 17405 2465 17417 2468
rect 17451 2465 17463 2499
rect 17405 2459 17463 2465
rect 18046 2456 18052 2508
rect 18104 2496 18110 2508
rect 18233 2499 18291 2505
rect 18233 2496 18245 2499
rect 18104 2468 18245 2496
rect 18104 2456 18110 2468
rect 18233 2465 18245 2468
rect 18279 2465 18291 2499
rect 18233 2459 18291 2465
rect 13780 2400 15056 2428
rect 16684 2428 16712 2456
rect 17129 2431 17187 2437
rect 17129 2428 17141 2431
rect 16684 2400 17141 2428
rect 13780 2388 13786 2400
rect 17129 2397 17141 2400
rect 17175 2397 17187 2431
rect 17129 2391 17187 2397
rect 17218 2388 17224 2440
rect 17276 2428 17282 2440
rect 17313 2431 17371 2437
rect 17313 2428 17325 2431
rect 17276 2400 17325 2428
rect 17276 2388 17282 2400
rect 17313 2397 17325 2400
rect 17359 2428 17371 2431
rect 17586 2428 17592 2440
rect 17359 2400 17592 2428
rect 17359 2397 17371 2400
rect 17313 2391 17371 2397
rect 17586 2388 17592 2400
rect 17644 2388 17650 2440
rect 17954 2388 17960 2440
rect 18012 2428 18018 2440
rect 18141 2431 18199 2437
rect 18141 2428 18153 2431
rect 18012 2400 18153 2428
rect 18012 2388 18018 2400
rect 18141 2397 18153 2400
rect 18187 2397 18199 2431
rect 18141 2391 18199 2397
rect 9493 2363 9551 2369
rect 9493 2360 9505 2363
rect 8996 2332 9260 2360
rect 9416 2332 9505 2360
rect 8996 2320 9002 2332
rect 4203 2264 4660 2292
rect 4203 2261 4215 2264
rect 4157 2255 4215 2261
rect 4798 2252 4804 2304
rect 4856 2292 4862 2304
rect 4893 2295 4951 2301
rect 4893 2292 4905 2295
rect 4856 2264 4905 2292
rect 4856 2252 4862 2264
rect 4893 2261 4905 2264
rect 4939 2261 4951 2295
rect 5442 2292 5448 2304
rect 5403 2264 5448 2292
rect 4893 2255 4951 2261
rect 5442 2252 5448 2264
rect 5500 2292 5506 2304
rect 6546 2292 6552 2304
rect 5500 2264 6552 2292
rect 5500 2252 5506 2264
rect 6546 2252 6552 2264
rect 6604 2252 6610 2304
rect 9232 2301 9260 2332
rect 9493 2329 9505 2332
rect 9539 2329 9551 2363
rect 9493 2323 9551 2329
rect 12250 2320 12256 2372
rect 12308 2320 12314 2372
rect 13814 2320 13820 2372
rect 13872 2360 13878 2372
rect 14274 2360 14280 2372
rect 13872 2332 14280 2360
rect 13872 2320 13878 2332
rect 14274 2320 14280 2332
rect 14332 2320 14338 2372
rect 14369 2363 14427 2369
rect 14369 2329 14381 2363
rect 14415 2360 14427 2363
rect 14415 2332 14964 2360
rect 14415 2329 14427 2332
rect 14369 2323 14427 2329
rect 9217 2295 9275 2301
rect 9217 2261 9229 2295
rect 9263 2261 9275 2295
rect 9217 2255 9275 2261
rect 9766 2252 9772 2304
rect 9824 2292 9830 2304
rect 9861 2295 9919 2301
rect 9861 2292 9873 2295
rect 9824 2264 9873 2292
rect 9824 2252 9830 2264
rect 9861 2261 9873 2264
rect 9907 2261 9919 2295
rect 9861 2255 9919 2261
rect 11885 2295 11943 2301
rect 11885 2261 11897 2295
rect 11931 2292 11943 2295
rect 11974 2292 11980 2304
rect 11931 2264 11980 2292
rect 11931 2261 11943 2264
rect 11885 2255 11943 2261
rect 11974 2252 11980 2264
rect 12032 2252 12038 2304
rect 12894 2252 12900 2304
rect 12952 2292 12958 2304
rect 14001 2295 14059 2301
rect 14001 2292 14013 2295
rect 12952 2264 14013 2292
rect 12952 2252 12958 2264
rect 14001 2261 14013 2264
rect 14047 2292 14059 2295
rect 14642 2292 14648 2304
rect 14047 2264 14648 2292
rect 14047 2261 14059 2264
rect 14001 2255 14059 2261
rect 14642 2252 14648 2264
rect 14700 2252 14706 2304
rect 14936 2292 14964 2332
rect 16666 2320 16672 2372
rect 16724 2360 16730 2372
rect 17865 2363 17923 2369
rect 17865 2360 17877 2363
rect 16724 2332 17877 2360
rect 16724 2320 16730 2332
rect 17865 2329 17877 2332
rect 17911 2329 17923 2363
rect 17865 2323 17923 2329
rect 16206 2292 16212 2304
rect 14936 2264 16212 2292
rect 16206 2252 16212 2264
rect 16264 2252 16270 2304
rect 16390 2252 16396 2304
rect 16448 2292 16454 2304
rect 16485 2295 16543 2301
rect 16485 2292 16497 2295
rect 16448 2264 16497 2292
rect 16448 2252 16454 2264
rect 16485 2261 16497 2264
rect 16531 2261 16543 2295
rect 17770 2292 17776 2304
rect 17731 2264 17776 2292
rect 16485 2255 16543 2261
rect 17770 2252 17776 2264
rect 17828 2252 17834 2304
rect 18046 2252 18052 2304
rect 18104 2292 18110 2304
rect 18414 2292 18420 2304
rect 18104 2264 18420 2292
rect 18104 2252 18110 2264
rect 18414 2252 18420 2264
rect 18472 2252 18478 2304
rect 184 2202 18924 2224
rect 184 2150 3110 2202
rect 3162 2150 3174 2202
rect 3226 2150 3238 2202
rect 3290 2150 3302 2202
rect 3354 2150 3366 2202
rect 3418 2150 6210 2202
rect 6262 2150 6274 2202
rect 6326 2150 6338 2202
rect 6390 2150 6402 2202
rect 6454 2150 6466 2202
rect 6518 2150 9310 2202
rect 9362 2150 9374 2202
rect 9426 2150 9438 2202
rect 9490 2150 9502 2202
rect 9554 2150 9566 2202
rect 9618 2150 12410 2202
rect 12462 2150 12474 2202
rect 12526 2150 12538 2202
rect 12590 2150 12602 2202
rect 12654 2150 12666 2202
rect 12718 2150 15510 2202
rect 15562 2150 15574 2202
rect 15626 2150 15638 2202
rect 15690 2150 15702 2202
rect 15754 2150 15766 2202
rect 15818 2150 18610 2202
rect 18662 2150 18674 2202
rect 18726 2150 18738 2202
rect 18790 2150 18802 2202
rect 18854 2150 18866 2202
rect 18918 2150 18924 2202
rect 184 2128 18924 2150
rect 4522 2048 4528 2100
rect 4580 2088 4586 2100
rect 4617 2091 4675 2097
rect 4617 2088 4629 2091
rect 4580 2060 4629 2088
rect 4580 2048 4586 2060
rect 4617 2057 4629 2060
rect 4663 2057 4675 2091
rect 4617 2051 4675 2057
rect 5997 2091 6055 2097
rect 5997 2057 6009 2091
rect 6043 2088 6055 2091
rect 7190 2088 7196 2100
rect 6043 2060 7196 2088
rect 6043 2057 6055 2060
rect 5997 2051 6055 2057
rect 7190 2048 7196 2060
rect 7248 2048 7254 2100
rect 7285 2091 7343 2097
rect 7285 2057 7297 2091
rect 7331 2088 7343 2091
rect 7650 2088 7656 2100
rect 7331 2060 7656 2088
rect 7331 2057 7343 2060
rect 7285 2051 7343 2057
rect 7650 2048 7656 2060
rect 7708 2048 7714 2100
rect 8202 2048 8208 2100
rect 8260 2088 8266 2100
rect 8297 2091 8355 2097
rect 8297 2088 8309 2091
rect 8260 2060 8309 2088
rect 8260 2048 8266 2060
rect 8297 2057 8309 2060
rect 8343 2057 8355 2091
rect 9214 2088 9220 2100
rect 8297 2051 8355 2057
rect 9048 2060 9220 2088
rect 5442 2020 5448 2032
rect 4264 1992 5448 2020
rect 2498 1844 2504 1896
rect 2556 1884 2562 1896
rect 4264 1893 4292 1992
rect 5442 1980 5448 1992
rect 5500 1980 5506 2032
rect 6086 1980 6092 2032
rect 6144 2020 6150 2032
rect 6144 1992 6500 2020
rect 6144 1980 6150 1992
rect 6472 1961 6500 1992
rect 6546 1980 6552 2032
rect 6604 2020 6610 2032
rect 9048 2020 9076 2060
rect 9214 2048 9220 2060
rect 9272 2048 9278 2100
rect 9401 2091 9459 2097
rect 9401 2057 9413 2091
rect 9447 2088 9459 2091
rect 9674 2088 9680 2100
rect 9447 2060 9680 2088
rect 9447 2057 9459 2060
rect 9401 2051 9459 2057
rect 9674 2048 9680 2060
rect 9732 2048 9738 2100
rect 9769 2091 9827 2097
rect 9769 2057 9781 2091
rect 9815 2088 9827 2091
rect 9858 2088 9864 2100
rect 9815 2060 9864 2088
rect 9815 2057 9827 2060
rect 9769 2051 9827 2057
rect 9858 2048 9864 2060
rect 9916 2048 9922 2100
rect 10781 2091 10839 2097
rect 10781 2088 10793 2091
rect 10152 2060 10793 2088
rect 6604 1992 9076 2020
rect 6604 1980 6610 1992
rect 5813 1955 5871 1961
rect 5813 1952 5825 1955
rect 4632 1924 5825 1952
rect 3053 1887 3111 1893
rect 3053 1884 3065 1887
rect 2556 1856 3065 1884
rect 2556 1844 2562 1856
rect 3053 1853 3065 1856
rect 3099 1853 3111 1887
rect 3053 1847 3111 1853
rect 4249 1887 4307 1893
rect 4249 1853 4261 1887
rect 4295 1853 4307 1887
rect 4249 1847 4307 1853
rect 4341 1887 4399 1893
rect 4341 1853 4353 1887
rect 4387 1853 4399 1887
rect 4341 1847 4399 1853
rect 2958 1816 2964 1828
rect 2919 1788 2964 1816
rect 2958 1776 2964 1788
rect 3016 1776 3022 1828
rect 4356 1816 4384 1847
rect 4430 1844 4436 1896
rect 4488 1884 4494 1896
rect 4488 1856 4533 1884
rect 4488 1844 4494 1856
rect 4522 1816 4528 1828
rect 4356 1788 4528 1816
rect 4522 1776 4528 1788
rect 4580 1776 4586 1828
rect 4065 1751 4123 1757
rect 4065 1717 4077 1751
rect 4111 1748 4123 1751
rect 4632 1748 4660 1924
rect 5813 1921 5825 1924
rect 5859 1921 5871 1955
rect 6273 1955 6331 1961
rect 6273 1952 6285 1955
rect 5813 1915 5871 1921
rect 5920 1924 6285 1952
rect 4798 1884 4804 1896
rect 4759 1856 4804 1884
rect 4798 1844 4804 1856
rect 4856 1844 4862 1896
rect 4982 1884 4988 1896
rect 4943 1856 4988 1884
rect 4982 1844 4988 1856
rect 5040 1844 5046 1896
rect 5077 1887 5135 1893
rect 5077 1853 5089 1887
rect 5123 1853 5135 1887
rect 5258 1884 5264 1896
rect 5219 1856 5264 1884
rect 5077 1847 5135 1853
rect 4111 1720 4660 1748
rect 5092 1748 5120 1847
rect 5258 1844 5264 1856
rect 5316 1844 5322 1896
rect 5718 1884 5724 1896
rect 5631 1856 5724 1884
rect 5718 1844 5724 1856
rect 5776 1884 5782 1896
rect 5920 1884 5948 1924
rect 6273 1921 6285 1924
rect 6319 1921 6331 1955
rect 6273 1915 6331 1921
rect 6457 1955 6515 1961
rect 6457 1921 6469 1955
rect 6503 1921 6515 1955
rect 6730 1952 6736 1964
rect 6691 1924 6736 1952
rect 6457 1915 6515 1921
rect 6730 1912 6736 1924
rect 6788 1912 6794 1964
rect 7006 1912 7012 1964
rect 7064 1952 7070 1964
rect 7101 1955 7159 1961
rect 7101 1952 7113 1955
rect 7064 1924 7113 1952
rect 7064 1912 7070 1924
rect 7101 1921 7113 1924
rect 7147 1952 7159 1955
rect 7561 1955 7619 1961
rect 7561 1952 7573 1955
rect 7147 1924 7573 1952
rect 7147 1921 7159 1924
rect 7101 1915 7159 1921
rect 7561 1921 7573 1924
rect 7607 1952 7619 1955
rect 7607 1924 8892 1952
rect 7607 1921 7619 1924
rect 7561 1915 7619 1921
rect 8864 1896 8892 1924
rect 5776 1856 5948 1884
rect 6089 1887 6147 1893
rect 5776 1844 5782 1856
rect 6089 1853 6101 1887
rect 6135 1853 6147 1887
rect 6089 1847 6147 1853
rect 5166 1776 5172 1828
rect 5224 1816 5230 1828
rect 6104 1816 6132 1847
rect 7650 1844 7656 1896
rect 7708 1884 7714 1896
rect 7745 1887 7803 1893
rect 7745 1884 7757 1887
rect 7708 1856 7757 1884
rect 7708 1844 7714 1856
rect 7745 1853 7757 1856
rect 7791 1853 7803 1887
rect 7745 1847 7803 1853
rect 8205 1881 8263 1887
rect 8846 1884 8852 1896
rect 8205 1847 8217 1881
rect 8251 1847 8263 1881
rect 8807 1856 8852 1884
rect 8205 1841 8263 1847
rect 8846 1844 8852 1856
rect 8904 1844 8910 1896
rect 9048 1893 9076 1992
rect 9582 1980 9588 2032
rect 9640 2020 9646 2032
rect 9640 1980 9674 2020
rect 9305 1960 9363 1961
rect 9232 1955 9363 1960
rect 9232 1952 9317 1955
rect 9140 1932 9317 1952
rect 9140 1924 9260 1932
rect 8941 1887 8999 1893
rect 8941 1853 8953 1887
rect 8987 1853 8999 1887
rect 8941 1847 8999 1853
rect 9029 1887 9087 1893
rect 9029 1853 9041 1887
rect 9075 1853 9087 1887
rect 9140 1884 9168 1924
rect 9305 1921 9317 1932
rect 9351 1921 9363 1955
rect 9646 1952 9674 1980
rect 10042 1952 10048 1964
rect 9646 1924 10048 1952
rect 9305 1915 9363 1921
rect 10042 1912 10048 1924
rect 10100 1912 10106 1964
rect 9217 1887 9275 1893
rect 9217 1884 9229 1887
rect 9140 1856 9229 1884
rect 9029 1847 9087 1853
rect 9217 1853 9229 1856
rect 9263 1853 9275 1887
rect 9217 1847 9275 1853
rect 5224 1788 6132 1816
rect 5224 1776 5230 1788
rect 5534 1748 5540 1760
rect 5092 1720 5540 1748
rect 4111 1717 4123 1720
rect 4065 1711 4123 1717
rect 5534 1708 5540 1720
rect 5592 1708 5598 1760
rect 5810 1748 5816 1760
rect 5771 1720 5816 1748
rect 5810 1708 5816 1720
rect 5868 1708 5874 1760
rect 7101 1751 7159 1757
rect 7101 1717 7113 1751
rect 7147 1748 7159 1751
rect 7190 1748 7196 1760
rect 7147 1720 7196 1748
rect 7147 1717 7159 1720
rect 7101 1711 7159 1717
rect 7190 1708 7196 1720
rect 7248 1708 7254 1760
rect 7466 1708 7472 1760
rect 7524 1748 7530 1760
rect 7653 1751 7711 1757
rect 7653 1748 7665 1751
rect 7524 1720 7665 1748
rect 7524 1708 7530 1720
rect 7653 1717 7665 1720
rect 7699 1717 7711 1751
rect 7653 1711 7711 1717
rect 8113 1751 8171 1757
rect 8113 1717 8125 1751
rect 8159 1748 8171 1751
rect 8220 1748 8248 1841
rect 8956 1816 8984 1847
rect 9398 1844 9404 1896
rect 9456 1884 9462 1896
rect 9493 1887 9551 1893
rect 9493 1884 9505 1887
rect 9456 1856 9505 1884
rect 9456 1844 9462 1856
rect 9493 1853 9505 1856
rect 9539 1853 9551 1887
rect 9493 1847 9551 1853
rect 9585 1887 9643 1893
rect 9585 1853 9597 1887
rect 9631 1884 9643 1887
rect 10152 1884 10180 2060
rect 10781 2057 10793 2060
rect 10827 2057 10839 2091
rect 12250 2088 12256 2100
rect 12211 2060 12256 2088
rect 10781 2051 10839 2057
rect 12250 2048 12256 2060
rect 12308 2048 12314 2100
rect 12621 2091 12679 2097
rect 12621 2057 12633 2091
rect 12667 2088 12679 2091
rect 16022 2088 16028 2100
rect 12667 2060 16028 2088
rect 12667 2057 12679 2060
rect 12621 2051 12679 2057
rect 16022 2048 16028 2060
rect 16080 2048 16086 2100
rect 16298 2048 16304 2100
rect 16356 2088 16362 2100
rect 16761 2091 16819 2097
rect 16761 2088 16773 2091
rect 16356 2060 16773 2088
rect 16356 2048 16362 2060
rect 16761 2057 16773 2060
rect 16807 2057 16819 2091
rect 16761 2051 16819 2057
rect 16853 2091 16911 2097
rect 16853 2057 16865 2091
rect 16899 2057 16911 2091
rect 17034 2088 17040 2100
rect 16995 2060 17040 2088
rect 16853 2051 16911 2057
rect 10597 2023 10655 2029
rect 10597 1989 10609 2023
rect 10643 1989 10655 2023
rect 10597 1983 10655 1989
rect 9631 1856 10180 1884
rect 10612 1884 10640 1983
rect 15838 1980 15844 2032
rect 15896 2020 15902 2032
rect 16316 2020 16344 2048
rect 15896 1992 16344 2020
rect 16868 2020 16896 2051
rect 17034 2048 17040 2060
rect 17092 2048 17098 2100
rect 18506 2088 18512 2100
rect 17604 2060 18092 2088
rect 18467 2060 18512 2088
rect 17604 2020 17632 2060
rect 17957 2023 18015 2029
rect 17957 2020 17969 2023
rect 16868 1992 17632 2020
rect 17789 1992 17969 2020
rect 15896 1980 15902 1992
rect 10778 1912 10784 1964
rect 10836 1952 10842 1964
rect 11609 1955 11667 1961
rect 11609 1952 11621 1955
rect 10836 1924 11621 1952
rect 10836 1912 10842 1924
rect 11609 1921 11621 1924
rect 11655 1921 11667 1955
rect 11609 1915 11667 1921
rect 12023 1955 12081 1961
rect 12023 1921 12035 1955
rect 12069 1952 12081 1955
rect 13265 1955 13323 1961
rect 13265 1952 13277 1955
rect 12069 1924 13277 1952
rect 12069 1921 12081 1924
rect 12023 1915 12081 1921
rect 13265 1921 13277 1924
rect 13311 1952 13323 1955
rect 13722 1952 13728 1964
rect 13311 1924 13728 1952
rect 13311 1921 13323 1924
rect 13265 1915 13323 1921
rect 13722 1912 13728 1924
rect 13780 1912 13786 1964
rect 13814 1912 13820 1964
rect 13872 1952 13878 1964
rect 13909 1955 13967 1961
rect 13909 1952 13921 1955
rect 13872 1924 13921 1952
rect 13872 1912 13878 1924
rect 13909 1921 13921 1924
rect 13955 1921 13967 1955
rect 13909 1915 13967 1921
rect 14093 1955 14151 1961
rect 14093 1921 14105 1955
rect 14139 1921 14151 1955
rect 14274 1952 14280 1964
rect 14235 1924 14280 1952
rect 14093 1915 14151 1921
rect 10689 1887 10747 1893
rect 10689 1884 10701 1887
rect 10612 1856 10701 1884
rect 9631 1853 9643 1856
rect 9585 1847 9643 1853
rect 10689 1853 10701 1856
rect 10735 1853 10747 1887
rect 11882 1884 11888 1896
rect 11843 1856 11888 1884
rect 10689 1847 10747 1853
rect 11882 1844 11888 1856
rect 11940 1844 11946 1896
rect 12158 1884 12164 1896
rect 12119 1856 12164 1884
rect 12158 1844 12164 1856
rect 12216 1844 12222 1896
rect 12342 1884 12348 1896
rect 12303 1856 12348 1884
rect 12342 1844 12348 1856
rect 12400 1844 12406 1896
rect 12802 1884 12808 1896
rect 12763 1856 12808 1884
rect 12802 1844 12808 1856
rect 12860 1844 12866 1896
rect 12986 1844 12992 1896
rect 13044 1884 13050 1896
rect 14108 1884 14136 1915
rect 14274 1912 14280 1924
rect 14332 1912 14338 1964
rect 16485 1955 16543 1961
rect 16485 1921 16497 1955
rect 16531 1952 16543 1955
rect 16758 1952 16764 1964
rect 16531 1924 16764 1952
rect 16531 1921 16543 1924
rect 16485 1915 16543 1921
rect 16758 1912 16764 1924
rect 16816 1912 16822 1964
rect 16850 1912 16856 1964
rect 16908 1941 16914 1964
rect 16945 1955 17003 1961
rect 16945 1941 16957 1955
rect 16908 1921 16957 1941
rect 16991 1921 17003 1955
rect 16908 1915 17003 1921
rect 16908 1913 16988 1915
rect 16908 1912 16914 1913
rect 17034 1912 17040 1964
rect 17092 1952 17098 1964
rect 17586 1952 17592 1964
rect 17092 1924 17448 1952
rect 17547 1924 17592 1952
rect 17092 1912 17098 1924
rect 14826 1884 14832 1896
rect 13044 1856 14044 1884
rect 14108 1856 14832 1884
rect 13044 1844 13050 1856
rect 9766 1816 9772 1828
rect 8956 1788 9772 1816
rect 9766 1776 9772 1788
rect 9824 1776 9830 1828
rect 10137 1819 10195 1825
rect 10137 1785 10149 1819
rect 10183 1816 10195 1819
rect 11517 1819 11575 1825
rect 11517 1816 11529 1819
rect 10183 1788 11529 1816
rect 10183 1785 10195 1788
rect 10137 1779 10195 1785
rect 11517 1785 11529 1788
rect 11563 1816 11575 1819
rect 13004 1816 13032 1844
rect 11563 1788 13032 1816
rect 11563 1785 11575 1788
rect 11517 1779 11575 1785
rect 8159 1720 8248 1748
rect 8159 1717 8171 1720
rect 8113 1711 8171 1717
rect 9030 1708 9036 1760
rect 9088 1748 9094 1760
rect 10152 1748 10180 1779
rect 13538 1776 13544 1828
rect 13596 1816 13602 1828
rect 13906 1816 13912 1828
rect 13596 1788 13912 1816
rect 13596 1776 13602 1788
rect 13906 1776 13912 1788
rect 13964 1776 13970 1828
rect 14016 1816 14044 1856
rect 14826 1844 14832 1856
rect 14884 1844 14890 1896
rect 16669 1887 16727 1893
rect 16669 1884 16681 1887
rect 14935 1856 16681 1884
rect 14544 1819 14602 1825
rect 14544 1816 14556 1819
rect 14016 1788 14556 1816
rect 14544 1785 14556 1788
rect 14590 1785 14602 1819
rect 14544 1779 14602 1785
rect 9088 1720 10180 1748
rect 10229 1751 10287 1757
rect 9088 1708 9094 1720
rect 10229 1717 10241 1751
rect 10275 1748 10287 1751
rect 11057 1751 11115 1757
rect 11057 1748 11069 1751
rect 10275 1720 11069 1748
rect 10275 1717 10287 1720
rect 10229 1711 10287 1717
rect 11057 1717 11069 1720
rect 11103 1717 11115 1751
rect 11422 1748 11428 1760
rect 11383 1720 11428 1748
rect 11057 1711 11115 1717
rect 11422 1708 11428 1720
rect 11480 1708 11486 1760
rect 13170 1708 13176 1760
rect 13228 1748 13234 1760
rect 13449 1751 13507 1757
rect 13449 1748 13461 1751
rect 13228 1720 13461 1748
rect 13228 1708 13234 1720
rect 13449 1717 13461 1720
rect 13495 1717 13507 1751
rect 13814 1748 13820 1760
rect 13775 1720 13820 1748
rect 13449 1711 13507 1717
rect 13814 1708 13820 1720
rect 13872 1708 13878 1760
rect 14559 1748 14587 1779
rect 14642 1776 14648 1828
rect 14700 1816 14706 1828
rect 14935 1816 14963 1856
rect 16669 1853 16681 1856
rect 16715 1884 16727 1887
rect 17126 1884 17132 1896
rect 16715 1856 17132 1884
rect 16715 1853 16727 1856
rect 16669 1847 16727 1853
rect 17126 1844 17132 1856
rect 17184 1844 17190 1896
rect 17420 1884 17448 1924
rect 17586 1912 17592 1924
rect 17644 1912 17650 1964
rect 17497 1887 17555 1893
rect 17497 1884 17509 1887
rect 17328 1856 17509 1884
rect 14700 1788 14963 1816
rect 14700 1776 14706 1788
rect 15470 1776 15476 1828
rect 15528 1816 15534 1828
rect 16298 1816 16304 1828
rect 15528 1788 16304 1816
rect 15528 1776 15534 1788
rect 16298 1776 16304 1788
rect 16356 1776 16362 1828
rect 16850 1776 16856 1828
rect 16908 1816 16914 1828
rect 17218 1816 17224 1828
rect 16908 1788 17224 1816
rect 16908 1776 16914 1788
rect 17218 1776 17224 1788
rect 17276 1776 17282 1828
rect 14734 1748 14740 1760
rect 14559 1720 14740 1748
rect 14734 1708 14740 1720
rect 14792 1708 14798 1760
rect 15654 1748 15660 1760
rect 15615 1720 15660 1748
rect 15654 1708 15660 1720
rect 15712 1708 15718 1760
rect 15838 1748 15844 1760
rect 15799 1720 15844 1748
rect 15838 1708 15844 1720
rect 15896 1708 15902 1760
rect 16206 1748 16212 1760
rect 16167 1720 16212 1748
rect 16206 1708 16212 1720
rect 16264 1708 16270 1760
rect 17328 1748 17356 1856
rect 17497 1853 17509 1856
rect 17543 1853 17555 1887
rect 17497 1847 17555 1853
rect 17405 1819 17463 1825
rect 17405 1785 17417 1819
rect 17451 1816 17463 1819
rect 17789 1816 17817 1992
rect 17957 1989 17969 1992
rect 18003 1989 18015 2023
rect 17957 1983 18015 1989
rect 17862 1844 17868 1896
rect 17920 1884 17926 1896
rect 18064 1893 18092 2060
rect 18506 2048 18512 2060
rect 18564 2048 18570 2100
rect 18049 1887 18107 1893
rect 17920 1856 17965 1884
rect 17920 1844 17926 1856
rect 18049 1853 18061 1887
rect 18095 1853 18107 1887
rect 18049 1847 18107 1853
rect 18325 1887 18383 1893
rect 18325 1853 18337 1887
rect 18371 1853 18383 1887
rect 18506 1884 18512 1896
rect 18467 1856 18512 1884
rect 18325 1847 18383 1853
rect 18340 1816 18368 1847
rect 18506 1844 18512 1856
rect 18564 1844 18570 1896
rect 17451 1788 17817 1816
rect 17880 1788 18368 1816
rect 17451 1785 17463 1788
rect 17405 1779 17463 1785
rect 17880 1748 17908 1788
rect 17328 1720 17908 1748
rect 184 1658 18860 1680
rect 184 1606 4660 1658
rect 4712 1606 4724 1658
rect 4776 1606 4788 1658
rect 4840 1606 4852 1658
rect 4904 1606 4916 1658
rect 4968 1606 7760 1658
rect 7812 1606 7824 1658
rect 7876 1606 7888 1658
rect 7940 1606 7952 1658
rect 8004 1606 8016 1658
rect 8068 1606 10860 1658
rect 10912 1606 10924 1658
rect 10976 1606 10988 1658
rect 11040 1606 11052 1658
rect 11104 1606 11116 1658
rect 11168 1606 13960 1658
rect 14012 1606 14024 1658
rect 14076 1606 14088 1658
rect 14140 1606 14152 1658
rect 14204 1606 14216 1658
rect 14268 1606 17060 1658
rect 17112 1606 17124 1658
rect 17176 1606 17188 1658
rect 17240 1606 17252 1658
rect 17304 1606 17316 1658
rect 17368 1606 18860 1658
rect 184 1584 18860 1606
rect 3510 1504 3516 1556
rect 3568 1504 3574 1556
rect 4522 1504 4528 1556
rect 4580 1544 4586 1556
rect 4663 1547 4721 1553
rect 4663 1544 4675 1547
rect 4580 1516 4675 1544
rect 4580 1504 4586 1516
rect 4663 1513 4675 1516
rect 4709 1544 4721 1547
rect 5166 1544 5172 1556
rect 4709 1516 5028 1544
rect 5127 1516 5172 1544
rect 4709 1513 4721 1516
rect 4663 1507 4721 1513
rect 3528 1476 3556 1504
rect 5000 1476 5028 1516
rect 5166 1504 5172 1516
rect 5224 1504 5230 1556
rect 5994 1504 6000 1556
rect 6052 1544 6058 1556
rect 6181 1547 6239 1553
rect 6181 1544 6193 1547
rect 6052 1516 6193 1544
rect 6052 1504 6058 1516
rect 6181 1513 6193 1516
rect 6227 1513 6239 1547
rect 6181 1507 6239 1513
rect 7469 1547 7527 1553
rect 7469 1513 7481 1547
rect 7515 1544 7527 1547
rect 7558 1544 7564 1556
rect 7515 1516 7564 1544
rect 7515 1513 7527 1516
rect 7469 1507 7527 1513
rect 7558 1504 7564 1516
rect 7616 1504 7622 1556
rect 7650 1504 7656 1556
rect 7708 1544 7714 1556
rect 7929 1547 7987 1553
rect 7929 1544 7941 1547
rect 7708 1516 7941 1544
rect 7708 1504 7714 1516
rect 7929 1513 7941 1516
rect 7975 1513 7987 1547
rect 7929 1507 7987 1513
rect 8294 1504 8300 1556
rect 8352 1544 8358 1556
rect 8757 1547 8815 1553
rect 8757 1544 8769 1547
rect 8352 1516 8769 1544
rect 8352 1504 8358 1516
rect 8757 1513 8769 1516
rect 8803 1513 8815 1547
rect 9858 1544 9864 1556
rect 8757 1507 8815 1513
rect 9416 1516 9864 1544
rect 7006 1476 7012 1488
rect 3528 1448 3634 1476
rect 5000 1448 7012 1476
rect 7006 1436 7012 1448
rect 7064 1476 7070 1488
rect 9416 1476 9444 1516
rect 9858 1504 9864 1516
rect 9916 1504 9922 1556
rect 10413 1547 10471 1553
rect 10413 1513 10425 1547
rect 10459 1544 10471 1547
rect 10778 1544 10784 1556
rect 10459 1516 10784 1544
rect 10459 1513 10471 1516
rect 10413 1507 10471 1513
rect 10428 1476 10456 1507
rect 10778 1504 10784 1516
rect 10836 1504 10842 1556
rect 11422 1544 11428 1556
rect 11383 1516 11428 1544
rect 11422 1504 11428 1516
rect 11480 1504 11486 1556
rect 11974 1544 11980 1556
rect 11935 1516 11980 1544
rect 11974 1504 11980 1516
rect 12032 1504 12038 1556
rect 12342 1504 12348 1556
rect 12400 1544 12406 1556
rect 12529 1547 12587 1553
rect 12529 1544 12541 1547
rect 12400 1516 12541 1544
rect 12400 1504 12406 1516
rect 12529 1513 12541 1516
rect 12575 1513 12587 1547
rect 12529 1507 12587 1513
rect 12897 1547 12955 1553
rect 12897 1513 12909 1547
rect 12943 1513 12955 1547
rect 13722 1544 13728 1556
rect 13683 1516 13728 1544
rect 12897 1507 12955 1513
rect 7064 1448 9444 1476
rect 7064 1436 7070 1448
rect 2869 1411 2927 1417
rect 2869 1377 2881 1411
rect 2915 1408 2927 1411
rect 2958 1408 2964 1420
rect 2915 1380 2964 1408
rect 2915 1377 2927 1380
rect 2869 1371 2927 1377
rect 2958 1368 2964 1380
rect 3016 1368 3022 1420
rect 5261 1411 5319 1417
rect 5261 1377 5273 1411
rect 5307 1408 5319 1411
rect 6086 1408 6092 1420
rect 5307 1380 5948 1408
rect 6047 1380 6092 1408
rect 5307 1377 5319 1380
rect 5261 1371 5319 1377
rect 3237 1343 3295 1349
rect 3237 1309 3249 1343
rect 3283 1340 3295 1343
rect 5810 1340 5816 1352
rect 3283 1312 5816 1340
rect 3283 1309 3295 1312
rect 3237 1303 3295 1309
rect 5810 1300 5816 1312
rect 5868 1300 5874 1352
rect 5721 1275 5779 1281
rect 5721 1241 5733 1275
rect 5767 1272 5779 1275
rect 5920 1272 5948 1380
rect 6086 1368 6092 1380
rect 6144 1368 6150 1420
rect 7745 1411 7803 1417
rect 7745 1377 7757 1411
rect 7791 1408 7803 1411
rect 8202 1408 8208 1420
rect 7791 1380 8208 1408
rect 7791 1377 7803 1380
rect 7745 1371 7803 1377
rect 8202 1368 8208 1380
rect 8260 1368 8266 1420
rect 8294 1368 8300 1420
rect 8352 1408 8358 1420
rect 9416 1417 9444 1448
rect 9646 1448 10456 1476
rect 9401 1411 9459 1417
rect 8352 1380 8397 1408
rect 8352 1368 8358 1380
rect 9401 1377 9413 1411
rect 9447 1377 9459 1411
rect 9646 1408 9674 1448
rect 10502 1436 10508 1488
rect 10560 1476 10566 1488
rect 11149 1479 11207 1485
rect 11149 1476 11161 1479
rect 10560 1448 11161 1476
rect 10560 1436 10566 1448
rect 11149 1445 11161 1448
rect 11195 1476 11207 1479
rect 12912 1476 12940 1507
rect 13722 1504 13728 1516
rect 13780 1504 13786 1556
rect 13814 1504 13820 1556
rect 13872 1544 13878 1556
rect 14093 1547 14151 1553
rect 14093 1544 14105 1547
rect 13872 1516 14105 1544
rect 13872 1504 13878 1516
rect 14093 1513 14105 1516
rect 14139 1513 14151 1547
rect 14458 1544 14464 1556
rect 14419 1516 14464 1544
rect 14093 1507 14151 1513
rect 14458 1504 14464 1516
rect 14516 1504 14522 1556
rect 14734 1504 14740 1556
rect 14792 1544 14798 1556
rect 16022 1544 16028 1556
rect 14792 1516 16028 1544
rect 14792 1504 14798 1516
rect 16022 1504 16028 1516
rect 16080 1504 16086 1556
rect 16301 1547 16359 1553
rect 16301 1513 16313 1547
rect 16347 1544 16359 1547
rect 16574 1544 16580 1556
rect 16347 1516 16580 1544
rect 16347 1513 16359 1516
rect 16301 1507 16359 1513
rect 16574 1504 16580 1516
rect 16632 1504 16638 1556
rect 17862 1544 17868 1556
rect 17308 1516 17868 1544
rect 16761 1479 16819 1485
rect 11195 1448 11928 1476
rect 12912 1448 16436 1476
rect 11195 1445 11207 1448
rect 11149 1439 11207 1445
rect 11900 1420 11928 1448
rect 9858 1408 9864 1420
rect 9401 1371 9459 1377
rect 9508 1380 9674 1408
rect 9819 1380 9864 1408
rect 6365 1343 6423 1349
rect 6365 1309 6377 1343
rect 6411 1340 6423 1343
rect 6914 1340 6920 1352
rect 6411 1312 6920 1340
rect 6411 1309 6423 1312
rect 6365 1303 6423 1309
rect 6914 1300 6920 1312
rect 6972 1300 6978 1352
rect 7098 1300 7104 1352
rect 7156 1340 7162 1352
rect 7469 1343 7527 1349
rect 7469 1340 7481 1343
rect 7156 1312 7481 1340
rect 7156 1300 7162 1312
rect 7469 1309 7481 1312
rect 7515 1309 7527 1343
rect 8386 1340 8392 1352
rect 8347 1312 8392 1340
rect 7469 1303 7527 1309
rect 8386 1300 8392 1312
rect 8444 1300 8450 1352
rect 8478 1300 8484 1352
rect 8536 1340 8542 1352
rect 9508 1340 9536 1380
rect 9858 1368 9864 1380
rect 9916 1368 9922 1420
rect 10137 1411 10195 1417
rect 10137 1377 10149 1411
rect 10183 1377 10195 1411
rect 10137 1371 10195 1377
rect 8536 1312 9536 1340
rect 9677 1343 9735 1349
rect 8536 1300 8542 1312
rect 9677 1309 9689 1343
rect 9723 1340 9735 1343
rect 9766 1340 9772 1352
rect 9723 1312 9772 1340
rect 9723 1309 9735 1312
rect 9677 1303 9735 1309
rect 9766 1300 9772 1312
rect 9824 1340 9830 1352
rect 10152 1340 10180 1371
rect 10226 1368 10232 1420
rect 10284 1408 10290 1420
rect 10689 1411 10747 1417
rect 10689 1408 10701 1411
rect 10284 1380 10701 1408
rect 10284 1368 10290 1380
rect 10689 1377 10701 1380
rect 10735 1377 10747 1411
rect 10689 1371 10747 1377
rect 11333 1411 11391 1417
rect 11333 1377 11345 1411
rect 11379 1377 11391 1411
rect 11514 1408 11520 1420
rect 11475 1380 11520 1408
rect 11333 1371 11391 1377
rect 9824 1312 10180 1340
rect 9824 1300 9830 1312
rect 5767 1244 5948 1272
rect 5767 1241 5779 1244
rect 5721 1235 5779 1241
rect 8754 1232 8760 1284
rect 8812 1272 8818 1284
rect 8938 1272 8944 1284
rect 8812 1244 8944 1272
rect 8812 1232 8818 1244
rect 8938 1232 8944 1244
rect 8996 1272 9002 1284
rect 9493 1275 9551 1281
rect 9493 1272 9505 1275
rect 8996 1244 9505 1272
rect 8996 1232 9002 1244
rect 9493 1241 9505 1244
rect 9539 1241 9551 1275
rect 9493 1235 9551 1241
rect 9585 1275 9643 1281
rect 9585 1241 9597 1275
rect 9631 1272 9643 1275
rect 11348 1272 11376 1371
rect 11514 1368 11520 1380
rect 11572 1368 11578 1420
rect 11882 1368 11888 1420
rect 11940 1408 11946 1420
rect 12253 1411 12311 1417
rect 12253 1408 12265 1411
rect 11940 1380 12265 1408
rect 11940 1368 11946 1380
rect 12253 1377 12265 1380
rect 12299 1408 12311 1411
rect 12802 1408 12808 1420
rect 12299 1380 12808 1408
rect 12299 1377 12311 1380
rect 12253 1371 12311 1377
rect 12802 1368 12808 1380
rect 12860 1368 12866 1420
rect 12894 1368 12900 1420
rect 12952 1408 12958 1420
rect 13173 1411 13231 1417
rect 13173 1408 13185 1411
rect 12952 1380 13185 1408
rect 12952 1368 12958 1380
rect 13173 1377 13185 1380
rect 13219 1377 13231 1411
rect 13173 1371 13231 1377
rect 13265 1411 13323 1417
rect 13265 1377 13277 1411
rect 13311 1408 13323 1411
rect 13354 1408 13360 1420
rect 13311 1380 13360 1408
rect 13311 1377 13323 1380
rect 13265 1371 13323 1377
rect 13354 1368 13360 1380
rect 13412 1368 13418 1420
rect 13630 1408 13636 1420
rect 13591 1380 13636 1408
rect 13630 1368 13636 1380
rect 13688 1368 13694 1420
rect 14918 1408 14924 1420
rect 14292 1380 14596 1408
rect 14879 1380 14924 1408
rect 12529 1343 12587 1349
rect 12529 1309 12541 1343
rect 12575 1340 12587 1343
rect 13078 1340 13084 1352
rect 12575 1312 13084 1340
rect 12575 1309 12587 1312
rect 12529 1303 12587 1309
rect 13078 1300 13084 1312
rect 13136 1300 13142 1352
rect 13449 1343 13507 1349
rect 13449 1309 13461 1343
rect 13495 1309 13507 1343
rect 13449 1303 13507 1309
rect 9631 1244 11376 1272
rect 9631 1241 9643 1244
rect 9585 1235 9643 1241
rect 12158 1232 12164 1284
rect 12216 1272 12222 1284
rect 12345 1275 12403 1281
rect 12345 1272 12357 1275
rect 12216 1244 12357 1272
rect 12216 1232 12222 1244
rect 12345 1241 12357 1244
rect 12391 1272 12403 1275
rect 12986 1272 12992 1284
rect 12391 1244 12992 1272
rect 12391 1241 12403 1244
rect 12345 1235 12403 1241
rect 12986 1232 12992 1244
rect 13044 1232 13050 1284
rect 13464 1272 13492 1303
rect 13814 1300 13820 1352
rect 13872 1340 13878 1352
rect 14292 1340 14320 1380
rect 13872 1312 14320 1340
rect 14568 1340 14596 1380
rect 14918 1368 14924 1380
rect 14976 1368 14982 1420
rect 15188 1411 15246 1417
rect 15188 1377 15200 1411
rect 15234 1408 15246 1411
rect 15470 1408 15476 1420
rect 15234 1380 15476 1408
rect 15234 1377 15246 1380
rect 15188 1371 15246 1377
rect 15470 1368 15476 1380
rect 15528 1368 15534 1420
rect 16408 1408 16436 1448
rect 16761 1445 16773 1479
rect 16807 1476 16819 1479
rect 16942 1476 16948 1488
rect 16807 1448 16948 1476
rect 16807 1445 16819 1448
rect 16761 1439 16819 1445
rect 16942 1436 16948 1448
rect 17000 1436 17006 1488
rect 17308 1408 17336 1516
rect 17862 1504 17868 1516
rect 17920 1504 17926 1556
rect 18049 1547 18107 1553
rect 18049 1513 18061 1547
rect 18095 1544 18107 1547
rect 18138 1544 18144 1556
rect 18095 1516 18144 1544
rect 18095 1513 18107 1516
rect 18049 1507 18107 1513
rect 18138 1504 18144 1516
rect 18196 1504 18202 1556
rect 17402 1436 17408 1488
rect 17460 1476 17466 1488
rect 17681 1479 17739 1485
rect 17681 1476 17693 1479
rect 17460 1448 17693 1476
rect 17460 1436 17466 1448
rect 17681 1445 17693 1448
rect 17727 1445 17739 1479
rect 17681 1439 17739 1445
rect 16408 1380 17336 1408
rect 17770 1368 17776 1420
rect 17828 1408 17834 1420
rect 17865 1411 17923 1417
rect 17865 1408 17877 1411
rect 17828 1380 17877 1408
rect 17828 1368 17834 1380
rect 17865 1377 17877 1380
rect 17911 1377 17923 1411
rect 17865 1371 17923 1377
rect 18046 1368 18052 1420
rect 18104 1408 18110 1420
rect 18141 1411 18199 1417
rect 18141 1408 18153 1411
rect 18104 1380 18153 1408
rect 18104 1368 18110 1380
rect 18141 1377 18153 1380
rect 18187 1377 18199 1411
rect 18325 1411 18383 1417
rect 18325 1408 18337 1411
rect 18141 1371 18199 1377
rect 18248 1380 18337 1408
rect 16390 1340 16396 1352
rect 14568 1312 14964 1340
rect 13872 1300 13878 1312
rect 14182 1272 14188 1284
rect 13464 1244 14188 1272
rect 14182 1232 14188 1244
rect 14240 1232 14246 1284
rect 14277 1275 14335 1281
rect 14277 1241 14289 1275
rect 14323 1272 14335 1275
rect 14550 1272 14556 1284
rect 14323 1244 14556 1272
rect 14323 1241 14335 1244
rect 14277 1235 14335 1241
rect 14550 1232 14556 1244
rect 14608 1232 14614 1284
rect 7190 1164 7196 1216
rect 7248 1204 7254 1216
rect 7653 1207 7711 1213
rect 7653 1204 7665 1207
rect 7248 1176 7665 1204
rect 7248 1164 7254 1176
rect 7653 1173 7665 1176
rect 7699 1204 7711 1207
rect 9398 1204 9404 1216
rect 7699 1176 9404 1204
rect 7699 1173 7711 1176
rect 7653 1167 7711 1173
rect 9398 1164 9404 1176
rect 9456 1164 9462 1216
rect 10042 1164 10048 1216
rect 10100 1204 10106 1216
rect 10873 1207 10931 1213
rect 10873 1204 10885 1207
rect 10100 1176 10885 1204
rect 10100 1164 10106 1176
rect 10873 1173 10885 1176
rect 10919 1173 10931 1207
rect 11882 1204 11888 1216
rect 11843 1176 11888 1204
rect 10873 1167 10931 1173
rect 11882 1164 11888 1176
rect 11940 1164 11946 1216
rect 11974 1164 11980 1216
rect 12032 1204 12038 1216
rect 12805 1207 12863 1213
rect 12805 1204 12817 1207
rect 12032 1176 12817 1204
rect 12032 1164 12038 1176
rect 12805 1173 12817 1176
rect 12851 1204 12863 1207
rect 12894 1204 12900 1216
rect 12851 1176 12900 1204
rect 12851 1173 12863 1176
rect 12805 1167 12863 1173
rect 12894 1164 12900 1176
rect 12952 1164 12958 1216
rect 13262 1204 13268 1216
rect 13223 1176 13268 1204
rect 13262 1164 13268 1176
rect 13320 1164 13326 1216
rect 13446 1164 13452 1216
rect 13504 1204 13510 1216
rect 14737 1207 14795 1213
rect 14737 1204 14749 1207
rect 13504 1176 14749 1204
rect 13504 1164 13510 1176
rect 14737 1173 14749 1176
rect 14783 1173 14795 1207
rect 14936 1204 14964 1312
rect 15948 1312 16396 1340
rect 15948 1204 15976 1312
rect 16390 1300 16396 1312
rect 16448 1340 16454 1352
rect 17037 1343 17095 1349
rect 17037 1340 17049 1343
rect 16448 1312 17049 1340
rect 16448 1300 16454 1312
rect 17037 1309 17049 1312
rect 17083 1309 17095 1343
rect 17402 1340 17408 1352
rect 17363 1312 17408 1340
rect 17037 1303 17095 1309
rect 17402 1300 17408 1312
rect 17460 1300 17466 1352
rect 16022 1232 16028 1284
rect 16080 1272 16086 1284
rect 16485 1275 16543 1281
rect 16485 1272 16497 1275
rect 16080 1244 16497 1272
rect 16080 1232 16086 1244
rect 16485 1241 16497 1244
rect 16531 1272 16543 1275
rect 16850 1272 16856 1284
rect 16531 1244 16856 1272
rect 16531 1241 16543 1244
rect 16485 1235 16543 1241
rect 16850 1232 16856 1244
rect 16908 1232 16914 1284
rect 17310 1272 17316 1284
rect 17052 1244 17316 1272
rect 14936 1176 15976 1204
rect 14737 1167 14795 1173
rect 16758 1164 16764 1216
rect 16816 1204 16822 1216
rect 17052 1204 17080 1244
rect 17310 1232 17316 1244
rect 17368 1272 17374 1284
rect 18248 1272 18276 1380
rect 18325 1377 18337 1380
rect 18371 1377 18383 1411
rect 18325 1371 18383 1377
rect 17368 1244 18276 1272
rect 17368 1232 17374 1244
rect 16816 1176 17080 1204
rect 16816 1164 16822 1176
rect 17126 1164 17132 1216
rect 17184 1204 17190 1216
rect 17494 1204 17500 1216
rect 17184 1176 17500 1204
rect 17184 1164 17190 1176
rect 17494 1164 17500 1176
rect 17552 1204 17558 1216
rect 18417 1207 18475 1213
rect 18417 1204 18429 1207
rect 17552 1176 18429 1204
rect 17552 1164 17558 1176
rect 18417 1173 18429 1176
rect 18463 1173 18475 1207
rect 18417 1167 18475 1173
rect 184 1114 18924 1136
rect 184 1062 3110 1114
rect 3162 1062 3174 1114
rect 3226 1062 3238 1114
rect 3290 1062 3302 1114
rect 3354 1062 3366 1114
rect 3418 1062 6210 1114
rect 6262 1062 6274 1114
rect 6326 1062 6338 1114
rect 6390 1062 6402 1114
rect 6454 1062 6466 1114
rect 6518 1062 9310 1114
rect 9362 1062 9374 1114
rect 9426 1062 9438 1114
rect 9490 1062 9502 1114
rect 9554 1062 9566 1114
rect 9618 1062 12410 1114
rect 12462 1062 12474 1114
rect 12526 1062 12538 1114
rect 12590 1062 12602 1114
rect 12654 1062 12666 1114
rect 12718 1062 15510 1114
rect 15562 1062 15574 1114
rect 15626 1062 15638 1114
rect 15690 1062 15702 1114
rect 15754 1062 15766 1114
rect 15818 1062 18610 1114
rect 18662 1062 18674 1114
rect 18726 1062 18738 1114
rect 18790 1062 18802 1114
rect 18854 1062 18866 1114
rect 18918 1062 18924 1114
rect 184 1040 18924 1062
rect 6086 960 6092 1012
rect 6144 1000 6150 1012
rect 7469 1003 7527 1009
rect 7469 1000 7481 1003
rect 6144 972 7481 1000
rect 6144 960 6150 972
rect 7469 969 7481 972
rect 7515 969 7527 1003
rect 7469 963 7527 969
rect 8294 960 8300 1012
rect 8352 1000 8358 1012
rect 8757 1003 8815 1009
rect 8757 1000 8769 1003
rect 8352 972 8769 1000
rect 8352 960 8358 972
rect 8757 969 8769 972
rect 8803 969 8815 1003
rect 8757 963 8815 969
rect 8938 960 8944 1012
rect 8996 1000 9002 1012
rect 9861 1003 9919 1009
rect 9861 1000 9873 1003
rect 8996 972 9873 1000
rect 8996 960 9002 972
rect 9861 969 9873 972
rect 9907 1000 9919 1003
rect 10134 1000 10140 1012
rect 9907 972 10140 1000
rect 9907 969 9919 972
rect 9861 963 9919 969
rect 10134 960 10140 972
rect 10192 960 10198 1012
rect 10229 1003 10287 1009
rect 10229 969 10241 1003
rect 10275 1000 10287 1003
rect 11514 1000 11520 1012
rect 10275 972 11520 1000
rect 10275 969 10287 972
rect 10229 963 10287 969
rect 11514 960 11520 972
rect 11572 960 11578 1012
rect 13538 1000 13544 1012
rect 13499 972 13544 1000
rect 13538 960 13544 972
rect 13596 960 13602 1012
rect 15378 960 15384 1012
rect 15436 1000 15442 1012
rect 15565 1003 15623 1009
rect 15565 1000 15577 1003
rect 15436 972 15577 1000
rect 15436 960 15442 972
rect 15565 969 15577 972
rect 15611 969 15623 1003
rect 15565 963 15623 969
rect 16206 960 16212 1012
rect 16264 1000 16270 1012
rect 16577 1003 16635 1009
rect 16577 1000 16589 1003
rect 16264 972 16589 1000
rect 16264 960 16270 972
rect 16577 969 16589 972
rect 16623 969 16635 1003
rect 17126 1000 17132 1012
rect 17087 972 17132 1000
rect 16577 963 16635 969
rect 17126 960 17132 972
rect 17184 960 17190 1012
rect 17310 960 17316 1012
rect 17368 1000 17374 1012
rect 17405 1003 17463 1009
rect 17405 1000 17417 1003
rect 17368 972 17417 1000
rect 17368 960 17374 972
rect 17405 969 17417 972
rect 17451 969 17463 1003
rect 17405 963 17463 969
rect 18230 960 18236 1012
rect 18288 1000 18294 1012
rect 18325 1003 18383 1009
rect 18325 1000 18337 1003
rect 18288 972 18337 1000
rect 18288 960 18294 972
rect 18325 969 18337 972
rect 18371 969 18383 1003
rect 18325 963 18383 969
rect 5994 892 6000 944
rect 6052 932 6058 944
rect 14090 932 14096 944
rect 6052 904 7972 932
rect 6052 892 6058 904
rect 6638 824 6644 876
rect 6696 864 6702 876
rect 7944 873 7972 904
rect 13556 904 14096 932
rect 6825 867 6883 873
rect 6825 864 6837 867
rect 6696 836 6837 864
rect 6696 824 6702 836
rect 6825 833 6837 836
rect 6871 864 6883 867
rect 7929 867 7987 873
rect 6871 836 7880 864
rect 6871 833 6883 836
rect 6825 827 6883 833
rect 6917 799 6975 805
rect 6917 765 6929 799
rect 6963 796 6975 799
rect 7006 796 7012 808
rect 6963 768 7012 796
rect 6963 765 6975 768
rect 6917 759 6975 765
rect 7006 756 7012 768
rect 7064 756 7070 808
rect 7852 796 7880 836
rect 7929 833 7941 867
rect 7975 833 7987 867
rect 7929 827 7987 833
rect 8113 867 8171 873
rect 8113 833 8125 867
rect 8159 864 8171 867
rect 8478 864 8484 876
rect 8159 836 8484 864
rect 8159 833 8171 836
rect 8113 827 8171 833
rect 8478 824 8484 836
rect 8536 824 8542 876
rect 9950 864 9956 876
rect 9911 836 9956 864
rect 9950 824 9956 836
rect 10008 824 10014 876
rect 12345 867 12403 873
rect 12345 833 12357 867
rect 12391 864 12403 867
rect 13170 864 13176 876
rect 12391 836 13176 864
rect 12391 833 12403 836
rect 12345 827 12403 833
rect 13170 824 13176 836
rect 13228 824 13234 876
rect 13262 824 13268 876
rect 13320 864 13326 876
rect 13320 836 13365 864
rect 13320 824 13326 836
rect 8754 796 8760 808
rect 7852 768 8760 796
rect 8754 756 8760 768
rect 8812 756 8818 808
rect 9766 756 9772 808
rect 9824 796 9830 808
rect 9861 799 9919 805
rect 9861 796 9873 799
rect 9824 768 9873 796
rect 9824 756 9830 768
rect 9861 765 9873 768
rect 9907 765 9919 799
rect 12802 796 12808 808
rect 12763 768 12808 796
rect 9861 759 9919 765
rect 12802 756 12808 768
rect 12860 756 12866 808
rect 12986 756 12992 808
rect 13044 796 13050 808
rect 13556 796 13584 904
rect 14090 892 14096 904
rect 14148 892 14154 944
rect 14185 935 14243 941
rect 14185 901 14197 935
rect 14231 932 14243 935
rect 14274 932 14280 944
rect 14231 904 14280 932
rect 14231 901 14243 904
rect 14185 895 14243 901
rect 14274 892 14280 904
rect 14332 892 14338 944
rect 14366 892 14372 944
rect 14424 932 14430 944
rect 14461 935 14519 941
rect 14461 932 14473 935
rect 14424 904 14473 932
rect 14424 892 14430 904
rect 14461 901 14473 904
rect 14507 901 14519 935
rect 14461 895 14519 901
rect 15473 935 15531 941
rect 15473 901 15485 935
rect 15519 932 15531 935
rect 16482 932 16488 944
rect 15519 904 16488 932
rect 15519 901 15531 904
rect 15473 895 15531 901
rect 16482 892 16488 904
rect 16540 892 16546 944
rect 14292 864 14320 892
rect 14292 836 15240 864
rect 13814 796 13820 808
rect 13044 768 13584 796
rect 13775 768 13820 796
rect 13044 756 13050 768
rect 13814 756 13820 768
rect 13872 756 13878 808
rect 14001 799 14059 805
rect 14001 765 14013 799
rect 14047 765 14059 799
rect 14274 796 14280 808
rect 14187 768 14280 796
rect 14001 759 14059 765
rect 7837 731 7895 737
rect 7837 728 7849 731
rect 7300 700 7849 728
rect 7300 669 7328 700
rect 7837 697 7849 700
rect 7883 697 7895 731
rect 14016 728 14044 759
rect 14274 756 14280 768
rect 14332 796 14338 808
rect 14734 796 14740 808
rect 14332 768 14740 796
rect 14332 756 14338 768
rect 14734 756 14740 768
rect 14792 756 14798 808
rect 14829 799 14887 805
rect 14829 765 14841 799
rect 14875 765 14887 799
rect 15010 796 15016 808
rect 14971 768 15016 796
rect 14829 759 14887 765
rect 14844 728 14872 759
rect 15010 756 15016 768
rect 15068 756 15074 808
rect 15212 805 15240 836
rect 16022 824 16028 876
rect 16080 864 16086 876
rect 17586 864 17592 876
rect 16080 836 17592 864
rect 16080 824 16086 836
rect 17586 824 17592 836
rect 17644 824 17650 876
rect 15197 799 15255 805
rect 15197 765 15209 799
rect 15243 765 15255 799
rect 17678 796 17684 808
rect 17639 768 17684 796
rect 15197 759 15255 765
rect 17678 756 17684 768
rect 17736 756 17742 808
rect 17862 756 17868 808
rect 17920 796 17926 808
rect 18506 796 18512 808
rect 17920 768 18013 796
rect 18467 768 18512 796
rect 17920 756 17926 768
rect 18506 756 18512 768
rect 18564 796 18570 808
rect 19058 796 19064 808
rect 18564 768 19064 796
rect 18564 756 18570 768
rect 19058 756 19064 768
rect 19116 756 19122 808
rect 16114 728 16120 740
rect 7837 691 7895 697
rect 13096 700 14044 728
rect 14108 700 14872 728
rect 16075 700 16120 728
rect 7285 663 7343 669
rect 7285 629 7297 663
rect 7331 629 7343 663
rect 12066 660 12072 672
rect 12027 632 12072 660
rect 7285 623 7343 629
rect 12066 620 12072 632
rect 12124 620 12130 672
rect 12526 660 12532 672
rect 12487 632 12532 660
rect 12526 620 12532 632
rect 12584 620 12590 672
rect 12710 660 12716 672
rect 12671 632 12716 660
rect 12710 620 12716 632
rect 12768 620 12774 672
rect 13096 669 13124 700
rect 13081 663 13139 669
rect 13081 629 13093 663
rect 13127 629 13139 663
rect 13081 623 13139 629
rect 13722 620 13728 672
rect 13780 660 13786 672
rect 14108 660 14136 700
rect 16114 688 16120 700
rect 16172 688 16178 740
rect 16209 731 16267 737
rect 16209 697 16221 731
rect 16255 728 16267 731
rect 16666 728 16672 740
rect 16255 700 16672 728
rect 16255 697 16267 700
rect 16209 691 16267 697
rect 16666 688 16672 700
rect 16724 688 16730 740
rect 16850 688 16856 740
rect 16908 728 16914 740
rect 17402 728 17408 740
rect 16908 700 17408 728
rect 16908 688 16914 700
rect 17402 688 17408 700
rect 17460 688 17466 740
rect 13780 632 14136 660
rect 13780 620 13786 632
rect 14182 620 14188 672
rect 14240 660 14246 672
rect 15197 663 15255 669
rect 15197 660 15209 663
rect 14240 632 15209 660
rect 14240 620 14246 632
rect 15197 629 15209 632
rect 15243 660 15255 663
rect 16022 660 16028 672
rect 15243 632 16028 660
rect 15243 629 15255 632
rect 15197 623 15255 629
rect 16022 620 16028 632
rect 16080 620 16086 672
rect 16482 620 16488 672
rect 16540 660 16546 672
rect 17880 660 17908 756
rect 16540 632 17908 660
rect 18049 663 18107 669
rect 16540 620 16546 632
rect 18049 629 18061 663
rect 18095 660 18107 663
rect 18322 660 18328 672
rect 18095 632 18328 660
rect 18095 629 18107 632
rect 18049 623 18107 629
rect 18322 620 18328 632
rect 18380 620 18386 672
rect 184 570 18860 592
rect 184 518 4660 570
rect 4712 518 4724 570
rect 4776 518 4788 570
rect 4840 518 4852 570
rect 4904 518 4916 570
rect 4968 518 7760 570
rect 7812 518 7824 570
rect 7876 518 7888 570
rect 7940 518 7952 570
rect 8004 518 8016 570
rect 8068 518 10860 570
rect 10912 518 10924 570
rect 10976 518 10988 570
rect 11040 518 11052 570
rect 11104 518 11116 570
rect 11168 518 13960 570
rect 14012 518 14024 570
rect 14076 518 14088 570
rect 14140 518 14152 570
rect 14204 518 14216 570
rect 14268 518 17060 570
rect 17112 518 17124 570
rect 17176 518 17188 570
rect 17240 518 17252 570
rect 17304 518 17316 570
rect 17368 518 18860 570
rect 184 496 18860 518
rect 12526 416 12532 468
rect 12584 456 12590 468
rect 15930 456 15936 468
rect 12584 428 15936 456
rect 12584 416 12590 428
rect 15930 416 15936 428
rect 15988 416 15994 468
rect 11882 348 11888 400
rect 11940 388 11946 400
rect 15286 388 15292 400
rect 11940 360 15292 388
rect 11940 348 11946 360
rect 15286 348 15292 360
rect 15344 348 15350 400
rect 12710 280 12716 332
rect 12768 320 12774 332
rect 15194 320 15200 332
rect 12768 292 15200 320
rect 12768 280 12774 292
rect 15194 280 15200 292
rect 15252 280 15258 332
rect 12894 212 12900 264
rect 12952 252 12958 264
rect 16850 252 16856 264
rect 12952 224 16856 252
rect 12952 212 12958 224
rect 16850 212 16856 224
rect 16908 212 16914 264
rect 13170 144 13176 196
rect 13228 184 13234 196
rect 16482 184 16488 196
rect 13228 156 16488 184
rect 13228 144 13234 156
rect 16482 144 16488 156
rect 16540 144 16546 196
rect 12066 76 12072 128
rect 12124 116 12130 128
rect 18506 116 18512 128
rect 12124 88 18512 116
rect 12124 76 12130 88
rect 18506 76 18512 88
rect 18564 76 18570 128
<< via1 >>
rect 7288 11364 7340 11416
rect 9680 11364 9732 11416
rect 17592 11364 17644 11416
rect 1308 11228 1360 11280
rect 4528 11228 4580 11280
rect 4620 11228 4672 11280
rect 6552 11228 6604 11280
rect 9772 11228 9824 11280
rect 4160 11160 4212 11212
rect 9128 11160 9180 11212
rect 12256 11160 12308 11212
rect 1952 11092 2004 11144
rect 8760 11092 8812 11144
rect 9220 11092 9272 11144
rect 12164 11092 12216 11144
rect 16120 11092 16172 11144
rect 17684 11092 17736 11144
rect 572 11024 624 11076
rect 2872 11024 2924 11076
rect 2964 11024 3016 11076
rect 4988 11024 5040 11076
rect 1860 10956 1912 11008
rect 6920 11024 6972 11076
rect 11888 11024 11940 11076
rect 16580 11024 16632 11076
rect 5264 10956 5316 11008
rect 7656 10956 7708 11008
rect 12072 10956 12124 11008
rect 18236 10956 18288 11008
rect 3110 10854 3162 10906
rect 3174 10854 3226 10906
rect 3238 10854 3290 10906
rect 3302 10854 3354 10906
rect 3366 10854 3418 10906
rect 6210 10854 6262 10906
rect 6274 10854 6326 10906
rect 6338 10854 6390 10906
rect 6402 10854 6454 10906
rect 6466 10854 6518 10906
rect 9310 10854 9362 10906
rect 9374 10854 9426 10906
rect 9438 10854 9490 10906
rect 9502 10854 9554 10906
rect 9566 10854 9618 10906
rect 12410 10854 12462 10906
rect 12474 10854 12526 10906
rect 12538 10854 12590 10906
rect 12602 10854 12654 10906
rect 12666 10854 12718 10906
rect 15510 10854 15562 10906
rect 15574 10854 15626 10906
rect 15638 10854 15690 10906
rect 15702 10854 15754 10906
rect 15766 10854 15818 10906
rect 18610 10854 18662 10906
rect 18674 10854 18726 10906
rect 18738 10854 18790 10906
rect 18802 10854 18854 10906
rect 18866 10854 18918 10906
rect 572 10795 624 10804
rect 572 10761 581 10795
rect 581 10761 615 10795
rect 615 10761 624 10795
rect 572 10752 624 10761
rect 1124 10659 1176 10668
rect 1124 10625 1133 10659
rect 1133 10625 1167 10659
rect 1167 10625 1176 10659
rect 1124 10616 1176 10625
rect 1952 10659 2004 10668
rect 1952 10625 1961 10659
rect 1961 10625 1995 10659
rect 1995 10625 2004 10659
rect 1952 10616 2004 10625
rect 4344 10752 4396 10804
rect 5264 10795 5316 10804
rect 5264 10761 5273 10795
rect 5273 10761 5307 10795
rect 5307 10761 5316 10795
rect 5264 10752 5316 10761
rect 2504 10727 2556 10736
rect 2504 10693 2513 10727
rect 2513 10693 2547 10727
rect 2547 10693 2556 10727
rect 2504 10684 2556 10693
rect 2964 10616 3016 10668
rect 4068 10616 4120 10668
rect 5816 10752 5868 10804
rect 756 10591 808 10600
rect 756 10557 765 10591
rect 765 10557 799 10591
rect 799 10557 808 10591
rect 756 10548 808 10557
rect 1400 10548 1452 10600
rect 1676 10591 1728 10600
rect 1676 10557 1685 10591
rect 1685 10557 1719 10591
rect 1719 10557 1728 10591
rect 1676 10548 1728 10557
rect 2780 10548 2832 10600
rect 4528 10591 4580 10600
rect 480 10480 532 10532
rect 2136 10455 2188 10464
rect 2136 10421 2145 10455
rect 2145 10421 2179 10455
rect 2179 10421 2188 10455
rect 2688 10455 2740 10464
rect 2136 10412 2188 10421
rect 2688 10421 2697 10455
rect 2697 10421 2731 10455
rect 2731 10421 2740 10455
rect 2688 10412 2740 10421
rect 3884 10412 3936 10464
rect 4068 10455 4120 10464
rect 4068 10421 4077 10455
rect 4077 10421 4111 10455
rect 4111 10421 4120 10455
rect 4068 10412 4120 10421
rect 4528 10557 4537 10591
rect 4537 10557 4571 10591
rect 4571 10557 4580 10591
rect 4528 10548 4580 10557
rect 4620 10591 4672 10600
rect 4620 10557 4629 10591
rect 4629 10557 4663 10591
rect 4663 10557 4672 10591
rect 9772 10752 9824 10804
rect 11888 10795 11940 10804
rect 5908 10659 5960 10668
rect 5908 10625 5917 10659
rect 5917 10625 5951 10659
rect 5951 10625 5960 10659
rect 5908 10616 5960 10625
rect 7012 10616 7064 10668
rect 9220 10684 9272 10736
rect 9680 10727 9732 10736
rect 9680 10693 9689 10727
rect 9689 10693 9723 10727
rect 9723 10693 9732 10727
rect 9680 10684 9732 10693
rect 7380 10616 7432 10668
rect 11888 10761 11897 10795
rect 11897 10761 11931 10795
rect 11931 10761 11940 10795
rect 11888 10752 11940 10761
rect 11980 10752 12032 10804
rect 14924 10752 14976 10804
rect 17960 10795 18012 10804
rect 17960 10761 17969 10795
rect 17969 10761 18003 10795
rect 18003 10761 18012 10795
rect 17960 10752 18012 10761
rect 18236 10795 18288 10804
rect 18236 10761 18245 10795
rect 18245 10761 18279 10795
rect 18279 10761 18288 10795
rect 18236 10752 18288 10761
rect 13452 10684 13504 10736
rect 17684 10727 17736 10736
rect 17684 10693 17693 10727
rect 17693 10693 17727 10727
rect 17727 10693 17736 10727
rect 17684 10684 17736 10693
rect 4620 10548 4672 10557
rect 7196 10548 7248 10600
rect 8116 10548 8168 10600
rect 8208 10548 8260 10600
rect 10140 10616 10192 10668
rect 10600 10659 10652 10668
rect 10600 10625 10609 10659
rect 10609 10625 10643 10659
rect 10643 10625 10652 10659
rect 10600 10616 10652 10625
rect 12164 10616 12216 10668
rect 12900 10616 12952 10668
rect 14464 10616 14516 10668
rect 14924 10659 14976 10668
rect 14924 10625 14933 10659
rect 14933 10625 14967 10659
rect 14967 10625 14976 10659
rect 14924 10616 14976 10625
rect 9220 10591 9272 10600
rect 9220 10557 9229 10591
rect 9229 10557 9263 10591
rect 9263 10557 9272 10591
rect 9220 10548 9272 10557
rect 9312 10548 9364 10600
rect 11520 10548 11572 10600
rect 11888 10591 11940 10600
rect 11888 10557 11897 10591
rect 11897 10557 11931 10591
rect 11931 10557 11940 10591
rect 11888 10548 11940 10557
rect 12072 10591 12124 10600
rect 12072 10557 12081 10591
rect 12081 10557 12115 10591
rect 12115 10557 12124 10591
rect 12072 10548 12124 10557
rect 12256 10591 12308 10600
rect 12256 10557 12265 10591
rect 12265 10557 12299 10591
rect 12299 10557 12308 10591
rect 12256 10548 12308 10557
rect 9772 10480 9824 10532
rect 5448 10412 5500 10464
rect 5540 10412 5592 10464
rect 6092 10412 6144 10464
rect 7288 10412 7340 10464
rect 7564 10412 7616 10464
rect 7656 10412 7708 10464
rect 8208 10412 8260 10464
rect 9128 10455 9180 10464
rect 9128 10421 9137 10455
rect 9137 10421 9171 10455
rect 9171 10421 9180 10455
rect 9496 10455 9548 10464
rect 9128 10412 9180 10421
rect 9496 10421 9505 10455
rect 9505 10421 9539 10455
rect 9539 10421 9548 10455
rect 9496 10412 9548 10421
rect 9956 10412 10008 10464
rect 10140 10412 10192 10464
rect 11336 10455 11388 10464
rect 11336 10421 11345 10455
rect 11345 10421 11379 10455
rect 11379 10421 11388 10455
rect 11336 10412 11388 10421
rect 12164 10480 12216 10532
rect 12808 10548 12860 10600
rect 14648 10591 14700 10600
rect 14648 10557 14657 10591
rect 14657 10557 14691 10591
rect 14691 10557 14700 10591
rect 14648 10548 14700 10557
rect 12440 10523 12492 10532
rect 12440 10489 12449 10523
rect 12449 10489 12483 10523
rect 12483 10489 12492 10523
rect 12440 10480 12492 10489
rect 13820 10480 13872 10532
rect 14832 10480 14884 10532
rect 12992 10455 13044 10464
rect 12992 10421 13001 10455
rect 13001 10421 13035 10455
rect 13035 10421 13044 10455
rect 12992 10412 13044 10421
rect 15660 10548 15712 10600
rect 18236 10616 18288 10668
rect 15292 10480 15344 10532
rect 16028 10523 16080 10532
rect 16028 10489 16037 10523
rect 16037 10489 16071 10523
rect 16071 10489 16080 10523
rect 16028 10480 16080 10489
rect 15200 10455 15252 10464
rect 15200 10421 15209 10455
rect 15209 10421 15243 10455
rect 15243 10421 15252 10455
rect 15200 10412 15252 10421
rect 15568 10455 15620 10464
rect 15568 10421 15577 10455
rect 15577 10421 15611 10455
rect 15611 10421 15620 10455
rect 15568 10412 15620 10421
rect 15936 10455 15988 10464
rect 15936 10421 15945 10455
rect 15945 10421 15979 10455
rect 15979 10421 15988 10455
rect 15936 10412 15988 10421
rect 16120 10455 16172 10464
rect 16120 10421 16129 10455
rect 16129 10421 16163 10455
rect 16163 10421 16172 10455
rect 16120 10412 16172 10421
rect 17776 10548 17828 10600
rect 17868 10591 17920 10600
rect 17868 10557 17877 10591
rect 17877 10557 17911 10591
rect 17911 10557 17920 10591
rect 17868 10548 17920 10557
rect 18144 10548 18196 10600
rect 18420 10591 18472 10600
rect 18420 10557 18429 10591
rect 18429 10557 18463 10591
rect 18463 10557 18472 10591
rect 18420 10548 18472 10557
rect 17592 10523 17644 10532
rect 16488 10455 16540 10464
rect 16488 10421 16497 10455
rect 16497 10421 16531 10455
rect 16531 10421 16540 10455
rect 16488 10412 16540 10421
rect 17592 10489 17601 10523
rect 17601 10489 17635 10523
rect 17635 10489 17644 10523
rect 17592 10480 17644 10489
rect 4660 10310 4712 10362
rect 4724 10310 4776 10362
rect 4788 10310 4840 10362
rect 4852 10310 4904 10362
rect 4916 10310 4968 10362
rect 7760 10310 7812 10362
rect 7824 10310 7876 10362
rect 7888 10310 7940 10362
rect 7952 10310 8004 10362
rect 8016 10310 8068 10362
rect 10860 10310 10912 10362
rect 10924 10310 10976 10362
rect 10988 10310 11040 10362
rect 11052 10310 11104 10362
rect 11116 10310 11168 10362
rect 13960 10310 14012 10362
rect 14024 10310 14076 10362
rect 14088 10310 14140 10362
rect 14152 10310 14204 10362
rect 14216 10310 14268 10362
rect 17060 10310 17112 10362
rect 17124 10310 17176 10362
rect 17188 10310 17240 10362
rect 17252 10310 17304 10362
rect 17316 10310 17368 10362
rect 2136 10208 2188 10260
rect 756 10140 808 10192
rect 2688 10140 2740 10192
rect 2872 10140 2924 10192
rect 4712 10140 4764 10192
rect 4988 10140 5040 10192
rect 4896 10115 4948 10124
rect 1860 10047 1912 10056
rect 1860 10013 1869 10047
rect 1869 10013 1903 10047
rect 1903 10013 1912 10047
rect 1860 10004 1912 10013
rect 2044 10047 2096 10056
rect 2044 10013 2053 10047
rect 2053 10013 2087 10047
rect 2087 10013 2096 10047
rect 2044 10004 2096 10013
rect 2964 9936 3016 9988
rect 3056 9936 3108 9988
rect 1400 9868 1452 9920
rect 1952 9868 2004 9920
rect 3148 9868 3200 9920
rect 4896 10081 4905 10115
rect 4905 10081 4939 10115
rect 4939 10081 4948 10115
rect 4896 10072 4948 10081
rect 5540 10140 5592 10192
rect 10140 10208 10192 10260
rect 5908 10072 5960 10124
rect 7288 10115 7340 10124
rect 7288 10081 7297 10115
rect 7297 10081 7331 10115
rect 7331 10081 7340 10115
rect 7288 10072 7340 10081
rect 8208 10140 8260 10192
rect 9496 10140 9548 10192
rect 9864 10115 9916 10124
rect 4160 10047 4212 10056
rect 4160 10013 4169 10047
rect 4169 10013 4203 10047
rect 4203 10013 4212 10047
rect 4160 10004 4212 10013
rect 4528 10047 4580 10056
rect 4528 10013 4537 10047
rect 4537 10013 4571 10047
rect 4571 10013 4580 10047
rect 4528 10004 4580 10013
rect 5172 10004 5224 10056
rect 7472 10047 7524 10056
rect 7472 10013 7481 10047
rect 7481 10013 7515 10047
rect 7515 10013 7524 10047
rect 7472 10004 7524 10013
rect 7840 10047 7892 10056
rect 7840 10013 7849 10047
rect 7849 10013 7883 10047
rect 7883 10013 7892 10047
rect 7840 10004 7892 10013
rect 9864 10081 9873 10115
rect 9873 10081 9907 10115
rect 9907 10081 9916 10115
rect 9864 10072 9916 10081
rect 12992 10208 13044 10260
rect 15568 10208 15620 10260
rect 17500 10251 17552 10260
rect 17500 10217 17509 10251
rect 17509 10217 17543 10251
rect 17543 10217 17552 10251
rect 17500 10208 17552 10217
rect 11888 10140 11940 10192
rect 14648 10140 14700 10192
rect 15936 10140 15988 10192
rect 16488 10140 16540 10192
rect 18144 10183 18196 10192
rect 12256 10072 12308 10124
rect 12440 10072 12492 10124
rect 9680 10004 9732 10056
rect 10140 10047 10192 10056
rect 10140 10013 10149 10047
rect 10149 10013 10183 10047
rect 10183 10013 10192 10047
rect 10140 10004 10192 10013
rect 4988 9936 5040 9988
rect 11336 10004 11388 10056
rect 12992 10047 13044 10056
rect 12992 10013 13001 10047
rect 13001 10013 13035 10047
rect 13035 10013 13044 10047
rect 12992 10004 13044 10013
rect 15016 10072 15068 10124
rect 15660 10072 15712 10124
rect 18144 10149 18153 10183
rect 18153 10149 18187 10183
rect 18187 10149 18196 10183
rect 18144 10140 18196 10149
rect 16212 10004 16264 10056
rect 11796 9936 11848 9988
rect 17500 10072 17552 10124
rect 17868 10072 17920 10124
rect 18236 10115 18288 10124
rect 18236 10081 18245 10115
rect 18245 10081 18279 10115
rect 18279 10081 18288 10115
rect 18236 10072 18288 10081
rect 18328 10115 18380 10124
rect 18328 10081 18337 10115
rect 18337 10081 18371 10115
rect 18371 10081 18380 10115
rect 18328 10072 18380 10081
rect 17868 9936 17920 9988
rect 18328 9936 18380 9988
rect 4620 9868 4672 9920
rect 5356 9868 5408 9920
rect 7840 9868 7892 9920
rect 8392 9868 8444 9920
rect 8668 9868 8720 9920
rect 9588 9911 9640 9920
rect 9588 9877 9597 9911
rect 9597 9877 9631 9911
rect 9631 9877 9640 9911
rect 9588 9868 9640 9877
rect 10232 9868 10284 9920
rect 10784 9868 10836 9920
rect 12164 9868 12216 9920
rect 12256 9911 12308 9920
rect 12256 9877 12265 9911
rect 12265 9877 12299 9911
rect 12299 9877 12308 9911
rect 12256 9868 12308 9877
rect 14924 9868 14976 9920
rect 15844 9868 15896 9920
rect 16764 9911 16816 9920
rect 16764 9877 16773 9911
rect 16773 9877 16807 9911
rect 16807 9877 16816 9911
rect 16764 9868 16816 9877
rect 16856 9868 16908 9920
rect 17960 9868 18012 9920
rect 18236 9868 18288 9920
rect 3110 9766 3162 9818
rect 3174 9766 3226 9818
rect 3238 9766 3290 9818
rect 3302 9766 3354 9818
rect 3366 9766 3418 9818
rect 6210 9766 6262 9818
rect 6274 9766 6326 9818
rect 6338 9766 6390 9818
rect 6402 9766 6454 9818
rect 6466 9766 6518 9818
rect 9310 9766 9362 9818
rect 9374 9766 9426 9818
rect 9438 9766 9490 9818
rect 9502 9766 9554 9818
rect 9566 9766 9618 9818
rect 12410 9766 12462 9818
rect 12474 9766 12526 9818
rect 12538 9766 12590 9818
rect 12602 9766 12654 9818
rect 12666 9766 12718 9818
rect 15510 9766 15562 9818
rect 15574 9766 15626 9818
rect 15638 9766 15690 9818
rect 15702 9766 15754 9818
rect 15766 9766 15818 9818
rect 18610 9766 18662 9818
rect 18674 9766 18726 9818
rect 18738 9766 18790 9818
rect 18802 9766 18854 9818
rect 18866 9766 18918 9818
rect 4160 9664 4212 9716
rect 4344 9707 4396 9716
rect 4344 9673 4353 9707
rect 4353 9673 4387 9707
rect 4387 9673 4396 9707
rect 4344 9664 4396 9673
rect 4528 9664 4580 9716
rect 4620 9664 4672 9716
rect 5080 9664 5132 9716
rect 6092 9664 6144 9716
rect 7288 9664 7340 9716
rect 13544 9664 13596 9716
rect 15292 9664 15344 9716
rect 1492 9596 1544 9648
rect 8392 9596 8444 9648
rect 8668 9639 8720 9648
rect 8668 9605 8677 9639
rect 8677 9605 8711 9639
rect 8711 9605 8720 9639
rect 8668 9596 8720 9605
rect 8760 9596 8812 9648
rect 10600 9639 10652 9648
rect 480 9503 532 9512
rect 480 9469 489 9503
rect 489 9469 523 9503
rect 523 9469 532 9503
rect 480 9460 532 9469
rect 1032 9503 1084 9512
rect 664 9392 716 9444
rect 1032 9469 1041 9503
rect 1041 9469 1075 9503
rect 1075 9469 1084 9503
rect 1032 9460 1084 9469
rect 1124 9497 1176 9512
rect 1124 9463 1133 9497
rect 1133 9463 1167 9497
rect 1167 9463 1176 9497
rect 1124 9460 1176 9463
rect 848 9367 900 9376
rect 848 9333 857 9367
rect 857 9333 891 9367
rect 891 9333 900 9367
rect 848 9324 900 9333
rect 940 9324 992 9376
rect 1400 9460 1452 9512
rect 3700 9528 3752 9580
rect 5724 9528 5776 9580
rect 8208 9528 8260 9580
rect 10600 9605 10609 9639
rect 10609 9605 10643 9639
rect 10643 9605 10652 9639
rect 10600 9596 10652 9605
rect 10784 9639 10836 9648
rect 10784 9605 10793 9639
rect 10793 9605 10827 9639
rect 10827 9605 10836 9639
rect 10784 9596 10836 9605
rect 12992 9596 13044 9648
rect 16120 9664 16172 9716
rect 16488 9664 16540 9716
rect 18236 9664 18288 9716
rect 17868 9596 17920 9648
rect 9496 9528 9548 9580
rect 9864 9528 9916 9580
rect 1768 9435 1820 9444
rect 1768 9401 1777 9435
rect 1777 9401 1811 9435
rect 1811 9401 1820 9435
rect 1768 9392 1820 9401
rect 3056 9392 3108 9444
rect 3792 9392 3844 9444
rect 4160 9503 4212 9512
rect 4160 9469 4169 9503
rect 4169 9469 4203 9503
rect 4203 9469 4212 9503
rect 4160 9460 4212 9469
rect 6552 9460 6604 9512
rect 7012 9503 7064 9512
rect 7012 9469 7021 9503
rect 7021 9469 7055 9503
rect 7055 9469 7064 9503
rect 7012 9460 7064 9469
rect 11336 9503 11388 9512
rect 5264 9392 5316 9444
rect 2136 9324 2188 9376
rect 3608 9324 3660 9376
rect 6644 9324 6696 9376
rect 6920 9324 6972 9376
rect 7380 9392 7432 9444
rect 10416 9392 10468 9444
rect 11336 9469 11345 9503
rect 11345 9469 11379 9503
rect 11379 9469 11388 9503
rect 11336 9460 11388 9469
rect 13452 9503 13504 9512
rect 13452 9469 13461 9503
rect 13461 9469 13495 9503
rect 13495 9469 13504 9503
rect 13452 9460 13504 9469
rect 11244 9392 11296 9444
rect 8300 9324 8352 9376
rect 9496 9324 9548 9376
rect 9864 9324 9916 9376
rect 10784 9324 10836 9376
rect 12256 9324 12308 9376
rect 14648 9392 14700 9444
rect 14832 9528 14884 9580
rect 16764 9528 16816 9580
rect 17592 9528 17644 9580
rect 17776 9528 17828 9580
rect 15200 9460 15252 9512
rect 16672 9460 16724 9512
rect 17408 9460 17460 9512
rect 14740 9367 14792 9376
rect 14740 9333 14749 9367
rect 14749 9333 14783 9367
rect 14783 9333 14792 9367
rect 14740 9324 14792 9333
rect 16028 9324 16080 9376
rect 17776 9392 17828 9444
rect 18052 9324 18104 9376
rect 4660 9222 4712 9274
rect 4724 9222 4776 9274
rect 4788 9222 4840 9274
rect 4852 9222 4904 9274
rect 4916 9222 4968 9274
rect 7760 9222 7812 9274
rect 7824 9222 7876 9274
rect 7888 9222 7940 9274
rect 7952 9222 8004 9274
rect 8016 9222 8068 9274
rect 10860 9222 10912 9274
rect 10924 9222 10976 9274
rect 10988 9222 11040 9274
rect 11052 9222 11104 9274
rect 11116 9222 11168 9274
rect 13960 9222 14012 9274
rect 14024 9222 14076 9274
rect 14088 9222 14140 9274
rect 14152 9222 14204 9274
rect 14216 9222 14268 9274
rect 17060 9222 17112 9274
rect 17124 9222 17176 9274
rect 17188 9222 17240 9274
rect 17252 9222 17304 9274
rect 17316 9222 17368 9274
rect 1676 9120 1728 9172
rect 3700 9120 3752 9172
rect 4436 9120 4488 9172
rect 8668 9120 8720 9172
rect 11428 9120 11480 9172
rect 13544 9163 13596 9172
rect 13544 9129 13553 9163
rect 13553 9129 13587 9163
rect 13587 9129 13596 9163
rect 13544 9120 13596 9129
rect 14648 9120 14700 9172
rect 2044 9052 2096 9104
rect 2872 9052 2924 9104
rect 3056 9052 3108 9104
rect 5264 9052 5316 9104
rect 6828 9052 6880 9104
rect 7472 9095 7524 9104
rect 572 8984 624 9036
rect 756 9027 808 9036
rect 756 8993 765 9027
rect 765 8993 799 9027
rect 799 8993 808 9027
rect 756 8984 808 8993
rect 1216 9027 1268 9036
rect 1216 8993 1225 9027
rect 1225 8993 1259 9027
rect 1259 8993 1268 9027
rect 1216 8984 1268 8993
rect 2136 9027 2188 9036
rect 2136 8993 2145 9027
rect 2145 8993 2179 9027
rect 2179 8993 2188 9027
rect 2136 8984 2188 8993
rect 2688 8984 2740 9036
rect 4436 9027 4488 9036
rect 4436 8993 4445 9027
rect 4445 8993 4479 9027
rect 4479 8993 4488 9027
rect 4436 8984 4488 8993
rect 1032 8916 1084 8968
rect 2320 8959 2372 8968
rect 2320 8925 2329 8959
rect 2329 8925 2363 8959
rect 2363 8925 2372 8959
rect 2320 8916 2372 8925
rect 3700 8916 3752 8968
rect 4988 8984 5040 9036
rect 7472 9061 7481 9095
rect 7481 9061 7515 9095
rect 7515 9061 7524 9095
rect 7472 9052 7524 9061
rect 9956 9052 10008 9104
rect 10784 9052 10836 9104
rect 11520 9052 11572 9104
rect 17776 9052 17828 9104
rect 4068 8848 4120 8900
rect 4160 8848 4212 8900
rect 7656 8984 7708 9036
rect 7840 9027 7892 9036
rect 7840 8993 7849 9027
rect 7849 8993 7883 9027
rect 7883 8993 7892 9027
rect 7840 8984 7892 8993
rect 7932 8959 7984 8968
rect 7932 8925 7941 8959
rect 7941 8925 7975 8959
rect 7975 8925 7984 8959
rect 7932 8916 7984 8925
rect 10232 8959 10284 8968
rect 10232 8925 10241 8959
rect 10241 8925 10275 8959
rect 10275 8925 10284 8959
rect 10232 8916 10284 8925
rect 11244 8916 11296 8968
rect 11888 8916 11940 8968
rect 12072 9027 12124 9036
rect 12072 8993 12081 9027
rect 12081 8993 12115 9027
rect 12115 8993 12124 9027
rect 12072 8984 12124 8993
rect 13728 8916 13780 8968
rect 16580 8984 16632 9036
rect 14832 8959 14884 8968
rect 14832 8925 14841 8959
rect 14841 8925 14875 8959
rect 14875 8925 14884 8959
rect 14832 8916 14884 8925
rect 16856 8916 16908 8968
rect 17500 8959 17552 8968
rect 17500 8925 17509 8959
rect 17509 8925 17543 8959
rect 17543 8925 17552 8959
rect 17500 8916 17552 8925
rect 4344 8780 4396 8832
rect 5724 8823 5776 8832
rect 5724 8789 5733 8823
rect 5733 8789 5767 8823
rect 5767 8789 5776 8823
rect 5724 8780 5776 8789
rect 16672 8848 16724 8900
rect 17592 8848 17644 8900
rect 9864 8780 9916 8832
rect 11980 8823 12032 8832
rect 11980 8789 11989 8823
rect 11989 8789 12023 8823
rect 12023 8789 12032 8823
rect 11980 8780 12032 8789
rect 15108 8780 15160 8832
rect 16764 8823 16816 8832
rect 16764 8789 16773 8823
rect 16773 8789 16807 8823
rect 16807 8789 16816 8823
rect 16764 8780 16816 8789
rect 3110 8678 3162 8730
rect 3174 8678 3226 8730
rect 3238 8678 3290 8730
rect 3302 8678 3354 8730
rect 3366 8678 3418 8730
rect 6210 8678 6262 8730
rect 6274 8678 6326 8730
rect 6338 8678 6390 8730
rect 6402 8678 6454 8730
rect 6466 8678 6518 8730
rect 9310 8678 9362 8730
rect 9374 8678 9426 8730
rect 9438 8678 9490 8730
rect 9502 8678 9554 8730
rect 9566 8678 9618 8730
rect 12410 8678 12462 8730
rect 12474 8678 12526 8730
rect 12538 8678 12590 8730
rect 12602 8678 12654 8730
rect 12666 8678 12718 8730
rect 15510 8678 15562 8730
rect 15574 8678 15626 8730
rect 15638 8678 15690 8730
rect 15702 8678 15754 8730
rect 15766 8678 15818 8730
rect 18610 8678 18662 8730
rect 18674 8678 18726 8730
rect 18738 8678 18790 8730
rect 18802 8678 18854 8730
rect 18866 8678 18918 8730
rect 756 8576 808 8628
rect 3424 8619 3476 8628
rect 572 8372 624 8424
rect 1308 8551 1360 8560
rect 1308 8517 1317 8551
rect 1317 8517 1351 8551
rect 1351 8517 1360 8551
rect 1308 8508 1360 8517
rect 3424 8585 3433 8619
rect 3433 8585 3467 8619
rect 3467 8585 3476 8619
rect 3424 8576 3476 8585
rect 3700 8619 3752 8628
rect 3700 8585 3709 8619
rect 3709 8585 3743 8619
rect 3743 8585 3752 8619
rect 3700 8576 3752 8585
rect 3976 8619 4028 8628
rect 3976 8585 3985 8619
rect 3985 8585 4019 8619
rect 4019 8585 4028 8619
rect 3976 8576 4028 8585
rect 4252 8619 4304 8628
rect 4252 8585 4261 8619
rect 4261 8585 4295 8619
rect 4295 8585 4304 8619
rect 4252 8576 4304 8585
rect 6552 8619 6604 8628
rect 6552 8585 6561 8619
rect 6561 8585 6595 8619
rect 6595 8585 6604 8619
rect 6552 8576 6604 8585
rect 9680 8576 9732 8628
rect 10600 8576 10652 8628
rect 3516 8508 3568 8560
rect 3608 8508 3660 8560
rect 1124 8440 1176 8492
rect 3424 8440 3476 8492
rect 8300 8508 8352 8560
rect 1400 8372 1452 8424
rect 2872 8372 2924 8424
rect 3056 8372 3108 8424
rect 3516 8415 3568 8424
rect 756 8304 808 8356
rect 3516 8381 3525 8415
rect 3525 8381 3559 8415
rect 3559 8381 3568 8415
rect 3516 8372 3568 8381
rect 5172 8440 5224 8492
rect 5540 8440 5592 8492
rect 3884 8415 3936 8424
rect 3884 8381 3893 8415
rect 3893 8381 3927 8415
rect 3927 8381 3936 8415
rect 3884 8372 3936 8381
rect 4252 8372 4304 8424
rect 7104 8440 7156 8492
rect 7840 8440 7892 8492
rect 12256 8508 12308 8560
rect 13820 8576 13872 8628
rect 15936 8576 15988 8628
rect 18328 8619 18380 8628
rect 18328 8585 18337 8619
rect 18337 8585 18371 8619
rect 18371 8585 18380 8619
rect 18328 8576 18380 8585
rect 6920 8372 6972 8424
rect 7932 8372 7984 8424
rect 9036 8372 9088 8424
rect 10600 8372 10652 8424
rect 12808 8440 12860 8492
rect 11428 8415 11480 8424
rect 572 8279 624 8288
rect 572 8245 581 8279
rect 581 8245 615 8279
rect 615 8245 624 8279
rect 572 8236 624 8245
rect 2596 8236 2648 8288
rect 4436 8304 4488 8356
rect 8852 8304 8904 8356
rect 10784 8304 10836 8356
rect 3424 8236 3476 8288
rect 5356 8236 5408 8288
rect 10140 8236 10192 8288
rect 11428 8381 11437 8415
rect 11437 8381 11471 8415
rect 11471 8381 11480 8415
rect 11428 8372 11480 8381
rect 12348 8372 12400 8424
rect 17592 8508 17644 8560
rect 13820 8440 13872 8492
rect 13544 8372 13596 8424
rect 13728 8372 13780 8424
rect 14372 8372 14424 8424
rect 17684 8440 17736 8492
rect 16764 8372 16816 8424
rect 16948 8372 17000 8424
rect 12164 8304 12216 8356
rect 15844 8347 15896 8356
rect 11520 8236 11572 8288
rect 12072 8236 12124 8288
rect 13084 8279 13136 8288
rect 13084 8245 13093 8279
rect 13093 8245 13127 8279
rect 13127 8245 13136 8279
rect 13084 8236 13136 8245
rect 13176 8236 13228 8288
rect 15844 8313 15853 8347
rect 15853 8313 15887 8347
rect 15887 8313 15896 8347
rect 15844 8304 15896 8313
rect 17500 8304 17552 8356
rect 18328 8372 18380 8424
rect 16856 8236 16908 8288
rect 17408 8236 17460 8288
rect 17960 8279 18012 8288
rect 17960 8245 17969 8279
rect 17969 8245 18003 8279
rect 18003 8245 18012 8279
rect 17960 8236 18012 8245
rect 4660 8134 4712 8186
rect 4724 8134 4776 8186
rect 4788 8134 4840 8186
rect 4852 8134 4904 8186
rect 4916 8134 4968 8186
rect 7760 8134 7812 8186
rect 7824 8134 7876 8186
rect 7888 8134 7940 8186
rect 7952 8134 8004 8186
rect 8016 8134 8068 8186
rect 10860 8134 10912 8186
rect 10924 8134 10976 8186
rect 10988 8134 11040 8186
rect 11052 8134 11104 8186
rect 11116 8134 11168 8186
rect 13960 8134 14012 8186
rect 14024 8134 14076 8186
rect 14088 8134 14140 8186
rect 14152 8134 14204 8186
rect 14216 8134 14268 8186
rect 17060 8134 17112 8186
rect 17124 8134 17176 8186
rect 17188 8134 17240 8186
rect 17252 8134 17304 8186
rect 17316 8134 17368 8186
rect 572 8032 624 8084
rect 2412 8032 2464 8084
rect 4160 8032 4212 8084
rect 5080 8032 5132 8084
rect 7196 8075 7248 8084
rect 7196 8041 7205 8075
rect 7205 8041 7239 8075
rect 7239 8041 7248 8075
rect 7196 8032 7248 8041
rect 9772 8032 9824 8084
rect 10048 8032 10100 8084
rect 14740 8032 14792 8084
rect 15016 8032 15068 8084
rect 16212 8032 16264 8084
rect 664 8007 716 8016
rect 664 7973 673 8007
rect 673 7973 707 8007
rect 707 7973 716 8007
rect 664 7964 716 7973
rect 2964 7964 3016 8016
rect 3884 7964 3936 8016
rect 4436 7964 4488 8016
rect 572 7896 624 7948
rect 1124 7896 1176 7948
rect 1216 7871 1268 7880
rect 1216 7837 1225 7871
rect 1225 7837 1259 7871
rect 1259 7837 1268 7871
rect 1216 7828 1268 7837
rect 2228 7871 2280 7880
rect 2228 7837 2237 7871
rect 2237 7837 2271 7871
rect 2271 7837 2280 7871
rect 2228 7828 2280 7837
rect 2412 7871 2464 7880
rect 2412 7837 2421 7871
rect 2421 7837 2455 7871
rect 2455 7837 2464 7871
rect 2412 7828 2464 7837
rect 2780 7828 2832 7880
rect 4068 7896 4120 7948
rect 8392 7964 8444 8016
rect 11704 7964 11756 8016
rect 11980 8007 12032 8016
rect 11980 7973 11989 8007
rect 11989 7973 12023 8007
rect 12023 7973 12032 8007
rect 11980 7964 12032 7973
rect 6092 7939 6144 7948
rect 6092 7905 6101 7939
rect 6101 7905 6135 7939
rect 6135 7905 6144 7939
rect 6092 7896 6144 7905
rect 6184 7896 6236 7948
rect 6644 7896 6696 7948
rect 6828 7939 6880 7948
rect 6828 7905 6837 7939
rect 6837 7905 6871 7939
rect 6871 7905 6880 7939
rect 6828 7896 6880 7905
rect 7012 7939 7064 7948
rect 7012 7905 7021 7939
rect 7021 7905 7055 7939
rect 7055 7905 7064 7939
rect 7012 7896 7064 7905
rect 7656 7896 7708 7948
rect 8300 7896 8352 7948
rect 9772 7896 9824 7948
rect 11796 7939 11848 7948
rect 11796 7905 11805 7939
rect 11805 7905 11839 7939
rect 11839 7905 11848 7939
rect 11796 7896 11848 7905
rect 12072 7939 12124 7948
rect 12072 7905 12081 7939
rect 12081 7905 12115 7939
rect 12115 7905 12124 7939
rect 12072 7896 12124 7905
rect 3516 7871 3568 7880
rect 3516 7837 3525 7871
rect 3525 7837 3559 7871
rect 3559 7837 3568 7871
rect 3516 7828 3568 7837
rect 4988 7828 5040 7880
rect 5724 7828 5776 7880
rect 6552 7828 6604 7880
rect 14372 7964 14424 8016
rect 16120 7964 16172 8016
rect 16488 7964 16540 8016
rect 16672 7964 16724 8016
rect 17316 8032 17368 8084
rect 17408 8032 17460 8084
rect 18144 8032 18196 8084
rect 13728 7896 13780 7948
rect 15016 7939 15068 7948
rect 15016 7905 15025 7939
rect 15025 7905 15059 7939
rect 15059 7905 15068 7939
rect 15016 7896 15068 7905
rect 16856 7939 16908 7948
rect 16856 7905 16865 7939
rect 16865 7905 16899 7939
rect 16899 7905 16908 7939
rect 16856 7896 16908 7905
rect 17224 7939 17276 7948
rect 17224 7905 17233 7939
rect 17233 7905 17267 7939
rect 17267 7905 17276 7939
rect 17224 7896 17276 7905
rect 17408 7896 17460 7948
rect 17684 7896 17736 7948
rect 18420 7939 18472 7948
rect 18420 7905 18429 7939
rect 18429 7905 18463 7939
rect 18463 7905 18472 7939
rect 18420 7896 18472 7905
rect 1492 7760 1544 7812
rect 2136 7760 2188 7812
rect 5172 7760 5224 7812
rect 9128 7760 9180 7812
rect 1676 7735 1728 7744
rect 1676 7701 1685 7735
rect 1685 7701 1719 7735
rect 1719 7701 1728 7735
rect 1676 7692 1728 7701
rect 2872 7692 2924 7744
rect 3056 7692 3108 7744
rect 3700 7692 3752 7744
rect 3884 7692 3936 7744
rect 5816 7692 5868 7744
rect 8484 7692 8536 7744
rect 9864 7692 9916 7744
rect 11888 7760 11940 7812
rect 13268 7760 13320 7812
rect 16120 7828 16172 7880
rect 17316 7828 17368 7880
rect 17868 7828 17920 7880
rect 11520 7692 11572 7744
rect 12256 7692 12308 7744
rect 13820 7692 13872 7744
rect 15292 7692 15344 7744
rect 18328 7760 18380 7812
rect 17408 7692 17460 7744
rect 3110 7590 3162 7642
rect 3174 7590 3226 7642
rect 3238 7590 3290 7642
rect 3302 7590 3354 7642
rect 3366 7590 3418 7642
rect 6210 7590 6262 7642
rect 6274 7590 6326 7642
rect 6338 7590 6390 7642
rect 6402 7590 6454 7642
rect 6466 7590 6518 7642
rect 9310 7590 9362 7642
rect 9374 7590 9426 7642
rect 9438 7590 9490 7642
rect 9502 7590 9554 7642
rect 9566 7590 9618 7642
rect 12410 7590 12462 7642
rect 12474 7590 12526 7642
rect 12538 7590 12590 7642
rect 12602 7590 12654 7642
rect 12666 7590 12718 7642
rect 15510 7590 15562 7642
rect 15574 7590 15626 7642
rect 15638 7590 15690 7642
rect 15702 7590 15754 7642
rect 15766 7590 15818 7642
rect 18610 7590 18662 7642
rect 18674 7590 18726 7642
rect 18738 7590 18790 7642
rect 18802 7590 18854 7642
rect 18866 7590 18918 7642
rect 756 7488 808 7540
rect 1216 7488 1268 7540
rect 3332 7488 3384 7540
rect 3608 7488 3660 7540
rect 940 7420 992 7472
rect 2780 7420 2832 7472
rect 3976 7420 4028 7472
rect 4068 7420 4120 7472
rect 848 7352 900 7404
rect 1308 7395 1360 7404
rect 1308 7361 1317 7395
rect 1317 7361 1351 7395
rect 1351 7361 1360 7395
rect 1308 7352 1360 7361
rect 2136 7352 2188 7404
rect 480 7327 532 7336
rect 480 7293 489 7327
rect 489 7293 523 7327
rect 523 7293 532 7327
rect 480 7284 532 7293
rect 1124 7284 1176 7336
rect 1216 7327 1268 7336
rect 1216 7293 1225 7327
rect 1225 7293 1259 7327
rect 1259 7293 1268 7327
rect 1216 7284 1268 7293
rect 1400 7284 1452 7336
rect 2872 7284 2924 7336
rect 3792 7352 3844 7404
rect 4068 7327 4120 7336
rect 1032 7148 1084 7200
rect 1768 7259 1820 7268
rect 1768 7225 1777 7259
rect 1777 7225 1811 7259
rect 1811 7225 1820 7259
rect 4068 7293 4077 7327
rect 4077 7293 4111 7327
rect 4111 7293 4120 7327
rect 4068 7284 4120 7293
rect 4252 7284 4304 7336
rect 4436 7284 4488 7336
rect 5356 7488 5408 7540
rect 5540 7327 5592 7336
rect 5540 7293 5549 7327
rect 5549 7293 5583 7327
rect 5583 7293 5592 7327
rect 5540 7284 5592 7293
rect 7012 7488 7064 7540
rect 7656 7488 7708 7540
rect 10140 7488 10192 7540
rect 11336 7531 11388 7540
rect 11336 7497 11345 7531
rect 11345 7497 11379 7531
rect 11379 7497 11388 7531
rect 11336 7488 11388 7497
rect 12992 7488 13044 7540
rect 16580 7488 16632 7540
rect 18512 7488 18564 7540
rect 6552 7352 6604 7404
rect 7656 7352 7708 7404
rect 8944 7420 8996 7472
rect 9404 7395 9456 7404
rect 9404 7361 9413 7395
rect 9413 7361 9447 7395
rect 9447 7361 9456 7395
rect 9404 7352 9456 7361
rect 9772 7420 9824 7472
rect 14372 7420 14424 7472
rect 15016 7420 15068 7472
rect 18328 7463 18380 7472
rect 11796 7352 11848 7404
rect 6644 7327 6696 7336
rect 6644 7293 6653 7327
rect 6653 7293 6687 7327
rect 6687 7293 6696 7327
rect 6644 7284 6696 7293
rect 8852 7284 8904 7336
rect 9036 7327 9088 7336
rect 9036 7293 9045 7327
rect 9045 7293 9079 7327
rect 9079 7293 9088 7327
rect 9036 7284 9088 7293
rect 10416 7327 10468 7336
rect 10416 7293 10425 7327
rect 10425 7293 10459 7327
rect 10459 7293 10468 7327
rect 10416 7284 10468 7293
rect 15844 7352 15896 7404
rect 18328 7429 18337 7463
rect 18337 7429 18371 7463
rect 18371 7429 18380 7463
rect 18328 7420 18380 7429
rect 13268 7327 13320 7336
rect 13268 7293 13277 7327
rect 13277 7293 13311 7327
rect 13311 7293 13320 7327
rect 13268 7284 13320 7293
rect 1768 7216 1820 7225
rect 2780 7148 2832 7200
rect 3424 7148 3476 7200
rect 5172 7216 5224 7268
rect 5816 7259 5868 7268
rect 5816 7225 5825 7259
rect 5825 7225 5859 7259
rect 5859 7225 5868 7259
rect 5816 7216 5868 7225
rect 3976 7191 4028 7200
rect 3976 7157 3985 7191
rect 3985 7157 4019 7191
rect 4019 7157 4028 7191
rect 3976 7148 4028 7157
rect 4988 7148 5040 7200
rect 5264 7148 5316 7200
rect 8300 7216 8352 7268
rect 9496 7216 9548 7268
rect 11704 7148 11756 7200
rect 13452 7259 13504 7268
rect 13452 7225 13461 7259
rect 13461 7225 13495 7259
rect 13495 7225 13504 7259
rect 15016 7284 15068 7336
rect 15936 7284 15988 7336
rect 17224 7352 17276 7404
rect 16212 7327 16264 7336
rect 16212 7293 16221 7327
rect 16221 7293 16255 7327
rect 16255 7293 16264 7327
rect 16212 7284 16264 7293
rect 18512 7327 18564 7336
rect 13452 7216 13504 7225
rect 18512 7293 18521 7327
rect 18521 7293 18555 7327
rect 18555 7293 18564 7327
rect 18512 7284 18564 7293
rect 16672 7216 16724 7268
rect 14740 7148 14792 7200
rect 15752 7148 15804 7200
rect 16212 7148 16264 7200
rect 16396 7148 16448 7200
rect 18328 7148 18380 7200
rect 4660 7046 4712 7098
rect 4724 7046 4776 7098
rect 4788 7046 4840 7098
rect 4852 7046 4904 7098
rect 4916 7046 4968 7098
rect 7760 7046 7812 7098
rect 7824 7046 7876 7098
rect 7888 7046 7940 7098
rect 7952 7046 8004 7098
rect 8016 7046 8068 7098
rect 10860 7046 10912 7098
rect 10924 7046 10976 7098
rect 10988 7046 11040 7098
rect 11052 7046 11104 7098
rect 11116 7046 11168 7098
rect 13960 7046 14012 7098
rect 14024 7046 14076 7098
rect 14088 7046 14140 7098
rect 14152 7046 14204 7098
rect 14216 7046 14268 7098
rect 17060 7046 17112 7098
rect 17124 7046 17176 7098
rect 17188 7046 17240 7098
rect 17252 7046 17304 7098
rect 17316 7046 17368 7098
rect 480 6944 532 6996
rect 2136 6944 2188 6996
rect 2412 6987 2464 6996
rect 2412 6953 2421 6987
rect 2421 6953 2455 6987
rect 2455 6953 2464 6987
rect 2412 6944 2464 6953
rect 3240 6944 3292 6996
rect 3332 6944 3384 6996
rect 4252 6944 4304 6996
rect 756 6851 808 6860
rect 756 6817 765 6851
rect 765 6817 799 6851
rect 799 6817 808 6851
rect 756 6808 808 6817
rect 848 6851 900 6860
rect 848 6817 857 6851
rect 857 6817 891 6851
rect 891 6817 900 6851
rect 848 6808 900 6817
rect 3056 6919 3108 6928
rect 3056 6885 3065 6919
rect 3065 6885 3099 6919
rect 3099 6885 3108 6919
rect 3056 6876 3108 6885
rect 4160 6876 4212 6928
rect 4988 6944 5040 6996
rect 6828 6944 6880 6996
rect 8760 6944 8812 6996
rect 9404 6944 9456 6996
rect 9680 6944 9732 6996
rect 10324 6944 10376 6996
rect 12900 6944 12952 6996
rect 13820 6944 13872 6996
rect 1492 6783 1544 6792
rect 1492 6749 1501 6783
rect 1501 6749 1535 6783
rect 1535 6749 1544 6783
rect 1492 6740 1544 6749
rect 1676 6783 1728 6792
rect 1676 6749 1685 6783
rect 1685 6749 1719 6783
rect 1719 6749 1728 6783
rect 1676 6740 1728 6749
rect 2964 6808 3016 6860
rect 3700 6808 3752 6860
rect 4252 6851 4304 6860
rect 4252 6817 4261 6851
rect 4261 6817 4295 6851
rect 4295 6817 4304 6851
rect 4252 6808 4304 6817
rect 6920 6808 6972 6860
rect 7196 6919 7248 6928
rect 7196 6885 7205 6919
rect 7205 6885 7239 6919
rect 7239 6885 7248 6919
rect 7196 6876 7248 6885
rect 8944 6876 8996 6928
rect 2688 6740 2740 6792
rect 4068 6740 4120 6792
rect 4528 6783 4580 6792
rect 4528 6749 4537 6783
rect 4537 6749 4571 6783
rect 4571 6749 4580 6783
rect 4528 6740 4580 6749
rect 5540 6740 5592 6792
rect 7288 6740 7340 6792
rect 7564 6808 7616 6860
rect 7840 6851 7892 6860
rect 7840 6817 7849 6851
rect 7849 6817 7883 6851
rect 7883 6817 7892 6851
rect 7840 6808 7892 6817
rect 7932 6851 7984 6860
rect 7932 6817 7941 6851
rect 7941 6817 7975 6851
rect 7975 6817 7984 6851
rect 7932 6808 7984 6817
rect 8392 6808 8444 6860
rect 8576 6851 8628 6860
rect 8576 6817 8585 6851
rect 8585 6817 8619 6851
rect 8619 6817 8628 6851
rect 8576 6808 8628 6817
rect 8852 6808 8904 6860
rect 9220 6808 9272 6860
rect 10140 6876 10192 6928
rect 12164 6876 12216 6928
rect 9496 6851 9548 6860
rect 9496 6817 9505 6851
rect 9505 6817 9539 6851
rect 9539 6817 9548 6851
rect 9496 6808 9548 6817
rect 9864 6851 9916 6860
rect 9864 6817 9873 6851
rect 9873 6817 9907 6851
rect 9907 6817 9916 6851
rect 9864 6808 9916 6817
rect 11888 6808 11940 6860
rect 14832 6944 14884 6996
rect 16212 6944 16264 6996
rect 15016 6876 15068 6928
rect 15108 6876 15160 6928
rect 15292 6876 15344 6928
rect 16396 6876 16448 6928
rect 3976 6672 4028 6724
rect 4620 6672 4672 6724
rect 1124 6604 1176 6656
rect 1860 6604 1912 6656
rect 2964 6604 3016 6656
rect 3240 6604 3292 6656
rect 4344 6604 4396 6656
rect 7012 6672 7064 6724
rect 5264 6604 5316 6656
rect 6920 6604 6972 6656
rect 7380 6672 7432 6724
rect 7656 6672 7708 6724
rect 7288 6604 7340 6656
rect 8760 6783 8812 6792
rect 8760 6749 8769 6783
rect 8769 6749 8803 6783
rect 8803 6749 8812 6783
rect 8760 6740 8812 6749
rect 9772 6740 9824 6792
rect 11704 6783 11756 6792
rect 11704 6749 11713 6783
rect 11713 6749 11747 6783
rect 11747 6749 11756 6783
rect 11704 6740 11756 6749
rect 11796 6740 11848 6792
rect 14648 6851 14700 6860
rect 12716 6740 12768 6792
rect 13452 6740 13504 6792
rect 13544 6740 13596 6792
rect 14648 6817 14657 6851
rect 14657 6817 14691 6851
rect 14691 6817 14700 6851
rect 14648 6808 14700 6817
rect 14832 6851 14884 6860
rect 14832 6817 14845 6851
rect 14845 6817 14884 6851
rect 14832 6808 14884 6817
rect 14924 6740 14976 6792
rect 14464 6672 14516 6724
rect 15016 6715 15068 6724
rect 15016 6681 15025 6715
rect 15025 6681 15059 6715
rect 15059 6681 15068 6715
rect 15016 6672 15068 6681
rect 8392 6604 8444 6656
rect 8852 6604 8904 6656
rect 8944 6604 8996 6656
rect 11980 6604 12032 6656
rect 12716 6604 12768 6656
rect 13728 6604 13780 6656
rect 13912 6604 13964 6656
rect 16120 6740 16172 6792
rect 16948 6808 17000 6860
rect 17132 6808 17184 6860
rect 16856 6604 16908 6656
rect 3110 6502 3162 6554
rect 3174 6502 3226 6554
rect 3238 6502 3290 6554
rect 3302 6502 3354 6554
rect 3366 6502 3418 6554
rect 6210 6502 6262 6554
rect 6274 6502 6326 6554
rect 6338 6502 6390 6554
rect 6402 6502 6454 6554
rect 6466 6502 6518 6554
rect 9310 6502 9362 6554
rect 9374 6502 9426 6554
rect 9438 6502 9490 6554
rect 9502 6502 9554 6554
rect 9566 6502 9618 6554
rect 12410 6502 12462 6554
rect 12474 6502 12526 6554
rect 12538 6502 12590 6554
rect 12602 6502 12654 6554
rect 12666 6502 12718 6554
rect 15510 6502 15562 6554
rect 15574 6502 15626 6554
rect 15638 6502 15690 6554
rect 15702 6502 15754 6554
rect 15766 6502 15818 6554
rect 18610 6502 18662 6554
rect 18674 6502 18726 6554
rect 18738 6502 18790 6554
rect 18802 6502 18854 6554
rect 18866 6502 18918 6554
rect 572 6443 624 6452
rect 572 6409 581 6443
rect 581 6409 615 6443
rect 615 6409 624 6443
rect 572 6400 624 6409
rect 1676 6400 1728 6452
rect 6000 6400 6052 6452
rect 6276 6400 6328 6452
rect 6828 6400 6880 6452
rect 9680 6400 9732 6452
rect 1124 6332 1176 6384
rect 2872 6332 2924 6384
rect 3056 6332 3108 6384
rect 3240 6375 3292 6384
rect 3240 6341 3249 6375
rect 3249 6341 3283 6375
rect 3283 6341 3292 6375
rect 3240 6332 3292 6341
rect 4528 6332 4580 6384
rect 1216 6264 1268 6316
rect 1860 6307 1912 6316
rect 848 6239 900 6248
rect 848 6205 857 6239
rect 857 6205 891 6239
rect 891 6205 900 6239
rect 848 6196 900 6205
rect 1032 6239 1084 6248
rect 1032 6205 1041 6239
rect 1041 6205 1075 6239
rect 1075 6205 1084 6239
rect 1032 6196 1084 6205
rect 1308 6239 1360 6248
rect 1308 6205 1317 6239
rect 1317 6205 1351 6239
rect 1351 6205 1360 6239
rect 1308 6196 1360 6205
rect 1492 6239 1544 6248
rect 1492 6205 1501 6239
rect 1501 6205 1535 6239
rect 1535 6205 1544 6239
rect 1492 6196 1544 6205
rect 1860 6273 1869 6307
rect 1869 6273 1903 6307
rect 1903 6273 1912 6307
rect 1860 6264 1912 6273
rect 2044 6264 2096 6316
rect 8668 6332 8720 6384
rect 8852 6332 8904 6384
rect 11888 6400 11940 6452
rect 12716 6400 12768 6452
rect 15384 6400 15436 6452
rect 15936 6400 15988 6452
rect 16488 6400 16540 6452
rect 16672 6400 16724 6452
rect 18052 6400 18104 6452
rect 5540 6264 5592 6316
rect 5908 6307 5960 6316
rect 5908 6273 5917 6307
rect 5917 6273 5951 6307
rect 5951 6273 5960 6307
rect 5908 6264 5960 6273
rect 3608 6196 3660 6248
rect 3976 6239 4028 6248
rect 3976 6205 3985 6239
rect 3985 6205 4019 6239
rect 4019 6205 4028 6239
rect 3976 6196 4028 6205
rect 7196 6264 7248 6316
rect 8208 6264 8260 6316
rect 6276 6239 6328 6248
rect 6276 6205 6285 6239
rect 6285 6205 6319 6239
rect 6319 6205 6328 6239
rect 6276 6196 6328 6205
rect 3884 6128 3936 6180
rect 4068 6060 4120 6112
rect 5632 6128 5684 6180
rect 6092 6128 6144 6180
rect 6552 6239 6604 6248
rect 6552 6205 6561 6239
rect 6561 6205 6595 6239
rect 6595 6205 6604 6239
rect 6552 6196 6604 6205
rect 6828 6196 6880 6248
rect 12900 6264 12952 6316
rect 8852 6239 8904 6248
rect 8852 6205 8861 6239
rect 8861 6205 8895 6239
rect 8895 6205 8904 6239
rect 8852 6196 8904 6205
rect 7656 6128 7708 6180
rect 9128 6171 9180 6180
rect 9128 6137 9137 6171
rect 9137 6137 9171 6171
rect 9171 6137 9180 6171
rect 9128 6128 9180 6137
rect 4988 6060 5040 6112
rect 5816 6103 5868 6112
rect 5816 6069 5825 6103
rect 5825 6069 5859 6103
rect 5859 6069 5868 6103
rect 5816 6060 5868 6069
rect 6000 6060 6052 6112
rect 7380 6060 7432 6112
rect 9220 6060 9272 6112
rect 11428 6128 11480 6180
rect 12072 6128 12124 6180
rect 13084 6171 13136 6180
rect 13084 6137 13093 6171
rect 13093 6137 13127 6171
rect 13127 6137 13136 6171
rect 13084 6128 13136 6137
rect 13452 6332 13504 6384
rect 13912 6307 13964 6316
rect 13912 6273 13921 6307
rect 13921 6273 13955 6307
rect 13955 6273 13964 6307
rect 13912 6264 13964 6273
rect 17868 6332 17920 6384
rect 18420 6332 18472 6384
rect 14556 6264 14608 6316
rect 12716 6060 12768 6112
rect 13544 6103 13596 6112
rect 13544 6069 13553 6103
rect 13553 6069 13587 6103
rect 13587 6069 13596 6103
rect 13544 6060 13596 6069
rect 14464 6128 14516 6180
rect 14924 6128 14976 6180
rect 16580 6264 16632 6316
rect 17776 6196 17828 6248
rect 17960 6196 18012 6248
rect 16120 6171 16172 6180
rect 16120 6137 16129 6171
rect 16129 6137 16163 6171
rect 16163 6137 16172 6171
rect 16120 6128 16172 6137
rect 18052 6171 18104 6180
rect 16212 6060 16264 6112
rect 16304 6060 16356 6112
rect 17684 6060 17736 6112
rect 18052 6137 18061 6171
rect 18061 6137 18095 6171
rect 18095 6137 18104 6171
rect 18052 6128 18104 6137
rect 18972 6196 19024 6248
rect 4660 5958 4712 6010
rect 4724 5958 4776 6010
rect 4788 5958 4840 6010
rect 4852 5958 4904 6010
rect 4916 5958 4968 6010
rect 7760 5958 7812 6010
rect 7824 5958 7876 6010
rect 7888 5958 7940 6010
rect 7952 5958 8004 6010
rect 8016 5958 8068 6010
rect 10860 5958 10912 6010
rect 10924 5958 10976 6010
rect 10988 5958 11040 6010
rect 11052 5958 11104 6010
rect 11116 5958 11168 6010
rect 13960 5958 14012 6010
rect 14024 5958 14076 6010
rect 14088 5958 14140 6010
rect 14152 5958 14204 6010
rect 14216 5958 14268 6010
rect 17060 5958 17112 6010
rect 17124 5958 17176 6010
rect 17188 5958 17240 6010
rect 17252 5958 17304 6010
rect 17316 5958 17368 6010
rect 1492 5856 1544 5908
rect 1584 5856 1636 5908
rect 3056 5856 3108 5908
rect 3516 5856 3568 5908
rect 3884 5856 3936 5908
rect 6920 5856 6972 5908
rect 8208 5856 8260 5908
rect 8576 5856 8628 5908
rect 9956 5856 10008 5908
rect 1492 5720 1544 5772
rect 2136 5763 2188 5772
rect 940 5652 992 5704
rect 2136 5729 2145 5763
rect 2145 5729 2179 5763
rect 2179 5729 2188 5763
rect 2136 5720 2188 5729
rect 3792 5788 3844 5840
rect 4068 5831 4120 5840
rect 4068 5797 4077 5831
rect 4077 5797 4111 5831
rect 4111 5797 4120 5831
rect 4068 5788 4120 5797
rect 2596 5720 2648 5772
rect 2780 5720 2832 5772
rect 4344 5788 4396 5840
rect 9128 5788 9180 5840
rect 2044 5695 2096 5704
rect 2044 5661 2053 5695
rect 2053 5661 2087 5695
rect 2087 5661 2096 5695
rect 2044 5652 2096 5661
rect 2228 5652 2280 5704
rect 4528 5652 4580 5704
rect 3700 5627 3752 5636
rect 3700 5593 3709 5627
rect 3709 5593 3743 5627
rect 3743 5593 3752 5627
rect 3700 5584 3752 5593
rect 5816 5720 5868 5772
rect 5908 5652 5960 5704
rect 6276 5652 6328 5704
rect 7380 5720 7432 5772
rect 7748 5720 7800 5772
rect 7932 5763 7984 5772
rect 7932 5729 7941 5763
rect 7941 5729 7975 5763
rect 7975 5729 7984 5763
rect 7932 5720 7984 5729
rect 8484 5720 8536 5772
rect 9680 5788 9732 5840
rect 10048 5788 10100 5840
rect 10692 5788 10744 5840
rect 11428 5788 11480 5840
rect 9404 5763 9456 5772
rect 9404 5729 9413 5763
rect 9413 5729 9447 5763
rect 9447 5729 9456 5763
rect 9404 5720 9456 5729
rect 11704 5763 11756 5772
rect 11704 5729 11713 5763
rect 11713 5729 11747 5763
rect 11747 5729 11756 5763
rect 11704 5720 11756 5729
rect 11888 5763 11940 5772
rect 11888 5729 11897 5763
rect 11897 5729 11931 5763
rect 11931 5729 11940 5763
rect 11888 5720 11940 5729
rect 12624 5788 12676 5840
rect 12992 5788 13044 5840
rect 14464 5856 14516 5908
rect 17132 5856 17184 5908
rect 17316 5856 17368 5908
rect 17500 5856 17552 5908
rect 18052 5856 18104 5908
rect 15108 5788 15160 5840
rect 16028 5788 16080 5840
rect 16396 5788 16448 5840
rect 8760 5695 8812 5704
rect 8760 5661 8769 5695
rect 8769 5661 8803 5695
rect 8803 5661 8812 5695
rect 8760 5652 8812 5661
rect 9036 5652 9088 5704
rect 5724 5584 5776 5636
rect 7012 5584 7064 5636
rect 7840 5627 7892 5636
rect 7840 5593 7849 5627
rect 7849 5593 7883 5627
rect 7883 5593 7892 5627
rect 7840 5584 7892 5593
rect 11612 5695 11664 5704
rect 11612 5661 11621 5695
rect 11621 5661 11655 5695
rect 11655 5661 11664 5695
rect 11612 5652 11664 5661
rect 14464 5720 14516 5772
rect 18144 5788 18196 5840
rect 16764 5720 16816 5772
rect 17224 5720 17276 5772
rect 18052 5763 18104 5772
rect 18052 5729 18061 5763
rect 18061 5729 18095 5763
rect 18095 5729 18104 5763
rect 18420 5788 18472 5840
rect 18052 5720 18104 5729
rect 12716 5652 12768 5704
rect 13084 5652 13136 5704
rect 1400 5516 1452 5568
rect 4436 5516 4488 5568
rect 5264 5516 5316 5568
rect 7656 5516 7708 5568
rect 8208 5559 8260 5568
rect 8208 5525 8217 5559
rect 8217 5525 8251 5559
rect 8251 5525 8260 5559
rect 8208 5516 8260 5525
rect 11704 5516 11756 5568
rect 12164 5516 12216 5568
rect 13452 5516 13504 5568
rect 13820 5516 13872 5568
rect 15108 5516 15160 5568
rect 16856 5652 16908 5704
rect 17500 5695 17552 5704
rect 17500 5661 17509 5695
rect 17509 5661 17543 5695
rect 17543 5661 17552 5695
rect 17500 5652 17552 5661
rect 16672 5584 16724 5636
rect 17224 5584 17276 5636
rect 16856 5516 16908 5568
rect 17040 5559 17092 5568
rect 17040 5525 17049 5559
rect 17049 5525 17083 5559
rect 17083 5525 17092 5559
rect 17040 5516 17092 5525
rect 17776 5652 17828 5704
rect 17684 5584 17736 5636
rect 18328 5584 18380 5636
rect 18236 5516 18288 5568
rect 3110 5414 3162 5466
rect 3174 5414 3226 5466
rect 3238 5414 3290 5466
rect 3302 5414 3354 5466
rect 3366 5414 3418 5466
rect 6210 5414 6262 5466
rect 6274 5414 6326 5466
rect 6338 5414 6390 5466
rect 6402 5414 6454 5466
rect 6466 5414 6518 5466
rect 9310 5414 9362 5466
rect 9374 5414 9426 5466
rect 9438 5414 9490 5466
rect 9502 5414 9554 5466
rect 9566 5414 9618 5466
rect 12410 5414 12462 5466
rect 12474 5414 12526 5466
rect 12538 5414 12590 5466
rect 12602 5414 12654 5466
rect 12666 5414 12718 5466
rect 15510 5414 15562 5466
rect 15574 5414 15626 5466
rect 15638 5414 15690 5466
rect 15702 5414 15754 5466
rect 15766 5414 15818 5466
rect 18610 5414 18662 5466
rect 18674 5414 18726 5466
rect 18738 5414 18790 5466
rect 18802 5414 18854 5466
rect 18866 5414 18918 5466
rect 1952 5312 2004 5364
rect 5632 5312 5684 5364
rect 6552 5312 6604 5364
rect 7196 5312 7248 5364
rect 7840 5312 7892 5364
rect 8484 5312 8536 5364
rect 8852 5355 8904 5364
rect 8852 5321 8861 5355
rect 8861 5321 8895 5355
rect 8895 5321 8904 5355
rect 8852 5312 8904 5321
rect 7748 5244 7800 5296
rect 10232 5312 10284 5364
rect 13176 5312 13228 5364
rect 1492 5176 1544 5228
rect 3884 5219 3936 5228
rect 3884 5185 3893 5219
rect 3893 5185 3927 5219
rect 3927 5185 3936 5219
rect 3884 5176 3936 5185
rect 4160 5176 4212 5228
rect 6736 5219 6788 5228
rect 4252 5151 4304 5160
rect 4252 5117 4261 5151
rect 4261 5117 4295 5151
rect 4295 5117 4304 5151
rect 4252 5108 4304 5117
rect 6736 5185 6745 5219
rect 6745 5185 6779 5219
rect 6779 5185 6788 5219
rect 6736 5176 6788 5185
rect 7012 5176 7064 5228
rect 6000 5151 6052 5160
rect 6000 5117 6009 5151
rect 6009 5117 6043 5151
rect 6043 5117 6052 5151
rect 6000 5108 6052 5117
rect 6092 5108 6144 5160
rect 7288 5108 7340 5160
rect 8116 5176 8168 5228
rect 8852 5176 8904 5228
rect 9220 5176 9272 5228
rect 9588 5176 9640 5228
rect 14740 5244 14792 5296
rect 9036 5151 9088 5160
rect 2964 5083 3016 5092
rect 2964 5049 2973 5083
rect 2973 5049 3007 5083
rect 3007 5049 3016 5083
rect 2964 5040 3016 5049
rect 5356 5040 5408 5092
rect 3608 4972 3660 5024
rect 5172 4972 5224 5024
rect 5540 5040 5592 5092
rect 7012 5040 7064 5092
rect 7104 5040 7156 5092
rect 8208 5083 8260 5092
rect 8208 5049 8217 5083
rect 8217 5049 8251 5083
rect 8251 5049 8260 5083
rect 8208 5040 8260 5049
rect 6828 4972 6880 5024
rect 7288 5015 7340 5024
rect 7288 4981 7297 5015
rect 7297 4981 7331 5015
rect 7331 4981 7340 5015
rect 7288 4972 7340 4981
rect 7380 4972 7432 5024
rect 7932 4972 7984 5024
rect 9036 5117 9045 5151
rect 9045 5117 9079 5151
rect 9079 5117 9088 5151
rect 9036 5108 9088 5117
rect 14372 5176 14424 5228
rect 14464 5176 14516 5228
rect 16120 5312 16172 5364
rect 16488 5244 16540 5296
rect 17132 5244 17184 5296
rect 17500 5312 17552 5364
rect 17868 5312 17920 5364
rect 12900 5151 12952 5160
rect 12900 5117 12909 5151
rect 12909 5117 12943 5151
rect 12943 5117 12952 5151
rect 12900 5108 12952 5117
rect 13084 5151 13136 5160
rect 13084 5117 13093 5151
rect 13093 5117 13127 5151
rect 13127 5117 13136 5151
rect 13452 5151 13504 5160
rect 13084 5108 13136 5117
rect 13452 5117 13461 5151
rect 13461 5117 13495 5151
rect 13495 5117 13504 5151
rect 13452 5108 13504 5117
rect 10692 5040 10744 5092
rect 12256 5040 12308 5092
rect 12440 5040 12492 5092
rect 13820 5040 13872 5092
rect 15200 5108 15252 5160
rect 15568 5151 15620 5160
rect 15568 5117 15577 5151
rect 15577 5117 15611 5151
rect 15611 5117 15620 5151
rect 15568 5108 15620 5117
rect 16672 5176 16724 5228
rect 16856 5151 16908 5160
rect 16856 5117 16865 5151
rect 16865 5117 16899 5151
rect 16899 5117 16908 5151
rect 16856 5108 16908 5117
rect 15016 5040 15068 5092
rect 15844 5040 15896 5092
rect 17040 5040 17092 5092
rect 17224 5151 17276 5160
rect 17224 5117 17233 5151
rect 17233 5117 17267 5151
rect 17267 5117 17276 5151
rect 17592 5176 17644 5228
rect 17776 5219 17828 5228
rect 17776 5185 17785 5219
rect 17785 5185 17819 5219
rect 17819 5185 17828 5219
rect 17776 5176 17828 5185
rect 17684 5151 17736 5160
rect 17224 5108 17276 5117
rect 17684 5117 17693 5151
rect 17693 5117 17727 5151
rect 17727 5117 17736 5151
rect 17684 5108 17736 5117
rect 18052 5108 18104 5160
rect 17316 5040 17368 5092
rect 17592 5040 17644 5092
rect 18144 5040 18196 5092
rect 19156 5040 19208 5092
rect 9864 4972 9916 5024
rect 10784 4972 10836 5024
rect 11428 4972 11480 5024
rect 12164 4972 12216 5024
rect 13360 4972 13412 5024
rect 15200 5015 15252 5024
rect 15200 4981 15209 5015
rect 15209 4981 15243 5015
rect 15243 4981 15252 5015
rect 15200 4972 15252 4981
rect 17408 4972 17460 5024
rect 18420 5015 18472 5024
rect 18420 4981 18429 5015
rect 18429 4981 18463 5015
rect 18463 4981 18472 5015
rect 18420 4972 18472 4981
rect 4660 4870 4712 4922
rect 4724 4870 4776 4922
rect 4788 4870 4840 4922
rect 4852 4870 4904 4922
rect 4916 4870 4968 4922
rect 7760 4870 7812 4922
rect 7824 4870 7876 4922
rect 7888 4870 7940 4922
rect 7952 4870 8004 4922
rect 8016 4870 8068 4922
rect 10860 4870 10912 4922
rect 10924 4870 10976 4922
rect 10988 4870 11040 4922
rect 11052 4870 11104 4922
rect 11116 4870 11168 4922
rect 13960 4870 14012 4922
rect 14024 4870 14076 4922
rect 14088 4870 14140 4922
rect 14152 4870 14204 4922
rect 14216 4870 14268 4922
rect 17060 4870 17112 4922
rect 17124 4870 17176 4922
rect 17188 4870 17240 4922
rect 17252 4870 17304 4922
rect 17316 4870 17368 4922
rect 2504 4768 2556 4820
rect 2964 4811 3016 4820
rect 2964 4777 2973 4811
rect 2973 4777 3007 4811
rect 3007 4777 3016 4811
rect 2964 4768 3016 4777
rect 4252 4768 4304 4820
rect 6552 4768 6604 4820
rect 2504 4632 2556 4684
rect 3516 4700 3568 4752
rect 4712 4700 4764 4752
rect 5356 4700 5408 4752
rect 6644 4700 6696 4752
rect 7012 4768 7064 4820
rect 7748 4768 7800 4820
rect 7656 4700 7708 4752
rect 7932 4743 7984 4752
rect 7932 4709 7941 4743
rect 7941 4709 7975 4743
rect 7975 4709 7984 4743
rect 7932 4700 7984 4709
rect 8668 4768 8720 4820
rect 9036 4768 9088 4820
rect 9956 4768 10008 4820
rect 11428 4768 11480 4820
rect 12440 4768 12492 4820
rect 12992 4768 13044 4820
rect 14648 4811 14700 4820
rect 4988 4564 5040 4616
rect 5264 4632 5316 4684
rect 5908 4632 5960 4684
rect 6092 4675 6144 4684
rect 6092 4641 6101 4675
rect 6101 4641 6135 4675
rect 6135 4641 6144 4675
rect 6092 4632 6144 4641
rect 6552 4632 6604 4684
rect 5264 4539 5316 4548
rect 2964 4428 3016 4480
rect 5264 4505 5273 4539
rect 5273 4505 5307 4539
rect 5307 4505 5316 4539
rect 5264 4496 5316 4505
rect 5448 4496 5500 4548
rect 5724 4539 5776 4548
rect 5724 4505 5733 4539
rect 5733 4505 5767 4539
rect 5767 4505 5776 4539
rect 5724 4496 5776 4505
rect 6000 4607 6052 4616
rect 6000 4573 6009 4607
rect 6009 4573 6043 4607
rect 6043 4573 6052 4607
rect 7196 4632 7248 4684
rect 8484 4700 8536 4752
rect 6000 4564 6052 4573
rect 7656 4496 7708 4548
rect 8484 4564 8536 4616
rect 8852 4632 8904 4684
rect 9220 4632 9272 4684
rect 9588 4632 9640 4684
rect 12256 4700 12308 4752
rect 10232 4675 10284 4684
rect 10232 4641 10241 4675
rect 10241 4641 10275 4675
rect 10275 4641 10284 4675
rect 10232 4632 10284 4641
rect 8576 4496 8628 4548
rect 9864 4607 9916 4616
rect 9864 4573 9873 4607
rect 9873 4573 9907 4607
rect 9907 4573 9916 4607
rect 9864 4564 9916 4573
rect 10324 4607 10376 4616
rect 10324 4573 10333 4607
rect 10333 4573 10367 4607
rect 10367 4573 10376 4607
rect 10324 4564 10376 4573
rect 10600 4607 10652 4616
rect 10600 4573 10609 4607
rect 10609 4573 10643 4607
rect 10643 4573 10652 4607
rect 10600 4564 10652 4573
rect 11060 4564 11112 4616
rect 12624 4675 12676 4684
rect 12624 4641 12633 4675
rect 12633 4641 12667 4675
rect 12667 4641 12676 4675
rect 12624 4632 12676 4641
rect 14648 4777 14657 4811
rect 14657 4777 14691 4811
rect 14691 4777 14700 4811
rect 14648 4768 14700 4777
rect 14556 4700 14608 4752
rect 16856 4768 16908 4820
rect 17592 4768 17644 4820
rect 17960 4768 18012 4820
rect 15752 4743 15804 4752
rect 15752 4709 15770 4743
rect 15770 4709 15804 4743
rect 16120 4743 16172 4752
rect 15752 4700 15804 4709
rect 16120 4709 16129 4743
rect 16129 4709 16163 4743
rect 16163 4709 16172 4743
rect 16120 4700 16172 4709
rect 14464 4632 14516 4684
rect 13728 4564 13780 4616
rect 16580 4632 16632 4684
rect 17224 4675 17276 4684
rect 17224 4641 17233 4675
rect 17233 4641 17267 4675
rect 17267 4641 17276 4675
rect 17224 4632 17276 4641
rect 16212 4564 16264 4616
rect 16672 4564 16724 4616
rect 18144 4675 18196 4684
rect 18144 4641 18153 4675
rect 18153 4641 18187 4675
rect 18187 4641 18196 4675
rect 18144 4632 18196 4641
rect 18328 4675 18380 4684
rect 18328 4641 18337 4675
rect 18337 4641 18371 4675
rect 18371 4641 18380 4675
rect 18328 4632 18380 4641
rect 19064 4564 19116 4616
rect 5816 4428 5868 4480
rect 6092 4428 6144 4480
rect 10140 4428 10192 4480
rect 11888 4428 11940 4480
rect 11980 4428 12032 4480
rect 13084 4428 13136 4480
rect 13728 4428 13780 4480
rect 14464 4471 14516 4480
rect 14464 4437 14473 4471
rect 14473 4437 14507 4471
rect 14507 4437 14516 4471
rect 14464 4428 14516 4437
rect 14648 4428 14700 4480
rect 14924 4428 14976 4480
rect 15844 4428 15896 4480
rect 17592 4496 17644 4548
rect 18236 4496 18288 4548
rect 17316 4471 17368 4480
rect 17316 4437 17325 4471
rect 17325 4437 17359 4471
rect 17359 4437 17368 4471
rect 17316 4428 17368 4437
rect 17408 4428 17460 4480
rect 3110 4326 3162 4378
rect 3174 4326 3226 4378
rect 3238 4326 3290 4378
rect 3302 4326 3354 4378
rect 3366 4326 3418 4378
rect 6210 4326 6262 4378
rect 6274 4326 6326 4378
rect 6338 4326 6390 4378
rect 6402 4326 6454 4378
rect 6466 4326 6518 4378
rect 9310 4326 9362 4378
rect 9374 4326 9426 4378
rect 9438 4326 9490 4378
rect 9502 4326 9554 4378
rect 9566 4326 9618 4378
rect 12410 4326 12462 4378
rect 12474 4326 12526 4378
rect 12538 4326 12590 4378
rect 12602 4326 12654 4378
rect 12666 4326 12718 4378
rect 15510 4326 15562 4378
rect 15574 4326 15626 4378
rect 15638 4326 15690 4378
rect 15702 4326 15754 4378
rect 15766 4326 15818 4378
rect 18610 4326 18662 4378
rect 18674 4326 18726 4378
rect 18738 4326 18790 4378
rect 18802 4326 18854 4378
rect 18866 4326 18918 4378
rect 1124 4224 1176 4276
rect 6000 4224 6052 4276
rect 6736 4224 6788 4276
rect 4712 4156 4764 4208
rect 3608 4020 3660 4072
rect 4344 4088 4396 4140
rect 4988 4131 5040 4140
rect 4988 4097 4997 4131
rect 4997 4097 5031 4131
rect 5031 4097 5040 4131
rect 4988 4088 5040 4097
rect 4160 4020 4212 4072
rect 5172 4020 5224 4072
rect 2228 3995 2280 4004
rect 2228 3961 2237 3995
rect 2237 3961 2271 3995
rect 2271 3961 2280 3995
rect 2228 3952 2280 3961
rect 5908 4088 5960 4140
rect 6184 4088 6236 4140
rect 2504 3884 2556 3936
rect 2596 3884 2648 3936
rect 4344 3927 4396 3936
rect 4344 3893 4353 3927
rect 4353 3893 4387 3927
rect 4387 3893 4396 3927
rect 4344 3884 4396 3893
rect 4528 3884 4580 3936
rect 5080 3884 5132 3936
rect 6092 3952 6144 4004
rect 5264 3884 5316 3936
rect 6644 4088 6696 4140
rect 6828 4088 6880 4140
rect 7196 4088 7248 4140
rect 6552 3952 6604 4004
rect 9220 4224 9272 4276
rect 8300 4156 8352 4208
rect 7748 4063 7800 4072
rect 7748 4029 7757 4063
rect 7757 4029 7791 4063
rect 7791 4029 7800 4063
rect 7748 4020 7800 4029
rect 7932 4063 7984 4072
rect 7932 4029 7941 4063
rect 7941 4029 7975 4063
rect 7975 4029 7984 4063
rect 7932 4020 7984 4029
rect 8024 4063 8076 4072
rect 8024 4029 8033 4063
rect 8033 4029 8067 4063
rect 8067 4029 8076 4063
rect 8024 4020 8076 4029
rect 8300 4063 8352 4072
rect 8300 4029 8309 4063
rect 8309 4029 8343 4063
rect 8343 4029 8352 4063
rect 8944 4088 8996 4140
rect 8300 4020 8352 4029
rect 8668 4063 8720 4072
rect 8668 4029 8677 4063
rect 8677 4029 8711 4063
rect 8711 4029 8720 4063
rect 8668 4020 8720 4029
rect 9036 4063 9088 4072
rect 9036 4029 9045 4063
rect 9045 4029 9079 4063
rect 9079 4029 9088 4063
rect 9036 4020 9088 4029
rect 10600 4224 10652 4276
rect 15844 4224 15896 4276
rect 17960 4224 18012 4276
rect 11428 4131 11480 4140
rect 11428 4097 11437 4131
rect 11437 4097 11471 4131
rect 11471 4097 11480 4131
rect 11428 4088 11480 4097
rect 13452 4131 13504 4140
rect 13452 4097 13461 4131
rect 13461 4097 13495 4131
rect 13495 4097 13504 4131
rect 13452 4088 13504 4097
rect 13728 4088 13780 4140
rect 17224 4156 17276 4208
rect 17776 4156 17828 4208
rect 18052 4199 18104 4208
rect 18052 4165 18061 4199
rect 18061 4165 18095 4199
rect 18095 4165 18104 4199
rect 18052 4156 18104 4165
rect 10784 4063 10836 4072
rect 10784 4029 10793 4063
rect 10793 4029 10827 4063
rect 10827 4029 10836 4063
rect 10784 4020 10836 4029
rect 11060 4063 11112 4072
rect 11060 4029 11069 4063
rect 11069 4029 11103 4063
rect 11103 4029 11112 4063
rect 11060 4020 11112 4029
rect 11336 4020 11388 4072
rect 11888 4020 11940 4072
rect 14924 4088 14976 4140
rect 16120 4088 16172 4140
rect 16580 4088 16632 4140
rect 16764 4088 16816 4140
rect 18236 4131 18288 4140
rect 6736 3884 6788 3936
rect 9772 3952 9824 4004
rect 8116 3884 8168 3936
rect 8208 3884 8260 3936
rect 8392 3927 8444 3936
rect 8392 3893 8401 3927
rect 8401 3893 8435 3927
rect 8435 3893 8444 3927
rect 8392 3884 8444 3893
rect 8576 3884 8628 3936
rect 12992 3952 13044 4004
rect 15016 3952 15068 4004
rect 15200 4020 15252 4072
rect 18236 4097 18245 4131
rect 18245 4097 18279 4131
rect 18279 4097 18288 4131
rect 18236 4088 18288 4097
rect 18604 4088 18656 4140
rect 16120 3952 16172 4004
rect 16580 3952 16632 4004
rect 18052 4020 18104 4072
rect 18512 4063 18564 4072
rect 18512 4029 18521 4063
rect 18521 4029 18555 4063
rect 18555 4029 18564 4063
rect 18512 4020 18564 4029
rect 10784 3884 10836 3936
rect 15200 3884 15252 3936
rect 15936 3884 15988 3936
rect 16488 3884 16540 3936
rect 17132 3884 17184 3936
rect 17684 3884 17736 3936
rect 18236 3927 18288 3936
rect 18236 3893 18245 3927
rect 18245 3893 18279 3927
rect 18279 3893 18288 3927
rect 18236 3884 18288 3893
rect 4660 3782 4712 3834
rect 4724 3782 4776 3834
rect 4788 3782 4840 3834
rect 4852 3782 4904 3834
rect 4916 3782 4968 3834
rect 7760 3782 7812 3834
rect 7824 3782 7876 3834
rect 7888 3782 7940 3834
rect 7952 3782 8004 3834
rect 8016 3782 8068 3834
rect 10860 3782 10912 3834
rect 10924 3782 10976 3834
rect 10988 3782 11040 3834
rect 11052 3782 11104 3834
rect 11116 3782 11168 3834
rect 13960 3782 14012 3834
rect 14024 3782 14076 3834
rect 14088 3782 14140 3834
rect 14152 3782 14204 3834
rect 14216 3782 14268 3834
rect 17060 3782 17112 3834
rect 17124 3782 17176 3834
rect 17188 3782 17240 3834
rect 17252 3782 17304 3834
rect 17316 3782 17368 3834
rect 2228 3680 2280 3732
rect 4252 3680 4304 3732
rect 5080 3680 5132 3732
rect 3608 3612 3660 3664
rect 4436 3612 4488 3664
rect 4988 3612 5040 3664
rect 5356 3612 5408 3664
rect 2596 3544 2648 3596
rect 4896 3587 4948 3596
rect 4896 3553 4905 3587
rect 4905 3553 4939 3587
rect 4939 3553 4948 3587
rect 4896 3544 4948 3553
rect 5172 3587 5224 3596
rect 5172 3553 5181 3587
rect 5181 3553 5215 3587
rect 5215 3553 5224 3587
rect 5172 3544 5224 3553
rect 5816 3544 5868 3596
rect 2504 3476 2556 3528
rect 2964 3519 3016 3528
rect 2964 3485 2973 3519
rect 2973 3485 3007 3519
rect 3007 3485 3016 3519
rect 2964 3476 3016 3485
rect 5540 3519 5592 3528
rect 5540 3485 5549 3519
rect 5549 3485 5583 3519
rect 5583 3485 5592 3519
rect 5540 3476 5592 3485
rect 6092 3476 6144 3528
rect 6552 3587 6604 3596
rect 6552 3553 6561 3587
rect 6561 3553 6595 3587
rect 6595 3553 6604 3587
rect 6552 3544 6604 3553
rect 6736 3544 6788 3596
rect 7196 3544 7248 3596
rect 7748 3587 7800 3596
rect 7748 3553 7757 3587
rect 7757 3553 7791 3587
rect 7791 3553 7800 3587
rect 7748 3544 7800 3553
rect 7932 3587 7984 3596
rect 7932 3553 7956 3587
rect 7956 3553 7984 3587
rect 7932 3544 7984 3553
rect 8116 3680 8168 3732
rect 8208 3680 8260 3732
rect 8300 3612 8352 3664
rect 8668 3680 8720 3732
rect 10048 3680 10100 3732
rect 13452 3680 13504 3732
rect 13820 3680 13872 3732
rect 14004 3680 14056 3732
rect 8760 3655 8812 3664
rect 8760 3621 8769 3655
rect 8769 3621 8803 3655
rect 8803 3621 8812 3655
rect 8760 3612 8812 3621
rect 9128 3612 9180 3664
rect 12900 3612 12952 3664
rect 14832 3723 14884 3732
rect 14832 3689 14841 3723
rect 14841 3689 14875 3723
rect 14875 3689 14884 3723
rect 14832 3680 14884 3689
rect 15200 3680 15252 3732
rect 8852 3587 8904 3596
rect 6644 3476 6696 3528
rect 7288 3476 7340 3528
rect 6000 3408 6052 3460
rect 7104 3408 7156 3460
rect 2872 3340 2924 3392
rect 4068 3340 4120 3392
rect 4620 3340 4672 3392
rect 4988 3340 5040 3392
rect 5264 3383 5316 3392
rect 5264 3349 5273 3383
rect 5273 3349 5307 3383
rect 5307 3349 5316 3383
rect 5264 3340 5316 3349
rect 5908 3383 5960 3392
rect 5908 3349 5917 3383
rect 5917 3349 5951 3383
rect 5951 3349 5960 3383
rect 5908 3340 5960 3349
rect 6828 3340 6880 3392
rect 7656 3340 7708 3392
rect 8024 3383 8076 3392
rect 8024 3349 8033 3383
rect 8033 3349 8067 3383
rect 8067 3349 8076 3383
rect 8024 3340 8076 3349
rect 8116 3340 8168 3392
rect 8852 3553 8861 3587
rect 8861 3553 8895 3587
rect 8895 3553 8904 3587
rect 8852 3544 8904 3553
rect 8944 3544 8996 3596
rect 9772 3544 9824 3596
rect 9956 3587 10008 3596
rect 9956 3553 9965 3587
rect 9965 3553 9999 3587
rect 9999 3553 10008 3587
rect 9956 3544 10008 3553
rect 11612 3544 11664 3596
rect 13084 3587 13136 3596
rect 13084 3553 13093 3587
rect 13093 3553 13127 3587
rect 13127 3553 13136 3587
rect 13084 3544 13136 3553
rect 17132 3612 17184 3664
rect 8760 3476 8812 3528
rect 10692 3476 10744 3528
rect 12164 3476 12216 3528
rect 12992 3476 13044 3528
rect 13544 3476 13596 3528
rect 13820 3587 13872 3596
rect 13820 3553 13829 3587
rect 13829 3553 13863 3587
rect 13863 3553 13872 3587
rect 13820 3544 13872 3553
rect 14188 3587 14240 3596
rect 14188 3553 14197 3587
rect 14197 3553 14231 3587
rect 14231 3553 14240 3587
rect 14188 3544 14240 3553
rect 14372 3476 14424 3528
rect 14648 3519 14700 3528
rect 14648 3485 14657 3519
rect 14657 3485 14691 3519
rect 14691 3485 14700 3519
rect 14648 3476 14700 3485
rect 8484 3383 8536 3392
rect 8484 3349 8493 3383
rect 8493 3349 8527 3383
rect 8527 3349 8536 3383
rect 8484 3340 8536 3349
rect 8576 3340 8628 3392
rect 13728 3408 13780 3460
rect 13820 3408 13872 3460
rect 15936 3587 15988 3596
rect 15936 3553 15954 3587
rect 15954 3553 15988 3587
rect 16212 3587 16264 3596
rect 15936 3544 15988 3553
rect 16212 3553 16221 3587
rect 16221 3553 16255 3587
rect 16255 3553 16264 3587
rect 16212 3544 16264 3553
rect 16488 3587 16540 3596
rect 16488 3553 16497 3587
rect 16497 3553 16531 3587
rect 16531 3553 16540 3587
rect 16488 3544 16540 3553
rect 19064 3680 19116 3732
rect 17684 3587 17736 3596
rect 17684 3553 17693 3587
rect 17693 3553 17727 3587
rect 17727 3553 17736 3587
rect 17684 3544 17736 3553
rect 18236 3612 18288 3664
rect 18420 3544 18472 3596
rect 18880 3544 18932 3596
rect 17224 3519 17276 3528
rect 17224 3485 17233 3519
rect 17233 3485 17267 3519
rect 17267 3485 17276 3519
rect 17224 3476 17276 3485
rect 17500 3476 17552 3528
rect 18604 3476 18656 3528
rect 16212 3408 16264 3460
rect 16304 3408 16356 3460
rect 16488 3408 16540 3460
rect 17960 3408 18012 3460
rect 18420 3408 18472 3460
rect 9128 3383 9180 3392
rect 9128 3349 9137 3383
rect 9137 3349 9171 3383
rect 9171 3349 9180 3383
rect 9128 3340 9180 3349
rect 9220 3340 9272 3392
rect 12072 3340 12124 3392
rect 12256 3340 12308 3392
rect 12992 3340 13044 3392
rect 13452 3340 13504 3392
rect 13912 3340 13964 3392
rect 14096 3340 14148 3392
rect 14832 3340 14884 3392
rect 16672 3340 16724 3392
rect 17776 3340 17828 3392
rect 3110 3238 3162 3290
rect 3174 3238 3226 3290
rect 3238 3238 3290 3290
rect 3302 3238 3354 3290
rect 3366 3238 3418 3290
rect 6210 3238 6262 3290
rect 6274 3238 6326 3290
rect 6338 3238 6390 3290
rect 6402 3238 6454 3290
rect 6466 3238 6518 3290
rect 9310 3238 9362 3290
rect 9374 3238 9426 3290
rect 9438 3238 9490 3290
rect 9502 3238 9554 3290
rect 9566 3238 9618 3290
rect 12410 3238 12462 3290
rect 12474 3238 12526 3290
rect 12538 3238 12590 3290
rect 12602 3238 12654 3290
rect 12666 3238 12718 3290
rect 15510 3238 15562 3290
rect 15574 3238 15626 3290
rect 15638 3238 15690 3290
rect 15702 3238 15754 3290
rect 15766 3238 15818 3290
rect 18610 3238 18662 3290
rect 18674 3238 18726 3290
rect 18738 3238 18790 3290
rect 18802 3238 18854 3290
rect 18866 3238 18918 3290
rect 2964 3136 3016 3188
rect 4068 3136 4120 3188
rect 2780 3000 2832 3052
rect 4344 3043 4396 3052
rect 4344 3009 4353 3043
rect 4353 3009 4387 3043
rect 4387 3009 4396 3043
rect 4344 3000 4396 3009
rect 7472 3179 7524 3188
rect 7472 3145 7481 3179
rect 7481 3145 7515 3179
rect 7515 3145 7524 3179
rect 7472 3136 7524 3145
rect 7564 3136 7616 3188
rect 6460 3068 6512 3120
rect 6736 3068 6788 3120
rect 6092 3000 6144 3052
rect 7380 3111 7432 3120
rect 7380 3077 7389 3111
rect 7389 3077 7423 3111
rect 7423 3077 7432 3111
rect 7380 3068 7432 3077
rect 1860 2975 1912 2984
rect 1860 2941 1869 2975
rect 1869 2941 1903 2975
rect 1903 2941 1912 2975
rect 1860 2932 1912 2941
rect 3608 2932 3660 2984
rect 4252 2975 4304 2984
rect 4252 2941 4261 2975
rect 4261 2941 4295 2975
rect 4295 2941 4304 2975
rect 4252 2932 4304 2941
rect 4620 2932 4672 2984
rect 6000 2932 6052 2984
rect 8484 3136 8536 3188
rect 9220 3136 9272 3188
rect 7932 3068 7984 3120
rect 8300 3068 8352 3120
rect 8116 3000 8168 3052
rect 8668 3000 8720 3052
rect 8944 3000 8996 3052
rect 9588 3000 9640 3052
rect 3700 2907 3752 2916
rect 3700 2873 3709 2907
rect 3709 2873 3743 2907
rect 3743 2873 3752 2907
rect 3700 2864 3752 2873
rect 1400 2796 1452 2848
rect 4804 2864 4856 2916
rect 4896 2864 4948 2916
rect 6092 2907 6144 2916
rect 4344 2796 4396 2848
rect 5080 2839 5132 2848
rect 5080 2805 5089 2839
rect 5089 2805 5123 2839
rect 5123 2805 5132 2839
rect 5080 2796 5132 2805
rect 5356 2796 5408 2848
rect 6092 2873 6101 2907
rect 6101 2873 6135 2907
rect 6135 2873 6144 2907
rect 6092 2864 6144 2873
rect 7012 2864 7064 2916
rect 7196 2864 7248 2916
rect 7472 2932 7524 2984
rect 7748 2975 7800 2984
rect 7748 2941 7757 2975
rect 7757 2941 7791 2975
rect 7791 2941 7800 2975
rect 7748 2932 7800 2941
rect 7840 2932 7892 2984
rect 8392 2975 8444 2984
rect 8392 2941 8401 2975
rect 8401 2941 8435 2975
rect 8435 2941 8444 2975
rect 8392 2932 8444 2941
rect 8576 2932 8628 2984
rect 8300 2864 8352 2916
rect 8852 2864 8904 2916
rect 9312 2932 9364 2984
rect 11244 3136 11296 3188
rect 11336 3136 11388 3188
rect 13452 3136 13504 3188
rect 14004 3136 14056 3188
rect 17132 3136 17184 3188
rect 17500 3136 17552 3188
rect 17868 3136 17920 3188
rect 18052 3179 18104 3188
rect 18052 3145 18061 3179
rect 18061 3145 18095 3179
rect 18095 3145 18104 3179
rect 18052 3136 18104 3145
rect 15292 3068 15344 3120
rect 15752 3068 15804 3120
rect 17316 3068 17368 3120
rect 10140 2932 10192 2984
rect 10508 3000 10560 3052
rect 12992 3000 13044 3052
rect 10784 2932 10836 2984
rect 11980 2932 12032 2984
rect 12716 2932 12768 2984
rect 6736 2796 6788 2848
rect 7472 2796 7524 2848
rect 7932 2796 7984 2848
rect 8668 2796 8720 2848
rect 12256 2864 12308 2916
rect 13452 2975 13504 2984
rect 13452 2941 13461 2975
rect 13461 2941 13495 2975
rect 13495 2941 13504 2975
rect 13452 2932 13504 2941
rect 14096 3000 14148 3052
rect 14924 3000 14976 3052
rect 17408 3000 17460 3052
rect 13820 2975 13872 2984
rect 13820 2941 13829 2975
rect 13829 2941 13863 2975
rect 13863 2941 13872 2975
rect 13820 2932 13872 2941
rect 14188 2975 14240 2984
rect 14188 2941 14197 2975
rect 14197 2941 14231 2975
rect 14231 2941 14240 2975
rect 14188 2932 14240 2941
rect 17592 2932 17644 2984
rect 17868 2975 17920 2984
rect 17868 2941 17877 2975
rect 17877 2941 17911 2975
rect 17911 2941 17920 2975
rect 17868 2932 17920 2941
rect 10600 2839 10652 2848
rect 10600 2805 10609 2839
rect 10609 2805 10643 2839
rect 10643 2805 10652 2839
rect 10600 2796 10652 2805
rect 11244 2796 11296 2848
rect 11612 2796 11664 2848
rect 13268 2864 13320 2916
rect 14556 2864 14608 2916
rect 18972 2932 19024 2984
rect 13912 2796 13964 2848
rect 15108 2796 15160 2848
rect 15844 2796 15896 2848
rect 15936 2796 15988 2848
rect 17776 2796 17828 2848
rect 4660 2694 4712 2746
rect 4724 2694 4776 2746
rect 4788 2694 4840 2746
rect 4852 2694 4904 2746
rect 4916 2694 4968 2746
rect 7760 2694 7812 2746
rect 7824 2694 7876 2746
rect 7888 2694 7940 2746
rect 7952 2694 8004 2746
rect 8016 2694 8068 2746
rect 10860 2694 10912 2746
rect 10924 2694 10976 2746
rect 10988 2694 11040 2746
rect 11052 2694 11104 2746
rect 11116 2694 11168 2746
rect 13960 2694 14012 2746
rect 14024 2694 14076 2746
rect 14088 2694 14140 2746
rect 14152 2694 14204 2746
rect 14216 2694 14268 2746
rect 17060 2694 17112 2746
rect 17124 2694 17176 2746
rect 17188 2694 17240 2746
rect 17252 2694 17304 2746
rect 17316 2694 17368 2746
rect 2780 2592 2832 2644
rect 4344 2592 4396 2644
rect 5540 2592 5592 2644
rect 6184 2592 6236 2644
rect 6460 2592 6512 2644
rect 7196 2592 7248 2644
rect 1860 2524 1912 2576
rect 2504 2456 2556 2508
rect 3700 2456 3752 2508
rect 3792 2431 3844 2440
rect 2872 2320 2924 2372
rect 3792 2397 3801 2431
rect 3801 2397 3835 2431
rect 3835 2397 3844 2431
rect 3792 2388 3844 2397
rect 4252 2456 4304 2508
rect 6000 2524 6052 2576
rect 5172 2456 5224 2508
rect 5724 2499 5776 2508
rect 5724 2465 5733 2499
rect 5733 2465 5767 2499
rect 5767 2465 5776 2499
rect 5724 2456 5776 2465
rect 6092 2499 6144 2508
rect 6092 2465 6101 2499
rect 6101 2465 6135 2499
rect 6135 2465 6144 2499
rect 6092 2456 6144 2465
rect 8760 2592 8812 2644
rect 9036 2592 9088 2644
rect 10600 2592 10652 2644
rect 12164 2592 12216 2644
rect 12256 2592 12308 2644
rect 14280 2592 14332 2644
rect 9772 2524 9824 2576
rect 13544 2524 13596 2576
rect 13912 2524 13964 2576
rect 14648 2567 14700 2576
rect 14648 2533 14657 2567
rect 14657 2533 14691 2567
rect 14691 2533 14700 2567
rect 14648 2524 14700 2533
rect 19156 2592 19208 2644
rect 16856 2524 16908 2576
rect 17132 2524 17184 2576
rect 9128 2456 9180 2508
rect 9588 2499 9640 2508
rect 7380 2388 7432 2440
rect 7748 2431 7800 2440
rect 5080 2320 5132 2372
rect 7288 2320 7340 2372
rect 7748 2397 7757 2431
rect 7757 2397 7791 2431
rect 7791 2397 7800 2431
rect 7748 2388 7800 2397
rect 8852 2320 8904 2372
rect 8944 2320 8996 2372
rect 9588 2465 9597 2499
rect 9597 2465 9631 2499
rect 9631 2465 9640 2499
rect 9588 2456 9640 2465
rect 11612 2499 11664 2508
rect 11612 2465 11621 2499
rect 11621 2465 11655 2499
rect 11655 2465 11664 2499
rect 11612 2456 11664 2465
rect 14188 2499 14240 2508
rect 14188 2465 14197 2499
rect 14197 2465 14231 2499
rect 14231 2465 14240 2499
rect 14188 2456 14240 2465
rect 14740 2456 14792 2508
rect 14924 2499 14976 2508
rect 14924 2465 14933 2499
rect 14933 2465 14967 2499
rect 14967 2465 14976 2499
rect 14924 2456 14976 2465
rect 15200 2499 15252 2508
rect 9680 2388 9732 2440
rect 13728 2388 13780 2440
rect 15200 2465 15223 2499
rect 15223 2465 15252 2499
rect 15200 2456 15252 2465
rect 16672 2456 16724 2508
rect 17040 2456 17092 2508
rect 18052 2456 18104 2508
rect 17224 2388 17276 2440
rect 17592 2388 17644 2440
rect 17960 2388 18012 2440
rect 4804 2252 4856 2304
rect 5448 2295 5500 2304
rect 5448 2261 5457 2295
rect 5457 2261 5491 2295
rect 5491 2261 5500 2295
rect 5448 2252 5500 2261
rect 6552 2252 6604 2304
rect 12256 2320 12308 2372
rect 13820 2320 13872 2372
rect 14280 2320 14332 2372
rect 9772 2252 9824 2304
rect 11980 2295 12032 2304
rect 11980 2261 11989 2295
rect 11989 2261 12023 2295
rect 12023 2261 12032 2295
rect 11980 2252 12032 2261
rect 12900 2252 12952 2304
rect 14648 2252 14700 2304
rect 16672 2320 16724 2372
rect 16212 2252 16264 2304
rect 16396 2252 16448 2304
rect 17776 2295 17828 2304
rect 17776 2261 17785 2295
rect 17785 2261 17819 2295
rect 17819 2261 17828 2295
rect 17776 2252 17828 2261
rect 18052 2252 18104 2304
rect 18420 2252 18472 2304
rect 3110 2150 3162 2202
rect 3174 2150 3226 2202
rect 3238 2150 3290 2202
rect 3302 2150 3354 2202
rect 3366 2150 3418 2202
rect 6210 2150 6262 2202
rect 6274 2150 6326 2202
rect 6338 2150 6390 2202
rect 6402 2150 6454 2202
rect 6466 2150 6518 2202
rect 9310 2150 9362 2202
rect 9374 2150 9426 2202
rect 9438 2150 9490 2202
rect 9502 2150 9554 2202
rect 9566 2150 9618 2202
rect 12410 2150 12462 2202
rect 12474 2150 12526 2202
rect 12538 2150 12590 2202
rect 12602 2150 12654 2202
rect 12666 2150 12718 2202
rect 15510 2150 15562 2202
rect 15574 2150 15626 2202
rect 15638 2150 15690 2202
rect 15702 2150 15754 2202
rect 15766 2150 15818 2202
rect 18610 2150 18662 2202
rect 18674 2150 18726 2202
rect 18738 2150 18790 2202
rect 18802 2150 18854 2202
rect 18866 2150 18918 2202
rect 4528 2048 4580 2100
rect 7196 2048 7248 2100
rect 7656 2048 7708 2100
rect 8208 2048 8260 2100
rect 2504 1844 2556 1896
rect 5448 1980 5500 2032
rect 6092 1980 6144 2032
rect 6552 1980 6604 2032
rect 9220 2048 9272 2100
rect 9680 2048 9732 2100
rect 9864 2048 9916 2100
rect 2964 1819 3016 1828
rect 2964 1785 2973 1819
rect 2973 1785 3007 1819
rect 3007 1785 3016 1819
rect 2964 1776 3016 1785
rect 4436 1887 4488 1896
rect 4436 1853 4445 1887
rect 4445 1853 4479 1887
rect 4479 1853 4488 1887
rect 4436 1844 4488 1853
rect 4528 1776 4580 1828
rect 4804 1887 4856 1896
rect 4804 1853 4813 1887
rect 4813 1853 4847 1887
rect 4847 1853 4856 1887
rect 4804 1844 4856 1853
rect 4988 1887 5040 1896
rect 4988 1853 4997 1887
rect 4997 1853 5031 1887
rect 5031 1853 5040 1887
rect 4988 1844 5040 1853
rect 5264 1887 5316 1896
rect 5264 1853 5273 1887
rect 5273 1853 5307 1887
rect 5307 1853 5316 1887
rect 5264 1844 5316 1853
rect 5724 1887 5776 1896
rect 5724 1853 5733 1887
rect 5733 1853 5767 1887
rect 5767 1853 5776 1887
rect 6736 1955 6788 1964
rect 6736 1921 6745 1955
rect 6745 1921 6779 1955
rect 6779 1921 6788 1955
rect 6736 1912 6788 1921
rect 7012 1912 7064 1964
rect 5724 1844 5776 1853
rect 5172 1776 5224 1828
rect 7656 1844 7708 1896
rect 8852 1887 8904 1896
rect 8852 1853 8861 1887
rect 8861 1853 8895 1887
rect 8895 1853 8904 1887
rect 8852 1844 8904 1853
rect 9588 1980 9640 2032
rect 10048 1955 10100 1964
rect 10048 1921 10057 1955
rect 10057 1921 10091 1955
rect 10091 1921 10100 1955
rect 10048 1912 10100 1921
rect 5540 1708 5592 1760
rect 5816 1751 5868 1760
rect 5816 1717 5825 1751
rect 5825 1717 5859 1751
rect 5859 1717 5868 1751
rect 5816 1708 5868 1717
rect 7196 1708 7248 1760
rect 7472 1708 7524 1760
rect 9404 1844 9456 1896
rect 12256 2091 12308 2100
rect 12256 2057 12265 2091
rect 12265 2057 12299 2091
rect 12299 2057 12308 2091
rect 12256 2048 12308 2057
rect 16028 2048 16080 2100
rect 16304 2048 16356 2100
rect 17040 2091 17092 2100
rect 15844 1980 15896 2032
rect 17040 2057 17049 2091
rect 17049 2057 17083 2091
rect 17083 2057 17092 2091
rect 17040 2048 17092 2057
rect 18512 2091 18564 2100
rect 10784 1912 10836 1964
rect 13728 1912 13780 1964
rect 13820 1912 13872 1964
rect 14280 1955 14332 1964
rect 11888 1887 11940 1896
rect 11888 1853 11897 1887
rect 11897 1853 11931 1887
rect 11931 1853 11940 1887
rect 11888 1844 11940 1853
rect 12164 1887 12216 1896
rect 12164 1853 12173 1887
rect 12173 1853 12207 1887
rect 12207 1853 12216 1887
rect 12164 1844 12216 1853
rect 12348 1887 12400 1896
rect 12348 1853 12357 1887
rect 12357 1853 12391 1887
rect 12391 1853 12400 1887
rect 12348 1844 12400 1853
rect 12808 1887 12860 1896
rect 12808 1853 12817 1887
rect 12817 1853 12851 1887
rect 12851 1853 12860 1887
rect 12808 1844 12860 1853
rect 12992 1844 13044 1896
rect 14280 1921 14289 1955
rect 14289 1921 14323 1955
rect 14323 1921 14332 1955
rect 14280 1912 14332 1921
rect 16764 1912 16816 1964
rect 16856 1912 16908 1964
rect 17040 1912 17092 1964
rect 17592 1955 17644 1964
rect 9772 1776 9824 1828
rect 9036 1708 9088 1760
rect 13544 1776 13596 1828
rect 13912 1776 13964 1828
rect 14832 1844 14884 1896
rect 11428 1751 11480 1760
rect 11428 1717 11437 1751
rect 11437 1717 11471 1751
rect 11471 1717 11480 1751
rect 11428 1708 11480 1717
rect 13176 1708 13228 1760
rect 13820 1751 13872 1760
rect 13820 1717 13829 1751
rect 13829 1717 13863 1751
rect 13863 1717 13872 1751
rect 13820 1708 13872 1717
rect 14648 1776 14700 1828
rect 17132 1844 17184 1896
rect 17592 1921 17601 1955
rect 17601 1921 17635 1955
rect 17635 1921 17644 1955
rect 17592 1912 17644 1921
rect 15476 1776 15528 1828
rect 16304 1819 16356 1828
rect 16304 1785 16313 1819
rect 16313 1785 16347 1819
rect 16347 1785 16356 1819
rect 16304 1776 16356 1785
rect 16856 1776 16908 1828
rect 17224 1776 17276 1828
rect 14740 1708 14792 1760
rect 15660 1751 15712 1760
rect 15660 1717 15669 1751
rect 15669 1717 15703 1751
rect 15703 1717 15712 1751
rect 15660 1708 15712 1717
rect 15844 1751 15896 1760
rect 15844 1717 15853 1751
rect 15853 1717 15887 1751
rect 15887 1717 15896 1751
rect 15844 1708 15896 1717
rect 16212 1751 16264 1760
rect 16212 1717 16221 1751
rect 16221 1717 16255 1751
rect 16255 1717 16264 1751
rect 16212 1708 16264 1717
rect 17868 1887 17920 1896
rect 17868 1853 17877 1887
rect 17877 1853 17911 1887
rect 17911 1853 17920 1887
rect 18512 2057 18521 2091
rect 18521 2057 18555 2091
rect 18555 2057 18564 2091
rect 18512 2048 18564 2057
rect 17868 1844 17920 1853
rect 18512 1887 18564 1896
rect 18512 1853 18521 1887
rect 18521 1853 18555 1887
rect 18555 1853 18564 1887
rect 18512 1844 18564 1853
rect 4660 1606 4712 1658
rect 4724 1606 4776 1658
rect 4788 1606 4840 1658
rect 4852 1606 4904 1658
rect 4916 1606 4968 1658
rect 7760 1606 7812 1658
rect 7824 1606 7876 1658
rect 7888 1606 7940 1658
rect 7952 1606 8004 1658
rect 8016 1606 8068 1658
rect 10860 1606 10912 1658
rect 10924 1606 10976 1658
rect 10988 1606 11040 1658
rect 11052 1606 11104 1658
rect 11116 1606 11168 1658
rect 13960 1606 14012 1658
rect 14024 1606 14076 1658
rect 14088 1606 14140 1658
rect 14152 1606 14204 1658
rect 14216 1606 14268 1658
rect 17060 1606 17112 1658
rect 17124 1606 17176 1658
rect 17188 1606 17240 1658
rect 17252 1606 17304 1658
rect 17316 1606 17368 1658
rect 3516 1504 3568 1556
rect 4528 1504 4580 1556
rect 5172 1547 5224 1556
rect 5172 1513 5181 1547
rect 5181 1513 5215 1547
rect 5215 1513 5224 1547
rect 5172 1504 5224 1513
rect 6000 1504 6052 1556
rect 7564 1504 7616 1556
rect 7656 1504 7708 1556
rect 8300 1504 8352 1556
rect 7012 1436 7064 1488
rect 9864 1504 9916 1556
rect 10784 1504 10836 1556
rect 11428 1547 11480 1556
rect 11428 1513 11437 1547
rect 11437 1513 11471 1547
rect 11471 1513 11480 1547
rect 11428 1504 11480 1513
rect 11980 1547 12032 1556
rect 11980 1513 11989 1547
rect 11989 1513 12023 1547
rect 12023 1513 12032 1547
rect 11980 1504 12032 1513
rect 12348 1504 12400 1556
rect 13728 1547 13780 1556
rect 2964 1368 3016 1420
rect 6092 1411 6144 1420
rect 5816 1300 5868 1352
rect 6092 1377 6101 1411
rect 6101 1377 6135 1411
rect 6135 1377 6144 1411
rect 6092 1368 6144 1377
rect 8208 1368 8260 1420
rect 8300 1411 8352 1420
rect 8300 1377 8309 1411
rect 8309 1377 8343 1411
rect 8343 1377 8352 1411
rect 8300 1368 8352 1377
rect 10508 1436 10560 1488
rect 13728 1513 13737 1547
rect 13737 1513 13771 1547
rect 13771 1513 13780 1547
rect 13728 1504 13780 1513
rect 13820 1504 13872 1556
rect 14464 1547 14516 1556
rect 14464 1513 14473 1547
rect 14473 1513 14507 1547
rect 14507 1513 14516 1547
rect 14464 1504 14516 1513
rect 14740 1504 14792 1556
rect 16028 1504 16080 1556
rect 16580 1504 16632 1556
rect 9864 1411 9916 1420
rect 6920 1300 6972 1352
rect 7104 1300 7156 1352
rect 8392 1343 8444 1352
rect 8392 1309 8401 1343
rect 8401 1309 8435 1343
rect 8435 1309 8444 1343
rect 8392 1300 8444 1309
rect 8484 1343 8536 1352
rect 8484 1309 8493 1343
rect 8493 1309 8527 1343
rect 8527 1309 8536 1343
rect 9864 1377 9873 1411
rect 9873 1377 9907 1411
rect 9907 1377 9916 1411
rect 9864 1368 9916 1377
rect 8484 1300 8536 1309
rect 9772 1300 9824 1352
rect 10232 1368 10284 1420
rect 11520 1411 11572 1420
rect 8760 1232 8812 1284
rect 8944 1232 8996 1284
rect 11520 1377 11529 1411
rect 11529 1377 11563 1411
rect 11563 1377 11572 1411
rect 11520 1368 11572 1377
rect 11888 1368 11940 1420
rect 12808 1368 12860 1420
rect 12900 1368 12952 1420
rect 13360 1368 13412 1420
rect 13636 1411 13688 1420
rect 13636 1377 13645 1411
rect 13645 1377 13679 1411
rect 13679 1377 13688 1411
rect 13636 1368 13688 1377
rect 14924 1411 14976 1420
rect 13084 1300 13136 1352
rect 12164 1232 12216 1284
rect 12992 1232 13044 1284
rect 13820 1300 13872 1352
rect 14924 1377 14933 1411
rect 14933 1377 14967 1411
rect 14967 1377 14976 1411
rect 14924 1368 14976 1377
rect 15476 1368 15528 1420
rect 16948 1436 17000 1488
rect 17868 1504 17920 1556
rect 18144 1504 18196 1556
rect 17408 1436 17460 1488
rect 17776 1368 17828 1420
rect 18052 1368 18104 1420
rect 14188 1232 14240 1284
rect 14556 1232 14608 1284
rect 7196 1164 7248 1216
rect 9404 1164 9456 1216
rect 10048 1164 10100 1216
rect 11888 1207 11940 1216
rect 11888 1173 11897 1207
rect 11897 1173 11931 1207
rect 11931 1173 11940 1207
rect 11888 1164 11940 1173
rect 11980 1164 12032 1216
rect 12900 1164 12952 1216
rect 13268 1207 13320 1216
rect 13268 1173 13277 1207
rect 13277 1173 13311 1207
rect 13311 1173 13320 1207
rect 13268 1164 13320 1173
rect 13452 1164 13504 1216
rect 16396 1300 16448 1352
rect 17408 1343 17460 1352
rect 17408 1309 17417 1343
rect 17417 1309 17451 1343
rect 17451 1309 17460 1343
rect 17408 1300 17460 1309
rect 16028 1232 16080 1284
rect 16856 1232 16908 1284
rect 16764 1164 16816 1216
rect 17316 1232 17368 1284
rect 17132 1164 17184 1216
rect 17500 1164 17552 1216
rect 3110 1062 3162 1114
rect 3174 1062 3226 1114
rect 3238 1062 3290 1114
rect 3302 1062 3354 1114
rect 3366 1062 3418 1114
rect 6210 1062 6262 1114
rect 6274 1062 6326 1114
rect 6338 1062 6390 1114
rect 6402 1062 6454 1114
rect 6466 1062 6518 1114
rect 9310 1062 9362 1114
rect 9374 1062 9426 1114
rect 9438 1062 9490 1114
rect 9502 1062 9554 1114
rect 9566 1062 9618 1114
rect 12410 1062 12462 1114
rect 12474 1062 12526 1114
rect 12538 1062 12590 1114
rect 12602 1062 12654 1114
rect 12666 1062 12718 1114
rect 15510 1062 15562 1114
rect 15574 1062 15626 1114
rect 15638 1062 15690 1114
rect 15702 1062 15754 1114
rect 15766 1062 15818 1114
rect 18610 1062 18662 1114
rect 18674 1062 18726 1114
rect 18738 1062 18790 1114
rect 18802 1062 18854 1114
rect 18866 1062 18918 1114
rect 6092 960 6144 1012
rect 8300 960 8352 1012
rect 8944 960 8996 1012
rect 10140 960 10192 1012
rect 11520 960 11572 1012
rect 13544 1003 13596 1012
rect 13544 969 13553 1003
rect 13553 969 13587 1003
rect 13587 969 13596 1003
rect 13544 960 13596 969
rect 15384 960 15436 1012
rect 16212 960 16264 1012
rect 17132 1003 17184 1012
rect 17132 969 17141 1003
rect 17141 969 17175 1003
rect 17175 969 17184 1003
rect 17132 960 17184 969
rect 17316 960 17368 1012
rect 18236 960 18288 1012
rect 6000 892 6052 944
rect 14096 935 14148 944
rect 6644 824 6696 876
rect 7012 756 7064 808
rect 8484 824 8536 876
rect 9956 867 10008 876
rect 9956 833 9965 867
rect 9965 833 9999 867
rect 9999 833 10008 867
rect 9956 824 10008 833
rect 13176 824 13228 876
rect 13268 867 13320 876
rect 13268 833 13277 867
rect 13277 833 13311 867
rect 13311 833 13320 867
rect 13268 824 13320 833
rect 8760 799 8812 808
rect 8760 765 8769 799
rect 8769 765 8803 799
rect 8803 765 8812 799
rect 8760 756 8812 765
rect 9772 756 9824 808
rect 12808 799 12860 808
rect 12808 765 12817 799
rect 12817 765 12851 799
rect 12851 765 12860 799
rect 12808 756 12860 765
rect 12992 799 13044 808
rect 12992 765 13001 799
rect 13001 765 13035 799
rect 13035 765 13044 799
rect 14096 901 14105 935
rect 14105 901 14139 935
rect 14139 901 14148 935
rect 14096 892 14148 901
rect 14280 892 14332 944
rect 14372 892 14424 944
rect 16488 892 16540 944
rect 13820 799 13872 808
rect 12992 756 13044 765
rect 13820 765 13829 799
rect 13829 765 13863 799
rect 13863 765 13872 799
rect 13820 756 13872 765
rect 14280 799 14332 808
rect 14280 765 14289 799
rect 14289 765 14323 799
rect 14323 765 14332 799
rect 14280 756 14332 765
rect 14740 756 14792 808
rect 15016 799 15068 808
rect 15016 765 15025 799
rect 15025 765 15059 799
rect 15059 765 15068 799
rect 15016 756 15068 765
rect 16028 867 16080 876
rect 16028 833 16037 867
rect 16037 833 16071 867
rect 16071 833 16080 867
rect 16028 824 16080 833
rect 17592 824 17644 876
rect 17684 799 17736 808
rect 17684 765 17693 799
rect 17693 765 17727 799
rect 17727 765 17736 799
rect 17684 756 17736 765
rect 17868 799 17920 808
rect 17868 765 17877 799
rect 17877 765 17911 799
rect 17911 765 17920 799
rect 18512 799 18564 808
rect 17868 756 17920 765
rect 18512 765 18521 799
rect 18521 765 18555 799
rect 18555 765 18564 799
rect 18512 756 18564 765
rect 19064 756 19116 808
rect 16120 731 16172 740
rect 12072 663 12124 672
rect 12072 629 12081 663
rect 12081 629 12115 663
rect 12115 629 12124 663
rect 12072 620 12124 629
rect 12532 663 12584 672
rect 12532 629 12541 663
rect 12541 629 12575 663
rect 12575 629 12584 663
rect 12532 620 12584 629
rect 12716 663 12768 672
rect 12716 629 12725 663
rect 12725 629 12759 663
rect 12759 629 12768 663
rect 12716 620 12768 629
rect 13728 620 13780 672
rect 16120 697 16129 731
rect 16129 697 16163 731
rect 16163 697 16172 731
rect 16120 688 16172 697
rect 16672 688 16724 740
rect 16856 731 16908 740
rect 16856 697 16865 731
rect 16865 697 16899 731
rect 16899 697 16908 731
rect 16856 688 16908 697
rect 17408 688 17460 740
rect 14188 620 14240 672
rect 16028 620 16080 672
rect 16488 620 16540 672
rect 18328 620 18380 672
rect 4660 518 4712 570
rect 4724 518 4776 570
rect 4788 518 4840 570
rect 4852 518 4904 570
rect 4916 518 4968 570
rect 7760 518 7812 570
rect 7824 518 7876 570
rect 7888 518 7940 570
rect 7952 518 8004 570
rect 8016 518 8068 570
rect 10860 518 10912 570
rect 10924 518 10976 570
rect 10988 518 11040 570
rect 11052 518 11104 570
rect 11116 518 11168 570
rect 13960 518 14012 570
rect 14024 518 14076 570
rect 14088 518 14140 570
rect 14152 518 14204 570
rect 14216 518 14268 570
rect 17060 518 17112 570
rect 17124 518 17176 570
rect 17188 518 17240 570
rect 17252 518 17304 570
rect 17316 518 17368 570
rect 12532 416 12584 468
rect 15936 416 15988 468
rect 11888 348 11940 400
rect 15292 348 15344 400
rect 12716 280 12768 332
rect 15200 280 15252 332
rect 12900 212 12952 264
rect 16856 212 16908 264
rect 13176 144 13228 196
rect 16488 144 16540 196
rect 12072 76 12124 128
rect 18512 76 18564 128
<< metal2 >>
rect 1308 11280 1360 11286
rect 1308 11222 1360 11228
rect 572 11076 624 11082
rect 572 11018 624 11024
rect 584 10810 612 11018
rect 572 10804 624 10810
rect 572 10746 624 10752
rect 1124 10668 1176 10674
rect 1124 10610 1176 10616
rect 756 10600 808 10606
rect 756 10542 808 10548
rect 480 10532 532 10538
rect 480 10474 532 10480
rect 492 9518 520 10474
rect 768 10198 796 10542
rect 756 10192 808 10198
rect 1136 10169 1164 10610
rect 756 10134 808 10140
rect 1122 10160 1178 10169
rect 1122 10095 1178 10104
rect 480 9512 532 9518
rect 1032 9512 1084 9518
rect 480 9454 532 9460
rect 662 9480 718 9489
rect 1032 9454 1084 9460
rect 1124 9512 1176 9518
rect 1124 9454 1176 9460
rect 662 9415 664 9424
rect 716 9415 718 9424
rect 664 9386 716 9392
rect 848 9376 900 9382
rect 848 9318 900 9324
rect 940 9376 992 9382
rect 940 9318 992 9324
rect 572 9036 624 9042
rect 756 9036 808 9042
rect 624 8996 704 9024
rect 572 8978 624 8984
rect 572 8424 624 8430
rect 570 8392 572 8401
rect 624 8392 626 8401
rect 570 8327 626 8336
rect 572 8288 624 8294
rect 572 8230 624 8236
rect 584 8090 612 8230
rect 572 8084 624 8090
rect 572 8026 624 8032
rect 676 8022 704 8996
rect 756 8978 808 8984
rect 768 8634 796 8978
rect 756 8628 808 8634
rect 756 8570 808 8576
rect 756 8356 808 8362
rect 756 8298 808 8304
rect 664 8016 716 8022
rect 662 7984 664 7993
rect 716 7984 718 7993
rect 572 7948 624 7954
rect 662 7919 718 7928
rect 572 7890 624 7896
rect 480 7336 532 7342
rect 584 7313 612 7890
rect 768 7546 796 8298
rect 756 7540 808 7546
rect 756 7482 808 7488
rect 860 7410 888 9318
rect 952 7478 980 9318
rect 1044 8974 1072 9454
rect 1032 8968 1084 8974
rect 1032 8910 1084 8916
rect 1044 8401 1072 8910
rect 1136 8498 1164 9454
rect 1216 9036 1268 9042
rect 1216 8978 1268 8984
rect 1124 8492 1176 8498
rect 1124 8434 1176 8440
rect 1030 8392 1086 8401
rect 1030 8327 1086 8336
rect 940 7472 992 7478
rect 938 7440 940 7449
rect 992 7440 994 7449
rect 848 7404 900 7410
rect 938 7375 994 7384
rect 848 7346 900 7352
rect 480 7278 532 7284
rect 570 7304 626 7313
rect 492 7002 520 7278
rect 1044 7290 1072 8327
rect 1228 7970 1256 8978
rect 1320 8566 1348 11222
rect 1398 11200 1454 12000
rect 1504 11206 2820 11234
rect 1504 11200 1532 11206
rect 1412 11172 1532 11200
rect 1952 11144 2004 11150
rect 1952 11086 2004 11092
rect 1860 11008 1912 11014
rect 1860 10950 1912 10956
rect 1400 10600 1452 10606
rect 1400 10542 1452 10548
rect 1676 10600 1728 10606
rect 1676 10542 1728 10548
rect 1412 9926 1440 10542
rect 1400 9920 1452 9926
rect 1400 9862 1452 9868
rect 1492 9648 1544 9654
rect 1492 9590 1544 9596
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 1308 8560 1360 8566
rect 1308 8502 1360 8508
rect 1412 8430 1440 9454
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1124 7948 1176 7954
rect 1228 7942 1348 7970
rect 1124 7890 1176 7896
rect 1136 7342 1164 7890
rect 1216 7880 1268 7886
rect 1216 7822 1268 7828
rect 1228 7546 1256 7822
rect 1216 7540 1268 7546
rect 1216 7482 1268 7488
rect 1320 7410 1348 7942
rect 1308 7404 1360 7410
rect 1308 7346 1360 7352
rect 1412 7342 1440 8366
rect 1504 7936 1532 9590
rect 1688 9178 1716 10542
rect 1872 10062 1900 10950
rect 1964 10674 1992 11086
rect 2504 10736 2556 10742
rect 2502 10704 2504 10713
rect 2556 10704 2558 10713
rect 1952 10668 2004 10674
rect 2502 10639 2558 10648
rect 1952 10610 2004 10616
rect 2792 10606 2820 11206
rect 4160 11212 4212 11218
rect 4250 11200 4306 12000
rect 4528 11280 4580 11286
rect 4528 11222 4580 11228
rect 4620 11280 4672 11286
rect 4620 11222 4672 11228
rect 6552 11280 6604 11286
rect 6552 11222 6604 11228
rect 4160 11154 4212 11160
rect 2872 11076 2924 11082
rect 2872 11018 2924 11024
rect 2964 11076 3016 11082
rect 2964 11018 3016 11024
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 2136 10464 2188 10470
rect 2136 10406 2188 10412
rect 2688 10464 2740 10470
rect 2688 10406 2740 10412
rect 2148 10266 2176 10406
rect 2136 10260 2188 10266
rect 2136 10202 2188 10208
rect 2700 10198 2728 10406
rect 2688 10192 2740 10198
rect 2688 10134 2740 10140
rect 1860 10056 1912 10062
rect 1860 9998 1912 10004
rect 2044 10056 2096 10062
rect 2044 9998 2096 10004
rect 1952 9920 2004 9926
rect 1952 9862 2004 9868
rect 1766 9480 1822 9489
rect 1766 9415 1768 9424
rect 1820 9415 1822 9424
rect 1768 9386 1820 9392
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 1504 7908 1624 7936
rect 1492 7812 1544 7818
rect 1492 7754 1544 7760
rect 570 7239 626 7248
rect 952 7262 1072 7290
rect 1124 7336 1176 7342
rect 1124 7278 1176 7284
rect 1216 7336 1268 7342
rect 1216 7278 1268 7284
rect 1400 7336 1452 7342
rect 1400 7278 1452 7284
rect 480 6996 532 7002
rect 480 6938 532 6944
rect 584 6458 612 7239
rect 846 7032 902 7041
rect 846 6967 902 6976
rect 754 6896 810 6905
rect 860 6866 888 6967
rect 754 6831 756 6840
rect 808 6831 810 6840
rect 848 6860 900 6866
rect 756 6802 808 6808
rect 848 6802 900 6808
rect 572 6452 624 6458
rect 572 6394 624 6400
rect 848 6248 900 6254
rect 846 6216 848 6225
rect 900 6216 902 6225
rect 846 6151 902 6160
rect 952 5710 980 7262
rect 1032 7200 1084 7206
rect 1228 7177 1256 7278
rect 1032 7142 1084 7148
rect 1214 7168 1270 7177
rect 1044 6254 1072 7142
rect 1214 7103 1270 7112
rect 1124 6656 1176 6662
rect 1124 6598 1176 6604
rect 1136 6390 1164 6598
rect 1124 6384 1176 6390
rect 1124 6326 1176 6332
rect 1032 6248 1084 6254
rect 1032 6190 1084 6196
rect 940 5704 992 5710
rect 940 5646 992 5652
rect 1136 4282 1164 6326
rect 1228 6322 1256 7103
rect 1306 6760 1362 6769
rect 1306 6695 1362 6704
rect 1216 6316 1268 6322
rect 1216 6258 1268 6264
rect 1320 6254 1348 6695
rect 1308 6248 1360 6254
rect 1308 6190 1360 6196
rect 1412 5794 1440 7278
rect 1504 6798 1532 7754
rect 1492 6792 1544 6798
rect 1492 6734 1544 6740
rect 1492 6248 1544 6254
rect 1492 6190 1544 6196
rect 1504 5914 1532 6190
rect 1596 5914 1624 7908
rect 1676 7744 1728 7750
rect 1676 7686 1728 7692
rect 1688 7256 1716 7686
rect 1768 7268 1820 7274
rect 1688 7228 1768 7256
rect 1768 7210 1820 7216
rect 1964 7154 1992 9862
rect 2056 9110 2084 9998
rect 2136 9376 2188 9382
rect 2188 9336 2360 9364
rect 2136 9318 2188 9324
rect 2044 9104 2096 9110
rect 2044 9046 2096 9052
rect 2136 9036 2188 9042
rect 2136 8978 2188 8984
rect 2148 7818 2176 8978
rect 2332 8974 2360 9336
rect 2688 9036 2740 9042
rect 2688 8978 2740 8984
rect 2320 8968 2372 8974
rect 2320 8910 2372 8916
rect 2332 7993 2360 8910
rect 2596 8288 2648 8294
rect 2596 8230 2648 8236
rect 2412 8084 2464 8090
rect 2412 8026 2464 8032
rect 2318 7984 2374 7993
rect 2318 7919 2374 7928
rect 2228 7880 2280 7886
rect 2332 7868 2360 7919
rect 2424 7886 2452 8026
rect 2280 7840 2360 7868
rect 2412 7880 2464 7886
rect 2228 7822 2280 7828
rect 2412 7822 2464 7828
rect 2136 7812 2188 7818
rect 2136 7754 2188 7760
rect 2136 7404 2188 7410
rect 2136 7346 2188 7352
rect 1780 7126 1992 7154
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 1688 6458 1716 6734
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 1780 6338 1808 7126
rect 2148 7002 2176 7346
rect 2136 6996 2188 7002
rect 2136 6938 2188 6944
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1688 6310 1808 6338
rect 1872 6322 1900 6598
rect 2148 6361 2176 6938
rect 2134 6352 2190 6361
rect 1860 6316 1912 6322
rect 1492 5908 1544 5914
rect 1492 5850 1544 5856
rect 1584 5908 1636 5914
rect 1584 5850 1636 5856
rect 1412 5778 1532 5794
rect 1412 5772 1544 5778
rect 1412 5766 1492 5772
rect 1492 5714 1544 5720
rect 1400 5568 1452 5574
rect 1400 5510 1452 5516
rect 1412 5114 1440 5510
rect 1504 5234 1532 5714
rect 1492 5228 1544 5234
rect 1492 5170 1544 5176
rect 1688 5114 1716 6310
rect 1860 6258 1912 6264
rect 2044 6316 2096 6322
rect 2134 6287 2190 6296
rect 2044 6258 2096 6264
rect 2056 5710 2084 6258
rect 2148 5778 2176 6287
rect 2136 5772 2188 5778
rect 2136 5714 2188 5720
rect 2240 5710 2268 7822
rect 2502 7304 2558 7313
rect 2502 7239 2558 7248
rect 2410 7032 2466 7041
rect 2410 6967 2412 6976
rect 2464 6967 2466 6976
rect 2412 6938 2464 6944
rect 2044 5704 2096 5710
rect 2044 5646 2096 5652
rect 2228 5704 2280 5710
rect 2228 5646 2280 5652
rect 1952 5364 2004 5370
rect 2056 5352 2084 5646
rect 2004 5324 2084 5352
rect 1952 5306 2004 5312
rect 1412 5086 1716 5114
rect 1124 4276 1176 4282
rect 1124 4218 1176 4224
rect 1412 2854 1440 5086
rect 2516 4826 2544 7239
rect 2608 5778 2636 8230
rect 2700 7868 2728 8978
rect 2792 8276 2820 10542
rect 2884 10198 2912 11018
rect 2976 10674 3004 11018
rect 3110 10908 3418 10917
rect 3110 10906 3116 10908
rect 3172 10906 3196 10908
rect 3252 10906 3276 10908
rect 3332 10906 3356 10908
rect 3412 10906 3418 10908
rect 3172 10854 3174 10906
rect 3354 10854 3356 10906
rect 3110 10852 3116 10854
rect 3172 10852 3196 10854
rect 3252 10852 3276 10854
rect 3332 10852 3356 10854
rect 3412 10852 3418 10854
rect 3110 10843 3418 10852
rect 4172 10690 4200 11154
rect 4080 10674 4200 10690
rect 2964 10668 3016 10674
rect 2964 10610 3016 10616
rect 4068 10668 4200 10674
rect 4120 10662 4200 10668
rect 4068 10610 4120 10616
rect 2872 10192 2924 10198
rect 2872 10134 2924 10140
rect 2884 9110 2912 10134
rect 2976 10112 3004 10610
rect 4066 10568 4122 10577
rect 4066 10503 4122 10512
rect 4080 10470 4108 10503
rect 3884 10464 3936 10470
rect 3884 10406 3936 10412
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 2976 10084 3096 10112
rect 3068 9994 3096 10084
rect 3146 10024 3202 10033
rect 2964 9988 3016 9994
rect 2964 9930 3016 9936
rect 3056 9988 3108 9994
rect 3146 9959 3202 9968
rect 3514 10024 3570 10033
rect 3514 9959 3570 9968
rect 3056 9930 3108 9936
rect 2872 9104 2924 9110
rect 2872 9046 2924 9052
rect 2884 8430 2912 9046
rect 2872 8424 2924 8430
rect 2872 8366 2924 8372
rect 2792 8248 2912 8276
rect 2780 7880 2832 7886
rect 2700 7840 2780 7868
rect 2884 7868 2912 8248
rect 2976 8022 3004 9930
rect 3160 9926 3188 9959
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 3110 9820 3418 9829
rect 3110 9818 3116 9820
rect 3172 9818 3196 9820
rect 3252 9818 3276 9820
rect 3332 9818 3356 9820
rect 3412 9818 3418 9820
rect 3172 9766 3174 9818
rect 3354 9766 3356 9818
rect 3110 9764 3116 9766
rect 3172 9764 3196 9766
rect 3252 9764 3276 9766
rect 3332 9764 3356 9766
rect 3412 9764 3418 9766
rect 3110 9755 3418 9764
rect 3056 9444 3108 9450
rect 3056 9386 3108 9392
rect 3068 9110 3096 9386
rect 3056 9104 3108 9110
rect 3056 9046 3108 9052
rect 3110 8732 3418 8741
rect 3110 8730 3116 8732
rect 3172 8730 3196 8732
rect 3252 8730 3276 8732
rect 3332 8730 3356 8732
rect 3412 8730 3418 8732
rect 3172 8678 3174 8730
rect 3354 8678 3356 8730
rect 3110 8676 3116 8678
rect 3172 8676 3196 8678
rect 3252 8676 3276 8678
rect 3332 8676 3356 8678
rect 3412 8676 3418 8678
rect 3110 8667 3418 8676
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 3436 8498 3464 8570
rect 3528 8566 3556 9959
rect 3700 9580 3752 9586
rect 3700 9522 3752 9528
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3620 8566 3648 9318
rect 3712 9178 3740 9522
rect 3792 9444 3844 9450
rect 3792 9386 3844 9392
rect 3700 9172 3752 9178
rect 3700 9114 3752 9120
rect 3700 8968 3752 8974
rect 3700 8910 3752 8916
rect 3712 8634 3740 8910
rect 3700 8628 3752 8634
rect 3700 8570 3752 8576
rect 3516 8560 3568 8566
rect 3516 8502 3568 8508
rect 3608 8560 3660 8566
rect 3608 8502 3660 8508
rect 3424 8492 3476 8498
rect 3424 8434 3476 8440
rect 3056 8424 3108 8430
rect 3056 8366 3108 8372
rect 2964 8016 3016 8022
rect 2964 7958 3016 7964
rect 2884 7840 3004 7868
rect 2780 7822 2832 7828
rect 2792 7478 2820 7822
rect 2872 7744 2924 7750
rect 2872 7686 2924 7692
rect 2780 7472 2832 7478
rect 2700 7432 2780 7460
rect 2700 6798 2728 7432
rect 2780 7414 2832 7420
rect 2884 7342 2912 7686
rect 2872 7336 2924 7342
rect 2872 7278 2924 7284
rect 2780 7200 2832 7206
rect 2976 7188 3004 7840
rect 3068 7750 3096 8366
rect 3436 8294 3464 8434
rect 3528 8430 3556 8502
rect 3516 8424 3568 8430
rect 3516 8366 3568 8372
rect 3528 8294 3556 8366
rect 3424 8288 3476 8294
rect 3528 8266 3648 8294
rect 3424 8230 3476 8236
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 3056 7744 3108 7750
rect 3056 7686 3108 7692
rect 3110 7644 3418 7653
rect 3110 7642 3116 7644
rect 3172 7642 3196 7644
rect 3252 7642 3276 7644
rect 3332 7642 3356 7644
rect 3412 7642 3418 7644
rect 3172 7590 3174 7642
rect 3354 7590 3356 7642
rect 3110 7588 3116 7590
rect 3172 7588 3196 7590
rect 3252 7588 3276 7590
rect 3332 7588 3356 7590
rect 3412 7588 3418 7590
rect 3110 7579 3418 7588
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 2780 7142 2832 7148
rect 2884 7160 3004 7188
rect 3054 7168 3110 7177
rect 2688 6792 2740 6798
rect 2688 6734 2740 6740
rect 2792 5778 2820 7142
rect 2884 6390 2912 7160
rect 3054 7103 3110 7112
rect 2962 7032 3018 7041
rect 2962 6967 3018 6976
rect 2976 6866 3004 6967
rect 3068 6934 3096 7103
rect 3344 7002 3372 7482
rect 3424 7200 3476 7206
rect 3424 7142 3476 7148
rect 3240 6996 3292 7002
rect 3240 6938 3292 6944
rect 3332 6996 3384 7002
rect 3332 6938 3384 6944
rect 3056 6928 3108 6934
rect 3056 6870 3108 6876
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 3252 6662 3280 6938
rect 3436 6769 3464 7142
rect 3422 6760 3478 6769
rect 3422 6695 3478 6704
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 2872 6384 2924 6390
rect 2872 6326 2924 6332
rect 2596 5772 2648 5778
rect 2596 5714 2648 5720
rect 2780 5772 2832 5778
rect 2780 5714 2832 5720
rect 2976 5098 3004 6598
rect 3110 6556 3418 6565
rect 3110 6554 3116 6556
rect 3172 6554 3196 6556
rect 3252 6554 3276 6556
rect 3332 6554 3356 6556
rect 3412 6554 3418 6556
rect 3172 6502 3174 6554
rect 3354 6502 3356 6554
rect 3110 6500 3116 6502
rect 3172 6500 3196 6502
rect 3252 6500 3276 6502
rect 3332 6500 3356 6502
rect 3412 6500 3418 6502
rect 3110 6491 3418 6500
rect 3056 6384 3108 6390
rect 3240 6384 3292 6390
rect 3056 6326 3108 6332
rect 3238 6352 3240 6361
rect 3292 6352 3294 6361
rect 3068 5914 3096 6326
rect 3238 6287 3294 6296
rect 3528 5914 3556 7822
rect 3620 7546 3648 8266
rect 3700 7744 3752 7750
rect 3700 7686 3752 7692
rect 3608 7540 3660 7546
rect 3608 7482 3660 7488
rect 3712 7018 3740 7686
rect 3804 7449 3832 9386
rect 3896 8430 3924 10406
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 4172 9722 4200 9998
rect 4160 9716 4212 9722
rect 4160 9658 4212 9664
rect 4160 9512 4212 9518
rect 3988 9460 4160 9466
rect 3988 9454 4212 9460
rect 3988 9438 4200 9454
rect 3988 8634 4016 9438
rect 4068 8900 4120 8906
rect 4068 8842 4120 8848
rect 4160 8900 4212 8906
rect 4160 8842 4212 8848
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 3884 8424 3936 8430
rect 3884 8366 3936 8372
rect 3884 8016 3936 8022
rect 3884 7958 3936 7964
rect 3896 7750 3924 7958
rect 4080 7954 4108 8842
rect 4172 8090 4200 8842
rect 4264 8634 4292 11200
rect 4344 10804 4396 10810
rect 4344 10746 4396 10752
rect 4356 9722 4384 10746
rect 4540 10606 4568 11222
rect 4632 10606 4660 11222
rect 4988 11076 5040 11082
rect 4988 11018 5040 11024
rect 4528 10600 4580 10606
rect 4528 10542 4580 10548
rect 4620 10600 4672 10606
rect 4620 10542 4672 10548
rect 4660 10364 4968 10373
rect 4660 10362 4666 10364
rect 4722 10362 4746 10364
rect 4802 10362 4826 10364
rect 4882 10362 4906 10364
rect 4962 10362 4968 10364
rect 4722 10310 4724 10362
rect 4904 10310 4906 10362
rect 4660 10308 4666 10310
rect 4722 10308 4746 10310
rect 4802 10308 4826 10310
rect 4882 10308 4906 10310
rect 4962 10308 4968 10310
rect 4660 10299 4968 10308
rect 5000 10198 5028 11018
rect 5264 11008 5316 11014
rect 5264 10950 5316 10956
rect 5276 10810 5304 10950
rect 6210 10908 6518 10917
rect 6210 10906 6216 10908
rect 6272 10906 6296 10908
rect 6352 10906 6376 10908
rect 6432 10906 6456 10908
rect 6512 10906 6518 10908
rect 6272 10854 6274 10906
rect 6454 10854 6456 10906
rect 6210 10852 6216 10854
rect 6272 10852 6296 10854
rect 6352 10852 6376 10854
rect 6432 10852 6456 10854
rect 6512 10852 6518 10854
rect 6210 10843 6518 10852
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 5538 10568 5594 10577
rect 5538 10503 5594 10512
rect 5552 10470 5580 10503
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 4712 10192 4764 10198
rect 4434 10160 4490 10169
rect 4712 10134 4764 10140
rect 4988 10192 5040 10198
rect 4988 10134 5040 10140
rect 4434 10095 4490 10104
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 4448 9178 4476 10095
rect 4528 10056 4580 10062
rect 4528 9998 4580 10004
rect 4540 9722 4568 9998
rect 4620 9920 4672 9926
rect 4620 9862 4672 9868
rect 4632 9722 4660 9862
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4620 9716 4672 9722
rect 4620 9658 4672 9664
rect 4724 9602 4752 10134
rect 4896 10124 4948 10130
rect 4896 10066 4948 10072
rect 4908 10033 4936 10066
rect 5172 10056 5224 10062
rect 4894 10024 4950 10033
rect 5172 9998 5224 10004
rect 4894 9959 4950 9968
rect 4988 9988 5040 9994
rect 4988 9930 5040 9936
rect 4540 9574 4752 9602
rect 4436 9172 4488 9178
rect 4436 9114 4488 9120
rect 4436 9036 4488 9042
rect 4436 8978 4488 8984
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 4252 8628 4304 8634
rect 4252 8570 4304 8576
rect 4264 8430 4292 8570
rect 4252 8424 4304 8430
rect 4252 8366 4304 8372
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 4068 7948 4120 7954
rect 4068 7890 4120 7896
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 4080 7478 4108 7890
rect 3976 7472 4028 7478
rect 3790 7440 3846 7449
rect 3976 7414 4028 7420
rect 4068 7472 4120 7478
rect 4068 7414 4120 7420
rect 3790 7375 3792 7384
rect 3844 7375 3846 7384
rect 3792 7346 3844 7352
rect 3804 7315 3832 7346
rect 3988 7206 4016 7414
rect 4068 7336 4120 7342
rect 4252 7336 4304 7342
rect 4068 7278 4120 7284
rect 4250 7304 4252 7313
rect 4304 7304 4306 7313
rect 3976 7200 4028 7206
rect 3976 7142 4028 7148
rect 3620 6990 3740 7018
rect 3620 6254 3648 6990
rect 3700 6860 3752 6866
rect 3700 6802 3752 6808
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3110 5468 3418 5477
rect 3110 5466 3116 5468
rect 3172 5466 3196 5468
rect 3252 5466 3276 5468
rect 3332 5466 3356 5468
rect 3412 5466 3418 5468
rect 3172 5414 3174 5466
rect 3354 5414 3356 5466
rect 3110 5412 3116 5414
rect 3172 5412 3196 5414
rect 3252 5412 3276 5414
rect 3332 5412 3356 5414
rect 3412 5412 3418 5414
rect 3110 5403 3418 5412
rect 2964 5092 3016 5098
rect 2964 5034 3016 5040
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 2964 4820 3016 4826
rect 2964 4762 3016 4768
rect 2504 4684 2556 4690
rect 2504 4626 2556 4632
rect 2228 4004 2280 4010
rect 2228 3946 2280 3952
rect 2240 3738 2268 3946
rect 2516 3942 2544 4626
rect 2976 4486 3004 4762
rect 3528 4758 3556 5850
rect 3620 5030 3648 6190
rect 3712 5642 3740 6802
rect 4080 6798 4108 7278
rect 4250 7239 4306 7248
rect 4158 7032 4214 7041
rect 4264 7002 4292 7239
rect 4158 6967 4214 6976
rect 4252 6996 4304 7002
rect 4172 6934 4200 6967
rect 4252 6938 4304 6944
rect 4160 6928 4212 6934
rect 4160 6870 4212 6876
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 3976 6724 4028 6730
rect 3976 6666 4028 6672
rect 3988 6254 4016 6666
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 3884 6180 3936 6186
rect 3884 6122 3936 6128
rect 3896 6066 3924 6122
rect 3804 6038 3924 6066
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 3804 5846 3832 6038
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 3792 5840 3844 5846
rect 3792 5782 3844 5788
rect 3700 5636 3752 5642
rect 3700 5578 3752 5584
rect 3896 5234 3924 5850
rect 4080 5846 4108 6054
rect 4068 5840 4120 5846
rect 4068 5782 4120 5788
rect 4172 5234 4200 6870
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 4264 6225 4292 6802
rect 4356 6662 4384 8774
rect 4448 8362 4476 8978
rect 4436 8356 4488 8362
rect 4436 8298 4488 8304
rect 4436 8016 4488 8022
rect 4436 7958 4488 7964
rect 4448 7342 4476 7958
rect 4436 7336 4488 7342
rect 4436 7278 4488 7284
rect 4344 6656 4396 6662
rect 4344 6598 4396 6604
rect 4250 6216 4306 6225
rect 4250 6151 4306 6160
rect 4356 5846 4384 6598
rect 4344 5840 4396 5846
rect 4344 5782 4396 5788
rect 3884 5228 3936 5234
rect 3884 5170 3936 5176
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 4252 5160 4304 5166
rect 4252 5102 4304 5108
rect 3608 5024 3660 5030
rect 3608 4966 3660 4972
rect 4264 4826 4292 5102
rect 4252 4820 4304 4826
rect 4252 4762 4304 4768
rect 3516 4752 3568 4758
rect 4356 4729 4384 5782
rect 4448 5574 4476 7278
rect 4540 6984 4568 9574
rect 4660 9276 4968 9285
rect 4660 9274 4666 9276
rect 4722 9274 4746 9276
rect 4802 9274 4826 9276
rect 4882 9274 4906 9276
rect 4962 9274 4968 9276
rect 4722 9222 4724 9274
rect 4904 9222 4906 9274
rect 4660 9220 4666 9222
rect 4722 9220 4746 9222
rect 4802 9220 4826 9222
rect 4882 9220 4906 9222
rect 4962 9220 4968 9222
rect 4660 9211 4968 9220
rect 5000 9042 5028 9930
rect 5080 9716 5132 9722
rect 5080 9658 5132 9664
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 4986 8392 5042 8401
rect 4986 8327 5042 8336
rect 4660 8188 4968 8197
rect 4660 8186 4666 8188
rect 4722 8186 4746 8188
rect 4802 8186 4826 8188
rect 4882 8186 4906 8188
rect 4962 8186 4968 8188
rect 4722 8134 4724 8186
rect 4904 8134 4906 8186
rect 4660 8132 4666 8134
rect 4722 8132 4746 8134
rect 4802 8132 4826 8134
rect 4882 8132 4906 8134
rect 4962 8132 4968 8134
rect 4660 8123 4968 8132
rect 5000 7886 5028 8327
rect 5092 8090 5120 9658
rect 5184 8498 5212 9998
rect 5356 9920 5408 9926
rect 5356 9862 5408 9868
rect 5264 9444 5316 9450
rect 5264 9386 5316 9392
rect 5276 9110 5304 9386
rect 5264 9104 5316 9110
rect 5264 9046 5316 9052
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 5172 7812 5224 7818
rect 5172 7754 5224 7760
rect 5184 7274 5212 7754
rect 5172 7268 5224 7274
rect 5172 7210 5224 7216
rect 5276 7206 5304 9046
rect 5368 8294 5396 9862
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 5368 7546 5396 8230
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 4660 7100 4968 7109
rect 4660 7098 4666 7100
rect 4722 7098 4746 7100
rect 4802 7098 4826 7100
rect 4882 7098 4906 7100
rect 4962 7098 4968 7100
rect 4722 7046 4724 7098
rect 4904 7046 4906 7098
rect 4660 7044 4666 7046
rect 4722 7044 4746 7046
rect 4802 7044 4826 7046
rect 4882 7044 4906 7046
rect 4962 7044 4968 7046
rect 4660 7035 4968 7044
rect 5000 7002 5028 7142
rect 4988 6996 5040 7002
rect 4540 6956 4660 6984
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 4540 6390 4568 6734
rect 4632 6730 4660 6956
rect 4988 6938 5040 6944
rect 5460 6905 5488 10406
rect 5552 10198 5580 10406
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5736 8838 5764 9522
rect 5724 8832 5776 8838
rect 5724 8774 5776 8780
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5552 7342 5580 8434
rect 5736 7886 5764 8774
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5828 7750 5856 10746
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 5920 10130 5948 10610
rect 6092 10464 6144 10470
rect 6092 10406 6144 10412
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 6104 9722 6132 10406
rect 6210 9820 6518 9829
rect 6210 9818 6216 9820
rect 6272 9818 6296 9820
rect 6352 9818 6376 9820
rect 6432 9818 6456 9820
rect 6512 9818 6518 9820
rect 6272 9766 6274 9818
rect 6454 9766 6456 9818
rect 6210 9764 6216 9766
rect 6272 9764 6296 9766
rect 6352 9764 6376 9766
rect 6432 9764 6456 9766
rect 6512 9764 6518 9766
rect 6210 9755 6518 9764
rect 6092 9716 6144 9722
rect 6092 9658 6144 9664
rect 6564 9674 6592 11222
rect 7102 11200 7158 12000
rect 7288 11416 7340 11422
rect 7288 11358 7340 11364
rect 9680 11416 9732 11422
rect 9680 11358 9732 11364
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 6104 7954 6132 9658
rect 6564 9646 6684 9674
rect 6552 9512 6604 9518
rect 6552 9454 6604 9460
rect 6210 8732 6518 8741
rect 6210 8730 6216 8732
rect 6272 8730 6296 8732
rect 6352 8730 6376 8732
rect 6432 8730 6456 8732
rect 6512 8730 6518 8732
rect 6272 8678 6274 8730
rect 6454 8678 6456 8730
rect 6210 8676 6216 8678
rect 6272 8676 6296 8678
rect 6352 8676 6376 8678
rect 6432 8676 6456 8678
rect 6512 8676 6518 8678
rect 6210 8667 6518 8676
rect 6564 8634 6592 9454
rect 6656 9382 6684 9646
rect 6932 9382 6960 11018
rect 7012 10668 7064 10674
rect 7012 10610 7064 10616
rect 7024 9518 7052 10610
rect 7012 9512 7064 9518
rect 7012 9454 7064 9460
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6552 8628 6604 8634
rect 6552 8570 6604 8576
rect 6656 7954 6684 9318
rect 6828 9104 6880 9110
rect 6828 9046 6880 9052
rect 6840 7954 6868 9046
rect 7116 8498 7144 11200
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 6092 7948 6144 7954
rect 6012 7908 6092 7936
rect 5816 7744 5868 7750
rect 5816 7686 5868 7692
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5828 7274 5856 7686
rect 5816 7268 5868 7274
rect 5816 7210 5868 7216
rect 5446 6896 5502 6905
rect 5446 6831 5502 6840
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 4620 6724 4672 6730
rect 4620 6666 4672 6672
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 4528 6384 4580 6390
rect 4528 6326 4580 6332
rect 4540 5710 4568 6326
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 4660 6012 4968 6021
rect 4660 6010 4666 6012
rect 4722 6010 4746 6012
rect 4802 6010 4826 6012
rect 4882 6010 4906 6012
rect 4962 6010 4968 6012
rect 4722 5958 4724 6010
rect 4904 5958 4906 6010
rect 4660 5956 4666 5958
rect 4722 5956 4746 5958
rect 4802 5956 4826 5958
rect 4882 5956 4906 5958
rect 4962 5956 4968 5958
rect 4660 5947 4968 5956
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4436 5568 4488 5574
rect 4436 5510 4488 5516
rect 4660 4924 4968 4933
rect 4660 4922 4666 4924
rect 4722 4922 4746 4924
rect 4802 4922 4826 4924
rect 4882 4922 4906 4924
rect 4962 4922 4968 4924
rect 4722 4870 4724 4922
rect 4904 4870 4906 4922
rect 4660 4868 4666 4870
rect 4722 4868 4746 4870
rect 4802 4868 4826 4870
rect 4882 4868 4906 4870
rect 4962 4868 4968 4870
rect 4660 4859 4968 4868
rect 4712 4752 4764 4758
rect 3516 4694 3568 4700
rect 4342 4720 4398 4729
rect 4712 4694 4764 4700
rect 4342 4655 4398 4664
rect 2964 4480 3016 4486
rect 2964 4422 3016 4428
rect 3110 4380 3418 4389
rect 3110 4378 3116 4380
rect 3172 4378 3196 4380
rect 3252 4378 3276 4380
rect 3332 4378 3356 4380
rect 3412 4378 3418 4380
rect 3172 4326 3174 4378
rect 3354 4326 3356 4378
rect 3110 4324 3116 4326
rect 3172 4324 3196 4326
rect 3252 4324 3276 4326
rect 3332 4324 3356 4326
rect 3412 4324 3418 4326
rect 3110 4315 3418 4324
rect 4356 4146 4384 4655
rect 4724 4214 4752 4694
rect 5000 4622 5028 6054
rect 5276 5574 5304 6598
rect 5552 6322 5580 6734
rect 6012 6458 6040 7908
rect 6092 7890 6144 7896
rect 6184 7948 6236 7954
rect 6184 7890 6236 7896
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6196 7800 6224 7890
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6104 7772 6224 7800
rect 6104 6905 6132 7772
rect 6210 7644 6518 7653
rect 6210 7642 6216 7644
rect 6272 7642 6296 7644
rect 6352 7642 6376 7644
rect 6432 7642 6456 7644
rect 6512 7642 6518 7644
rect 6272 7590 6274 7642
rect 6454 7590 6456 7642
rect 6210 7588 6216 7590
rect 6272 7588 6296 7590
rect 6352 7588 6376 7590
rect 6432 7588 6456 7590
rect 6512 7588 6518 7590
rect 6210 7579 6518 7588
rect 6564 7410 6592 7822
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6644 7336 6696 7342
rect 6644 7278 6696 7284
rect 6090 6896 6146 6905
rect 6090 6831 6146 6840
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5908 6316 5960 6322
rect 5908 6258 5960 6264
rect 5446 5672 5502 5681
rect 5446 5607 5502 5616
rect 5264 5568 5316 5574
rect 5264 5510 5316 5516
rect 5172 5024 5224 5030
rect 5276 5012 5304 5510
rect 5356 5092 5408 5098
rect 5356 5034 5408 5040
rect 5224 4984 5304 5012
rect 5172 4966 5224 4972
rect 5276 4690 5304 4984
rect 5368 4758 5396 5034
rect 5356 4752 5408 4758
rect 5356 4694 5408 4700
rect 5264 4684 5316 4690
rect 5264 4626 5316 4632
rect 4988 4616 5040 4622
rect 4988 4558 5040 4564
rect 5460 4554 5488 5607
rect 5552 5250 5580 6258
rect 5632 6180 5684 6186
rect 5632 6122 5684 6128
rect 5644 5370 5672 6122
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 5828 5778 5856 6054
rect 5920 5817 5948 6258
rect 6104 6186 6132 6831
rect 6210 6556 6518 6565
rect 6210 6554 6216 6556
rect 6272 6554 6296 6556
rect 6352 6554 6376 6556
rect 6432 6554 6456 6556
rect 6512 6554 6518 6556
rect 6272 6502 6274 6554
rect 6454 6502 6456 6554
rect 6210 6500 6216 6502
rect 6272 6500 6296 6502
rect 6352 6500 6376 6502
rect 6432 6500 6456 6502
rect 6512 6500 6518 6502
rect 6210 6491 6518 6500
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6288 6254 6316 6394
rect 6276 6248 6328 6254
rect 6276 6190 6328 6196
rect 6552 6248 6604 6254
rect 6552 6190 6604 6196
rect 6092 6180 6144 6186
rect 6092 6122 6144 6128
rect 6000 6112 6052 6118
rect 6000 6054 6052 6060
rect 5906 5808 5962 5817
rect 5816 5772 5868 5778
rect 5906 5743 5962 5752
rect 5816 5714 5868 5720
rect 5724 5636 5776 5642
rect 5724 5578 5776 5584
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5552 5222 5672 5250
rect 5540 5092 5592 5098
rect 5540 5034 5592 5040
rect 5264 4548 5316 4554
rect 5448 4548 5500 4554
rect 5316 4508 5396 4536
rect 5264 4490 5316 4496
rect 4712 4208 4764 4214
rect 4712 4150 4764 4156
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 3608 4072 3660 4078
rect 3608 4014 3660 4020
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 2504 3936 2556 3942
rect 2504 3878 2556 3884
rect 2596 3936 2648 3942
rect 2596 3878 2648 3884
rect 2228 3732 2280 3738
rect 2228 3674 2280 3680
rect 2516 3534 2544 3878
rect 2608 3602 2636 3878
rect 3620 3670 3648 4014
rect 4172 3720 4200 4014
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 4528 3936 4580 3942
rect 4528 3878 4580 3884
rect 4252 3732 4304 3738
rect 4172 3692 4252 3720
rect 3608 3664 3660 3670
rect 3608 3606 3660 3612
rect 2596 3596 2648 3602
rect 2596 3538 2648 3544
rect 2504 3528 2556 3534
rect 2504 3470 2556 3476
rect 2964 3528 3016 3534
rect 2964 3470 3016 3476
rect 1860 2984 1912 2990
rect 1860 2926 1912 2932
rect 1400 2848 1452 2854
rect 1400 2790 1452 2796
rect 1872 2582 1900 2926
rect 1860 2576 1912 2582
rect 1860 2518 1912 2524
rect 2516 2514 2544 3470
rect 2872 3392 2924 3398
rect 2872 3334 2924 3340
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2792 2650 2820 2994
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 2504 2508 2556 2514
rect 2504 2450 2556 2456
rect 2516 1902 2544 2450
rect 2884 2378 2912 3334
rect 2976 3194 3004 3470
rect 3110 3292 3418 3301
rect 3110 3290 3116 3292
rect 3172 3290 3196 3292
rect 3252 3290 3276 3292
rect 3332 3290 3356 3292
rect 3412 3290 3418 3292
rect 3172 3238 3174 3290
rect 3354 3238 3356 3290
rect 3110 3236 3116 3238
rect 3172 3236 3196 3238
rect 3252 3236 3276 3238
rect 3332 3236 3356 3238
rect 3412 3236 3418 3238
rect 3110 3227 3418 3236
rect 2964 3188 3016 3194
rect 2964 3130 3016 3136
rect 3620 2990 3648 3606
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 4080 3194 4108 3334
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 3608 2984 3660 2990
rect 3608 2926 3660 2932
rect 3620 2774 3648 2926
rect 3700 2916 3752 2922
rect 3700 2858 3752 2864
rect 3528 2746 3648 2774
rect 2872 2372 2924 2378
rect 2872 2314 2924 2320
rect 3110 2204 3418 2213
rect 3110 2202 3116 2204
rect 3172 2202 3196 2204
rect 3252 2202 3276 2204
rect 3332 2202 3356 2204
rect 3412 2202 3418 2204
rect 3172 2150 3174 2202
rect 3354 2150 3356 2202
rect 3110 2148 3116 2150
rect 3172 2148 3196 2150
rect 3252 2148 3276 2150
rect 3332 2148 3356 2150
rect 3412 2148 3418 2150
rect 3110 2139 3418 2148
rect 2504 1896 2556 1902
rect 2504 1838 2556 1844
rect 2964 1828 3016 1834
rect 2964 1770 3016 1776
rect 2976 1426 3004 1770
rect 3528 1562 3556 2746
rect 3712 2514 3740 2858
rect 4172 2774 4200 3692
rect 4252 3674 4304 3680
rect 4356 3058 4384 3878
rect 4436 3664 4488 3670
rect 4436 3606 4488 3612
rect 4344 3052 4396 3058
rect 4344 2994 4396 3000
rect 4252 2984 4304 2990
rect 4252 2926 4304 2932
rect 3804 2746 4200 2774
rect 3700 2508 3752 2514
rect 3700 2450 3752 2456
rect 3804 2446 3832 2746
rect 4264 2514 4292 2926
rect 4344 2848 4396 2854
rect 4344 2790 4396 2796
rect 4356 2650 4384 2790
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 4252 2508 4304 2514
rect 4252 2450 4304 2456
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 4448 1902 4476 3606
rect 4540 2106 4568 3878
rect 4660 3836 4968 3845
rect 4660 3834 4666 3836
rect 4722 3834 4746 3836
rect 4802 3834 4826 3836
rect 4882 3834 4906 3836
rect 4962 3834 4968 3836
rect 4722 3782 4724 3834
rect 4904 3782 4906 3834
rect 4660 3780 4666 3782
rect 4722 3780 4746 3782
rect 4802 3780 4826 3782
rect 4882 3780 4906 3782
rect 4962 3780 4968 3782
rect 4660 3771 4968 3780
rect 5000 3670 5028 4082
rect 5172 4072 5224 4078
rect 5172 4014 5224 4020
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 5092 3738 5120 3878
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 4988 3664 5040 3670
rect 4988 3606 5040 3612
rect 5184 3602 5212 4014
rect 5264 3936 5316 3942
rect 5264 3878 5316 3884
rect 4896 3596 4948 3602
rect 4896 3538 4948 3544
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 4802 3496 4858 3505
rect 4802 3431 4858 3440
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4632 2990 4660 3334
rect 4620 2984 4672 2990
rect 4620 2926 4672 2932
rect 4816 2922 4844 3431
rect 4908 2922 4936 3538
rect 5276 3398 5304 3878
rect 5368 3670 5396 4508
rect 5448 4490 5500 4496
rect 5356 3664 5408 3670
rect 5356 3606 5408 3612
rect 5552 3534 5580 5034
rect 5644 3641 5672 5222
rect 5736 4554 5764 5578
rect 5724 4548 5776 4554
rect 5724 4490 5776 4496
rect 5828 4486 5856 5714
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 5920 5012 5948 5646
rect 6012 5166 6040 6054
rect 6104 5166 6132 6122
rect 6288 5710 6316 6190
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 6210 5468 6518 5477
rect 6210 5466 6216 5468
rect 6272 5466 6296 5468
rect 6352 5466 6376 5468
rect 6432 5466 6456 5468
rect 6512 5466 6518 5468
rect 6272 5414 6274 5466
rect 6454 5414 6456 5466
rect 6210 5412 6216 5414
rect 6272 5412 6296 5414
rect 6352 5412 6376 5414
rect 6432 5412 6456 5414
rect 6512 5412 6518 5414
rect 6210 5403 6518 5412
rect 6564 5370 6592 6190
rect 6552 5364 6604 5370
rect 6552 5306 6604 5312
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 6092 5160 6144 5166
rect 6092 5102 6144 5108
rect 5920 4984 6040 5012
rect 5906 4856 5962 4865
rect 5906 4791 5962 4800
rect 5920 4690 5948 4791
rect 5908 4684 5960 4690
rect 5908 4626 5960 4632
rect 5816 4480 5868 4486
rect 5816 4422 5868 4428
rect 5630 3632 5686 3641
rect 5828 3602 5856 4422
rect 5920 4146 5948 4626
rect 6012 4622 6040 4984
rect 6104 4729 6132 5102
rect 6564 4826 6592 5306
rect 6552 4820 6604 4826
rect 6552 4762 6604 4768
rect 6656 4758 6684 7278
rect 6840 7002 6868 7890
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6734 6760 6790 6769
rect 6734 6695 6790 6704
rect 6748 5234 6776 6695
rect 6840 6458 6868 6938
rect 6932 6866 6960 8366
rect 7012 7948 7064 7954
rect 7012 7890 7064 7896
rect 7024 7546 7052 7890
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 7012 6724 7064 6730
rect 7116 6712 7144 8434
rect 7208 8090 7236 10542
rect 7300 10470 7328 11358
rect 9128 11212 9180 11218
rect 9128 11154 9180 11160
rect 8760 11144 8812 11150
rect 8760 11086 8812 11092
rect 7656 11008 7708 11014
rect 7656 10950 7708 10956
rect 7380 10668 7432 10674
rect 7380 10610 7432 10616
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7300 9722 7328 10066
rect 7288 9716 7340 9722
rect 7288 9658 7340 9664
rect 7392 9568 7420 10610
rect 7668 10470 7696 10950
rect 8116 10600 8168 10606
rect 8116 10542 8168 10548
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7656 10464 7708 10470
rect 7656 10406 7708 10412
rect 7472 10056 7524 10062
rect 7472 9998 7524 10004
rect 7300 9540 7420 9568
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7196 6928 7248 6934
rect 7194 6896 7196 6905
rect 7248 6896 7250 6905
rect 7194 6831 7250 6840
rect 7300 6798 7328 9540
rect 7380 9444 7432 9450
rect 7380 9386 7432 9392
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 7392 6730 7420 9386
rect 7484 9110 7512 9998
rect 7472 9104 7524 9110
rect 7472 9046 7524 9052
rect 7576 7018 7604 10406
rect 7668 9042 7696 10406
rect 7760 10364 8068 10373
rect 7760 10362 7766 10364
rect 7822 10362 7846 10364
rect 7902 10362 7926 10364
rect 7982 10362 8006 10364
rect 8062 10362 8068 10364
rect 7822 10310 7824 10362
rect 8004 10310 8006 10362
rect 7760 10308 7766 10310
rect 7822 10308 7846 10310
rect 7902 10308 7926 10310
rect 7982 10308 8006 10310
rect 8062 10308 8068 10310
rect 7760 10299 8068 10308
rect 7840 10056 7892 10062
rect 7840 9998 7892 10004
rect 7852 9926 7880 9998
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7760 9276 8068 9285
rect 7760 9274 7766 9276
rect 7822 9274 7846 9276
rect 7902 9274 7926 9276
rect 7982 9274 8006 9276
rect 8062 9274 8068 9276
rect 7822 9222 7824 9274
rect 8004 9222 8006 9274
rect 7760 9220 7766 9222
rect 7822 9220 7846 9222
rect 7902 9220 7926 9222
rect 7982 9220 8006 9222
rect 8062 9220 8068 9222
rect 7760 9211 8068 9220
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 7852 8498 7880 8978
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 7944 8430 7972 8910
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 7760 8188 8068 8197
rect 7760 8186 7766 8188
rect 7822 8186 7846 8188
rect 7902 8186 7926 8188
rect 7982 8186 8006 8188
rect 8062 8186 8068 8188
rect 7822 8134 7824 8186
rect 8004 8134 8006 8186
rect 7760 8132 7766 8134
rect 7822 8132 7846 8134
rect 7902 8132 7926 8134
rect 7982 8132 8006 8134
rect 8062 8132 8068 8134
rect 7760 8123 8068 8132
rect 7656 7948 7708 7954
rect 7656 7890 7708 7896
rect 7668 7546 7696 7890
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7484 6990 7604 7018
rect 7064 6684 7144 6712
rect 7380 6724 7432 6730
rect 7012 6666 7064 6672
rect 7380 6666 7432 6672
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 6840 6254 6868 6394
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6932 6066 6960 6598
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 6840 6038 6960 6066
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6748 4865 6776 5170
rect 6840 5030 6868 6038
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6734 4856 6790 4865
rect 6734 4791 6790 4800
rect 6644 4752 6696 4758
rect 6090 4720 6146 4729
rect 6644 4694 6696 4700
rect 6090 4655 6092 4664
rect 6144 4655 6146 4664
rect 6552 4684 6604 4690
rect 6092 4626 6144 4632
rect 6552 4626 6604 4632
rect 6000 4616 6052 4622
rect 6000 4558 6052 4564
rect 6012 4282 6040 4558
rect 6104 4486 6132 4626
rect 6092 4480 6144 4486
rect 6092 4422 6144 4428
rect 6210 4380 6518 4389
rect 6210 4378 6216 4380
rect 6272 4378 6296 4380
rect 6352 4378 6376 4380
rect 6432 4378 6456 4380
rect 6512 4378 6518 4380
rect 6272 4326 6274 4378
rect 6454 4326 6456 4378
rect 6210 4324 6216 4326
rect 6272 4324 6296 4326
rect 6352 4324 6376 4326
rect 6432 4324 6456 4326
rect 6512 4324 6518 4326
rect 6210 4315 6518 4324
rect 6000 4276 6052 4282
rect 6000 4218 6052 4224
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 6196 4049 6224 4082
rect 6182 4040 6238 4049
rect 6092 4004 6144 4010
rect 6564 4010 6592 4626
rect 6642 4312 6698 4321
rect 6642 4247 6698 4256
rect 6736 4276 6788 4282
rect 6656 4146 6684 4247
rect 6736 4218 6788 4224
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 6182 3975 6238 3984
rect 6552 4004 6604 4010
rect 6092 3946 6144 3952
rect 6552 3946 6604 3952
rect 5906 3768 5962 3777
rect 5906 3703 5962 3712
rect 5630 3567 5686 3576
rect 5816 3596 5868 3602
rect 5816 3538 5868 3544
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5920 3398 5948 3703
rect 6104 3534 6132 3946
rect 6748 3942 6776 4218
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6748 3602 6776 3878
rect 6552 3596 6604 3602
rect 6552 3538 6604 3544
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6092 3528 6144 3534
rect 6092 3470 6144 3476
rect 6000 3460 6052 3466
rect 6000 3402 6052 3408
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 5264 3392 5316 3398
rect 5264 3334 5316 3340
rect 5908 3392 5960 3398
rect 5908 3334 5960 3340
rect 4804 2916 4856 2922
rect 4804 2858 4856 2864
rect 4896 2916 4948 2922
rect 4896 2858 4948 2864
rect 4660 2748 4968 2757
rect 4660 2746 4666 2748
rect 4722 2746 4746 2748
rect 4802 2746 4826 2748
rect 4882 2746 4906 2748
rect 4962 2746 4968 2748
rect 4722 2694 4724 2746
rect 4904 2694 4906 2746
rect 4660 2692 4666 2694
rect 4722 2692 4746 2694
rect 4802 2692 4826 2694
rect 4882 2692 4906 2694
rect 4962 2692 4968 2694
rect 4660 2683 4968 2692
rect 4804 2304 4856 2310
rect 4804 2246 4856 2252
rect 4528 2100 4580 2106
rect 4528 2042 4580 2048
rect 4816 1902 4844 2246
rect 5000 1902 5028 3334
rect 6012 2990 6040 3402
rect 6104 3058 6132 3470
rect 6210 3292 6518 3301
rect 6210 3290 6216 3292
rect 6272 3290 6296 3292
rect 6352 3290 6376 3292
rect 6432 3290 6456 3292
rect 6512 3290 6518 3292
rect 6272 3238 6274 3290
rect 6454 3238 6456 3290
rect 6210 3236 6216 3238
rect 6272 3236 6296 3238
rect 6352 3236 6376 3238
rect 6432 3236 6456 3238
rect 6512 3236 6518 3238
rect 6210 3227 6518 3236
rect 6460 3120 6512 3126
rect 6182 3088 6238 3097
rect 6092 3052 6144 3058
rect 6460 3062 6512 3068
rect 6182 3023 6238 3032
rect 6092 2994 6144 3000
rect 6000 2984 6052 2990
rect 6000 2926 6052 2932
rect 6092 2916 6144 2922
rect 6092 2858 6144 2864
rect 5080 2848 5132 2854
rect 5080 2790 5132 2796
rect 5356 2848 5408 2854
rect 5356 2790 5408 2796
rect 5092 2378 5120 2790
rect 5368 2553 5396 2790
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 5354 2544 5410 2553
rect 5172 2508 5224 2514
rect 5224 2468 5304 2496
rect 5354 2479 5410 2488
rect 5172 2450 5224 2456
rect 5080 2372 5132 2378
rect 5080 2314 5132 2320
rect 5276 1902 5304 2468
rect 5448 2304 5500 2310
rect 5448 2246 5500 2252
rect 5460 2038 5488 2246
rect 5448 2032 5500 2038
rect 5448 1974 5500 1980
rect 4436 1896 4488 1902
rect 4436 1838 4488 1844
rect 4804 1896 4856 1902
rect 4804 1838 4856 1844
rect 4988 1896 5040 1902
rect 4988 1838 5040 1844
rect 5264 1896 5316 1902
rect 5264 1838 5316 1844
rect 4528 1828 4580 1834
rect 4528 1770 4580 1776
rect 5172 1828 5224 1834
rect 5172 1770 5224 1776
rect 4540 1562 4568 1770
rect 4660 1660 4968 1669
rect 4660 1658 4666 1660
rect 4722 1658 4746 1660
rect 4802 1658 4826 1660
rect 4882 1658 4906 1660
rect 4962 1658 4968 1660
rect 4722 1606 4724 1658
rect 4904 1606 4906 1658
rect 4660 1604 4666 1606
rect 4722 1604 4746 1606
rect 4802 1604 4826 1606
rect 4882 1604 4906 1606
rect 4962 1604 4968 1606
rect 4660 1595 4968 1604
rect 5184 1562 5212 1770
rect 5552 1766 5580 2586
rect 6000 2576 6052 2582
rect 6000 2518 6052 2524
rect 5724 2508 5776 2514
rect 5724 2450 5776 2456
rect 5736 1902 5764 2450
rect 5724 1896 5776 1902
rect 5724 1838 5776 1844
rect 5540 1760 5592 1766
rect 5540 1702 5592 1708
rect 5816 1760 5868 1766
rect 5816 1702 5868 1708
rect 3516 1556 3568 1562
rect 3516 1498 3568 1504
rect 4528 1556 4580 1562
rect 4528 1498 4580 1504
rect 5172 1556 5224 1562
rect 5172 1498 5224 1504
rect 2964 1420 3016 1426
rect 2964 1362 3016 1368
rect 5828 1358 5856 1702
rect 6012 1562 6040 2518
rect 6104 2514 6132 2858
rect 6196 2650 6224 3023
rect 6472 2650 6500 3062
rect 6184 2644 6236 2650
rect 6184 2586 6236 2592
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 6092 2508 6144 2514
rect 6092 2450 6144 2456
rect 6104 2038 6132 2450
rect 6564 2310 6592 3538
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 6552 2304 6604 2310
rect 6552 2246 6604 2252
rect 6210 2204 6518 2213
rect 6210 2202 6216 2204
rect 6272 2202 6296 2204
rect 6352 2202 6376 2204
rect 6432 2202 6456 2204
rect 6512 2202 6518 2204
rect 6272 2150 6274 2202
rect 6454 2150 6456 2202
rect 6210 2148 6216 2150
rect 6272 2148 6296 2150
rect 6352 2148 6376 2150
rect 6432 2148 6456 2150
rect 6512 2148 6518 2150
rect 6210 2139 6518 2148
rect 6564 2038 6592 2246
rect 6092 2032 6144 2038
rect 6092 1974 6144 1980
rect 6552 2032 6604 2038
rect 6552 1974 6604 1980
rect 6000 1556 6052 1562
rect 6000 1498 6052 1504
rect 5816 1352 5868 1358
rect 5816 1294 5868 1300
rect 3110 1116 3418 1125
rect 3110 1114 3116 1116
rect 3172 1114 3196 1116
rect 3252 1114 3276 1116
rect 3332 1114 3356 1116
rect 3412 1114 3418 1116
rect 3172 1062 3174 1114
rect 3354 1062 3356 1114
rect 3110 1060 3116 1062
rect 3172 1060 3196 1062
rect 3252 1060 3276 1062
rect 3332 1060 3356 1062
rect 3412 1060 3418 1062
rect 3110 1051 3418 1060
rect 6012 950 6040 1498
rect 6092 1420 6144 1426
rect 6092 1362 6144 1368
rect 6104 1018 6132 1362
rect 6210 1116 6518 1125
rect 6210 1114 6216 1116
rect 6272 1114 6296 1116
rect 6352 1114 6376 1116
rect 6432 1114 6456 1116
rect 6512 1114 6518 1116
rect 6272 1062 6274 1114
rect 6454 1062 6456 1114
rect 6210 1060 6216 1062
rect 6272 1060 6296 1062
rect 6352 1060 6376 1062
rect 6432 1060 6456 1062
rect 6512 1060 6518 1062
rect 6210 1051 6518 1060
rect 6092 1012 6144 1018
rect 6092 954 6144 960
rect 6000 944 6052 950
rect 6000 886 6052 892
rect 6656 882 6684 3470
rect 6748 3126 6776 3538
rect 6840 3398 6868 4082
rect 6828 3392 6880 3398
rect 6826 3360 6828 3369
rect 6880 3360 6882 3369
rect 6826 3295 6882 3304
rect 6736 3120 6788 3126
rect 6736 3062 6788 3068
rect 6734 2952 6790 2961
rect 6734 2887 6790 2896
rect 6748 2854 6776 2887
rect 6736 2848 6788 2854
rect 6736 2790 6788 2796
rect 6748 1970 6776 2790
rect 6932 2774 6960 5850
rect 7102 5808 7158 5817
rect 7102 5743 7158 5752
rect 7012 5636 7064 5642
rect 7012 5578 7064 5584
rect 7024 5234 7052 5578
rect 7012 5228 7064 5234
rect 7116 5216 7144 5743
rect 7208 5370 7236 6258
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 7116 5188 7236 5216
rect 7012 5170 7064 5176
rect 7024 5098 7052 5170
rect 7012 5092 7064 5098
rect 7012 5034 7064 5040
rect 7104 5092 7156 5098
rect 7104 5034 7156 5040
rect 7024 4826 7052 5034
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 7116 3584 7144 5034
rect 7208 4690 7236 5188
rect 7300 5166 7328 6598
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7392 5778 7420 6054
rect 7380 5772 7432 5778
rect 7380 5714 7432 5720
rect 7288 5160 7340 5166
rect 7288 5102 7340 5108
rect 7288 5024 7340 5030
rect 7288 4966 7340 4972
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7196 4684 7248 4690
rect 7196 4626 7248 4632
rect 7208 4146 7236 4626
rect 7196 4140 7248 4146
rect 7196 4082 7248 4088
rect 7196 3596 7248 3602
rect 7116 3556 7196 3584
rect 7196 3538 7248 3544
rect 7104 3460 7156 3466
rect 7104 3402 7156 3408
rect 7012 2916 7064 2922
rect 7012 2858 7064 2864
rect 6840 2746 6960 2774
rect 6840 2689 6868 2746
rect 6826 2680 6882 2689
rect 6826 2615 6882 2624
rect 7024 1970 7052 2858
rect 6736 1964 6788 1970
rect 7012 1964 7064 1970
rect 6736 1906 6788 1912
rect 6932 1924 7012 1952
rect 6932 1358 6960 1924
rect 7012 1906 7064 1912
rect 7012 1488 7064 1494
rect 7012 1430 7064 1436
rect 6920 1352 6972 1358
rect 6920 1294 6972 1300
rect 6644 876 6696 882
rect 6644 818 6696 824
rect 7024 814 7052 1430
rect 7116 1358 7144 3402
rect 7208 2922 7236 3538
rect 7300 3534 7328 4966
rect 7392 3777 7420 4966
rect 7378 3768 7434 3777
rect 7378 3703 7434 3712
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 7378 3224 7434 3233
rect 7484 3194 7512 6990
rect 7668 6882 7696 7346
rect 7760 7100 8068 7109
rect 7760 7098 7766 7100
rect 7822 7098 7846 7100
rect 7902 7098 7926 7100
rect 7982 7098 8006 7100
rect 8062 7098 8068 7100
rect 7822 7046 7824 7098
rect 8004 7046 8006 7098
rect 7760 7044 7766 7046
rect 7822 7044 7846 7046
rect 7902 7044 7926 7046
rect 7982 7044 8006 7046
rect 8062 7044 8068 7046
rect 7760 7035 8068 7044
rect 7564 6860 7616 6866
rect 7668 6854 7788 6882
rect 7760 6848 7788 6854
rect 7840 6860 7892 6866
rect 7760 6820 7840 6848
rect 7564 6802 7616 6808
rect 7840 6802 7892 6808
rect 7932 6860 7984 6866
rect 7932 6802 7984 6808
rect 7576 3194 7604 6802
rect 7944 6769 7972 6802
rect 7930 6760 7986 6769
rect 7656 6724 7708 6730
rect 7930 6695 7986 6704
rect 7656 6666 7708 6672
rect 7668 6186 7696 6666
rect 7656 6180 7708 6186
rect 7656 6122 7708 6128
rect 7760 6012 8068 6021
rect 7760 6010 7766 6012
rect 7822 6010 7846 6012
rect 7902 6010 7926 6012
rect 7982 6010 8006 6012
rect 8062 6010 8068 6012
rect 7822 5958 7824 6010
rect 8004 5958 8006 6010
rect 7760 5956 7766 5958
rect 7822 5956 7846 5958
rect 7902 5956 7926 5958
rect 7982 5956 8006 5958
rect 8062 5956 8068 5958
rect 7760 5947 8068 5956
rect 7930 5808 7986 5817
rect 7748 5772 7800 5778
rect 7930 5743 7932 5752
rect 7748 5714 7800 5720
rect 7984 5743 7986 5752
rect 7932 5714 7984 5720
rect 7656 5568 7708 5574
rect 7656 5510 7708 5516
rect 7668 4758 7696 5510
rect 7760 5302 7788 5714
rect 7840 5636 7892 5642
rect 7840 5578 7892 5584
rect 7852 5370 7880 5578
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 7748 5296 7800 5302
rect 7748 5238 7800 5244
rect 7944 5030 7972 5714
rect 8128 5658 8156 10542
rect 8220 10470 8248 10542
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8208 10192 8260 10198
rect 8260 10152 8340 10180
rect 8208 10134 8260 10140
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8220 6322 8248 9522
rect 8312 9382 8340 10152
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8404 9654 8432 9862
rect 8680 9654 8708 9862
rect 8772 9654 8800 11086
rect 9140 10470 9168 11154
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 9232 10742 9260 11086
rect 9310 10908 9618 10917
rect 9310 10906 9316 10908
rect 9372 10906 9396 10908
rect 9452 10906 9476 10908
rect 9532 10906 9556 10908
rect 9612 10906 9618 10908
rect 9372 10854 9374 10906
rect 9554 10854 9556 10906
rect 9310 10852 9316 10854
rect 9372 10852 9396 10854
rect 9452 10852 9476 10854
rect 9532 10852 9556 10854
rect 9612 10852 9618 10854
rect 9310 10843 9618 10852
rect 9692 10742 9720 11358
rect 9772 11280 9824 11286
rect 9772 11222 9824 11228
rect 9784 10810 9812 11222
rect 9954 11200 10010 12000
rect 12256 11212 12308 11218
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9220 10736 9272 10742
rect 9680 10736 9732 10742
rect 9220 10678 9272 10684
rect 9310 10704 9366 10713
rect 9232 10606 9260 10678
rect 9680 10678 9732 10684
rect 9310 10639 9366 10648
rect 9324 10606 9352 10639
rect 9220 10600 9272 10606
rect 9220 10542 9272 10548
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 9968 10554 9996 11200
rect 12806 11200 12862 12000
rect 12912 11206 13216 11234
rect 12256 11154 12308 11160
rect 12164 11144 12216 11150
rect 12164 11086 12216 11092
rect 11888 11076 11940 11082
rect 11888 11018 11940 11024
rect 11900 10810 11928 11018
rect 12072 11008 12124 11014
rect 12072 10950 12124 10956
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 11980 10804 12032 10810
rect 11980 10746 12032 10752
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 10152 10577 10180 10610
rect 10138 10568 10194 10577
rect 9772 10532 9824 10538
rect 9968 10526 10088 10554
rect 9772 10474 9824 10480
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 8392 9648 8444 9654
rect 8392 9590 8444 9596
rect 8668 9648 8720 9654
rect 8668 9590 8720 9596
rect 8760 9648 8812 9654
rect 8760 9590 8812 9596
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 8680 9178 8708 9590
rect 8668 9172 8720 9178
rect 8668 9114 8720 9120
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 8312 7954 8340 8502
rect 9036 8424 9088 8430
rect 9036 8366 9088 8372
rect 8852 8356 8904 8362
rect 8852 8298 8904 8304
rect 8392 8016 8444 8022
rect 8392 7958 8444 7964
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8300 7268 8352 7274
rect 8300 7210 8352 7216
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 8220 5914 8248 6258
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 8128 5630 8248 5658
rect 8220 5574 8248 5630
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 7760 4924 8068 4933
rect 7760 4922 7766 4924
rect 7822 4922 7846 4924
rect 7902 4922 7926 4924
rect 7982 4922 8006 4924
rect 8062 4922 8068 4924
rect 7822 4870 7824 4922
rect 8004 4870 8006 4922
rect 7760 4868 7766 4870
rect 7822 4868 7846 4870
rect 7902 4868 7926 4870
rect 7982 4868 8006 4870
rect 8062 4868 8068 4870
rect 7760 4859 8068 4868
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 7656 4752 7708 4758
rect 7656 4694 7708 4700
rect 7656 4548 7708 4554
rect 7656 4490 7708 4496
rect 7668 3398 7696 4490
rect 7760 4078 7788 4762
rect 7932 4752 7984 4758
rect 7932 4694 7984 4700
rect 7944 4078 7972 4694
rect 7748 4072 7800 4078
rect 7748 4014 7800 4020
rect 7932 4072 7984 4078
rect 8024 4072 8076 4078
rect 7932 4014 7984 4020
rect 8022 4040 8024 4049
rect 8076 4040 8078 4049
rect 8022 3975 8078 3984
rect 8128 3942 8156 5170
rect 8208 5092 8260 5098
rect 8208 5034 8260 5040
rect 8220 4321 8248 5034
rect 8206 4312 8262 4321
rect 8206 4247 8262 4256
rect 8312 4214 8340 7210
rect 8404 6866 8432 7958
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8300 4208 8352 4214
rect 8300 4150 8352 4156
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 7760 3836 8068 3845
rect 7760 3834 7766 3836
rect 7822 3834 7846 3836
rect 7902 3834 7926 3836
rect 7982 3834 8006 3836
rect 8062 3834 8068 3836
rect 7822 3782 7824 3834
rect 8004 3782 8006 3834
rect 7760 3780 7766 3782
rect 7822 3780 7846 3782
rect 7902 3780 7926 3782
rect 7982 3780 8006 3782
rect 8062 3780 8068 3782
rect 7760 3771 8068 3780
rect 8220 3738 8248 3878
rect 8116 3732 8168 3738
rect 7760 3692 8116 3720
rect 7760 3602 7788 3692
rect 8116 3674 8168 3680
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 8312 3670 8340 4014
rect 8404 3942 8432 6598
rect 8496 5778 8524 7686
rect 8864 7342 8892 8298
rect 8944 7472 8996 7478
rect 8944 7414 8996 7420
rect 8852 7336 8904 7342
rect 8852 7278 8904 7284
rect 8760 6996 8812 7002
rect 8760 6938 8812 6944
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 8588 5914 8616 6802
rect 8772 6798 8800 6938
rect 8864 6866 8892 7278
rect 8956 6934 8984 7414
rect 9048 7342 9076 8366
rect 9140 7818 9168 10406
rect 9508 10198 9536 10406
rect 9496 10192 9548 10198
rect 9496 10134 9548 10140
rect 9680 10056 9732 10062
rect 9586 10024 9642 10033
rect 9680 9998 9732 10004
rect 9586 9959 9642 9968
rect 9600 9926 9628 9959
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 9310 9820 9618 9829
rect 9310 9818 9316 9820
rect 9372 9818 9396 9820
rect 9452 9818 9476 9820
rect 9532 9818 9556 9820
rect 9612 9818 9618 9820
rect 9372 9766 9374 9818
rect 9554 9766 9556 9818
rect 9310 9764 9316 9766
rect 9372 9764 9396 9766
rect 9452 9764 9476 9766
rect 9532 9764 9556 9766
rect 9612 9764 9618 9766
rect 9310 9755 9618 9764
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9508 9382 9536 9522
rect 9496 9376 9548 9382
rect 9496 9318 9548 9324
rect 9310 8732 9618 8741
rect 9310 8730 9316 8732
rect 9372 8730 9396 8732
rect 9452 8730 9476 8732
rect 9532 8730 9556 8732
rect 9612 8730 9618 8732
rect 9372 8678 9374 8730
rect 9554 8678 9556 8730
rect 9310 8676 9316 8678
rect 9372 8676 9396 8678
rect 9452 8676 9476 8678
rect 9532 8676 9556 8678
rect 9612 8676 9618 8678
rect 9310 8667 9618 8676
rect 9692 8634 9720 9998
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9784 8106 9812 10474
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 9864 10124 9916 10130
rect 9864 10066 9916 10072
rect 9876 9586 9904 10066
rect 9864 9580 9916 9586
rect 9864 9522 9916 9528
rect 9864 9376 9916 9382
rect 9864 9318 9916 9324
rect 9876 8922 9904 9318
rect 9968 9110 9996 10406
rect 9956 9104 10008 9110
rect 9956 9046 10008 9052
rect 9876 8894 9996 8922
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 9692 8090 9812 8106
rect 9692 8084 9824 8090
rect 9692 8078 9772 8084
rect 9128 7812 9180 7818
rect 9128 7754 9180 7760
rect 9310 7644 9618 7653
rect 9310 7642 9316 7644
rect 9372 7642 9396 7644
rect 9452 7642 9476 7644
rect 9532 7642 9556 7644
rect 9612 7642 9618 7644
rect 9372 7590 9374 7642
rect 9554 7590 9556 7642
rect 9310 7588 9316 7590
rect 9372 7588 9396 7590
rect 9452 7588 9476 7590
rect 9532 7588 9556 7590
rect 9612 7588 9618 7590
rect 9310 7579 9618 7588
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 8944 6928 8996 6934
rect 8944 6870 8996 6876
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 8668 6384 8720 6390
rect 8668 6326 8720 6332
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8484 5772 8536 5778
rect 8484 5714 8536 5720
rect 8484 5364 8536 5370
rect 8484 5306 8536 5312
rect 8496 4758 8524 5306
rect 8680 4826 8708 6326
rect 8772 5710 8800 6734
rect 8852 6656 8904 6662
rect 8852 6598 8904 6604
rect 8944 6656 8996 6662
rect 8944 6598 8996 6604
rect 8864 6390 8892 6598
rect 8852 6384 8904 6390
rect 8852 6326 8904 6332
rect 8852 6248 8904 6254
rect 8852 6190 8904 6196
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 8864 5370 8892 6190
rect 8852 5364 8904 5370
rect 8852 5306 8904 5312
rect 8852 5228 8904 5234
rect 8852 5170 8904 5176
rect 8668 4820 8720 4826
rect 8668 4762 8720 4768
rect 8484 4752 8536 4758
rect 8484 4694 8536 4700
rect 8864 4690 8892 5170
rect 8852 4684 8904 4690
rect 8852 4626 8904 4632
rect 8484 4616 8536 4622
rect 8484 4558 8536 4564
rect 8392 3936 8444 3942
rect 8392 3878 8444 3884
rect 8496 3754 8524 4558
rect 8576 4548 8628 4554
rect 8576 4490 8628 4496
rect 8588 3942 8616 4490
rect 8956 4146 8984 6598
rect 9048 5710 9076 7278
rect 9416 7002 9444 7346
rect 9496 7268 9548 7274
rect 9496 7210 9548 7216
rect 9404 6996 9456 7002
rect 9404 6938 9456 6944
rect 9508 6866 9536 7210
rect 9692 7002 9720 8078
rect 9772 8026 9824 8032
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 9784 7478 9812 7890
rect 9876 7750 9904 8774
rect 9864 7744 9916 7750
rect 9864 7686 9916 7692
rect 9772 7472 9824 7478
rect 9772 7414 9824 7420
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9876 6866 9904 7686
rect 9220 6860 9272 6866
rect 9220 6802 9272 6808
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9232 6440 9260 6802
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9310 6556 9618 6565
rect 9310 6554 9316 6556
rect 9372 6554 9396 6556
rect 9452 6554 9476 6556
rect 9532 6554 9556 6556
rect 9612 6554 9618 6556
rect 9372 6502 9374 6554
rect 9554 6502 9556 6554
rect 9310 6500 9316 6502
rect 9372 6500 9396 6502
rect 9452 6500 9476 6502
rect 9532 6500 9556 6502
rect 9612 6500 9618 6502
rect 9310 6491 9618 6500
rect 9680 6452 9732 6458
rect 9232 6412 9444 6440
rect 9128 6180 9180 6186
rect 9128 6122 9180 6128
rect 9140 5846 9168 6122
rect 9220 6112 9272 6118
rect 9220 6054 9272 6060
rect 9128 5840 9180 5846
rect 9128 5782 9180 5788
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 9036 5160 9088 5166
rect 9036 5102 9088 5108
rect 9048 4826 9076 5102
rect 9036 4820 9088 4826
rect 9036 4762 9088 4768
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 9036 4072 9088 4078
rect 9036 4014 9088 4020
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 8496 3726 8616 3754
rect 8680 3738 8708 4014
rect 8300 3664 8352 3670
rect 7838 3632 7894 3641
rect 7748 3596 7800 3602
rect 8114 3632 8170 3641
rect 7838 3567 7894 3576
rect 7932 3596 7984 3602
rect 7748 3538 7800 3544
rect 7656 3392 7708 3398
rect 7656 3334 7708 3340
rect 7378 3159 7434 3168
rect 7472 3188 7524 3194
rect 7392 3126 7420 3159
rect 7472 3130 7524 3136
rect 7564 3188 7616 3194
rect 7564 3130 7616 3136
rect 7380 3120 7432 3126
rect 7380 3062 7432 3068
rect 7760 2990 7788 3538
rect 7852 2990 7880 3567
rect 7984 3576 8114 3584
rect 8352 3624 8432 3652
rect 8300 3606 8352 3612
rect 7984 3567 8170 3576
rect 7984 3556 8156 3567
rect 7932 3538 7984 3544
rect 8128 3516 8156 3556
rect 8128 3488 8248 3516
rect 8024 3392 8076 3398
rect 7930 3360 7986 3369
rect 8024 3334 8076 3340
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 7930 3295 7986 3304
rect 7944 3126 7972 3295
rect 7932 3120 7984 3126
rect 7932 3062 7984 3068
rect 7472 2984 7524 2990
rect 7748 2984 7800 2990
rect 7472 2926 7524 2932
rect 7668 2944 7748 2972
rect 7196 2916 7248 2922
rect 7196 2858 7248 2864
rect 7208 2650 7236 2858
rect 7484 2854 7512 2926
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 7286 2680 7342 2689
rect 7196 2644 7248 2650
rect 7286 2615 7342 2624
rect 7196 2586 7248 2592
rect 7300 2378 7328 2615
rect 7380 2440 7432 2446
rect 7484 2428 7512 2790
rect 7432 2400 7512 2428
rect 7380 2382 7432 2388
rect 7288 2372 7340 2378
rect 7288 2314 7340 2320
rect 7196 2100 7248 2106
rect 7196 2042 7248 2048
rect 7208 1766 7236 2042
rect 7484 1766 7512 2400
rect 7668 2106 7696 2944
rect 7748 2926 7800 2932
rect 7840 2984 7892 2990
rect 7840 2926 7892 2932
rect 7944 2854 7972 3062
rect 8036 2904 8064 3334
rect 8128 3233 8156 3334
rect 8114 3224 8170 3233
rect 8114 3159 8170 3168
rect 8114 3088 8170 3097
rect 8114 3023 8116 3032
rect 8168 3023 8170 3032
rect 8116 2994 8168 3000
rect 8036 2876 8156 2904
rect 7932 2848 7984 2854
rect 7932 2790 7984 2796
rect 7760 2748 8068 2757
rect 7760 2746 7766 2748
rect 7822 2746 7846 2748
rect 7902 2746 7926 2748
rect 7982 2746 8006 2748
rect 8062 2746 8068 2748
rect 7822 2694 7824 2746
rect 8004 2694 8006 2746
rect 7760 2692 7766 2694
rect 7822 2692 7846 2694
rect 7902 2692 7926 2694
rect 7982 2692 8006 2694
rect 8062 2692 8068 2694
rect 7760 2683 8068 2692
rect 8128 2553 8156 2876
rect 8220 2802 8248 3488
rect 8300 3120 8352 3126
rect 8404 3097 8432 3624
rect 8588 3398 8616 3726
rect 8668 3732 8720 3738
rect 8668 3674 8720 3680
rect 8760 3664 8812 3670
rect 8680 3612 8760 3618
rect 8680 3606 8812 3612
rect 8680 3590 8800 3606
rect 8852 3596 8904 3602
rect 8484 3392 8536 3398
rect 8484 3334 8536 3340
rect 8576 3392 8628 3398
rect 8576 3334 8628 3340
rect 8496 3194 8524 3334
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8300 3062 8352 3068
rect 8390 3088 8446 3097
rect 8312 2922 8340 3062
rect 8390 3023 8446 3032
rect 8588 2990 8616 3334
rect 8680 3058 8708 3590
rect 8852 3538 8904 3544
rect 8944 3596 8996 3602
rect 8944 3538 8996 3544
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 8392 2984 8444 2990
rect 8392 2926 8444 2932
rect 8576 2984 8628 2990
rect 8576 2926 8628 2932
rect 8300 2916 8352 2922
rect 8300 2858 8352 2864
rect 8220 2774 8340 2802
rect 8114 2544 8170 2553
rect 8114 2479 8170 2488
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 7656 2100 7708 2106
rect 7656 2042 7708 2048
rect 7760 1986 7788 2382
rect 8208 2100 8260 2106
rect 8208 2042 8260 2048
rect 7576 1958 7788 1986
rect 7196 1760 7248 1766
rect 7196 1702 7248 1708
rect 7472 1760 7524 1766
rect 7472 1702 7524 1708
rect 7104 1352 7156 1358
rect 7104 1294 7156 1300
rect 7208 1222 7236 1702
rect 7576 1562 7604 1958
rect 7656 1896 7708 1902
rect 7656 1838 7708 1844
rect 7668 1562 7696 1838
rect 7760 1660 8068 1669
rect 7760 1658 7766 1660
rect 7822 1658 7846 1660
rect 7902 1658 7926 1660
rect 7982 1658 8006 1660
rect 8062 1658 8068 1660
rect 7822 1606 7824 1658
rect 8004 1606 8006 1658
rect 7760 1604 7766 1606
rect 7822 1604 7846 1606
rect 7902 1604 7926 1606
rect 7982 1604 8006 1606
rect 8062 1604 8068 1606
rect 7760 1595 8068 1604
rect 7564 1556 7616 1562
rect 7564 1498 7616 1504
rect 7656 1556 7708 1562
rect 7656 1498 7708 1504
rect 8220 1426 8248 2042
rect 8312 1562 8340 2774
rect 8300 1556 8352 1562
rect 8300 1498 8352 1504
rect 8208 1420 8260 1426
rect 8208 1362 8260 1368
rect 8300 1420 8352 1426
rect 8300 1362 8352 1368
rect 7196 1216 7248 1222
rect 7196 1158 7248 1164
rect 8312 1018 8340 1362
rect 8404 1358 8432 2926
rect 8668 2848 8720 2854
rect 8668 2790 8720 2796
rect 8482 2680 8538 2689
rect 8482 2615 8538 2624
rect 8496 1358 8524 2615
rect 8680 2394 8708 2790
rect 8772 2650 8800 3470
rect 8864 3346 8892 3538
rect 8956 3505 8984 3538
rect 8942 3496 8998 3505
rect 8942 3431 8998 3440
rect 8864 3318 8984 3346
rect 8956 3058 8984 3318
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 8850 2952 8906 2961
rect 8850 2887 8852 2896
rect 8904 2887 8906 2896
rect 8852 2858 8904 2864
rect 8956 2689 8984 2994
rect 8942 2680 8998 2689
rect 8760 2644 8812 2650
rect 9048 2650 9076 4014
rect 9140 3670 9168 5782
rect 9232 5234 9260 6054
rect 9416 5778 9444 6412
rect 9680 6394 9732 6400
rect 9692 5846 9720 6394
rect 9680 5840 9732 5846
rect 9680 5782 9732 5788
rect 9404 5772 9456 5778
rect 9404 5714 9456 5720
rect 9416 5681 9444 5714
rect 9402 5672 9458 5681
rect 9402 5607 9458 5616
rect 9310 5468 9618 5477
rect 9310 5466 9316 5468
rect 9372 5466 9396 5468
rect 9452 5466 9476 5468
rect 9532 5466 9556 5468
rect 9612 5466 9618 5468
rect 9372 5414 9374 5466
rect 9554 5414 9556 5466
rect 9310 5412 9316 5414
rect 9372 5412 9396 5414
rect 9452 5412 9476 5414
rect 9532 5412 9556 5414
rect 9612 5412 9618 5414
rect 9310 5403 9618 5412
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 9600 4690 9628 5170
rect 9220 4684 9272 4690
rect 9220 4626 9272 4632
rect 9588 4684 9640 4690
rect 9588 4626 9640 4632
rect 9232 4282 9260 4626
rect 9310 4380 9618 4389
rect 9310 4378 9316 4380
rect 9372 4378 9396 4380
rect 9452 4378 9476 4380
rect 9532 4378 9556 4380
rect 9612 4378 9618 4380
rect 9372 4326 9374 4378
rect 9554 4326 9556 4378
rect 9310 4324 9316 4326
rect 9372 4324 9396 4326
rect 9452 4324 9476 4326
rect 9532 4324 9556 4326
rect 9612 4324 9618 4326
rect 9310 4315 9618 4324
rect 9220 4276 9272 4282
rect 9220 4218 9272 4224
rect 9784 4010 9812 6734
rect 9968 5914 9996 8894
rect 10060 8090 10088 10526
rect 10138 10503 10194 10512
rect 10140 10464 10192 10470
rect 10140 10406 10192 10412
rect 10152 10266 10180 10406
rect 10140 10260 10192 10266
rect 10140 10202 10192 10208
rect 10138 10160 10194 10169
rect 10138 10095 10194 10104
rect 10152 10062 10180 10095
rect 10140 10056 10192 10062
rect 10140 9998 10192 10004
rect 10414 10024 10470 10033
rect 10414 9959 10470 9968
rect 10232 9920 10284 9926
rect 10232 9862 10284 9868
rect 10244 8974 10272 9862
rect 10428 9450 10456 9959
rect 10612 9654 10640 10610
rect 11520 10600 11572 10606
rect 11520 10542 11572 10548
rect 11888 10600 11940 10606
rect 11888 10542 11940 10548
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 10860 10364 11168 10373
rect 10860 10362 10866 10364
rect 10922 10362 10946 10364
rect 11002 10362 11026 10364
rect 11082 10362 11106 10364
rect 11162 10362 11168 10364
rect 10922 10310 10924 10362
rect 11104 10310 11106 10362
rect 10860 10308 10866 10310
rect 10922 10308 10946 10310
rect 11002 10308 11026 10310
rect 11082 10308 11106 10310
rect 11162 10308 11168 10310
rect 10860 10299 11168 10308
rect 11348 10062 11376 10406
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 10784 9920 10836 9926
rect 10784 9862 10836 9868
rect 10796 9654 10824 9862
rect 10600 9648 10652 9654
rect 10600 9590 10652 9596
rect 10784 9648 10836 9654
rect 10784 9590 10836 9596
rect 11348 9518 11376 9998
rect 11336 9512 11388 9518
rect 11336 9454 11388 9460
rect 10416 9444 10468 9450
rect 10416 9386 10468 9392
rect 11244 9444 11296 9450
rect 11244 9386 11296 9392
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10796 9110 10824 9318
rect 10860 9276 11168 9285
rect 10860 9274 10866 9276
rect 10922 9274 10946 9276
rect 11002 9274 11026 9276
rect 11082 9274 11106 9276
rect 11162 9274 11168 9276
rect 10922 9222 10924 9274
rect 11104 9222 11106 9274
rect 10860 9220 10866 9222
rect 10922 9220 10946 9222
rect 11002 9220 11026 9222
rect 11082 9220 11106 9222
rect 11162 9220 11168 9222
rect 10860 9211 11168 9220
rect 10784 9104 10836 9110
rect 10784 9046 10836 9052
rect 11256 8974 11284 9386
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10612 8430 10640 8570
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10782 8392 10838 8401
rect 10782 8327 10784 8336
rect 10836 8327 10838 8336
rect 10784 8298 10836 8304
rect 10140 8288 10192 8294
rect 10140 8230 10192 8236
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 10152 7546 10180 8230
rect 10860 8188 11168 8197
rect 10860 8186 10866 8188
rect 10922 8186 10946 8188
rect 11002 8186 11026 8188
rect 11082 8186 11106 8188
rect 11162 8186 11168 8188
rect 10922 8134 10924 8186
rect 11104 8134 11106 8186
rect 10860 8132 10866 8134
rect 10922 8132 10946 8134
rect 11002 8132 11026 8134
rect 11082 8132 11106 8134
rect 11162 8132 11168 8134
rect 10860 8123 11168 8132
rect 11348 7546 11376 9454
rect 11428 9172 11480 9178
rect 11428 9114 11480 9120
rect 11440 8430 11468 9114
rect 11532 9110 11560 10542
rect 11900 10198 11928 10542
rect 11888 10192 11940 10198
rect 11992 10169 12020 10746
rect 12084 10606 12112 10950
rect 12176 10674 12204 11086
rect 12164 10668 12216 10674
rect 12164 10610 12216 10616
rect 12268 10606 12296 11154
rect 12820 11132 12848 11200
rect 12912 11132 12940 11206
rect 12820 11104 12940 11132
rect 12410 10908 12718 10917
rect 12410 10906 12416 10908
rect 12472 10906 12496 10908
rect 12552 10906 12576 10908
rect 12632 10906 12656 10908
rect 12712 10906 12718 10908
rect 12472 10854 12474 10906
rect 12654 10854 12656 10906
rect 12410 10852 12416 10854
rect 12472 10852 12496 10854
rect 12552 10852 12576 10854
rect 12632 10852 12656 10854
rect 12712 10852 12718 10854
rect 12410 10843 12718 10852
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 12072 10600 12124 10606
rect 12072 10542 12124 10548
rect 12256 10600 12308 10606
rect 12256 10542 12308 10548
rect 12808 10600 12860 10606
rect 12808 10542 12860 10548
rect 12164 10532 12216 10538
rect 12164 10474 12216 10480
rect 12440 10532 12492 10538
rect 12440 10474 12492 10480
rect 11888 10134 11940 10140
rect 11978 10160 12034 10169
rect 11978 10095 12034 10104
rect 11796 9988 11848 9994
rect 11796 9930 11848 9936
rect 11520 9104 11572 9110
rect 11520 9046 11572 9052
rect 11428 8424 11480 8430
rect 11428 8366 11480 8372
rect 11520 8288 11572 8294
rect 11520 8230 11572 8236
rect 11532 7750 11560 8230
rect 11704 8016 11756 8022
rect 11702 7984 11704 7993
rect 11756 7984 11758 7993
rect 11808 7954 11836 9930
rect 12176 9926 12204 10474
rect 12452 10130 12480 10474
rect 12256 10124 12308 10130
rect 12256 10066 12308 10072
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12268 9926 12296 10066
rect 12164 9920 12216 9926
rect 12164 9862 12216 9868
rect 12256 9920 12308 9926
rect 12256 9862 12308 9868
rect 12268 9382 12296 9862
rect 12410 9820 12718 9829
rect 12410 9818 12416 9820
rect 12472 9818 12496 9820
rect 12552 9818 12576 9820
rect 12632 9818 12656 9820
rect 12712 9818 12718 9820
rect 12472 9766 12474 9818
rect 12654 9766 12656 9818
rect 12410 9764 12416 9766
rect 12472 9764 12496 9766
rect 12552 9764 12576 9766
rect 12632 9764 12656 9766
rect 12712 9764 12718 9766
rect 12410 9755 12718 9764
rect 12256 9376 12308 9382
rect 12176 9324 12256 9330
rect 12176 9318 12308 9324
rect 12176 9302 12296 9318
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 11888 8968 11940 8974
rect 11888 8910 11940 8916
rect 11702 7919 11758 7928
rect 11796 7948 11848 7954
rect 11796 7890 11848 7896
rect 11520 7744 11572 7750
rect 11520 7686 11572 7692
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 11336 7540 11388 7546
rect 11336 7482 11388 7488
rect 10152 6934 10180 7482
rect 11808 7410 11836 7890
rect 11900 7818 11928 8910
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 11992 8022 12020 8774
rect 12084 8294 12112 8978
rect 12176 8362 12204 9302
rect 12410 8732 12718 8741
rect 12410 8730 12416 8732
rect 12472 8730 12496 8732
rect 12552 8730 12576 8732
rect 12632 8730 12656 8732
rect 12712 8730 12718 8732
rect 12472 8678 12474 8730
rect 12654 8678 12656 8730
rect 12410 8676 12416 8678
rect 12472 8676 12496 8678
rect 12552 8676 12576 8678
rect 12632 8676 12656 8678
rect 12712 8676 12718 8678
rect 12410 8667 12718 8676
rect 12256 8560 12308 8566
rect 12256 8502 12308 8508
rect 12164 8356 12216 8362
rect 12164 8298 12216 8304
rect 12072 8288 12124 8294
rect 12072 8230 12124 8236
rect 11980 8016 12032 8022
rect 11980 7958 12032 7964
rect 12084 7954 12112 8230
rect 12176 7993 12204 8298
rect 12162 7984 12218 7993
rect 12072 7948 12124 7954
rect 12162 7919 12218 7928
rect 12072 7890 12124 7896
rect 11888 7812 11940 7818
rect 11888 7754 11940 7760
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 10416 7336 10468 7342
rect 10414 7304 10416 7313
rect 10468 7304 10470 7313
rect 10414 7239 10470 7248
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 10860 7100 11168 7109
rect 10860 7098 10866 7100
rect 10922 7098 10946 7100
rect 11002 7098 11026 7100
rect 11082 7098 11106 7100
rect 11162 7098 11168 7100
rect 10922 7046 10924 7098
rect 11104 7046 11106 7098
rect 10860 7044 10866 7046
rect 10922 7044 10946 7046
rect 11002 7044 11026 7046
rect 11082 7044 11106 7046
rect 11162 7044 11168 7046
rect 10860 7035 11168 7044
rect 10324 6996 10376 7002
rect 10324 6938 10376 6944
rect 10140 6928 10192 6934
rect 10046 6896 10102 6905
rect 10140 6870 10192 6876
rect 10046 6831 10102 6840
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 10060 5846 10088 6831
rect 10048 5840 10100 5846
rect 10048 5782 10100 5788
rect 10232 5364 10284 5370
rect 10232 5306 10284 5312
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 9876 4622 9904 4966
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 9864 4616 9916 4622
rect 9864 4558 9916 4564
rect 9772 4004 9824 4010
rect 9772 3946 9824 3952
rect 9784 3720 9812 3946
rect 9692 3692 9812 3720
rect 9128 3664 9180 3670
rect 9128 3606 9180 3612
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 9220 3392 9272 3398
rect 9220 3334 9272 3340
rect 8942 2615 8998 2624
rect 9036 2644 9088 2650
rect 8760 2586 8812 2592
rect 9036 2586 9088 2592
rect 8772 2530 8800 2586
rect 8772 2502 9076 2530
rect 9140 2514 9168 3334
rect 9232 3194 9260 3334
rect 9310 3292 9618 3301
rect 9310 3290 9316 3292
rect 9372 3290 9396 3292
rect 9452 3290 9476 3292
rect 9532 3290 9556 3292
rect 9612 3290 9618 3292
rect 9372 3238 9374 3290
rect 9554 3238 9556 3290
rect 9310 3236 9316 3238
rect 9372 3236 9396 3238
rect 9452 3236 9476 3238
rect 9532 3236 9556 3238
rect 9612 3236 9618 3238
rect 9310 3227 9618 3236
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9312 2984 9364 2990
rect 9232 2944 9312 2972
rect 8680 2378 8892 2394
rect 8680 2372 8904 2378
rect 8680 2366 8852 2372
rect 8852 2314 8904 2320
rect 8944 2372 8996 2378
rect 8944 2314 8996 2320
rect 8850 2000 8906 2009
rect 8850 1935 8906 1944
rect 8864 1902 8892 1935
rect 8852 1896 8904 1902
rect 8852 1838 8904 1844
rect 8392 1352 8444 1358
rect 8392 1294 8444 1300
rect 8484 1352 8536 1358
rect 8484 1294 8536 1300
rect 8300 1012 8352 1018
rect 8300 954 8352 960
rect 8496 882 8524 1294
rect 8956 1290 8984 2314
rect 9048 1766 9076 2502
rect 9128 2508 9180 2514
rect 9128 2450 9180 2456
rect 9232 2106 9260 2944
rect 9312 2926 9364 2932
rect 9600 2514 9628 2994
rect 9692 2774 9720 3692
rect 9968 3602 9996 4762
rect 10244 4690 10272 5306
rect 10232 4684 10284 4690
rect 10232 4626 10284 4632
rect 10336 4622 10364 6938
rect 11716 6798 11744 7142
rect 11808 6798 11836 7346
rect 12176 6934 12204 7919
rect 12268 7750 12296 8502
rect 12820 8498 12848 10542
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 12348 8424 12400 8430
rect 12346 8392 12348 8401
rect 12400 8392 12402 8401
rect 12346 8327 12402 8336
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 12410 7644 12718 7653
rect 12410 7642 12416 7644
rect 12472 7642 12496 7644
rect 12552 7642 12576 7644
rect 12632 7642 12656 7644
rect 12712 7642 12718 7644
rect 12472 7590 12474 7642
rect 12654 7590 12656 7642
rect 12410 7588 12416 7590
rect 12472 7588 12496 7590
rect 12552 7588 12576 7590
rect 12632 7588 12656 7590
rect 12712 7588 12718 7590
rect 12410 7579 12718 7588
rect 12912 7528 12940 10610
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 13004 10266 13032 10406
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 12992 10056 13044 10062
rect 12992 9998 13044 10004
rect 13004 9654 13032 9998
rect 12992 9648 13044 9654
rect 12992 9590 13044 9596
rect 13188 8294 13216 11206
rect 15396 11206 15608 11234
rect 14924 10804 14976 10810
rect 14924 10746 14976 10752
rect 13452 10736 13504 10742
rect 13452 10678 13504 10684
rect 13464 9518 13492 10678
rect 14936 10674 14964 10746
rect 14464 10668 14516 10674
rect 14464 10610 14516 10616
rect 14924 10668 14976 10674
rect 14924 10610 14976 10616
rect 13820 10532 13872 10538
rect 13820 10474 13872 10480
rect 13544 9716 13596 9722
rect 13544 9658 13596 9664
rect 13452 9512 13504 9518
rect 13452 9454 13504 9460
rect 13556 9178 13584 9658
rect 13544 9172 13596 9178
rect 13544 9114 13596 9120
rect 13556 8430 13584 9114
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13740 8430 13768 8910
rect 13832 8634 13860 10474
rect 13960 10364 14268 10373
rect 13960 10362 13966 10364
rect 14022 10362 14046 10364
rect 14102 10362 14126 10364
rect 14182 10362 14206 10364
rect 14262 10362 14268 10364
rect 14022 10310 14024 10362
rect 14204 10310 14206 10362
rect 13960 10308 13966 10310
rect 14022 10308 14046 10310
rect 14102 10308 14126 10310
rect 14182 10308 14206 10310
rect 14262 10308 14268 10310
rect 13960 10299 14268 10308
rect 13960 9276 14268 9285
rect 13960 9274 13966 9276
rect 14022 9274 14046 9276
rect 14102 9274 14126 9276
rect 14182 9274 14206 9276
rect 14262 9274 14268 9276
rect 14022 9222 14024 9274
rect 14204 9222 14206 9274
rect 13960 9220 13966 9222
rect 14022 9220 14046 9222
rect 14102 9220 14126 9222
rect 14182 9220 14206 9222
rect 14262 9220 14268 9222
rect 13960 9211 14268 9220
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13728 8424 13780 8430
rect 13728 8366 13780 8372
rect 13084 8288 13136 8294
rect 13084 8230 13136 8236
rect 13176 8288 13228 8294
rect 13176 8230 13228 8236
rect 12728 7500 12940 7528
rect 12992 7540 13044 7546
rect 12164 6928 12216 6934
rect 12164 6870 12216 6876
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 11900 6458 11928 6802
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11992 6225 12020 6598
rect 11978 6216 12034 6225
rect 11428 6180 11480 6186
rect 11978 6151 12034 6160
rect 12072 6180 12124 6186
rect 11428 6122 11480 6128
rect 12176 6168 12204 6870
rect 12728 6798 12756 7500
rect 12992 7482 13044 7488
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 12716 6792 12768 6798
rect 12716 6734 12768 6740
rect 12728 6662 12756 6734
rect 12716 6656 12768 6662
rect 12716 6598 12768 6604
rect 12410 6556 12718 6565
rect 12410 6554 12416 6556
rect 12472 6554 12496 6556
rect 12552 6554 12576 6556
rect 12632 6554 12656 6556
rect 12712 6554 12718 6556
rect 12472 6502 12474 6554
rect 12654 6502 12656 6554
rect 12410 6500 12416 6502
rect 12472 6500 12496 6502
rect 12552 6500 12576 6502
rect 12632 6500 12656 6502
rect 12712 6500 12718 6502
rect 12410 6491 12718 6500
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 12124 6140 12204 6168
rect 12072 6122 12124 6128
rect 10860 6012 11168 6021
rect 10860 6010 10866 6012
rect 10922 6010 10946 6012
rect 11002 6010 11026 6012
rect 11082 6010 11106 6012
rect 11162 6010 11168 6012
rect 10922 5958 10924 6010
rect 11104 5958 11106 6010
rect 10860 5956 10866 5958
rect 10922 5956 10946 5958
rect 11002 5956 11026 5958
rect 11082 5956 11106 5958
rect 11162 5956 11168 5958
rect 10860 5947 11168 5956
rect 11440 5846 11468 6122
rect 10692 5840 10744 5846
rect 10692 5782 10744 5788
rect 11428 5840 11480 5846
rect 11428 5782 11480 5788
rect 10704 5098 10732 5782
rect 11704 5772 11756 5778
rect 11704 5714 11756 5720
rect 11888 5772 11940 5778
rect 11888 5714 11940 5720
rect 11612 5704 11664 5710
rect 11612 5646 11664 5652
rect 10692 5092 10744 5098
rect 10692 5034 10744 5040
rect 10324 4616 10376 4622
rect 10324 4558 10376 4564
rect 10600 4616 10652 4622
rect 10600 4558 10652 4564
rect 10140 4480 10192 4486
rect 10140 4422 10192 4428
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 9772 3596 9824 3602
rect 9956 3596 10008 3602
rect 9824 3556 9904 3584
rect 9772 3538 9824 3544
rect 9876 3482 9904 3556
rect 9956 3538 10008 3544
rect 10060 3482 10088 3674
rect 9876 3454 10088 3482
rect 9692 2746 9812 2774
rect 9784 2582 9812 2746
rect 9772 2576 9824 2582
rect 9772 2518 9824 2524
rect 9588 2508 9640 2514
rect 9588 2450 9640 2456
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 9310 2204 9618 2213
rect 9310 2202 9316 2204
rect 9372 2202 9396 2204
rect 9452 2202 9476 2204
rect 9532 2202 9556 2204
rect 9612 2202 9618 2204
rect 9372 2150 9374 2202
rect 9554 2150 9556 2202
rect 9310 2148 9316 2150
rect 9372 2148 9396 2150
rect 9452 2148 9476 2150
rect 9532 2148 9556 2150
rect 9612 2148 9618 2150
rect 9310 2139 9618 2148
rect 9692 2106 9720 2382
rect 9772 2304 9824 2310
rect 9772 2246 9824 2252
rect 9220 2100 9272 2106
rect 9220 2042 9272 2048
rect 9680 2100 9732 2106
rect 9680 2042 9732 2048
rect 9588 2032 9640 2038
rect 9586 2000 9588 2009
rect 9640 2000 9642 2009
rect 9586 1935 9642 1944
rect 9404 1896 9456 1902
rect 9404 1838 9456 1844
rect 9036 1760 9088 1766
rect 9036 1702 9088 1708
rect 8760 1284 8812 1290
rect 8760 1226 8812 1232
rect 8944 1284 8996 1290
rect 8944 1226 8996 1232
rect 8484 876 8536 882
rect 8484 818 8536 824
rect 8772 814 8800 1226
rect 8956 1018 8984 1226
rect 9416 1222 9444 1838
rect 9784 1834 9812 2246
rect 9876 2106 9904 3454
rect 10152 2990 10180 4422
rect 10612 4282 10640 4558
rect 10600 4276 10652 4282
rect 10600 4218 10652 4224
rect 10704 3534 10732 5034
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 11428 5024 11480 5030
rect 11428 4966 11480 4972
rect 10796 4078 10824 4966
rect 10860 4924 11168 4933
rect 10860 4922 10866 4924
rect 10922 4922 10946 4924
rect 11002 4922 11026 4924
rect 11082 4922 11106 4924
rect 11162 4922 11168 4924
rect 10922 4870 10924 4922
rect 11104 4870 11106 4922
rect 10860 4868 10866 4870
rect 10922 4868 10946 4870
rect 11002 4868 11026 4870
rect 11082 4868 11106 4870
rect 11162 4868 11168 4870
rect 10860 4859 11168 4868
rect 11440 4826 11468 4966
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 11334 4584 11390 4593
rect 11072 4078 11100 4558
rect 11334 4519 11390 4528
rect 11348 4078 11376 4519
rect 11440 4146 11468 4762
rect 11428 4140 11480 4146
rect 11428 4082 11480 4088
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 11060 4072 11112 4078
rect 11060 4014 11112 4020
rect 11336 4072 11388 4078
rect 11336 4014 11388 4020
rect 10784 3936 10836 3942
rect 11072 3924 11100 4014
rect 11072 3896 11284 3924
rect 10784 3878 10836 3884
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 9864 2100 9916 2106
rect 9864 2042 9916 2048
rect 10048 1964 10100 1970
rect 10048 1906 10100 1912
rect 9772 1828 9824 1834
rect 9772 1770 9824 1776
rect 9784 1358 9812 1770
rect 9864 1556 9916 1562
rect 9864 1498 9916 1504
rect 9876 1426 9904 1498
rect 9864 1420 9916 1426
rect 9916 1380 9996 1408
rect 9864 1362 9916 1368
rect 9772 1352 9824 1358
rect 9772 1294 9824 1300
rect 9404 1216 9456 1222
rect 9404 1158 9456 1164
rect 9310 1116 9618 1125
rect 9310 1114 9316 1116
rect 9372 1114 9396 1116
rect 9452 1114 9476 1116
rect 9532 1114 9556 1116
rect 9612 1114 9618 1116
rect 9372 1062 9374 1114
rect 9554 1062 9556 1114
rect 9310 1060 9316 1062
rect 9372 1060 9396 1062
rect 9452 1060 9476 1062
rect 9532 1060 9556 1062
rect 9612 1060 9618 1062
rect 9310 1051 9618 1060
rect 8944 1012 8996 1018
rect 8944 954 8996 960
rect 9784 814 9812 1294
rect 9968 882 9996 1380
rect 10060 1222 10088 1906
rect 10520 1494 10548 2994
rect 10796 2990 10824 3878
rect 10860 3836 11168 3845
rect 10860 3834 10866 3836
rect 10922 3834 10946 3836
rect 11002 3834 11026 3836
rect 11082 3834 11106 3836
rect 11162 3834 11168 3836
rect 10922 3782 10924 3834
rect 11104 3782 11106 3834
rect 10860 3780 10866 3782
rect 10922 3780 10946 3782
rect 11002 3780 11026 3782
rect 11082 3780 11106 3782
rect 11162 3780 11168 3782
rect 10860 3771 11168 3780
rect 11256 3194 11284 3896
rect 11348 3194 11376 4014
rect 11624 3602 11652 5646
rect 11716 5574 11744 5714
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 11900 4486 11928 5714
rect 12176 5574 12204 6140
rect 12728 6118 12756 6394
rect 12912 6322 12940 6938
rect 12900 6316 12952 6322
rect 12900 6258 12952 6264
rect 12716 6112 12768 6118
rect 12716 6054 12768 6060
rect 13004 5930 13032 7482
rect 13096 6338 13124 8230
rect 13740 7954 13768 8366
rect 13728 7948 13780 7954
rect 13728 7890 13780 7896
rect 13268 7812 13320 7818
rect 13268 7754 13320 7760
rect 13280 7342 13308 7754
rect 13832 7750 13860 8434
rect 14372 8424 14424 8430
rect 14372 8366 14424 8372
rect 13960 8188 14268 8197
rect 13960 8186 13966 8188
rect 14022 8186 14046 8188
rect 14102 8186 14126 8188
rect 14182 8186 14206 8188
rect 14262 8186 14268 8188
rect 14022 8134 14024 8186
rect 14204 8134 14206 8186
rect 13960 8132 13966 8134
rect 14022 8132 14046 8134
rect 14102 8132 14126 8134
rect 14182 8132 14206 8134
rect 14262 8132 14268 8134
rect 13960 8123 14268 8132
rect 14384 8022 14412 8366
rect 14372 8016 14424 8022
rect 14372 7958 14424 7964
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 13268 7336 13320 7342
rect 13268 7278 13320 7284
rect 13452 7268 13504 7274
rect 13452 7210 13504 7216
rect 13464 6882 13492 7210
rect 13832 7002 13860 7686
rect 14372 7472 14424 7478
rect 14372 7414 14424 7420
rect 13960 7100 14268 7109
rect 13960 7098 13966 7100
rect 14022 7098 14046 7100
rect 14102 7098 14126 7100
rect 14182 7098 14206 7100
rect 14262 7098 14268 7100
rect 14022 7046 14024 7098
rect 14204 7046 14206 7098
rect 13960 7044 13966 7046
rect 14022 7044 14046 7046
rect 14102 7044 14126 7046
rect 14182 7044 14206 7046
rect 14262 7044 14268 7046
rect 13960 7035 14268 7044
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 13280 6854 13492 6882
rect 13096 6310 13216 6338
rect 13084 6180 13136 6186
rect 13084 6122 13136 6128
rect 12820 5902 13032 5930
rect 12624 5840 12676 5846
rect 12676 5788 12756 5794
rect 12624 5782 12756 5788
rect 12636 5766 12756 5782
rect 12728 5710 12756 5766
rect 12716 5704 12768 5710
rect 12716 5646 12768 5652
rect 12164 5568 12216 5574
rect 12164 5510 12216 5516
rect 12176 5030 12204 5510
rect 12410 5468 12718 5477
rect 12410 5466 12416 5468
rect 12472 5466 12496 5468
rect 12552 5466 12576 5468
rect 12632 5466 12656 5468
rect 12712 5466 12718 5468
rect 12472 5414 12474 5466
rect 12654 5414 12656 5466
rect 12410 5412 12416 5414
rect 12472 5412 12496 5414
rect 12552 5412 12576 5414
rect 12632 5412 12656 5414
rect 12712 5412 12718 5414
rect 12410 5403 12718 5412
rect 12256 5092 12308 5098
rect 12256 5034 12308 5040
rect 12440 5092 12492 5098
rect 12440 5034 12492 5040
rect 12164 5024 12216 5030
rect 12164 4966 12216 4972
rect 12268 4758 12296 5034
rect 12452 4826 12480 5034
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12256 4752 12308 4758
rect 12256 4694 12308 4700
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 11980 4480 12032 4486
rect 11980 4422 12032 4428
rect 11888 4072 11940 4078
rect 11888 4014 11940 4020
rect 11900 3641 11928 4014
rect 11886 3632 11942 3641
rect 11612 3596 11664 3602
rect 11886 3567 11942 3576
rect 11612 3538 11664 3544
rect 11244 3188 11296 3194
rect 11244 3130 11296 3136
rect 11336 3188 11388 3194
rect 11336 3130 11388 3136
rect 11242 3088 11298 3097
rect 11242 3023 11298 3032
rect 10784 2984 10836 2990
rect 10784 2926 10836 2932
rect 11256 2854 11284 3023
rect 11624 2854 11652 3538
rect 11992 2990 12020 4422
rect 12164 3528 12216 3534
rect 12164 3470 12216 3476
rect 12072 3392 12124 3398
rect 12072 3334 12124 3340
rect 11980 2984 12032 2990
rect 11980 2926 12032 2932
rect 10600 2848 10652 2854
rect 10600 2790 10652 2796
rect 11244 2848 11296 2854
rect 11244 2790 11296 2796
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 10612 2650 10640 2790
rect 10860 2748 11168 2757
rect 10860 2746 10866 2748
rect 10922 2746 10946 2748
rect 11002 2746 11026 2748
rect 11082 2746 11106 2748
rect 11162 2746 11168 2748
rect 10922 2694 10924 2746
rect 11104 2694 11106 2746
rect 10860 2692 10866 2694
rect 10922 2692 10946 2694
rect 11002 2692 11026 2694
rect 11082 2692 11106 2694
rect 11162 2692 11168 2694
rect 10860 2683 11168 2692
rect 10600 2644 10652 2650
rect 10600 2586 10652 2592
rect 11256 2553 11284 2790
rect 11242 2544 11298 2553
rect 11624 2514 11652 2790
rect 11242 2479 11298 2488
rect 11612 2508 11664 2514
rect 11612 2450 11664 2456
rect 11980 2304 12032 2310
rect 11980 2246 12032 2252
rect 10784 1964 10836 1970
rect 10784 1906 10836 1912
rect 10796 1562 10824 1906
rect 11888 1896 11940 1902
rect 11888 1838 11940 1844
rect 11428 1760 11480 1766
rect 11428 1702 11480 1708
rect 10860 1660 11168 1669
rect 10860 1658 10866 1660
rect 10922 1658 10946 1660
rect 11002 1658 11026 1660
rect 11082 1658 11106 1660
rect 11162 1658 11168 1660
rect 10922 1606 10924 1658
rect 11104 1606 11106 1658
rect 10860 1604 10866 1606
rect 10922 1604 10946 1606
rect 11002 1604 11026 1606
rect 11082 1604 11106 1606
rect 11162 1604 11168 1606
rect 10860 1595 11168 1604
rect 11440 1562 11468 1702
rect 10784 1556 10836 1562
rect 10784 1498 10836 1504
rect 11428 1556 11480 1562
rect 11428 1498 11480 1504
rect 10508 1488 10560 1494
rect 10508 1430 10560 1436
rect 11900 1426 11928 1838
rect 11992 1562 12020 2246
rect 12084 1873 12112 3334
rect 12176 2650 12204 3470
rect 12268 3398 12296 4694
rect 12624 4684 12676 4690
rect 12624 4626 12676 4632
rect 12636 4593 12664 4626
rect 12622 4584 12678 4593
rect 12622 4519 12678 4528
rect 12410 4380 12718 4389
rect 12410 4378 12416 4380
rect 12472 4378 12496 4380
rect 12552 4378 12576 4380
rect 12632 4378 12656 4380
rect 12712 4378 12718 4380
rect 12472 4326 12474 4378
rect 12654 4326 12656 4378
rect 12410 4324 12416 4326
rect 12472 4324 12496 4326
rect 12552 4324 12576 4326
rect 12632 4324 12656 4326
rect 12712 4324 12718 4326
rect 12410 4315 12718 4324
rect 12820 3777 12848 5902
rect 12992 5840 13044 5846
rect 12992 5782 13044 5788
rect 13004 5250 13032 5782
rect 13096 5710 13124 6122
rect 13084 5704 13136 5710
rect 13084 5646 13136 5652
rect 13188 5370 13216 6310
rect 13176 5364 13228 5370
rect 13176 5306 13228 5312
rect 13004 5222 13216 5250
rect 12900 5160 12952 5166
rect 12900 5102 12952 5108
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 12806 3768 12862 3777
rect 12806 3703 12862 3712
rect 12912 3670 12940 5102
rect 12992 4820 13044 4826
rect 12992 4762 13044 4768
rect 13004 4010 13032 4762
rect 13096 4486 13124 5102
rect 13084 4480 13136 4486
rect 13084 4422 13136 4428
rect 12992 4004 13044 4010
rect 12992 3946 13044 3952
rect 12900 3664 12952 3670
rect 12900 3606 12952 3612
rect 12256 3392 12308 3398
rect 12256 3334 12308 3340
rect 12268 2922 12296 3334
rect 12410 3292 12718 3301
rect 12410 3290 12416 3292
rect 12472 3290 12496 3292
rect 12552 3290 12576 3292
rect 12632 3290 12656 3292
rect 12712 3290 12718 3292
rect 12472 3238 12474 3290
rect 12654 3238 12656 3290
rect 12410 3236 12416 3238
rect 12472 3236 12496 3238
rect 12552 3236 12576 3238
rect 12632 3236 12656 3238
rect 12712 3236 12718 3238
rect 12410 3227 12718 3236
rect 12716 2984 12768 2990
rect 12714 2952 12716 2961
rect 12768 2952 12770 2961
rect 12256 2916 12308 2922
rect 12912 2938 12940 3606
rect 13004 3534 13032 3946
rect 13096 3602 13124 4422
rect 13084 3596 13136 3602
rect 13084 3538 13136 3544
rect 12992 3528 13044 3534
rect 13188 3505 13216 5222
rect 12992 3470 13044 3476
rect 13174 3496 13230 3505
rect 13004 3398 13032 3470
rect 13174 3431 13230 3440
rect 12992 3392 13044 3398
rect 12992 3334 13044 3340
rect 13280 3074 13308 6854
rect 13452 6792 13504 6798
rect 13452 6734 13504 6740
rect 13544 6792 13596 6798
rect 13596 6752 13676 6780
rect 13544 6734 13596 6740
rect 13464 6390 13492 6734
rect 13452 6384 13504 6390
rect 13452 6326 13504 6332
rect 13542 6216 13598 6225
rect 13542 6151 13598 6160
rect 13556 6118 13584 6151
rect 13544 6112 13596 6118
rect 13544 6054 13596 6060
rect 13452 5568 13504 5574
rect 13452 5510 13504 5516
rect 13464 5166 13492 5510
rect 13556 5273 13584 6054
rect 13542 5264 13598 5273
rect 13542 5199 13598 5208
rect 13452 5160 13504 5166
rect 13452 5102 13504 5108
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 13004 3058 13308 3074
rect 12992 3052 13308 3058
rect 13044 3046 13308 3052
rect 12992 2994 13044 3000
rect 13266 2952 13322 2961
rect 12912 2910 13032 2938
rect 12714 2887 12770 2896
rect 12256 2858 12308 2864
rect 12268 2650 12296 2858
rect 12164 2644 12216 2650
rect 12164 2586 12216 2592
rect 12256 2644 12308 2650
rect 12256 2586 12308 2592
rect 12176 1902 12204 2586
rect 12256 2372 12308 2378
rect 12256 2314 12308 2320
rect 12268 2106 12296 2314
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 12410 2204 12718 2213
rect 12410 2202 12416 2204
rect 12472 2202 12496 2204
rect 12552 2202 12576 2204
rect 12632 2202 12656 2204
rect 12712 2202 12718 2204
rect 12472 2150 12474 2202
rect 12654 2150 12656 2202
rect 12410 2148 12416 2150
rect 12472 2148 12496 2150
rect 12552 2148 12576 2150
rect 12632 2148 12656 2150
rect 12712 2148 12718 2150
rect 12410 2139 12718 2148
rect 12256 2100 12308 2106
rect 12256 2042 12308 2048
rect 12164 1896 12216 1902
rect 12070 1864 12126 1873
rect 12164 1838 12216 1844
rect 12348 1896 12400 1902
rect 12348 1838 12400 1844
rect 12808 1896 12860 1902
rect 12912 1884 12940 2246
rect 13004 1902 13032 2910
rect 13266 2887 13268 2896
rect 13320 2887 13322 2896
rect 13268 2858 13320 2864
rect 13372 2836 13400 4966
rect 13464 4146 13492 5102
rect 13452 4140 13504 4146
rect 13452 4082 13504 4088
rect 13648 3890 13676 6752
rect 13728 6656 13780 6662
rect 13728 6598 13780 6604
rect 13912 6656 13964 6662
rect 13912 6598 13964 6604
rect 13740 4622 13768 6598
rect 13924 6322 13952 6598
rect 13912 6316 13964 6322
rect 13912 6258 13964 6264
rect 13960 6012 14268 6021
rect 13960 6010 13966 6012
rect 14022 6010 14046 6012
rect 14102 6010 14126 6012
rect 14182 6010 14206 6012
rect 14262 6010 14268 6012
rect 14022 5958 14024 6010
rect 14204 5958 14206 6010
rect 13960 5956 13966 5958
rect 14022 5956 14046 5958
rect 14102 5956 14126 5958
rect 14182 5956 14206 5958
rect 14262 5956 14268 5958
rect 13960 5947 14268 5956
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 13832 5098 13860 5510
rect 14384 5234 14412 7414
rect 14476 6730 14504 10610
rect 14648 10600 14700 10606
rect 14648 10542 14700 10548
rect 15198 10568 15254 10577
rect 14660 10198 14688 10542
rect 14832 10532 14884 10538
rect 15198 10503 15254 10512
rect 15292 10532 15344 10538
rect 14832 10474 14884 10480
rect 14648 10192 14700 10198
rect 14648 10134 14700 10140
rect 14660 9450 14688 10134
rect 14844 9586 14872 10474
rect 15212 10470 15240 10503
rect 15292 10474 15344 10480
rect 15200 10464 15252 10470
rect 15120 10424 15200 10452
rect 15016 10124 15068 10130
rect 15016 10066 15068 10072
rect 14924 9920 14976 9926
rect 14924 9862 14976 9868
rect 14832 9580 14884 9586
rect 14832 9522 14884 9528
rect 14648 9444 14700 9450
rect 14648 9386 14700 9392
rect 14660 9178 14688 9386
rect 14740 9376 14792 9382
rect 14740 9318 14792 9324
rect 14648 9172 14700 9178
rect 14648 9114 14700 9120
rect 14752 8090 14780 9318
rect 14844 8974 14872 9522
rect 14832 8968 14884 8974
rect 14832 8910 14884 8916
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 14646 6896 14702 6905
rect 14646 6831 14648 6840
rect 14700 6831 14702 6840
rect 14648 6802 14700 6808
rect 14464 6724 14516 6730
rect 14464 6666 14516 6672
rect 14556 6316 14608 6322
rect 14556 6258 14608 6264
rect 14464 6180 14516 6186
rect 14464 6122 14516 6128
rect 14476 5914 14504 6122
rect 14464 5908 14516 5914
rect 14464 5850 14516 5856
rect 14464 5772 14516 5778
rect 14464 5714 14516 5720
rect 14476 5234 14504 5714
rect 14372 5228 14424 5234
rect 14372 5170 14424 5176
rect 14464 5228 14516 5234
rect 14464 5170 14516 5176
rect 13820 5092 13872 5098
rect 13820 5034 13872 5040
rect 13960 4924 14268 4933
rect 13960 4922 13966 4924
rect 14022 4922 14046 4924
rect 14102 4922 14126 4924
rect 14182 4922 14206 4924
rect 14262 4922 14268 4924
rect 14022 4870 14024 4922
rect 14204 4870 14206 4922
rect 13960 4868 13966 4870
rect 14022 4868 14046 4870
rect 14102 4868 14126 4870
rect 14182 4868 14206 4870
rect 14262 4868 14268 4870
rect 13960 4859 14268 4868
rect 14476 4690 14504 5170
rect 14568 4758 14596 6258
rect 14752 5794 14780 7142
rect 14844 7002 14872 8910
rect 14936 7936 14964 9862
rect 15028 8090 15056 10066
rect 15120 8838 15148 10424
rect 15200 10406 15252 10412
rect 15198 10024 15254 10033
rect 15198 9959 15254 9968
rect 15212 9518 15240 9959
rect 15304 9722 15332 10474
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15200 9512 15252 9518
rect 15200 9454 15252 9460
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 15016 8084 15068 8090
rect 15016 8026 15068 8032
rect 15016 7948 15068 7954
rect 14936 7908 15016 7936
rect 15016 7890 15068 7896
rect 15028 7478 15056 7890
rect 15016 7472 15068 7478
rect 15016 7414 15068 7420
rect 15016 7336 15068 7342
rect 15016 7278 15068 7284
rect 14832 6996 14884 7002
rect 14832 6938 14884 6944
rect 15028 6934 15056 7278
rect 15120 6934 15148 8774
rect 15016 6928 15068 6934
rect 15016 6870 15068 6876
rect 15108 6928 15160 6934
rect 15108 6870 15160 6876
rect 14832 6860 14884 6866
rect 14832 6802 14884 6808
rect 14660 5766 14780 5794
rect 14660 4826 14688 5766
rect 14740 5296 14792 5302
rect 14740 5238 14792 5244
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 14556 4752 14608 4758
rect 14556 4694 14608 4700
rect 14464 4684 14516 4690
rect 14464 4626 14516 4632
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 14462 4584 14518 4593
rect 14462 4519 14518 4528
rect 14476 4486 14504 4519
rect 13728 4480 13780 4486
rect 13728 4422 13780 4428
rect 14464 4480 14516 4486
rect 14464 4422 14516 4428
rect 13740 4146 13768 4422
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 13648 3862 13860 3890
rect 13726 3768 13782 3777
rect 13452 3732 13504 3738
rect 13832 3738 13860 3862
rect 13960 3836 14268 3845
rect 13960 3834 13966 3836
rect 14022 3834 14046 3836
rect 14102 3834 14126 3836
rect 14182 3834 14206 3836
rect 14262 3834 14268 3836
rect 14022 3782 14024 3834
rect 14204 3782 14206 3834
rect 13960 3780 13966 3782
rect 14022 3780 14046 3782
rect 14102 3780 14126 3782
rect 14182 3780 14206 3782
rect 14262 3780 14268 3782
rect 13960 3771 14268 3780
rect 13726 3703 13782 3712
rect 13820 3732 13872 3738
rect 13452 3674 13504 3680
rect 13464 3398 13492 3674
rect 13740 3584 13768 3703
rect 13820 3674 13872 3680
rect 14004 3732 14056 3738
rect 14004 3674 14056 3680
rect 13820 3596 13872 3602
rect 13740 3556 13820 3584
rect 13820 3538 13872 3544
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13452 3392 13504 3398
rect 13452 3334 13504 3340
rect 13450 3224 13506 3233
rect 13450 3159 13452 3168
rect 13504 3159 13506 3168
rect 13452 3130 13504 3136
rect 13464 2990 13492 3130
rect 13452 2984 13504 2990
rect 13452 2926 13504 2932
rect 13372 2808 13492 2836
rect 13358 2000 13414 2009
rect 13358 1935 13414 1944
rect 12860 1856 12940 1884
rect 12808 1838 12860 1844
rect 12070 1799 12126 1808
rect 11980 1556 12032 1562
rect 11980 1498 12032 1504
rect 10232 1420 10284 1426
rect 10152 1380 10232 1408
rect 10048 1216 10100 1222
rect 10048 1158 10100 1164
rect 10152 1018 10180 1380
rect 10232 1362 10284 1368
rect 11520 1420 11572 1426
rect 11520 1362 11572 1368
rect 11888 1420 11940 1426
rect 11888 1362 11940 1368
rect 11532 1018 11560 1362
rect 11992 1222 12020 1498
rect 12176 1290 12204 1838
rect 12360 1562 12388 1838
rect 12348 1556 12400 1562
rect 12348 1498 12400 1504
rect 12912 1426 12940 1856
rect 12992 1896 13044 1902
rect 12992 1838 13044 1844
rect 13176 1760 13228 1766
rect 13176 1702 13228 1708
rect 13188 1442 13216 1702
rect 12808 1420 12860 1426
rect 12808 1362 12860 1368
rect 12900 1420 12952 1426
rect 12900 1362 12952 1368
rect 13096 1414 13216 1442
rect 13372 1426 13400 1935
rect 13360 1420 13412 1426
rect 12164 1284 12216 1290
rect 12164 1226 12216 1232
rect 11888 1216 11940 1222
rect 11888 1158 11940 1164
rect 11980 1216 12032 1222
rect 11980 1158 12032 1164
rect 10140 1012 10192 1018
rect 10140 954 10192 960
rect 11520 1012 11572 1018
rect 11520 954 11572 960
rect 9956 876 10008 882
rect 9956 818 10008 824
rect 7012 808 7064 814
rect 7012 750 7064 756
rect 8760 808 8812 814
rect 8760 750 8812 756
rect 9772 808 9824 814
rect 9772 750 9824 756
rect 4660 572 4968 581
rect 4660 570 4666 572
rect 4722 570 4746 572
rect 4802 570 4826 572
rect 4882 570 4906 572
rect 4962 570 4968 572
rect 4722 518 4724 570
rect 4904 518 4906 570
rect 4660 516 4666 518
rect 4722 516 4746 518
rect 4802 516 4826 518
rect 4882 516 4906 518
rect 4962 516 4968 518
rect 4660 507 4968 516
rect 7760 572 8068 581
rect 7760 570 7766 572
rect 7822 570 7846 572
rect 7902 570 7926 572
rect 7982 570 8006 572
rect 8062 570 8068 572
rect 7822 518 7824 570
rect 8004 518 8006 570
rect 7760 516 7766 518
rect 7822 516 7846 518
rect 7902 516 7926 518
rect 7982 516 8006 518
rect 8062 516 8068 518
rect 7760 507 8068 516
rect 10860 572 11168 581
rect 10860 570 10866 572
rect 10922 570 10946 572
rect 11002 570 11026 572
rect 11082 570 11106 572
rect 11162 570 11168 572
rect 10922 518 10924 570
rect 11104 518 11106 570
rect 10860 516 10866 518
rect 10922 516 10946 518
rect 11002 516 11026 518
rect 11082 516 11106 518
rect 11162 516 11168 518
rect 10860 507 11168 516
rect 11900 406 11928 1158
rect 12410 1116 12718 1125
rect 12410 1114 12416 1116
rect 12472 1114 12496 1116
rect 12552 1114 12576 1116
rect 12632 1114 12656 1116
rect 12712 1114 12718 1116
rect 12472 1062 12474 1114
rect 12654 1062 12656 1114
rect 12410 1060 12416 1062
rect 12472 1060 12496 1062
rect 12552 1060 12576 1062
rect 12632 1060 12656 1062
rect 12712 1060 12718 1062
rect 12410 1051 12718 1060
rect 12820 814 12848 1362
rect 13096 1358 13124 1414
rect 13360 1362 13412 1368
rect 13084 1352 13136 1358
rect 13084 1294 13136 1300
rect 12992 1284 13044 1290
rect 12992 1226 13044 1232
rect 12900 1216 12952 1222
rect 12900 1158 12952 1164
rect 12808 808 12860 814
rect 12806 776 12808 785
rect 12860 776 12862 785
rect 12806 711 12862 720
rect 12072 672 12124 678
rect 12072 614 12124 620
rect 12532 672 12584 678
rect 12532 614 12584 620
rect 12716 672 12768 678
rect 12716 614 12768 620
rect 11888 400 11940 406
rect 11888 342 11940 348
rect 12084 134 12112 614
rect 12544 474 12572 614
rect 12532 468 12584 474
rect 12532 410 12584 416
rect 12728 338 12756 614
rect 12716 332 12768 338
rect 12716 274 12768 280
rect 12912 270 12940 1158
rect 13004 814 13032 1226
rect 13464 1222 13492 2808
rect 13556 2582 13584 3470
rect 13728 3460 13780 3466
rect 13728 3402 13780 3408
rect 13820 3460 13872 3466
rect 13820 3402 13872 3408
rect 13544 2576 13596 2582
rect 13544 2518 13596 2524
rect 13740 2446 13768 3402
rect 13832 3369 13860 3402
rect 13912 3392 13964 3398
rect 13818 3360 13874 3369
rect 13912 3334 13964 3340
rect 13818 3295 13874 3304
rect 13820 2984 13872 2990
rect 13820 2926 13872 2932
rect 13728 2440 13780 2446
rect 13728 2382 13780 2388
rect 13740 2088 13768 2382
rect 13832 2378 13860 2926
rect 13924 2854 13952 3334
rect 14016 3194 14044 3674
rect 14188 3596 14240 3602
rect 14188 3538 14240 3544
rect 14096 3392 14148 3398
rect 14096 3334 14148 3340
rect 14004 3188 14056 3194
rect 14004 3130 14056 3136
rect 14108 3058 14136 3334
rect 14200 3233 14228 3538
rect 14372 3528 14424 3534
rect 14568 3516 14596 4694
rect 14648 4480 14700 4486
rect 14648 4422 14700 4428
rect 14660 3534 14688 4422
rect 14424 3488 14596 3516
rect 14648 3528 14700 3534
rect 14372 3470 14424 3476
rect 14186 3224 14242 3233
rect 14186 3159 14242 3168
rect 14096 3052 14148 3058
rect 14096 2994 14148 3000
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 13912 2848 13964 2854
rect 14200 2836 14228 2926
rect 14200 2808 14412 2836
rect 13912 2790 13964 2796
rect 13960 2748 14268 2757
rect 13960 2746 13966 2748
rect 14022 2746 14046 2748
rect 14102 2746 14126 2748
rect 14182 2746 14206 2748
rect 14262 2746 14268 2748
rect 14022 2694 14024 2746
rect 14204 2694 14206 2746
rect 13960 2692 13966 2694
rect 14022 2692 14046 2694
rect 14102 2692 14126 2694
rect 14182 2692 14206 2694
rect 14262 2692 14268 2694
rect 13960 2683 14268 2692
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 13912 2576 13964 2582
rect 13910 2544 13912 2553
rect 13964 2544 13966 2553
rect 13910 2479 13966 2488
rect 14186 2544 14242 2553
rect 14186 2479 14188 2488
rect 13820 2372 13872 2378
rect 13820 2314 13872 2320
rect 13648 2060 13860 2088
rect 13544 1828 13596 1834
rect 13544 1770 13596 1776
rect 13268 1216 13320 1222
rect 13268 1158 13320 1164
rect 13452 1216 13504 1222
rect 13452 1158 13504 1164
rect 13280 1057 13308 1158
rect 13266 1048 13322 1057
rect 13556 1018 13584 1770
rect 13648 1426 13676 2060
rect 13832 1970 13860 2060
rect 13728 1964 13780 1970
rect 13728 1906 13780 1912
rect 13820 1964 13872 1970
rect 13820 1906 13872 1912
rect 13740 1562 13768 1906
rect 13924 1834 13952 2479
rect 14240 2479 14242 2488
rect 14188 2450 14240 2456
rect 14292 2378 14320 2586
rect 14280 2372 14332 2378
rect 14280 2314 14332 2320
rect 14292 1970 14320 2314
rect 14280 1964 14332 1970
rect 14280 1906 14332 1912
rect 13912 1828 13964 1834
rect 13912 1770 13964 1776
rect 13820 1760 13872 1766
rect 13820 1702 13872 1708
rect 13832 1562 13860 1702
rect 13960 1660 14268 1669
rect 13960 1658 13966 1660
rect 14022 1658 14046 1660
rect 14102 1658 14126 1660
rect 14182 1658 14206 1660
rect 14262 1658 14268 1660
rect 14022 1606 14024 1658
rect 14204 1606 14206 1658
rect 13960 1604 13966 1606
rect 14022 1604 14046 1606
rect 14102 1604 14126 1606
rect 14182 1604 14206 1606
rect 14262 1604 14268 1606
rect 13960 1595 14268 1604
rect 13728 1556 13780 1562
rect 13728 1498 13780 1504
rect 13820 1556 13872 1562
rect 13820 1498 13872 1504
rect 13636 1420 13688 1426
rect 13636 1362 13688 1368
rect 13266 983 13322 992
rect 13544 1012 13596 1018
rect 13544 954 13596 960
rect 13266 912 13322 921
rect 13176 876 13228 882
rect 13266 847 13268 856
rect 13176 818 13228 824
rect 13320 847 13322 856
rect 13268 818 13320 824
rect 12992 808 13044 814
rect 12992 750 13044 756
rect 12900 264 12952 270
rect 12900 206 12952 212
rect 13188 202 13216 818
rect 13740 678 13768 1498
rect 14094 1456 14150 1465
rect 14094 1391 14150 1400
rect 13820 1352 13872 1358
rect 13820 1294 13872 1300
rect 13832 814 13860 1294
rect 14108 950 14136 1391
rect 14188 1284 14240 1290
rect 14188 1226 14240 1232
rect 14096 944 14148 950
rect 14096 886 14148 892
rect 13820 808 13872 814
rect 13820 750 13872 756
rect 14200 678 14228 1226
rect 14278 1048 14334 1057
rect 14278 983 14334 992
rect 14292 950 14320 983
rect 14384 950 14412 2808
rect 14476 1562 14504 3488
rect 14648 3470 14700 3476
rect 14556 2916 14608 2922
rect 14556 2858 14608 2864
rect 14464 1556 14516 1562
rect 14464 1498 14516 1504
rect 14568 1290 14596 2858
rect 14660 2582 14688 3470
rect 14752 3369 14780 5238
rect 14844 3738 14872 6802
rect 14924 6792 14976 6798
rect 14922 6760 14924 6769
rect 15212 6780 15240 9454
rect 15292 7744 15344 7750
rect 15292 7686 15344 7692
rect 15304 6934 15332 7686
rect 15292 6928 15344 6934
rect 15292 6870 15344 6876
rect 14976 6760 14978 6769
rect 15212 6752 15332 6780
rect 14922 6695 14978 6704
rect 15016 6724 15068 6730
rect 15068 6684 15240 6712
rect 15016 6666 15068 6672
rect 15106 6216 15162 6225
rect 14924 6180 14976 6186
rect 14976 6160 15106 6168
rect 14976 6151 15162 6160
rect 14976 6140 15148 6151
rect 14924 6122 14976 6128
rect 15120 5846 15148 6140
rect 15108 5840 15160 5846
rect 15108 5782 15160 5788
rect 15120 5574 15148 5782
rect 15108 5568 15160 5574
rect 15108 5510 15160 5516
rect 14922 5264 14978 5273
rect 14922 5199 14978 5208
rect 14936 4486 14964 5199
rect 15016 5092 15068 5098
rect 15016 5034 15068 5040
rect 14924 4480 14976 4486
rect 14924 4422 14976 4428
rect 14924 4140 14976 4146
rect 14924 4082 14976 4088
rect 14832 3732 14884 3738
rect 14832 3674 14884 3680
rect 14832 3392 14884 3398
rect 14738 3360 14794 3369
rect 14832 3334 14884 3340
rect 14738 3295 14794 3304
rect 14648 2576 14700 2582
rect 14648 2518 14700 2524
rect 14740 2508 14792 2514
rect 14740 2450 14792 2456
rect 14648 2304 14700 2310
rect 14648 2246 14700 2252
rect 14660 1834 14688 2246
rect 14752 2009 14780 2450
rect 14738 2000 14794 2009
rect 14738 1935 14794 1944
rect 14844 1902 14872 3334
rect 14936 3058 14964 4082
rect 15028 4049 15056 5034
rect 15120 4865 15148 5510
rect 15212 5166 15240 6684
rect 15200 5160 15252 5166
rect 15200 5102 15252 5108
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 15106 4856 15162 4865
rect 15106 4791 15162 4800
rect 15014 4040 15070 4049
rect 15014 3975 15016 3984
rect 15068 3975 15070 3984
rect 15016 3946 15068 3952
rect 14924 3052 14976 3058
rect 14924 2994 14976 3000
rect 14936 2514 14964 2994
rect 15120 2854 15148 4791
rect 15212 4078 15240 4966
rect 15200 4072 15252 4078
rect 15200 4014 15252 4020
rect 15304 4026 15332 6752
rect 15396 6458 15424 11206
rect 15580 11132 15608 11206
rect 15658 11200 15714 12000
rect 17592 11416 17644 11422
rect 17592 11358 17644 11364
rect 15672 11132 15700 11200
rect 15580 11104 15700 11132
rect 16120 11144 16172 11150
rect 16120 11086 16172 11092
rect 15510 10908 15818 10917
rect 15510 10906 15516 10908
rect 15572 10906 15596 10908
rect 15652 10906 15676 10908
rect 15732 10906 15756 10908
rect 15812 10906 15818 10908
rect 15572 10854 15574 10906
rect 15754 10854 15756 10906
rect 15510 10852 15516 10854
rect 15572 10852 15596 10854
rect 15652 10852 15676 10854
rect 15732 10852 15756 10854
rect 15812 10852 15818 10854
rect 15510 10843 15818 10852
rect 15660 10600 15712 10606
rect 15660 10542 15712 10548
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 15580 10266 15608 10406
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 15672 10130 15700 10542
rect 16028 10532 16080 10538
rect 16028 10474 16080 10480
rect 15936 10464 15988 10470
rect 15936 10406 15988 10412
rect 15948 10198 15976 10406
rect 15936 10192 15988 10198
rect 15936 10134 15988 10140
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 15844 9920 15896 9926
rect 15844 9862 15896 9868
rect 15510 9820 15818 9829
rect 15510 9818 15516 9820
rect 15572 9818 15596 9820
rect 15652 9818 15676 9820
rect 15732 9818 15756 9820
rect 15812 9818 15818 9820
rect 15572 9766 15574 9818
rect 15754 9766 15756 9818
rect 15510 9764 15516 9766
rect 15572 9764 15596 9766
rect 15652 9764 15676 9766
rect 15732 9764 15756 9766
rect 15812 9764 15818 9766
rect 15510 9755 15818 9764
rect 15510 8732 15818 8741
rect 15510 8730 15516 8732
rect 15572 8730 15596 8732
rect 15652 8730 15676 8732
rect 15732 8730 15756 8732
rect 15812 8730 15818 8732
rect 15572 8678 15574 8730
rect 15754 8678 15756 8730
rect 15510 8676 15516 8678
rect 15572 8676 15596 8678
rect 15652 8676 15676 8678
rect 15732 8676 15756 8678
rect 15812 8676 15818 8678
rect 15510 8667 15818 8676
rect 15856 8362 15884 9862
rect 16040 9466 16068 10474
rect 16132 10470 16160 11086
rect 16580 11076 16632 11082
rect 16580 11018 16632 11024
rect 16302 10568 16358 10577
rect 16302 10503 16358 10512
rect 16120 10464 16172 10470
rect 16172 10424 16252 10452
rect 16120 10406 16172 10412
rect 16224 10062 16252 10424
rect 16212 10056 16264 10062
rect 16212 9998 16264 10004
rect 16120 9716 16172 9722
rect 16120 9658 16172 9664
rect 15948 9438 16068 9466
rect 15948 8634 15976 9438
rect 16028 9376 16080 9382
rect 16028 9318 16080 9324
rect 15936 8628 15988 8634
rect 15936 8570 15988 8576
rect 15844 8356 15896 8362
rect 15844 8298 15896 8304
rect 15510 7644 15818 7653
rect 15510 7642 15516 7644
rect 15572 7642 15596 7644
rect 15652 7642 15676 7644
rect 15732 7642 15756 7644
rect 15812 7642 15818 7644
rect 15572 7590 15574 7642
rect 15754 7590 15756 7642
rect 15510 7588 15516 7590
rect 15572 7588 15596 7590
rect 15652 7588 15676 7590
rect 15732 7588 15756 7590
rect 15812 7588 15818 7590
rect 15510 7579 15818 7588
rect 15856 7410 15884 8298
rect 15844 7404 15896 7410
rect 15844 7346 15896 7352
rect 15936 7336 15988 7342
rect 15936 7278 15988 7284
rect 15752 7200 15804 7206
rect 15752 7142 15804 7148
rect 15764 6712 15792 7142
rect 15764 6684 15884 6712
rect 15510 6556 15818 6565
rect 15510 6554 15516 6556
rect 15572 6554 15596 6556
rect 15652 6554 15676 6556
rect 15732 6554 15756 6556
rect 15812 6554 15818 6556
rect 15572 6502 15574 6554
rect 15754 6502 15756 6554
rect 15510 6500 15516 6502
rect 15572 6500 15596 6502
rect 15652 6500 15676 6502
rect 15732 6500 15756 6502
rect 15812 6500 15818 6502
rect 15510 6491 15818 6500
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 15510 5468 15818 5477
rect 15510 5466 15516 5468
rect 15572 5466 15596 5468
rect 15652 5466 15676 5468
rect 15732 5466 15756 5468
rect 15812 5466 15818 5468
rect 15572 5414 15574 5466
rect 15754 5414 15756 5466
rect 15510 5412 15516 5414
rect 15572 5412 15596 5414
rect 15652 5412 15676 5414
rect 15732 5412 15756 5414
rect 15812 5412 15818 5414
rect 15510 5403 15818 5412
rect 15566 5264 15622 5273
rect 15566 5199 15622 5208
rect 15580 5166 15608 5199
rect 15568 5160 15620 5166
rect 15568 5102 15620 5108
rect 15856 5098 15884 6684
rect 15948 6458 15976 7278
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 15934 6352 15990 6361
rect 15934 6287 15990 6296
rect 15844 5092 15896 5098
rect 15844 5034 15896 5040
rect 15752 4752 15804 4758
rect 15750 4720 15752 4729
rect 15804 4720 15806 4729
rect 15750 4655 15806 4664
rect 15844 4480 15896 4486
rect 15844 4422 15896 4428
rect 15510 4380 15818 4389
rect 15510 4378 15516 4380
rect 15572 4378 15596 4380
rect 15652 4378 15676 4380
rect 15732 4378 15756 4380
rect 15812 4378 15818 4380
rect 15572 4326 15574 4378
rect 15754 4326 15756 4378
rect 15510 4324 15516 4326
rect 15572 4324 15596 4326
rect 15652 4324 15676 4326
rect 15732 4324 15756 4326
rect 15812 4324 15818 4326
rect 15510 4315 15818 4324
rect 15856 4282 15884 4422
rect 15844 4276 15896 4282
rect 15844 4218 15896 4224
rect 15948 4162 15976 6287
rect 16040 5846 16068 9318
rect 16132 8022 16160 9658
rect 16224 8090 16252 9998
rect 16212 8084 16264 8090
rect 16212 8026 16264 8032
rect 16120 8016 16172 8022
rect 16120 7958 16172 7964
rect 16120 7880 16172 7886
rect 16120 7822 16172 7828
rect 16132 7290 16160 7822
rect 16224 7449 16252 8026
rect 16210 7440 16266 7449
rect 16210 7375 16266 7384
rect 16212 7336 16264 7342
rect 16132 7284 16212 7290
rect 16132 7278 16264 7284
rect 16132 7262 16252 7278
rect 16132 6798 16160 7262
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 16224 7002 16252 7142
rect 16212 6996 16264 7002
rect 16212 6938 16264 6944
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 16120 6180 16172 6186
rect 16120 6122 16172 6128
rect 16028 5840 16080 5846
rect 16028 5782 16080 5788
rect 16026 5672 16082 5681
rect 16026 5607 16082 5616
rect 15856 4134 15976 4162
rect 15304 3998 15516 4026
rect 15200 3936 15252 3942
rect 15200 3878 15252 3884
rect 15212 3738 15240 3878
rect 15200 3732 15252 3738
rect 15200 3674 15252 3680
rect 15108 2848 15160 2854
rect 15108 2790 15160 2796
rect 15212 2514 15240 3674
rect 15488 3618 15516 3998
rect 15396 3590 15516 3618
rect 15292 3120 15344 3126
rect 15292 3062 15344 3068
rect 14924 2508 14976 2514
rect 14924 2450 14976 2456
rect 15200 2508 15252 2514
rect 15200 2450 15252 2456
rect 14832 1896 14884 1902
rect 14832 1838 14884 1844
rect 14648 1828 14700 1834
rect 14648 1770 14700 1776
rect 14740 1760 14792 1766
rect 14740 1702 14792 1708
rect 14752 1562 14780 1702
rect 14740 1556 14792 1562
rect 14740 1498 14792 1504
rect 14556 1284 14608 1290
rect 14556 1226 14608 1232
rect 14280 944 14332 950
rect 14280 886 14332 892
rect 14372 944 14424 950
rect 14372 886 14424 892
rect 14280 808 14332 814
rect 14278 776 14280 785
rect 14740 808 14792 814
rect 14332 776 14334 785
rect 14844 796 14872 1838
rect 14936 1426 14964 2450
rect 15198 2408 15254 2417
rect 15198 2343 15254 2352
rect 15014 2000 15070 2009
rect 15014 1935 15070 1944
rect 14924 1420 14976 1426
rect 14924 1362 14976 1368
rect 15028 814 15056 1935
rect 14792 768 14872 796
rect 15016 808 15068 814
rect 14740 750 14792 756
rect 15016 750 15068 756
rect 14278 711 14334 720
rect 13728 672 13780 678
rect 13728 614 13780 620
rect 14188 672 14240 678
rect 14188 614 14240 620
rect 13960 572 14268 581
rect 13960 570 13966 572
rect 14022 570 14046 572
rect 14102 570 14126 572
rect 14182 570 14206 572
rect 14262 570 14268 572
rect 14022 518 14024 570
rect 14204 518 14206 570
rect 13960 516 13966 518
rect 14022 516 14046 518
rect 14102 516 14126 518
rect 14182 516 14206 518
rect 14262 516 14268 518
rect 13960 507 14268 516
rect 15212 338 15240 2343
rect 15304 406 15332 3062
rect 15396 1018 15424 3590
rect 15510 3292 15818 3301
rect 15510 3290 15516 3292
rect 15572 3290 15596 3292
rect 15652 3290 15676 3292
rect 15732 3290 15756 3292
rect 15812 3290 15818 3292
rect 15572 3238 15574 3290
rect 15754 3238 15756 3290
rect 15510 3236 15516 3238
rect 15572 3236 15596 3238
rect 15652 3236 15676 3238
rect 15732 3236 15756 3238
rect 15812 3236 15818 3238
rect 15510 3227 15818 3236
rect 15752 3120 15804 3126
rect 15856 3074 15884 4134
rect 15936 3936 15988 3942
rect 15936 3878 15988 3884
rect 15948 3602 15976 3878
rect 15936 3596 15988 3602
rect 15936 3538 15988 3544
rect 15804 3068 15884 3074
rect 15752 3062 15884 3068
rect 15764 3046 15884 3062
rect 15844 2848 15896 2854
rect 15844 2790 15896 2796
rect 15936 2848 15988 2854
rect 15936 2790 15988 2796
rect 15856 2553 15884 2790
rect 15842 2544 15898 2553
rect 15842 2479 15898 2488
rect 15510 2204 15818 2213
rect 15510 2202 15516 2204
rect 15572 2202 15596 2204
rect 15652 2202 15676 2204
rect 15732 2202 15756 2204
rect 15812 2202 15818 2204
rect 15572 2150 15574 2202
rect 15754 2150 15756 2202
rect 15510 2148 15516 2150
rect 15572 2148 15596 2150
rect 15652 2148 15676 2150
rect 15732 2148 15756 2150
rect 15812 2148 15818 2150
rect 15510 2139 15818 2148
rect 15856 2038 15884 2479
rect 15844 2032 15896 2038
rect 15844 1974 15896 1980
rect 15474 1864 15530 1873
rect 15474 1799 15476 1808
rect 15528 1799 15530 1808
rect 15658 1864 15714 1873
rect 15658 1799 15714 1808
rect 15476 1770 15528 1776
rect 15488 1426 15516 1770
rect 15672 1766 15700 1799
rect 15660 1760 15712 1766
rect 15660 1702 15712 1708
rect 15844 1760 15896 1766
rect 15844 1702 15896 1708
rect 15476 1420 15528 1426
rect 15476 1362 15528 1368
rect 15510 1116 15818 1125
rect 15510 1114 15516 1116
rect 15572 1114 15596 1116
rect 15652 1114 15676 1116
rect 15732 1114 15756 1116
rect 15812 1114 15818 1116
rect 15572 1062 15574 1114
rect 15754 1062 15756 1114
rect 15510 1060 15516 1062
rect 15572 1060 15596 1062
rect 15652 1060 15676 1062
rect 15732 1060 15756 1062
rect 15812 1060 15818 1062
rect 15510 1051 15818 1060
rect 15384 1012 15436 1018
rect 15384 954 15436 960
rect 15856 921 15884 1702
rect 15842 912 15898 921
rect 15842 847 15898 856
rect 15948 474 15976 2790
rect 16040 2106 16068 5607
rect 16132 5370 16160 6122
rect 16224 6118 16252 6938
rect 16316 6361 16344 10503
rect 16488 10464 16540 10470
rect 16488 10406 16540 10412
rect 16500 10198 16528 10406
rect 16488 10192 16540 10198
rect 16488 10134 16540 10140
rect 16500 9722 16528 10134
rect 16488 9716 16540 9722
rect 16488 9658 16540 9664
rect 16592 9042 16620 11018
rect 17604 10538 17632 11358
rect 18510 11200 18566 12000
rect 17684 11144 17736 11150
rect 17684 11086 17736 11092
rect 18418 11112 18474 11121
rect 17696 10742 17724 11086
rect 18418 11047 18474 11056
rect 18236 11008 18288 11014
rect 18236 10950 18288 10956
rect 18248 10810 18276 10950
rect 17960 10804 18012 10810
rect 17960 10746 18012 10752
rect 18236 10804 18288 10810
rect 18236 10746 18288 10752
rect 17684 10736 17736 10742
rect 17684 10678 17736 10684
rect 17776 10600 17828 10606
rect 17776 10542 17828 10548
rect 17868 10600 17920 10606
rect 17868 10542 17920 10548
rect 17592 10532 17644 10538
rect 17592 10474 17644 10480
rect 17060 10364 17368 10373
rect 17060 10362 17066 10364
rect 17122 10362 17146 10364
rect 17202 10362 17226 10364
rect 17282 10362 17306 10364
rect 17362 10362 17368 10364
rect 17122 10310 17124 10362
rect 17304 10310 17306 10362
rect 17060 10308 17066 10310
rect 17122 10308 17146 10310
rect 17202 10308 17226 10310
rect 17282 10308 17306 10310
rect 17362 10308 17368 10310
rect 17060 10299 17368 10308
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17512 10130 17540 10202
rect 17500 10124 17552 10130
rect 17500 10066 17552 10072
rect 16764 9920 16816 9926
rect 16764 9862 16816 9868
rect 16856 9920 16908 9926
rect 16856 9862 16908 9868
rect 16776 9586 16804 9862
rect 16764 9580 16816 9586
rect 16764 9522 16816 9528
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 16580 9036 16632 9042
rect 16580 8978 16632 8984
rect 16684 8906 16712 9454
rect 16868 8974 16896 9862
rect 17408 9512 17460 9518
rect 17408 9454 17460 9460
rect 17060 9276 17368 9285
rect 17060 9274 17066 9276
rect 17122 9274 17146 9276
rect 17202 9274 17226 9276
rect 17282 9274 17306 9276
rect 17362 9274 17368 9276
rect 17122 9222 17124 9274
rect 17304 9222 17306 9274
rect 17060 9220 17066 9222
rect 17122 9220 17146 9222
rect 17202 9220 17226 9222
rect 17282 9220 17306 9222
rect 17362 9220 17368 9222
rect 17060 9211 17368 9220
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 16672 8900 16724 8906
rect 16672 8842 16724 8848
rect 16764 8832 16816 8838
rect 16764 8774 16816 8780
rect 16776 8430 16804 8774
rect 16764 8424 16816 8430
rect 16764 8366 16816 8372
rect 16948 8424 17000 8430
rect 16948 8366 17000 8372
rect 16488 8016 16540 8022
rect 16408 7976 16488 8004
rect 16408 7206 16436 7976
rect 16488 7958 16540 7964
rect 16672 8016 16724 8022
rect 16776 8004 16804 8366
rect 16856 8288 16908 8294
rect 16856 8230 16908 8236
rect 16724 7976 16804 8004
rect 16672 7958 16724 7964
rect 16580 7540 16632 7546
rect 16580 7482 16632 7488
rect 16396 7200 16448 7206
rect 16396 7142 16448 7148
rect 16408 6934 16436 7142
rect 16396 6928 16448 6934
rect 16396 6870 16448 6876
rect 16302 6352 16358 6361
rect 16302 6287 16358 6296
rect 16408 6225 16436 6870
rect 16488 6452 16540 6458
rect 16488 6394 16540 6400
rect 16394 6216 16450 6225
rect 16394 6151 16450 6160
rect 16212 6112 16264 6118
rect 16212 6054 16264 6060
rect 16304 6112 16356 6118
rect 16304 6054 16356 6060
rect 16120 5364 16172 5370
rect 16120 5306 16172 5312
rect 16118 4856 16174 4865
rect 16118 4791 16174 4800
rect 16132 4758 16160 4791
rect 16120 4752 16172 4758
rect 16120 4694 16172 4700
rect 16224 4622 16252 6054
rect 16212 4616 16264 4622
rect 16212 4558 16264 4564
rect 16120 4140 16172 4146
rect 16120 4082 16172 4088
rect 16132 4010 16160 4082
rect 16120 4004 16172 4010
rect 16120 3946 16172 3952
rect 16028 2100 16080 2106
rect 16028 2042 16080 2048
rect 16028 1556 16080 1562
rect 16028 1498 16080 1504
rect 16040 1290 16068 1498
rect 16028 1284 16080 1290
rect 16028 1226 16080 1232
rect 16028 876 16080 882
rect 16028 818 16080 824
rect 16040 678 16068 818
rect 16132 746 16160 3946
rect 16224 3602 16252 4558
rect 16212 3596 16264 3602
rect 16212 3538 16264 3544
rect 16316 3466 16344 6054
rect 16396 5840 16448 5846
rect 16396 5782 16448 5788
rect 16408 4457 16436 5782
rect 16500 5302 16528 6394
rect 16592 6322 16620 7482
rect 16672 7268 16724 7274
rect 16672 7210 16724 7216
rect 16684 6458 16712 7210
rect 16776 6905 16804 7976
rect 16868 7954 16896 8230
rect 16856 7948 16908 7954
rect 16856 7890 16908 7896
rect 16762 6896 16818 6905
rect 16762 6831 16818 6840
rect 16672 6452 16724 6458
rect 16672 6394 16724 6400
rect 16776 6338 16804 6831
rect 16868 6662 16896 7890
rect 16960 6866 16988 8366
rect 17420 8294 17448 9454
rect 17512 9058 17540 10066
rect 17604 9586 17632 10474
rect 17788 9586 17816 10542
rect 17880 10130 17908 10542
rect 17868 10124 17920 10130
rect 17868 10066 17920 10072
rect 17868 9988 17920 9994
rect 17868 9930 17920 9936
rect 17880 9654 17908 9930
rect 17972 9926 18000 10746
rect 18236 10668 18288 10674
rect 18236 10610 18288 10616
rect 18144 10600 18196 10606
rect 18144 10542 18196 10548
rect 18156 10198 18184 10542
rect 18144 10192 18196 10198
rect 18144 10134 18196 10140
rect 17960 9920 18012 9926
rect 17960 9862 18012 9868
rect 17868 9648 17920 9654
rect 17868 9590 17920 9596
rect 17592 9580 17644 9586
rect 17592 9522 17644 9528
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 17776 9444 17828 9450
rect 17776 9386 17828 9392
rect 17788 9110 17816 9386
rect 18052 9376 18104 9382
rect 18052 9318 18104 9324
rect 17776 9104 17828 9110
rect 17512 9030 17632 9058
rect 17776 9046 17828 9052
rect 17500 8968 17552 8974
rect 17500 8910 17552 8916
rect 17512 8362 17540 8910
rect 17604 8906 17632 9030
rect 17592 8900 17644 8906
rect 17592 8842 17644 8848
rect 17604 8566 17632 8842
rect 17592 8560 17644 8566
rect 17592 8502 17644 8508
rect 17500 8356 17552 8362
rect 17500 8298 17552 8304
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17060 8188 17368 8197
rect 17060 8186 17066 8188
rect 17122 8186 17146 8188
rect 17202 8186 17226 8188
rect 17282 8186 17306 8188
rect 17362 8186 17368 8188
rect 17122 8134 17124 8186
rect 17304 8134 17306 8186
rect 17060 8132 17066 8134
rect 17122 8132 17146 8134
rect 17202 8132 17226 8134
rect 17282 8132 17306 8134
rect 17362 8132 17368 8134
rect 17060 8123 17368 8132
rect 17420 8090 17448 8230
rect 17316 8084 17368 8090
rect 17316 8026 17368 8032
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 17224 7948 17276 7954
rect 17224 7890 17276 7896
rect 17236 7410 17264 7890
rect 17328 7886 17356 8026
rect 17408 7948 17460 7954
rect 17460 7908 17540 7936
rect 17408 7890 17460 7896
rect 17316 7880 17368 7886
rect 17316 7822 17368 7828
rect 17408 7744 17460 7750
rect 17408 7686 17460 7692
rect 17224 7404 17276 7410
rect 17224 7346 17276 7352
rect 17060 7100 17368 7109
rect 17060 7098 17066 7100
rect 17122 7098 17146 7100
rect 17202 7098 17226 7100
rect 17282 7098 17306 7100
rect 17362 7098 17368 7100
rect 17122 7046 17124 7098
rect 17304 7046 17306 7098
rect 17060 7044 17066 7046
rect 17122 7044 17146 7046
rect 17202 7044 17226 7046
rect 17282 7044 17306 7046
rect 17362 7044 17368 7046
rect 17060 7035 17368 7044
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 17132 6860 17184 6866
rect 17132 6802 17184 6808
rect 16856 6656 16908 6662
rect 16856 6598 16908 6604
rect 16580 6316 16632 6322
rect 16580 6258 16632 6264
rect 16684 6310 16804 6338
rect 16684 5642 16712 6310
rect 16764 5772 16816 5778
rect 16764 5714 16816 5720
rect 16672 5636 16724 5642
rect 16672 5578 16724 5584
rect 16488 5296 16540 5302
rect 16488 5238 16540 5244
rect 16670 5264 16726 5273
rect 16394 4448 16450 4457
rect 16394 4383 16450 4392
rect 16394 4176 16450 4185
rect 16394 4111 16450 4120
rect 16212 3460 16264 3466
rect 16212 3402 16264 3408
rect 16304 3460 16356 3466
rect 16304 3402 16356 3408
rect 16224 2310 16252 3402
rect 16302 3360 16358 3369
rect 16302 3295 16358 3304
rect 16212 2304 16264 2310
rect 16316 2292 16344 3295
rect 16408 2417 16436 4111
rect 16500 3942 16528 5238
rect 16670 5199 16672 5208
rect 16724 5199 16726 5208
rect 16672 5170 16724 5176
rect 16684 4729 16712 5170
rect 16670 4720 16726 4729
rect 16580 4684 16632 4690
rect 16670 4655 16726 4664
rect 16580 4626 16632 4632
rect 16592 4146 16620 4626
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 16580 4140 16632 4146
rect 16580 4082 16632 4088
rect 16578 4040 16634 4049
rect 16578 3975 16580 3984
rect 16632 3975 16634 3984
rect 16580 3946 16632 3952
rect 16488 3936 16540 3942
rect 16488 3878 16540 3884
rect 16500 3602 16528 3878
rect 16488 3596 16540 3602
rect 16488 3538 16540 3544
rect 16488 3460 16540 3466
rect 16488 3402 16540 3408
rect 16394 2408 16450 2417
rect 16394 2343 16450 2352
rect 16396 2304 16448 2310
rect 16316 2264 16396 2292
rect 16212 2246 16264 2252
rect 16396 2246 16448 2252
rect 16302 2136 16358 2145
rect 16302 2071 16304 2080
rect 16356 2071 16358 2080
rect 16304 2042 16356 2048
rect 16302 2000 16358 2009
rect 16302 1935 16358 1944
rect 16316 1834 16344 1935
rect 16304 1828 16356 1834
rect 16304 1770 16356 1776
rect 16212 1760 16264 1766
rect 16212 1702 16264 1708
rect 16224 1018 16252 1702
rect 16408 1358 16436 2246
rect 16396 1352 16448 1358
rect 16396 1294 16448 1300
rect 16212 1012 16264 1018
rect 16212 954 16264 960
rect 16500 950 16528 3402
rect 16684 3398 16712 4558
rect 16776 4146 16804 5714
rect 16868 5710 16896 6598
rect 16856 5704 16908 5710
rect 16856 5646 16908 5652
rect 16856 5568 16908 5574
rect 16856 5510 16908 5516
rect 16868 5166 16896 5510
rect 16856 5160 16908 5166
rect 16856 5102 16908 5108
rect 16856 4820 16908 4826
rect 16856 4762 16908 4768
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 16672 3392 16724 3398
rect 16672 3334 16724 3340
rect 16578 2680 16634 2689
rect 16578 2615 16634 2624
rect 16592 1562 16620 2615
rect 16684 2514 16712 3334
rect 16776 2825 16804 4082
rect 16762 2816 16818 2825
rect 16762 2751 16818 2760
rect 16868 2582 16896 4762
rect 16960 3652 16988 6802
rect 17144 6769 17172 6802
rect 17130 6760 17186 6769
rect 17130 6695 17186 6704
rect 17060 6012 17368 6021
rect 17060 6010 17066 6012
rect 17122 6010 17146 6012
rect 17202 6010 17226 6012
rect 17282 6010 17306 6012
rect 17362 6010 17368 6012
rect 17122 5958 17124 6010
rect 17304 5958 17306 6010
rect 17060 5956 17066 5958
rect 17122 5956 17146 5958
rect 17202 5956 17226 5958
rect 17282 5956 17306 5958
rect 17362 5956 17368 5958
rect 17060 5947 17368 5956
rect 17132 5908 17184 5914
rect 17132 5850 17184 5856
rect 17316 5908 17368 5914
rect 17316 5850 17368 5856
rect 17144 5817 17172 5850
rect 17130 5808 17186 5817
rect 17130 5743 17186 5752
rect 17224 5772 17276 5778
rect 17224 5714 17276 5720
rect 17236 5642 17264 5714
rect 17224 5636 17276 5642
rect 17224 5578 17276 5584
rect 17040 5568 17092 5574
rect 17040 5510 17092 5516
rect 17052 5098 17080 5510
rect 17132 5296 17184 5302
rect 17236 5273 17264 5578
rect 17132 5238 17184 5244
rect 17222 5264 17278 5273
rect 17144 5148 17172 5238
rect 17222 5199 17278 5208
rect 17224 5160 17276 5166
rect 17144 5120 17224 5148
rect 17224 5102 17276 5108
rect 17328 5098 17356 5850
rect 17040 5092 17092 5098
rect 17040 5034 17092 5040
rect 17316 5092 17368 5098
rect 17316 5034 17368 5040
rect 17420 5030 17448 7686
rect 17512 5914 17540 7908
rect 17500 5908 17552 5914
rect 17500 5850 17552 5856
rect 17500 5704 17552 5710
rect 17500 5646 17552 5652
rect 17512 5370 17540 5646
rect 17500 5364 17552 5370
rect 17500 5306 17552 5312
rect 17604 5234 17632 8502
rect 17684 8492 17736 8498
rect 17684 8434 17736 8440
rect 17696 7954 17724 8434
rect 17684 7948 17736 7954
rect 17684 7890 17736 7896
rect 17696 6118 17724 7890
rect 17788 6254 17816 9046
rect 17960 8288 18012 8294
rect 17960 8230 18012 8236
rect 17868 7880 17920 7886
rect 17868 7822 17920 7828
rect 17880 6390 17908 7822
rect 17868 6384 17920 6390
rect 17868 6326 17920 6332
rect 17972 6254 18000 8230
rect 18064 6458 18092 9318
rect 18156 8090 18184 10134
rect 18248 10130 18276 10610
rect 18432 10606 18460 11047
rect 18420 10600 18472 10606
rect 18418 10568 18420 10577
rect 18472 10568 18474 10577
rect 18418 10503 18474 10512
rect 18236 10124 18288 10130
rect 18236 10066 18288 10072
rect 18328 10124 18380 10130
rect 18328 10066 18380 10072
rect 18340 9994 18368 10066
rect 18328 9988 18380 9994
rect 18328 9930 18380 9936
rect 18236 9920 18288 9926
rect 18236 9862 18288 9868
rect 18248 9722 18276 9862
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 18052 6452 18104 6458
rect 18052 6394 18104 6400
rect 17776 6248 17828 6254
rect 17960 6248 18012 6254
rect 17828 6208 17908 6236
rect 17776 6190 17828 6196
rect 17684 6112 17736 6118
rect 17684 6054 17736 6060
rect 17696 5642 17724 6054
rect 17776 5704 17828 5710
rect 17776 5646 17828 5652
rect 17684 5636 17736 5642
rect 17684 5578 17736 5584
rect 17592 5228 17644 5234
rect 17592 5170 17644 5176
rect 17696 5166 17724 5578
rect 17788 5234 17816 5646
rect 17880 5370 17908 6208
rect 17960 6190 18012 6196
rect 18052 6180 18104 6186
rect 18052 6122 18104 6128
rect 18064 5914 18092 6122
rect 18052 5908 18104 5914
rect 18052 5850 18104 5856
rect 18144 5840 18196 5846
rect 17958 5808 18014 5817
rect 18144 5782 18196 5788
rect 17958 5743 18014 5752
rect 18052 5772 18104 5778
rect 17868 5364 17920 5370
rect 17868 5306 17920 5312
rect 17866 5264 17922 5273
rect 17776 5228 17828 5234
rect 17866 5199 17922 5208
rect 17776 5170 17828 5176
rect 17684 5160 17736 5166
rect 17684 5102 17736 5108
rect 17592 5092 17644 5098
rect 17592 5034 17644 5040
rect 17408 5024 17460 5030
rect 17408 4966 17460 4972
rect 17060 4924 17368 4933
rect 17060 4922 17066 4924
rect 17122 4922 17146 4924
rect 17202 4922 17226 4924
rect 17282 4922 17306 4924
rect 17362 4922 17368 4924
rect 17122 4870 17124 4922
rect 17304 4870 17306 4922
rect 17060 4868 17066 4870
rect 17122 4868 17146 4870
rect 17202 4868 17226 4870
rect 17282 4868 17306 4870
rect 17362 4868 17368 4870
rect 17060 4859 17368 4868
rect 17604 4826 17632 5034
rect 17592 4820 17644 4826
rect 17592 4762 17644 4768
rect 17224 4684 17276 4690
rect 17224 4626 17276 4632
rect 17130 4448 17186 4457
rect 17130 4383 17186 4392
rect 17144 3942 17172 4383
rect 17236 4214 17264 4626
rect 17498 4584 17554 4593
rect 17498 4519 17554 4528
rect 17592 4548 17644 4554
rect 17316 4480 17368 4486
rect 17314 4448 17316 4457
rect 17408 4480 17460 4486
rect 17368 4448 17370 4457
rect 17408 4422 17460 4428
rect 17314 4383 17370 4392
rect 17224 4208 17276 4214
rect 17224 4150 17276 4156
rect 17132 3936 17184 3942
rect 17132 3878 17184 3884
rect 17060 3836 17368 3845
rect 17060 3834 17066 3836
rect 17122 3834 17146 3836
rect 17202 3834 17226 3836
rect 17282 3834 17306 3836
rect 17362 3834 17368 3836
rect 17122 3782 17124 3834
rect 17304 3782 17306 3834
rect 17060 3780 17066 3782
rect 17122 3780 17146 3782
rect 17202 3780 17226 3782
rect 17282 3780 17306 3782
rect 17362 3780 17368 3782
rect 17060 3771 17368 3780
rect 17132 3664 17184 3670
rect 16960 3624 17080 3652
rect 16946 3360 17002 3369
rect 16946 3295 17002 3304
rect 16856 2576 16908 2582
rect 16856 2518 16908 2524
rect 16672 2508 16724 2514
rect 16724 2468 16804 2496
rect 16672 2450 16724 2456
rect 16672 2372 16724 2378
rect 16672 2314 16724 2320
rect 16580 1556 16632 1562
rect 16580 1498 16632 1504
rect 16488 944 16540 950
rect 16488 886 16540 892
rect 16684 746 16712 2314
rect 16776 1970 16804 2468
rect 16854 2408 16910 2417
rect 16854 2343 16910 2352
rect 16868 1970 16896 2343
rect 16764 1964 16816 1970
rect 16764 1906 16816 1912
rect 16856 1964 16908 1970
rect 16856 1906 16908 1912
rect 16960 1952 16988 3295
rect 17052 2938 17080 3624
rect 17132 3606 17184 3612
rect 17314 3632 17370 3641
rect 17144 3194 17172 3606
rect 17314 3567 17370 3576
rect 17224 3528 17276 3534
rect 17224 3470 17276 3476
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 17236 3097 17264 3470
rect 17328 3126 17356 3567
rect 17316 3120 17368 3126
rect 17222 3088 17278 3097
rect 17316 3062 17368 3068
rect 17420 3058 17448 4422
rect 17512 3534 17540 4519
rect 17592 4490 17644 4496
rect 17500 3528 17552 3534
rect 17500 3470 17552 3476
rect 17512 3369 17540 3470
rect 17498 3360 17554 3369
rect 17498 3295 17554 3304
rect 17500 3188 17552 3194
rect 17604 3176 17632 4490
rect 17776 4208 17828 4214
rect 17776 4150 17828 4156
rect 17684 3936 17736 3942
rect 17684 3878 17736 3884
rect 17696 3602 17724 3878
rect 17684 3596 17736 3602
rect 17684 3538 17736 3544
rect 17696 3369 17724 3538
rect 17788 3398 17816 4150
rect 17776 3392 17828 3398
rect 17682 3360 17738 3369
rect 17776 3334 17828 3340
rect 17682 3295 17738 3304
rect 17880 3194 17908 5199
rect 17972 4826 18000 5743
rect 18052 5714 18104 5720
rect 18064 5545 18092 5714
rect 18050 5536 18106 5545
rect 18050 5471 18106 5480
rect 18052 5160 18104 5166
rect 18052 5102 18104 5108
rect 17960 4820 18012 4826
rect 17960 4762 18012 4768
rect 17960 4276 18012 4282
rect 17960 4218 18012 4224
rect 17972 3466 18000 4218
rect 18064 4214 18092 5102
rect 18156 5098 18184 5782
rect 18248 5574 18276 9658
rect 18340 8634 18368 9930
rect 18328 8628 18380 8634
rect 18328 8570 18380 8576
rect 18340 8537 18368 8570
rect 18326 8528 18382 8537
rect 18326 8463 18382 8472
rect 18328 8424 18380 8430
rect 18380 8384 18460 8412
rect 18328 8366 18380 8372
rect 18432 7954 18460 8384
rect 18420 7948 18472 7954
rect 18420 7890 18472 7896
rect 18328 7812 18380 7818
rect 18328 7754 18380 7760
rect 18340 7478 18368 7754
rect 18328 7472 18380 7478
rect 18328 7414 18380 7420
rect 18432 7290 18460 7890
rect 18524 7546 18552 11200
rect 18610 10908 18918 10917
rect 18610 10906 18616 10908
rect 18672 10906 18696 10908
rect 18752 10906 18776 10908
rect 18832 10906 18856 10908
rect 18912 10906 18918 10908
rect 18672 10854 18674 10906
rect 18854 10854 18856 10906
rect 18610 10852 18616 10854
rect 18672 10852 18696 10854
rect 18752 10852 18776 10854
rect 18832 10852 18856 10854
rect 18912 10852 18918 10854
rect 18610 10843 18918 10852
rect 18610 9820 18918 9829
rect 18610 9818 18616 9820
rect 18672 9818 18696 9820
rect 18752 9818 18776 9820
rect 18832 9818 18856 9820
rect 18912 9818 18918 9820
rect 18672 9766 18674 9818
rect 18854 9766 18856 9818
rect 18610 9764 18616 9766
rect 18672 9764 18696 9766
rect 18752 9764 18776 9766
rect 18832 9764 18856 9766
rect 18912 9764 18918 9766
rect 18610 9755 18918 9764
rect 18610 8732 18918 8741
rect 18610 8730 18616 8732
rect 18672 8730 18696 8732
rect 18752 8730 18776 8732
rect 18832 8730 18856 8732
rect 18912 8730 18918 8732
rect 18672 8678 18674 8730
rect 18854 8678 18856 8730
rect 18610 8676 18616 8678
rect 18672 8676 18696 8678
rect 18752 8676 18776 8678
rect 18832 8676 18856 8678
rect 18912 8676 18918 8678
rect 18610 8667 18918 8676
rect 18970 8256 19026 8265
rect 18970 8191 19026 8200
rect 18610 7644 18918 7653
rect 18610 7642 18616 7644
rect 18672 7642 18696 7644
rect 18752 7642 18776 7644
rect 18832 7642 18856 7644
rect 18912 7642 18918 7644
rect 18672 7590 18674 7642
rect 18854 7590 18856 7642
rect 18610 7588 18616 7590
rect 18672 7588 18696 7590
rect 18752 7588 18776 7590
rect 18832 7588 18856 7590
rect 18912 7588 18918 7590
rect 18610 7579 18918 7588
rect 18512 7540 18564 7546
rect 18512 7482 18564 7488
rect 18340 7262 18460 7290
rect 18512 7336 18564 7342
rect 18512 7278 18564 7284
rect 18340 7206 18368 7262
rect 18328 7200 18380 7206
rect 18328 7142 18380 7148
rect 18340 5642 18368 7142
rect 18524 6769 18552 7278
rect 18510 6760 18566 6769
rect 18510 6695 18566 6704
rect 18420 6384 18472 6390
rect 18420 6326 18472 6332
rect 18432 5846 18460 6326
rect 18420 5840 18472 5846
rect 18420 5782 18472 5788
rect 18524 5681 18552 6695
rect 18610 6556 18918 6565
rect 18610 6554 18616 6556
rect 18672 6554 18696 6556
rect 18752 6554 18776 6556
rect 18832 6554 18856 6556
rect 18912 6554 18918 6556
rect 18672 6502 18674 6554
rect 18854 6502 18856 6554
rect 18610 6500 18616 6502
rect 18672 6500 18696 6502
rect 18752 6500 18776 6502
rect 18832 6500 18856 6502
rect 18912 6500 18918 6502
rect 18610 6491 18918 6500
rect 18984 6254 19012 8191
rect 18972 6248 19024 6254
rect 18972 6190 19024 6196
rect 18510 5672 18566 5681
rect 18328 5636 18380 5642
rect 18510 5607 18566 5616
rect 18328 5578 18380 5584
rect 18236 5568 18288 5574
rect 18236 5510 18288 5516
rect 18610 5468 18918 5477
rect 18610 5466 18616 5468
rect 18672 5466 18696 5468
rect 18752 5466 18776 5468
rect 18832 5466 18856 5468
rect 18912 5466 18918 5468
rect 18672 5414 18674 5466
rect 18854 5414 18856 5466
rect 18610 5412 18616 5414
rect 18672 5412 18696 5414
rect 18752 5412 18776 5414
rect 18832 5412 18856 5414
rect 18912 5412 18918 5414
rect 18610 5403 18918 5412
rect 18970 5264 19026 5273
rect 18970 5199 19026 5208
rect 18144 5092 18196 5098
rect 18144 5034 18196 5040
rect 18420 5024 18472 5030
rect 18420 4966 18472 4972
rect 18144 4684 18196 4690
rect 18144 4626 18196 4632
rect 18328 4684 18380 4690
rect 18328 4626 18380 4632
rect 18052 4208 18104 4214
rect 18052 4150 18104 4156
rect 18052 4072 18104 4078
rect 18052 4014 18104 4020
rect 17960 3460 18012 3466
rect 17960 3402 18012 3408
rect 18064 3194 18092 4014
rect 17868 3188 17920 3194
rect 17604 3148 17816 3176
rect 17500 3130 17552 3136
rect 17222 3023 17278 3032
rect 17408 3052 17460 3058
rect 17408 2994 17460 3000
rect 17052 2910 17448 2938
rect 17060 2748 17368 2757
rect 17060 2746 17066 2748
rect 17122 2746 17146 2748
rect 17202 2746 17226 2748
rect 17282 2746 17306 2748
rect 17362 2746 17368 2748
rect 17122 2694 17124 2746
rect 17304 2694 17306 2746
rect 17060 2692 17066 2694
rect 17122 2692 17146 2694
rect 17202 2692 17226 2694
rect 17282 2692 17306 2694
rect 17362 2692 17368 2694
rect 17060 2683 17368 2692
rect 17132 2576 17184 2582
rect 17132 2518 17184 2524
rect 17040 2508 17092 2514
rect 17040 2450 17092 2456
rect 17052 2106 17080 2450
rect 17040 2100 17092 2106
rect 17040 2042 17092 2048
rect 17040 1964 17092 1970
rect 16960 1924 17040 1952
rect 16776 1222 16804 1906
rect 16856 1828 16908 1834
rect 16856 1770 16908 1776
rect 16868 1290 16896 1770
rect 16960 1494 16988 1924
rect 17040 1906 17092 1912
rect 17144 1902 17172 2518
rect 17224 2440 17276 2446
rect 17224 2382 17276 2388
rect 17132 1896 17184 1902
rect 17132 1838 17184 1844
rect 17236 1834 17264 2382
rect 17224 1828 17276 1834
rect 17224 1770 17276 1776
rect 17060 1660 17368 1669
rect 17060 1658 17066 1660
rect 17122 1658 17146 1660
rect 17202 1658 17226 1660
rect 17282 1658 17306 1660
rect 17362 1658 17368 1660
rect 17122 1606 17124 1658
rect 17304 1606 17306 1658
rect 17060 1604 17066 1606
rect 17122 1604 17146 1606
rect 17202 1604 17226 1606
rect 17282 1604 17306 1606
rect 17362 1604 17368 1606
rect 17060 1595 17368 1604
rect 17420 1494 17448 2910
rect 16948 1488 17000 1494
rect 16948 1430 17000 1436
rect 17408 1488 17460 1494
rect 17408 1430 17460 1436
rect 17408 1352 17460 1358
rect 17406 1320 17408 1329
rect 17460 1320 17462 1329
rect 16856 1284 16908 1290
rect 16856 1226 16908 1232
rect 17316 1284 17368 1290
rect 17406 1255 17462 1264
rect 17316 1226 17368 1232
rect 16764 1216 16816 1222
rect 16764 1158 16816 1164
rect 17132 1216 17184 1222
rect 17132 1158 17184 1164
rect 17144 1018 17172 1158
rect 17328 1018 17356 1226
rect 17132 1012 17184 1018
rect 17132 954 17184 960
rect 17316 1012 17368 1018
rect 17316 954 17368 960
rect 17420 746 17448 1255
rect 17512 1222 17540 3130
rect 17682 3088 17738 3097
rect 17682 3023 17738 3032
rect 17592 2984 17644 2990
rect 17592 2926 17644 2932
rect 17604 2446 17632 2926
rect 17592 2440 17644 2446
rect 17592 2382 17644 2388
rect 17592 1964 17644 1970
rect 17592 1906 17644 1912
rect 17500 1216 17552 1222
rect 17500 1158 17552 1164
rect 17604 882 17632 1906
rect 17592 876 17644 882
rect 17592 818 17644 824
rect 17696 814 17724 3023
rect 17788 2854 17816 3148
rect 17868 3130 17920 3136
rect 18052 3188 18104 3194
rect 18052 3130 18104 3136
rect 17868 2984 17920 2990
rect 17868 2926 17920 2932
rect 18050 2952 18106 2961
rect 17776 2848 17828 2854
rect 17776 2790 17828 2796
rect 17788 2417 17816 2790
rect 17774 2408 17830 2417
rect 17774 2343 17830 2352
rect 17776 2304 17828 2310
rect 17776 2246 17828 2252
rect 17788 1426 17816 2246
rect 17880 2009 17908 2926
rect 18050 2887 18106 2896
rect 18064 2514 18092 2887
rect 18052 2508 18104 2514
rect 18052 2450 18104 2456
rect 17960 2440 18012 2446
rect 17960 2382 18012 2388
rect 17972 2145 18000 2382
rect 18052 2304 18104 2310
rect 18052 2246 18104 2252
rect 17958 2136 18014 2145
rect 17958 2071 18014 2080
rect 17866 2000 17922 2009
rect 17866 1935 17922 1944
rect 17868 1896 17920 1902
rect 17868 1838 17920 1844
rect 17880 1562 17908 1838
rect 17868 1556 17920 1562
rect 17868 1498 17920 1504
rect 18064 1465 18092 2246
rect 18156 1562 18184 4626
rect 18236 4548 18288 4554
rect 18236 4490 18288 4496
rect 18248 4146 18276 4490
rect 18236 4140 18288 4146
rect 18236 4082 18288 4088
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 18248 3670 18276 3878
rect 18236 3664 18288 3670
rect 18236 3606 18288 3612
rect 18234 3496 18290 3505
rect 18234 3431 18290 3440
rect 18144 1556 18196 1562
rect 18144 1498 18196 1504
rect 18050 1456 18106 1465
rect 17776 1420 17828 1426
rect 18050 1391 18052 1400
rect 17776 1362 17828 1368
rect 18104 1391 18106 1400
rect 18052 1362 18104 1368
rect 18064 1331 18092 1362
rect 18248 1018 18276 3431
rect 18236 1012 18288 1018
rect 18236 954 18288 960
rect 17684 808 17736 814
rect 17868 808 17920 814
rect 17684 750 17736 756
rect 17866 776 17868 785
rect 17920 776 17922 785
rect 16120 740 16172 746
rect 16120 682 16172 688
rect 16672 740 16724 746
rect 16672 682 16724 688
rect 16856 740 16908 746
rect 16856 682 16908 688
rect 17408 740 17460 746
rect 17866 711 17922 720
rect 17408 682 17460 688
rect 16028 672 16080 678
rect 16028 614 16080 620
rect 16488 672 16540 678
rect 16488 614 16540 620
rect 15936 468 15988 474
rect 15936 410 15988 416
rect 15292 400 15344 406
rect 15292 342 15344 348
rect 15200 332 15252 338
rect 15200 274 15252 280
rect 16500 202 16528 614
rect 16868 270 16896 682
rect 18340 678 18368 4626
rect 18432 3602 18460 4966
rect 18610 4380 18918 4389
rect 18610 4378 18616 4380
rect 18672 4378 18696 4380
rect 18752 4378 18776 4380
rect 18832 4378 18856 4380
rect 18912 4378 18918 4380
rect 18672 4326 18674 4378
rect 18854 4326 18856 4378
rect 18610 4324 18616 4326
rect 18672 4324 18696 4326
rect 18752 4324 18776 4326
rect 18832 4324 18856 4326
rect 18912 4324 18918 4326
rect 18610 4315 18918 4324
rect 18984 4185 19012 5199
rect 19156 5092 19208 5098
rect 19156 5034 19208 5040
rect 19064 4616 19116 4622
rect 19064 4558 19116 4564
rect 18970 4176 19026 4185
rect 18604 4140 18656 4146
rect 18970 4111 19026 4120
rect 18604 4082 18656 4088
rect 18512 4072 18564 4078
rect 18512 4014 18564 4020
rect 18420 3596 18472 3602
rect 18420 3538 18472 3544
rect 18420 3460 18472 3466
rect 18420 3402 18472 3408
rect 18432 2310 18460 3402
rect 18420 2304 18472 2310
rect 18420 2246 18472 2252
rect 18524 2106 18552 4014
rect 18616 3534 18644 4082
rect 18984 3890 19012 4111
rect 18892 3862 19012 3890
rect 18892 3602 18920 3862
rect 18970 3768 19026 3777
rect 19076 3738 19104 4558
rect 18970 3703 19026 3712
rect 19064 3732 19116 3738
rect 18880 3596 18932 3602
rect 18880 3538 18932 3544
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 18610 3292 18918 3301
rect 18610 3290 18616 3292
rect 18672 3290 18696 3292
rect 18752 3290 18776 3292
rect 18832 3290 18856 3292
rect 18912 3290 18918 3292
rect 18672 3238 18674 3290
rect 18854 3238 18856 3290
rect 18610 3236 18616 3238
rect 18672 3236 18696 3238
rect 18752 3236 18776 3238
rect 18832 3236 18856 3238
rect 18912 3236 18918 3238
rect 18610 3227 18918 3236
rect 18984 2990 19012 3703
rect 19064 3674 19116 3680
rect 18972 2984 19024 2990
rect 18972 2926 19024 2932
rect 19168 2650 19196 5034
rect 19156 2644 19208 2650
rect 19156 2586 19208 2592
rect 19062 2272 19118 2281
rect 18610 2204 18918 2213
rect 19062 2207 19118 2216
rect 18610 2202 18616 2204
rect 18672 2202 18696 2204
rect 18752 2202 18776 2204
rect 18832 2202 18856 2204
rect 18912 2202 18918 2204
rect 18672 2150 18674 2202
rect 18854 2150 18856 2202
rect 18610 2148 18616 2150
rect 18672 2148 18696 2150
rect 18752 2148 18776 2150
rect 18832 2148 18856 2150
rect 18912 2148 18918 2150
rect 18610 2139 18918 2148
rect 18512 2100 18564 2106
rect 18512 2042 18564 2048
rect 18510 2000 18566 2009
rect 18510 1935 18566 1944
rect 18524 1902 18552 1935
rect 18512 1896 18564 1902
rect 18512 1838 18564 1844
rect 18610 1116 18918 1125
rect 18610 1114 18616 1116
rect 18672 1114 18696 1116
rect 18752 1114 18776 1116
rect 18832 1114 18856 1116
rect 18912 1114 18918 1116
rect 18672 1062 18674 1114
rect 18854 1062 18856 1114
rect 18610 1060 18616 1062
rect 18672 1060 18696 1062
rect 18752 1060 18776 1062
rect 18832 1060 18856 1062
rect 18912 1060 18918 1062
rect 18610 1051 18918 1060
rect 19076 814 19104 2207
rect 18512 808 18564 814
rect 18512 750 18564 756
rect 19064 808 19116 814
rect 19064 750 19116 756
rect 18328 672 18380 678
rect 18328 614 18380 620
rect 17060 572 17368 581
rect 17060 570 17066 572
rect 17122 570 17146 572
rect 17202 570 17226 572
rect 17282 570 17306 572
rect 17362 570 17368 572
rect 17122 518 17124 570
rect 17304 518 17306 570
rect 17060 516 17066 518
rect 17122 516 17146 518
rect 17202 516 17226 518
rect 17282 516 17306 518
rect 17362 516 17368 518
rect 17060 507 17368 516
rect 16856 264 16908 270
rect 16856 206 16908 212
rect 13176 196 13228 202
rect 13176 138 13228 144
rect 16488 196 16540 202
rect 16488 138 16540 144
rect 18524 134 18552 750
rect 12072 128 12124 134
rect 12072 70 12124 76
rect 18512 128 18564 134
rect 18512 70 18564 76
<< via2 >>
rect 1122 10104 1178 10160
rect 662 9444 718 9480
rect 662 9424 664 9444
rect 664 9424 716 9444
rect 716 9424 718 9444
rect 570 8372 572 8392
rect 572 8372 624 8392
rect 624 8372 626 8392
rect 570 8336 626 8372
rect 662 7964 664 7984
rect 664 7964 716 7984
rect 716 7964 718 7984
rect 662 7928 718 7964
rect 1030 8336 1086 8392
rect 938 7420 940 7440
rect 940 7420 992 7440
rect 992 7420 994 7440
rect 938 7384 994 7420
rect 570 7248 626 7304
rect 2502 10684 2504 10704
rect 2504 10684 2556 10704
rect 2556 10684 2558 10704
rect 2502 10648 2558 10684
rect 1766 9444 1822 9480
rect 1766 9424 1768 9444
rect 1768 9424 1820 9444
rect 1820 9424 1822 9444
rect 846 6976 902 7032
rect 754 6860 810 6896
rect 754 6840 756 6860
rect 756 6840 808 6860
rect 808 6840 810 6860
rect 846 6196 848 6216
rect 848 6196 900 6216
rect 900 6196 902 6216
rect 846 6160 902 6196
rect 1214 7112 1270 7168
rect 1306 6704 1362 6760
rect 2318 7928 2374 7984
rect 2134 6296 2190 6352
rect 2502 7248 2558 7304
rect 2410 6996 2466 7032
rect 2410 6976 2412 6996
rect 2412 6976 2464 6996
rect 2464 6976 2466 6996
rect 3116 10906 3172 10908
rect 3196 10906 3252 10908
rect 3276 10906 3332 10908
rect 3356 10906 3412 10908
rect 3116 10854 3162 10906
rect 3162 10854 3172 10906
rect 3196 10854 3226 10906
rect 3226 10854 3238 10906
rect 3238 10854 3252 10906
rect 3276 10854 3290 10906
rect 3290 10854 3302 10906
rect 3302 10854 3332 10906
rect 3356 10854 3366 10906
rect 3366 10854 3412 10906
rect 3116 10852 3172 10854
rect 3196 10852 3252 10854
rect 3276 10852 3332 10854
rect 3356 10852 3412 10854
rect 4066 10512 4122 10568
rect 3146 9968 3202 10024
rect 3514 9968 3570 10024
rect 3116 9818 3172 9820
rect 3196 9818 3252 9820
rect 3276 9818 3332 9820
rect 3356 9818 3412 9820
rect 3116 9766 3162 9818
rect 3162 9766 3172 9818
rect 3196 9766 3226 9818
rect 3226 9766 3238 9818
rect 3238 9766 3252 9818
rect 3276 9766 3290 9818
rect 3290 9766 3302 9818
rect 3302 9766 3332 9818
rect 3356 9766 3366 9818
rect 3366 9766 3412 9818
rect 3116 9764 3172 9766
rect 3196 9764 3252 9766
rect 3276 9764 3332 9766
rect 3356 9764 3412 9766
rect 3116 8730 3172 8732
rect 3196 8730 3252 8732
rect 3276 8730 3332 8732
rect 3356 8730 3412 8732
rect 3116 8678 3162 8730
rect 3162 8678 3172 8730
rect 3196 8678 3226 8730
rect 3226 8678 3238 8730
rect 3238 8678 3252 8730
rect 3276 8678 3290 8730
rect 3290 8678 3302 8730
rect 3302 8678 3332 8730
rect 3356 8678 3366 8730
rect 3366 8678 3412 8730
rect 3116 8676 3172 8678
rect 3196 8676 3252 8678
rect 3276 8676 3332 8678
rect 3356 8676 3412 8678
rect 3116 7642 3172 7644
rect 3196 7642 3252 7644
rect 3276 7642 3332 7644
rect 3356 7642 3412 7644
rect 3116 7590 3162 7642
rect 3162 7590 3172 7642
rect 3196 7590 3226 7642
rect 3226 7590 3238 7642
rect 3238 7590 3252 7642
rect 3276 7590 3290 7642
rect 3290 7590 3302 7642
rect 3302 7590 3332 7642
rect 3356 7590 3366 7642
rect 3366 7590 3412 7642
rect 3116 7588 3172 7590
rect 3196 7588 3252 7590
rect 3276 7588 3332 7590
rect 3356 7588 3412 7590
rect 3054 7112 3110 7168
rect 2962 6976 3018 7032
rect 3422 6704 3478 6760
rect 3116 6554 3172 6556
rect 3196 6554 3252 6556
rect 3276 6554 3332 6556
rect 3356 6554 3412 6556
rect 3116 6502 3162 6554
rect 3162 6502 3172 6554
rect 3196 6502 3226 6554
rect 3226 6502 3238 6554
rect 3238 6502 3252 6554
rect 3276 6502 3290 6554
rect 3290 6502 3302 6554
rect 3302 6502 3332 6554
rect 3356 6502 3366 6554
rect 3366 6502 3412 6554
rect 3116 6500 3172 6502
rect 3196 6500 3252 6502
rect 3276 6500 3332 6502
rect 3356 6500 3412 6502
rect 3238 6332 3240 6352
rect 3240 6332 3292 6352
rect 3292 6332 3294 6352
rect 3238 6296 3294 6332
rect 4666 10362 4722 10364
rect 4746 10362 4802 10364
rect 4826 10362 4882 10364
rect 4906 10362 4962 10364
rect 4666 10310 4712 10362
rect 4712 10310 4722 10362
rect 4746 10310 4776 10362
rect 4776 10310 4788 10362
rect 4788 10310 4802 10362
rect 4826 10310 4840 10362
rect 4840 10310 4852 10362
rect 4852 10310 4882 10362
rect 4906 10310 4916 10362
rect 4916 10310 4962 10362
rect 4666 10308 4722 10310
rect 4746 10308 4802 10310
rect 4826 10308 4882 10310
rect 4906 10308 4962 10310
rect 6216 10906 6272 10908
rect 6296 10906 6352 10908
rect 6376 10906 6432 10908
rect 6456 10906 6512 10908
rect 6216 10854 6262 10906
rect 6262 10854 6272 10906
rect 6296 10854 6326 10906
rect 6326 10854 6338 10906
rect 6338 10854 6352 10906
rect 6376 10854 6390 10906
rect 6390 10854 6402 10906
rect 6402 10854 6432 10906
rect 6456 10854 6466 10906
rect 6466 10854 6512 10906
rect 6216 10852 6272 10854
rect 6296 10852 6352 10854
rect 6376 10852 6432 10854
rect 6456 10852 6512 10854
rect 5538 10512 5594 10568
rect 4434 10104 4490 10160
rect 4894 9968 4950 10024
rect 3790 7404 3846 7440
rect 3790 7384 3792 7404
rect 3792 7384 3844 7404
rect 3844 7384 3846 7404
rect 4250 7284 4252 7304
rect 4252 7284 4304 7304
rect 4304 7284 4306 7304
rect 3116 5466 3172 5468
rect 3196 5466 3252 5468
rect 3276 5466 3332 5468
rect 3356 5466 3412 5468
rect 3116 5414 3162 5466
rect 3162 5414 3172 5466
rect 3196 5414 3226 5466
rect 3226 5414 3238 5466
rect 3238 5414 3252 5466
rect 3276 5414 3290 5466
rect 3290 5414 3302 5466
rect 3302 5414 3332 5466
rect 3356 5414 3366 5466
rect 3366 5414 3412 5466
rect 3116 5412 3172 5414
rect 3196 5412 3252 5414
rect 3276 5412 3332 5414
rect 3356 5412 3412 5414
rect 4250 7248 4306 7284
rect 4158 6976 4214 7032
rect 4250 6160 4306 6216
rect 4666 9274 4722 9276
rect 4746 9274 4802 9276
rect 4826 9274 4882 9276
rect 4906 9274 4962 9276
rect 4666 9222 4712 9274
rect 4712 9222 4722 9274
rect 4746 9222 4776 9274
rect 4776 9222 4788 9274
rect 4788 9222 4802 9274
rect 4826 9222 4840 9274
rect 4840 9222 4852 9274
rect 4852 9222 4882 9274
rect 4906 9222 4916 9274
rect 4916 9222 4962 9274
rect 4666 9220 4722 9222
rect 4746 9220 4802 9222
rect 4826 9220 4882 9222
rect 4906 9220 4962 9222
rect 4986 8336 5042 8392
rect 4666 8186 4722 8188
rect 4746 8186 4802 8188
rect 4826 8186 4882 8188
rect 4906 8186 4962 8188
rect 4666 8134 4712 8186
rect 4712 8134 4722 8186
rect 4746 8134 4776 8186
rect 4776 8134 4788 8186
rect 4788 8134 4802 8186
rect 4826 8134 4840 8186
rect 4840 8134 4852 8186
rect 4852 8134 4882 8186
rect 4906 8134 4916 8186
rect 4916 8134 4962 8186
rect 4666 8132 4722 8134
rect 4746 8132 4802 8134
rect 4826 8132 4882 8134
rect 4906 8132 4962 8134
rect 4666 7098 4722 7100
rect 4746 7098 4802 7100
rect 4826 7098 4882 7100
rect 4906 7098 4962 7100
rect 4666 7046 4712 7098
rect 4712 7046 4722 7098
rect 4746 7046 4776 7098
rect 4776 7046 4788 7098
rect 4788 7046 4802 7098
rect 4826 7046 4840 7098
rect 4840 7046 4852 7098
rect 4852 7046 4882 7098
rect 4906 7046 4916 7098
rect 4916 7046 4962 7098
rect 4666 7044 4722 7046
rect 4746 7044 4802 7046
rect 4826 7044 4882 7046
rect 4906 7044 4962 7046
rect 6216 9818 6272 9820
rect 6296 9818 6352 9820
rect 6376 9818 6432 9820
rect 6456 9818 6512 9820
rect 6216 9766 6262 9818
rect 6262 9766 6272 9818
rect 6296 9766 6326 9818
rect 6326 9766 6338 9818
rect 6338 9766 6352 9818
rect 6376 9766 6390 9818
rect 6390 9766 6402 9818
rect 6402 9766 6432 9818
rect 6456 9766 6466 9818
rect 6466 9766 6512 9818
rect 6216 9764 6272 9766
rect 6296 9764 6352 9766
rect 6376 9764 6432 9766
rect 6456 9764 6512 9766
rect 6216 8730 6272 8732
rect 6296 8730 6352 8732
rect 6376 8730 6432 8732
rect 6456 8730 6512 8732
rect 6216 8678 6262 8730
rect 6262 8678 6272 8730
rect 6296 8678 6326 8730
rect 6326 8678 6338 8730
rect 6338 8678 6352 8730
rect 6376 8678 6390 8730
rect 6390 8678 6402 8730
rect 6402 8678 6432 8730
rect 6456 8678 6466 8730
rect 6466 8678 6512 8730
rect 6216 8676 6272 8678
rect 6296 8676 6352 8678
rect 6376 8676 6432 8678
rect 6456 8676 6512 8678
rect 5446 6840 5502 6896
rect 4666 6010 4722 6012
rect 4746 6010 4802 6012
rect 4826 6010 4882 6012
rect 4906 6010 4962 6012
rect 4666 5958 4712 6010
rect 4712 5958 4722 6010
rect 4746 5958 4776 6010
rect 4776 5958 4788 6010
rect 4788 5958 4802 6010
rect 4826 5958 4840 6010
rect 4840 5958 4852 6010
rect 4852 5958 4882 6010
rect 4906 5958 4916 6010
rect 4916 5958 4962 6010
rect 4666 5956 4722 5958
rect 4746 5956 4802 5958
rect 4826 5956 4882 5958
rect 4906 5956 4962 5958
rect 4666 4922 4722 4924
rect 4746 4922 4802 4924
rect 4826 4922 4882 4924
rect 4906 4922 4962 4924
rect 4666 4870 4712 4922
rect 4712 4870 4722 4922
rect 4746 4870 4776 4922
rect 4776 4870 4788 4922
rect 4788 4870 4802 4922
rect 4826 4870 4840 4922
rect 4840 4870 4852 4922
rect 4852 4870 4882 4922
rect 4906 4870 4916 4922
rect 4916 4870 4962 4922
rect 4666 4868 4722 4870
rect 4746 4868 4802 4870
rect 4826 4868 4882 4870
rect 4906 4868 4962 4870
rect 4342 4664 4398 4720
rect 3116 4378 3172 4380
rect 3196 4378 3252 4380
rect 3276 4378 3332 4380
rect 3356 4378 3412 4380
rect 3116 4326 3162 4378
rect 3162 4326 3172 4378
rect 3196 4326 3226 4378
rect 3226 4326 3238 4378
rect 3238 4326 3252 4378
rect 3276 4326 3290 4378
rect 3290 4326 3302 4378
rect 3302 4326 3332 4378
rect 3356 4326 3366 4378
rect 3366 4326 3412 4378
rect 3116 4324 3172 4326
rect 3196 4324 3252 4326
rect 3276 4324 3332 4326
rect 3356 4324 3412 4326
rect 6216 7642 6272 7644
rect 6296 7642 6352 7644
rect 6376 7642 6432 7644
rect 6456 7642 6512 7644
rect 6216 7590 6262 7642
rect 6262 7590 6272 7642
rect 6296 7590 6326 7642
rect 6326 7590 6338 7642
rect 6338 7590 6352 7642
rect 6376 7590 6390 7642
rect 6390 7590 6402 7642
rect 6402 7590 6432 7642
rect 6456 7590 6466 7642
rect 6466 7590 6512 7642
rect 6216 7588 6272 7590
rect 6296 7588 6352 7590
rect 6376 7588 6432 7590
rect 6456 7588 6512 7590
rect 6090 6840 6146 6896
rect 5446 5616 5502 5672
rect 6216 6554 6272 6556
rect 6296 6554 6352 6556
rect 6376 6554 6432 6556
rect 6456 6554 6512 6556
rect 6216 6502 6262 6554
rect 6262 6502 6272 6554
rect 6296 6502 6326 6554
rect 6326 6502 6338 6554
rect 6338 6502 6352 6554
rect 6376 6502 6390 6554
rect 6390 6502 6402 6554
rect 6402 6502 6432 6554
rect 6456 6502 6466 6554
rect 6466 6502 6512 6554
rect 6216 6500 6272 6502
rect 6296 6500 6352 6502
rect 6376 6500 6432 6502
rect 6456 6500 6512 6502
rect 5906 5752 5962 5808
rect 3116 3290 3172 3292
rect 3196 3290 3252 3292
rect 3276 3290 3332 3292
rect 3356 3290 3412 3292
rect 3116 3238 3162 3290
rect 3162 3238 3172 3290
rect 3196 3238 3226 3290
rect 3226 3238 3238 3290
rect 3238 3238 3252 3290
rect 3276 3238 3290 3290
rect 3290 3238 3302 3290
rect 3302 3238 3332 3290
rect 3356 3238 3366 3290
rect 3366 3238 3412 3290
rect 3116 3236 3172 3238
rect 3196 3236 3252 3238
rect 3276 3236 3332 3238
rect 3356 3236 3412 3238
rect 3116 2202 3172 2204
rect 3196 2202 3252 2204
rect 3276 2202 3332 2204
rect 3356 2202 3412 2204
rect 3116 2150 3162 2202
rect 3162 2150 3172 2202
rect 3196 2150 3226 2202
rect 3226 2150 3238 2202
rect 3238 2150 3252 2202
rect 3276 2150 3290 2202
rect 3290 2150 3302 2202
rect 3302 2150 3332 2202
rect 3356 2150 3366 2202
rect 3366 2150 3412 2202
rect 3116 2148 3172 2150
rect 3196 2148 3252 2150
rect 3276 2148 3332 2150
rect 3356 2148 3412 2150
rect 4666 3834 4722 3836
rect 4746 3834 4802 3836
rect 4826 3834 4882 3836
rect 4906 3834 4962 3836
rect 4666 3782 4712 3834
rect 4712 3782 4722 3834
rect 4746 3782 4776 3834
rect 4776 3782 4788 3834
rect 4788 3782 4802 3834
rect 4826 3782 4840 3834
rect 4840 3782 4852 3834
rect 4852 3782 4882 3834
rect 4906 3782 4916 3834
rect 4916 3782 4962 3834
rect 4666 3780 4722 3782
rect 4746 3780 4802 3782
rect 4826 3780 4882 3782
rect 4906 3780 4962 3782
rect 4802 3440 4858 3496
rect 6216 5466 6272 5468
rect 6296 5466 6352 5468
rect 6376 5466 6432 5468
rect 6456 5466 6512 5468
rect 6216 5414 6262 5466
rect 6262 5414 6272 5466
rect 6296 5414 6326 5466
rect 6326 5414 6338 5466
rect 6338 5414 6352 5466
rect 6376 5414 6390 5466
rect 6390 5414 6402 5466
rect 6402 5414 6432 5466
rect 6456 5414 6466 5466
rect 6466 5414 6512 5466
rect 6216 5412 6272 5414
rect 6296 5412 6352 5414
rect 6376 5412 6432 5414
rect 6456 5412 6512 5414
rect 5906 4800 5962 4856
rect 5630 3576 5686 3632
rect 6734 6704 6790 6760
rect 7194 6876 7196 6896
rect 7196 6876 7248 6896
rect 7248 6876 7250 6896
rect 7194 6840 7250 6876
rect 7766 10362 7822 10364
rect 7846 10362 7902 10364
rect 7926 10362 7982 10364
rect 8006 10362 8062 10364
rect 7766 10310 7812 10362
rect 7812 10310 7822 10362
rect 7846 10310 7876 10362
rect 7876 10310 7888 10362
rect 7888 10310 7902 10362
rect 7926 10310 7940 10362
rect 7940 10310 7952 10362
rect 7952 10310 7982 10362
rect 8006 10310 8016 10362
rect 8016 10310 8062 10362
rect 7766 10308 7822 10310
rect 7846 10308 7902 10310
rect 7926 10308 7982 10310
rect 8006 10308 8062 10310
rect 7766 9274 7822 9276
rect 7846 9274 7902 9276
rect 7926 9274 7982 9276
rect 8006 9274 8062 9276
rect 7766 9222 7812 9274
rect 7812 9222 7822 9274
rect 7846 9222 7876 9274
rect 7876 9222 7888 9274
rect 7888 9222 7902 9274
rect 7926 9222 7940 9274
rect 7940 9222 7952 9274
rect 7952 9222 7982 9274
rect 8006 9222 8016 9274
rect 8016 9222 8062 9274
rect 7766 9220 7822 9222
rect 7846 9220 7902 9222
rect 7926 9220 7982 9222
rect 8006 9220 8062 9222
rect 7766 8186 7822 8188
rect 7846 8186 7902 8188
rect 7926 8186 7982 8188
rect 8006 8186 8062 8188
rect 7766 8134 7812 8186
rect 7812 8134 7822 8186
rect 7846 8134 7876 8186
rect 7876 8134 7888 8186
rect 7888 8134 7902 8186
rect 7926 8134 7940 8186
rect 7940 8134 7952 8186
rect 7952 8134 7982 8186
rect 8006 8134 8016 8186
rect 8016 8134 8062 8186
rect 7766 8132 7822 8134
rect 7846 8132 7902 8134
rect 7926 8132 7982 8134
rect 8006 8132 8062 8134
rect 6734 4800 6790 4856
rect 6090 4684 6146 4720
rect 6090 4664 6092 4684
rect 6092 4664 6144 4684
rect 6144 4664 6146 4684
rect 6216 4378 6272 4380
rect 6296 4378 6352 4380
rect 6376 4378 6432 4380
rect 6456 4378 6512 4380
rect 6216 4326 6262 4378
rect 6262 4326 6272 4378
rect 6296 4326 6326 4378
rect 6326 4326 6338 4378
rect 6338 4326 6352 4378
rect 6376 4326 6390 4378
rect 6390 4326 6402 4378
rect 6402 4326 6432 4378
rect 6456 4326 6466 4378
rect 6466 4326 6512 4378
rect 6216 4324 6272 4326
rect 6296 4324 6352 4326
rect 6376 4324 6432 4326
rect 6456 4324 6512 4326
rect 6182 3984 6238 4040
rect 6642 4256 6698 4312
rect 5906 3712 5962 3768
rect 4666 2746 4722 2748
rect 4746 2746 4802 2748
rect 4826 2746 4882 2748
rect 4906 2746 4962 2748
rect 4666 2694 4712 2746
rect 4712 2694 4722 2746
rect 4746 2694 4776 2746
rect 4776 2694 4788 2746
rect 4788 2694 4802 2746
rect 4826 2694 4840 2746
rect 4840 2694 4852 2746
rect 4852 2694 4882 2746
rect 4906 2694 4916 2746
rect 4916 2694 4962 2746
rect 4666 2692 4722 2694
rect 4746 2692 4802 2694
rect 4826 2692 4882 2694
rect 4906 2692 4962 2694
rect 6216 3290 6272 3292
rect 6296 3290 6352 3292
rect 6376 3290 6432 3292
rect 6456 3290 6512 3292
rect 6216 3238 6262 3290
rect 6262 3238 6272 3290
rect 6296 3238 6326 3290
rect 6326 3238 6338 3290
rect 6338 3238 6352 3290
rect 6376 3238 6390 3290
rect 6390 3238 6402 3290
rect 6402 3238 6432 3290
rect 6456 3238 6466 3290
rect 6466 3238 6512 3290
rect 6216 3236 6272 3238
rect 6296 3236 6352 3238
rect 6376 3236 6432 3238
rect 6456 3236 6512 3238
rect 6182 3032 6238 3088
rect 5354 2488 5410 2544
rect 4666 1658 4722 1660
rect 4746 1658 4802 1660
rect 4826 1658 4882 1660
rect 4906 1658 4962 1660
rect 4666 1606 4712 1658
rect 4712 1606 4722 1658
rect 4746 1606 4776 1658
rect 4776 1606 4788 1658
rect 4788 1606 4802 1658
rect 4826 1606 4840 1658
rect 4840 1606 4852 1658
rect 4852 1606 4882 1658
rect 4906 1606 4916 1658
rect 4916 1606 4962 1658
rect 4666 1604 4722 1606
rect 4746 1604 4802 1606
rect 4826 1604 4882 1606
rect 4906 1604 4962 1606
rect 6216 2202 6272 2204
rect 6296 2202 6352 2204
rect 6376 2202 6432 2204
rect 6456 2202 6512 2204
rect 6216 2150 6262 2202
rect 6262 2150 6272 2202
rect 6296 2150 6326 2202
rect 6326 2150 6338 2202
rect 6338 2150 6352 2202
rect 6376 2150 6390 2202
rect 6390 2150 6402 2202
rect 6402 2150 6432 2202
rect 6456 2150 6466 2202
rect 6466 2150 6512 2202
rect 6216 2148 6272 2150
rect 6296 2148 6352 2150
rect 6376 2148 6432 2150
rect 6456 2148 6512 2150
rect 3116 1114 3172 1116
rect 3196 1114 3252 1116
rect 3276 1114 3332 1116
rect 3356 1114 3412 1116
rect 3116 1062 3162 1114
rect 3162 1062 3172 1114
rect 3196 1062 3226 1114
rect 3226 1062 3238 1114
rect 3238 1062 3252 1114
rect 3276 1062 3290 1114
rect 3290 1062 3302 1114
rect 3302 1062 3332 1114
rect 3356 1062 3366 1114
rect 3366 1062 3412 1114
rect 3116 1060 3172 1062
rect 3196 1060 3252 1062
rect 3276 1060 3332 1062
rect 3356 1060 3412 1062
rect 6216 1114 6272 1116
rect 6296 1114 6352 1116
rect 6376 1114 6432 1116
rect 6456 1114 6512 1116
rect 6216 1062 6262 1114
rect 6262 1062 6272 1114
rect 6296 1062 6326 1114
rect 6326 1062 6338 1114
rect 6338 1062 6352 1114
rect 6376 1062 6390 1114
rect 6390 1062 6402 1114
rect 6402 1062 6432 1114
rect 6456 1062 6466 1114
rect 6466 1062 6512 1114
rect 6216 1060 6272 1062
rect 6296 1060 6352 1062
rect 6376 1060 6432 1062
rect 6456 1060 6512 1062
rect 6826 3340 6828 3360
rect 6828 3340 6880 3360
rect 6880 3340 6882 3360
rect 6826 3304 6882 3340
rect 6734 2896 6790 2952
rect 7102 5752 7158 5808
rect 6826 2624 6882 2680
rect 7378 3712 7434 3768
rect 7378 3168 7434 3224
rect 7766 7098 7822 7100
rect 7846 7098 7902 7100
rect 7926 7098 7982 7100
rect 8006 7098 8062 7100
rect 7766 7046 7812 7098
rect 7812 7046 7822 7098
rect 7846 7046 7876 7098
rect 7876 7046 7888 7098
rect 7888 7046 7902 7098
rect 7926 7046 7940 7098
rect 7940 7046 7952 7098
rect 7952 7046 7982 7098
rect 8006 7046 8016 7098
rect 8016 7046 8062 7098
rect 7766 7044 7822 7046
rect 7846 7044 7902 7046
rect 7926 7044 7982 7046
rect 8006 7044 8062 7046
rect 7930 6704 7986 6760
rect 7766 6010 7822 6012
rect 7846 6010 7902 6012
rect 7926 6010 7982 6012
rect 8006 6010 8062 6012
rect 7766 5958 7812 6010
rect 7812 5958 7822 6010
rect 7846 5958 7876 6010
rect 7876 5958 7888 6010
rect 7888 5958 7902 6010
rect 7926 5958 7940 6010
rect 7940 5958 7952 6010
rect 7952 5958 7982 6010
rect 8006 5958 8016 6010
rect 8016 5958 8062 6010
rect 7766 5956 7822 5958
rect 7846 5956 7902 5958
rect 7926 5956 7982 5958
rect 8006 5956 8062 5958
rect 7930 5772 7986 5808
rect 7930 5752 7932 5772
rect 7932 5752 7984 5772
rect 7984 5752 7986 5772
rect 9316 10906 9372 10908
rect 9396 10906 9452 10908
rect 9476 10906 9532 10908
rect 9556 10906 9612 10908
rect 9316 10854 9362 10906
rect 9362 10854 9372 10906
rect 9396 10854 9426 10906
rect 9426 10854 9438 10906
rect 9438 10854 9452 10906
rect 9476 10854 9490 10906
rect 9490 10854 9502 10906
rect 9502 10854 9532 10906
rect 9556 10854 9566 10906
rect 9566 10854 9612 10906
rect 9316 10852 9372 10854
rect 9396 10852 9452 10854
rect 9476 10852 9532 10854
rect 9556 10852 9612 10854
rect 9310 10648 9366 10704
rect 7766 4922 7822 4924
rect 7846 4922 7902 4924
rect 7926 4922 7982 4924
rect 8006 4922 8062 4924
rect 7766 4870 7812 4922
rect 7812 4870 7822 4922
rect 7846 4870 7876 4922
rect 7876 4870 7888 4922
rect 7888 4870 7902 4922
rect 7926 4870 7940 4922
rect 7940 4870 7952 4922
rect 7952 4870 7982 4922
rect 8006 4870 8016 4922
rect 8016 4870 8062 4922
rect 7766 4868 7822 4870
rect 7846 4868 7902 4870
rect 7926 4868 7982 4870
rect 8006 4868 8062 4870
rect 8022 4020 8024 4040
rect 8024 4020 8076 4040
rect 8076 4020 8078 4040
rect 8022 3984 8078 4020
rect 8206 4256 8262 4312
rect 7766 3834 7822 3836
rect 7846 3834 7902 3836
rect 7926 3834 7982 3836
rect 8006 3834 8062 3836
rect 7766 3782 7812 3834
rect 7812 3782 7822 3834
rect 7846 3782 7876 3834
rect 7876 3782 7888 3834
rect 7888 3782 7902 3834
rect 7926 3782 7940 3834
rect 7940 3782 7952 3834
rect 7952 3782 7982 3834
rect 8006 3782 8016 3834
rect 8016 3782 8062 3834
rect 7766 3780 7822 3782
rect 7846 3780 7902 3782
rect 7926 3780 7982 3782
rect 8006 3780 8062 3782
rect 9586 9968 9642 10024
rect 9316 9818 9372 9820
rect 9396 9818 9452 9820
rect 9476 9818 9532 9820
rect 9556 9818 9612 9820
rect 9316 9766 9362 9818
rect 9362 9766 9372 9818
rect 9396 9766 9426 9818
rect 9426 9766 9438 9818
rect 9438 9766 9452 9818
rect 9476 9766 9490 9818
rect 9490 9766 9502 9818
rect 9502 9766 9532 9818
rect 9556 9766 9566 9818
rect 9566 9766 9612 9818
rect 9316 9764 9372 9766
rect 9396 9764 9452 9766
rect 9476 9764 9532 9766
rect 9556 9764 9612 9766
rect 9316 8730 9372 8732
rect 9396 8730 9452 8732
rect 9476 8730 9532 8732
rect 9556 8730 9612 8732
rect 9316 8678 9362 8730
rect 9362 8678 9372 8730
rect 9396 8678 9426 8730
rect 9426 8678 9438 8730
rect 9438 8678 9452 8730
rect 9476 8678 9490 8730
rect 9490 8678 9502 8730
rect 9502 8678 9532 8730
rect 9556 8678 9566 8730
rect 9566 8678 9612 8730
rect 9316 8676 9372 8678
rect 9396 8676 9452 8678
rect 9476 8676 9532 8678
rect 9556 8676 9612 8678
rect 9316 7642 9372 7644
rect 9396 7642 9452 7644
rect 9476 7642 9532 7644
rect 9556 7642 9612 7644
rect 9316 7590 9362 7642
rect 9362 7590 9372 7642
rect 9396 7590 9426 7642
rect 9426 7590 9438 7642
rect 9438 7590 9452 7642
rect 9476 7590 9490 7642
rect 9490 7590 9502 7642
rect 9502 7590 9532 7642
rect 9556 7590 9566 7642
rect 9566 7590 9612 7642
rect 9316 7588 9372 7590
rect 9396 7588 9452 7590
rect 9476 7588 9532 7590
rect 9556 7588 9612 7590
rect 9316 6554 9372 6556
rect 9396 6554 9452 6556
rect 9476 6554 9532 6556
rect 9556 6554 9612 6556
rect 9316 6502 9362 6554
rect 9362 6502 9372 6554
rect 9396 6502 9426 6554
rect 9426 6502 9438 6554
rect 9438 6502 9452 6554
rect 9476 6502 9490 6554
rect 9490 6502 9502 6554
rect 9502 6502 9532 6554
rect 9556 6502 9566 6554
rect 9566 6502 9612 6554
rect 9316 6500 9372 6502
rect 9396 6500 9452 6502
rect 9476 6500 9532 6502
rect 9556 6500 9612 6502
rect 7838 3576 7894 3632
rect 8114 3576 8170 3632
rect 7930 3304 7986 3360
rect 7286 2624 7342 2680
rect 8114 3168 8170 3224
rect 8114 3052 8170 3088
rect 8114 3032 8116 3052
rect 8116 3032 8168 3052
rect 8168 3032 8170 3052
rect 7766 2746 7822 2748
rect 7846 2746 7902 2748
rect 7926 2746 7982 2748
rect 8006 2746 8062 2748
rect 7766 2694 7812 2746
rect 7812 2694 7822 2746
rect 7846 2694 7876 2746
rect 7876 2694 7888 2746
rect 7888 2694 7902 2746
rect 7926 2694 7940 2746
rect 7940 2694 7952 2746
rect 7952 2694 7982 2746
rect 8006 2694 8016 2746
rect 8016 2694 8062 2746
rect 7766 2692 7822 2694
rect 7846 2692 7902 2694
rect 7926 2692 7982 2694
rect 8006 2692 8062 2694
rect 8390 3032 8446 3088
rect 8114 2488 8170 2544
rect 7766 1658 7822 1660
rect 7846 1658 7902 1660
rect 7926 1658 7982 1660
rect 8006 1658 8062 1660
rect 7766 1606 7812 1658
rect 7812 1606 7822 1658
rect 7846 1606 7876 1658
rect 7876 1606 7888 1658
rect 7888 1606 7902 1658
rect 7926 1606 7940 1658
rect 7940 1606 7952 1658
rect 7952 1606 7982 1658
rect 8006 1606 8016 1658
rect 8016 1606 8062 1658
rect 7766 1604 7822 1606
rect 7846 1604 7902 1606
rect 7926 1604 7982 1606
rect 8006 1604 8062 1606
rect 8482 2624 8538 2680
rect 8942 3440 8998 3496
rect 8850 2916 8906 2952
rect 8850 2896 8852 2916
rect 8852 2896 8904 2916
rect 8904 2896 8906 2916
rect 8942 2624 8998 2680
rect 9402 5616 9458 5672
rect 9316 5466 9372 5468
rect 9396 5466 9452 5468
rect 9476 5466 9532 5468
rect 9556 5466 9612 5468
rect 9316 5414 9362 5466
rect 9362 5414 9372 5466
rect 9396 5414 9426 5466
rect 9426 5414 9438 5466
rect 9438 5414 9452 5466
rect 9476 5414 9490 5466
rect 9490 5414 9502 5466
rect 9502 5414 9532 5466
rect 9556 5414 9566 5466
rect 9566 5414 9612 5466
rect 9316 5412 9372 5414
rect 9396 5412 9452 5414
rect 9476 5412 9532 5414
rect 9556 5412 9612 5414
rect 9316 4378 9372 4380
rect 9396 4378 9452 4380
rect 9476 4378 9532 4380
rect 9556 4378 9612 4380
rect 9316 4326 9362 4378
rect 9362 4326 9372 4378
rect 9396 4326 9426 4378
rect 9426 4326 9438 4378
rect 9438 4326 9452 4378
rect 9476 4326 9490 4378
rect 9490 4326 9502 4378
rect 9502 4326 9532 4378
rect 9556 4326 9566 4378
rect 9566 4326 9612 4378
rect 9316 4324 9372 4326
rect 9396 4324 9452 4326
rect 9476 4324 9532 4326
rect 9556 4324 9612 4326
rect 10138 10512 10194 10568
rect 10138 10104 10194 10160
rect 10414 9968 10470 10024
rect 10866 10362 10922 10364
rect 10946 10362 11002 10364
rect 11026 10362 11082 10364
rect 11106 10362 11162 10364
rect 10866 10310 10912 10362
rect 10912 10310 10922 10362
rect 10946 10310 10976 10362
rect 10976 10310 10988 10362
rect 10988 10310 11002 10362
rect 11026 10310 11040 10362
rect 11040 10310 11052 10362
rect 11052 10310 11082 10362
rect 11106 10310 11116 10362
rect 11116 10310 11162 10362
rect 10866 10308 10922 10310
rect 10946 10308 11002 10310
rect 11026 10308 11082 10310
rect 11106 10308 11162 10310
rect 10866 9274 10922 9276
rect 10946 9274 11002 9276
rect 11026 9274 11082 9276
rect 11106 9274 11162 9276
rect 10866 9222 10912 9274
rect 10912 9222 10922 9274
rect 10946 9222 10976 9274
rect 10976 9222 10988 9274
rect 10988 9222 11002 9274
rect 11026 9222 11040 9274
rect 11040 9222 11052 9274
rect 11052 9222 11082 9274
rect 11106 9222 11116 9274
rect 11116 9222 11162 9274
rect 10866 9220 10922 9222
rect 10946 9220 11002 9222
rect 11026 9220 11082 9222
rect 11106 9220 11162 9222
rect 10782 8356 10838 8392
rect 10782 8336 10784 8356
rect 10784 8336 10836 8356
rect 10836 8336 10838 8356
rect 10866 8186 10922 8188
rect 10946 8186 11002 8188
rect 11026 8186 11082 8188
rect 11106 8186 11162 8188
rect 10866 8134 10912 8186
rect 10912 8134 10922 8186
rect 10946 8134 10976 8186
rect 10976 8134 10988 8186
rect 10988 8134 11002 8186
rect 11026 8134 11040 8186
rect 11040 8134 11052 8186
rect 11052 8134 11082 8186
rect 11106 8134 11116 8186
rect 11116 8134 11162 8186
rect 10866 8132 10922 8134
rect 10946 8132 11002 8134
rect 11026 8132 11082 8134
rect 11106 8132 11162 8134
rect 12416 10906 12472 10908
rect 12496 10906 12552 10908
rect 12576 10906 12632 10908
rect 12656 10906 12712 10908
rect 12416 10854 12462 10906
rect 12462 10854 12472 10906
rect 12496 10854 12526 10906
rect 12526 10854 12538 10906
rect 12538 10854 12552 10906
rect 12576 10854 12590 10906
rect 12590 10854 12602 10906
rect 12602 10854 12632 10906
rect 12656 10854 12666 10906
rect 12666 10854 12712 10906
rect 12416 10852 12472 10854
rect 12496 10852 12552 10854
rect 12576 10852 12632 10854
rect 12656 10852 12712 10854
rect 11978 10104 12034 10160
rect 11702 7964 11704 7984
rect 11704 7964 11756 7984
rect 11756 7964 11758 7984
rect 11702 7928 11758 7964
rect 12416 9818 12472 9820
rect 12496 9818 12552 9820
rect 12576 9818 12632 9820
rect 12656 9818 12712 9820
rect 12416 9766 12462 9818
rect 12462 9766 12472 9818
rect 12496 9766 12526 9818
rect 12526 9766 12538 9818
rect 12538 9766 12552 9818
rect 12576 9766 12590 9818
rect 12590 9766 12602 9818
rect 12602 9766 12632 9818
rect 12656 9766 12666 9818
rect 12666 9766 12712 9818
rect 12416 9764 12472 9766
rect 12496 9764 12552 9766
rect 12576 9764 12632 9766
rect 12656 9764 12712 9766
rect 12416 8730 12472 8732
rect 12496 8730 12552 8732
rect 12576 8730 12632 8732
rect 12656 8730 12712 8732
rect 12416 8678 12462 8730
rect 12462 8678 12472 8730
rect 12496 8678 12526 8730
rect 12526 8678 12538 8730
rect 12538 8678 12552 8730
rect 12576 8678 12590 8730
rect 12590 8678 12602 8730
rect 12602 8678 12632 8730
rect 12656 8678 12666 8730
rect 12666 8678 12712 8730
rect 12416 8676 12472 8678
rect 12496 8676 12552 8678
rect 12576 8676 12632 8678
rect 12656 8676 12712 8678
rect 12162 7928 12218 7984
rect 10414 7284 10416 7304
rect 10416 7284 10468 7304
rect 10468 7284 10470 7304
rect 10414 7248 10470 7284
rect 10866 7098 10922 7100
rect 10946 7098 11002 7100
rect 11026 7098 11082 7100
rect 11106 7098 11162 7100
rect 10866 7046 10912 7098
rect 10912 7046 10922 7098
rect 10946 7046 10976 7098
rect 10976 7046 10988 7098
rect 10988 7046 11002 7098
rect 11026 7046 11040 7098
rect 11040 7046 11052 7098
rect 11052 7046 11082 7098
rect 11106 7046 11116 7098
rect 11116 7046 11162 7098
rect 10866 7044 10922 7046
rect 10946 7044 11002 7046
rect 11026 7044 11082 7046
rect 11106 7044 11162 7046
rect 10046 6840 10102 6896
rect 9316 3290 9372 3292
rect 9396 3290 9452 3292
rect 9476 3290 9532 3292
rect 9556 3290 9612 3292
rect 9316 3238 9362 3290
rect 9362 3238 9372 3290
rect 9396 3238 9426 3290
rect 9426 3238 9438 3290
rect 9438 3238 9452 3290
rect 9476 3238 9490 3290
rect 9490 3238 9502 3290
rect 9502 3238 9532 3290
rect 9556 3238 9566 3290
rect 9566 3238 9612 3290
rect 9316 3236 9372 3238
rect 9396 3236 9452 3238
rect 9476 3236 9532 3238
rect 9556 3236 9612 3238
rect 8850 1944 8906 2000
rect 12346 8372 12348 8392
rect 12348 8372 12400 8392
rect 12400 8372 12402 8392
rect 12346 8336 12402 8372
rect 12416 7642 12472 7644
rect 12496 7642 12552 7644
rect 12576 7642 12632 7644
rect 12656 7642 12712 7644
rect 12416 7590 12462 7642
rect 12462 7590 12472 7642
rect 12496 7590 12526 7642
rect 12526 7590 12538 7642
rect 12538 7590 12552 7642
rect 12576 7590 12590 7642
rect 12590 7590 12602 7642
rect 12602 7590 12632 7642
rect 12656 7590 12666 7642
rect 12666 7590 12712 7642
rect 12416 7588 12472 7590
rect 12496 7588 12552 7590
rect 12576 7588 12632 7590
rect 12656 7588 12712 7590
rect 13966 10362 14022 10364
rect 14046 10362 14102 10364
rect 14126 10362 14182 10364
rect 14206 10362 14262 10364
rect 13966 10310 14012 10362
rect 14012 10310 14022 10362
rect 14046 10310 14076 10362
rect 14076 10310 14088 10362
rect 14088 10310 14102 10362
rect 14126 10310 14140 10362
rect 14140 10310 14152 10362
rect 14152 10310 14182 10362
rect 14206 10310 14216 10362
rect 14216 10310 14262 10362
rect 13966 10308 14022 10310
rect 14046 10308 14102 10310
rect 14126 10308 14182 10310
rect 14206 10308 14262 10310
rect 13966 9274 14022 9276
rect 14046 9274 14102 9276
rect 14126 9274 14182 9276
rect 14206 9274 14262 9276
rect 13966 9222 14012 9274
rect 14012 9222 14022 9274
rect 14046 9222 14076 9274
rect 14076 9222 14088 9274
rect 14088 9222 14102 9274
rect 14126 9222 14140 9274
rect 14140 9222 14152 9274
rect 14152 9222 14182 9274
rect 14206 9222 14216 9274
rect 14216 9222 14262 9274
rect 13966 9220 14022 9222
rect 14046 9220 14102 9222
rect 14126 9220 14182 9222
rect 14206 9220 14262 9222
rect 11978 6160 12034 6216
rect 12416 6554 12472 6556
rect 12496 6554 12552 6556
rect 12576 6554 12632 6556
rect 12656 6554 12712 6556
rect 12416 6502 12462 6554
rect 12462 6502 12472 6554
rect 12496 6502 12526 6554
rect 12526 6502 12538 6554
rect 12538 6502 12552 6554
rect 12576 6502 12590 6554
rect 12590 6502 12602 6554
rect 12602 6502 12632 6554
rect 12656 6502 12666 6554
rect 12666 6502 12712 6554
rect 12416 6500 12472 6502
rect 12496 6500 12552 6502
rect 12576 6500 12632 6502
rect 12656 6500 12712 6502
rect 10866 6010 10922 6012
rect 10946 6010 11002 6012
rect 11026 6010 11082 6012
rect 11106 6010 11162 6012
rect 10866 5958 10912 6010
rect 10912 5958 10922 6010
rect 10946 5958 10976 6010
rect 10976 5958 10988 6010
rect 10988 5958 11002 6010
rect 11026 5958 11040 6010
rect 11040 5958 11052 6010
rect 11052 5958 11082 6010
rect 11106 5958 11116 6010
rect 11116 5958 11162 6010
rect 10866 5956 10922 5958
rect 10946 5956 11002 5958
rect 11026 5956 11082 5958
rect 11106 5956 11162 5958
rect 9316 2202 9372 2204
rect 9396 2202 9452 2204
rect 9476 2202 9532 2204
rect 9556 2202 9612 2204
rect 9316 2150 9362 2202
rect 9362 2150 9372 2202
rect 9396 2150 9426 2202
rect 9426 2150 9438 2202
rect 9438 2150 9452 2202
rect 9476 2150 9490 2202
rect 9490 2150 9502 2202
rect 9502 2150 9532 2202
rect 9556 2150 9566 2202
rect 9566 2150 9612 2202
rect 9316 2148 9372 2150
rect 9396 2148 9452 2150
rect 9476 2148 9532 2150
rect 9556 2148 9612 2150
rect 9586 1980 9588 2000
rect 9588 1980 9640 2000
rect 9640 1980 9642 2000
rect 9586 1944 9642 1980
rect 10866 4922 10922 4924
rect 10946 4922 11002 4924
rect 11026 4922 11082 4924
rect 11106 4922 11162 4924
rect 10866 4870 10912 4922
rect 10912 4870 10922 4922
rect 10946 4870 10976 4922
rect 10976 4870 10988 4922
rect 10988 4870 11002 4922
rect 11026 4870 11040 4922
rect 11040 4870 11052 4922
rect 11052 4870 11082 4922
rect 11106 4870 11116 4922
rect 11116 4870 11162 4922
rect 10866 4868 10922 4870
rect 10946 4868 11002 4870
rect 11026 4868 11082 4870
rect 11106 4868 11162 4870
rect 11334 4528 11390 4584
rect 9316 1114 9372 1116
rect 9396 1114 9452 1116
rect 9476 1114 9532 1116
rect 9556 1114 9612 1116
rect 9316 1062 9362 1114
rect 9362 1062 9372 1114
rect 9396 1062 9426 1114
rect 9426 1062 9438 1114
rect 9438 1062 9452 1114
rect 9476 1062 9490 1114
rect 9490 1062 9502 1114
rect 9502 1062 9532 1114
rect 9556 1062 9566 1114
rect 9566 1062 9612 1114
rect 9316 1060 9372 1062
rect 9396 1060 9452 1062
rect 9476 1060 9532 1062
rect 9556 1060 9612 1062
rect 10866 3834 10922 3836
rect 10946 3834 11002 3836
rect 11026 3834 11082 3836
rect 11106 3834 11162 3836
rect 10866 3782 10912 3834
rect 10912 3782 10922 3834
rect 10946 3782 10976 3834
rect 10976 3782 10988 3834
rect 10988 3782 11002 3834
rect 11026 3782 11040 3834
rect 11040 3782 11052 3834
rect 11052 3782 11082 3834
rect 11106 3782 11116 3834
rect 11116 3782 11162 3834
rect 10866 3780 10922 3782
rect 10946 3780 11002 3782
rect 11026 3780 11082 3782
rect 11106 3780 11162 3782
rect 13966 8186 14022 8188
rect 14046 8186 14102 8188
rect 14126 8186 14182 8188
rect 14206 8186 14262 8188
rect 13966 8134 14012 8186
rect 14012 8134 14022 8186
rect 14046 8134 14076 8186
rect 14076 8134 14088 8186
rect 14088 8134 14102 8186
rect 14126 8134 14140 8186
rect 14140 8134 14152 8186
rect 14152 8134 14182 8186
rect 14206 8134 14216 8186
rect 14216 8134 14262 8186
rect 13966 8132 14022 8134
rect 14046 8132 14102 8134
rect 14126 8132 14182 8134
rect 14206 8132 14262 8134
rect 13966 7098 14022 7100
rect 14046 7098 14102 7100
rect 14126 7098 14182 7100
rect 14206 7098 14262 7100
rect 13966 7046 14012 7098
rect 14012 7046 14022 7098
rect 14046 7046 14076 7098
rect 14076 7046 14088 7098
rect 14088 7046 14102 7098
rect 14126 7046 14140 7098
rect 14140 7046 14152 7098
rect 14152 7046 14182 7098
rect 14206 7046 14216 7098
rect 14216 7046 14262 7098
rect 13966 7044 14022 7046
rect 14046 7044 14102 7046
rect 14126 7044 14182 7046
rect 14206 7044 14262 7046
rect 12416 5466 12472 5468
rect 12496 5466 12552 5468
rect 12576 5466 12632 5468
rect 12656 5466 12712 5468
rect 12416 5414 12462 5466
rect 12462 5414 12472 5466
rect 12496 5414 12526 5466
rect 12526 5414 12538 5466
rect 12538 5414 12552 5466
rect 12576 5414 12590 5466
rect 12590 5414 12602 5466
rect 12602 5414 12632 5466
rect 12656 5414 12666 5466
rect 12666 5414 12712 5466
rect 12416 5412 12472 5414
rect 12496 5412 12552 5414
rect 12576 5412 12632 5414
rect 12656 5412 12712 5414
rect 11886 3576 11942 3632
rect 11242 3032 11298 3088
rect 10866 2746 10922 2748
rect 10946 2746 11002 2748
rect 11026 2746 11082 2748
rect 11106 2746 11162 2748
rect 10866 2694 10912 2746
rect 10912 2694 10922 2746
rect 10946 2694 10976 2746
rect 10976 2694 10988 2746
rect 10988 2694 11002 2746
rect 11026 2694 11040 2746
rect 11040 2694 11052 2746
rect 11052 2694 11082 2746
rect 11106 2694 11116 2746
rect 11116 2694 11162 2746
rect 10866 2692 10922 2694
rect 10946 2692 11002 2694
rect 11026 2692 11082 2694
rect 11106 2692 11162 2694
rect 11242 2488 11298 2544
rect 10866 1658 10922 1660
rect 10946 1658 11002 1660
rect 11026 1658 11082 1660
rect 11106 1658 11162 1660
rect 10866 1606 10912 1658
rect 10912 1606 10922 1658
rect 10946 1606 10976 1658
rect 10976 1606 10988 1658
rect 10988 1606 11002 1658
rect 11026 1606 11040 1658
rect 11040 1606 11052 1658
rect 11052 1606 11082 1658
rect 11106 1606 11116 1658
rect 11116 1606 11162 1658
rect 10866 1604 10922 1606
rect 10946 1604 11002 1606
rect 11026 1604 11082 1606
rect 11106 1604 11162 1606
rect 12622 4528 12678 4584
rect 12416 4378 12472 4380
rect 12496 4378 12552 4380
rect 12576 4378 12632 4380
rect 12656 4378 12712 4380
rect 12416 4326 12462 4378
rect 12462 4326 12472 4378
rect 12496 4326 12526 4378
rect 12526 4326 12538 4378
rect 12538 4326 12552 4378
rect 12576 4326 12590 4378
rect 12590 4326 12602 4378
rect 12602 4326 12632 4378
rect 12656 4326 12666 4378
rect 12666 4326 12712 4378
rect 12416 4324 12472 4326
rect 12496 4324 12552 4326
rect 12576 4324 12632 4326
rect 12656 4324 12712 4326
rect 12806 3712 12862 3768
rect 12416 3290 12472 3292
rect 12496 3290 12552 3292
rect 12576 3290 12632 3292
rect 12656 3290 12712 3292
rect 12416 3238 12462 3290
rect 12462 3238 12472 3290
rect 12496 3238 12526 3290
rect 12526 3238 12538 3290
rect 12538 3238 12552 3290
rect 12576 3238 12590 3290
rect 12590 3238 12602 3290
rect 12602 3238 12632 3290
rect 12656 3238 12666 3290
rect 12666 3238 12712 3290
rect 12416 3236 12472 3238
rect 12496 3236 12552 3238
rect 12576 3236 12632 3238
rect 12656 3236 12712 3238
rect 12714 2932 12716 2952
rect 12716 2932 12768 2952
rect 12768 2932 12770 2952
rect 12714 2896 12770 2932
rect 13174 3440 13230 3496
rect 13542 6160 13598 6216
rect 13542 5208 13598 5264
rect 12416 2202 12472 2204
rect 12496 2202 12552 2204
rect 12576 2202 12632 2204
rect 12656 2202 12712 2204
rect 12416 2150 12462 2202
rect 12462 2150 12472 2202
rect 12496 2150 12526 2202
rect 12526 2150 12538 2202
rect 12538 2150 12552 2202
rect 12576 2150 12590 2202
rect 12590 2150 12602 2202
rect 12602 2150 12632 2202
rect 12656 2150 12666 2202
rect 12666 2150 12712 2202
rect 12416 2148 12472 2150
rect 12496 2148 12552 2150
rect 12576 2148 12632 2150
rect 12656 2148 12712 2150
rect 12070 1808 12126 1864
rect 13266 2916 13322 2952
rect 13266 2896 13268 2916
rect 13268 2896 13320 2916
rect 13320 2896 13322 2916
rect 13966 6010 14022 6012
rect 14046 6010 14102 6012
rect 14126 6010 14182 6012
rect 14206 6010 14262 6012
rect 13966 5958 14012 6010
rect 14012 5958 14022 6010
rect 14046 5958 14076 6010
rect 14076 5958 14088 6010
rect 14088 5958 14102 6010
rect 14126 5958 14140 6010
rect 14140 5958 14152 6010
rect 14152 5958 14182 6010
rect 14206 5958 14216 6010
rect 14216 5958 14262 6010
rect 13966 5956 14022 5958
rect 14046 5956 14102 5958
rect 14126 5956 14182 5958
rect 14206 5956 14262 5958
rect 15198 10512 15254 10568
rect 14646 6860 14702 6896
rect 14646 6840 14648 6860
rect 14648 6840 14700 6860
rect 14700 6840 14702 6860
rect 13966 4922 14022 4924
rect 14046 4922 14102 4924
rect 14126 4922 14182 4924
rect 14206 4922 14262 4924
rect 13966 4870 14012 4922
rect 14012 4870 14022 4922
rect 14046 4870 14076 4922
rect 14076 4870 14088 4922
rect 14088 4870 14102 4922
rect 14126 4870 14140 4922
rect 14140 4870 14152 4922
rect 14152 4870 14182 4922
rect 14206 4870 14216 4922
rect 14216 4870 14262 4922
rect 13966 4868 14022 4870
rect 14046 4868 14102 4870
rect 14126 4868 14182 4870
rect 14206 4868 14262 4870
rect 15198 9968 15254 10024
rect 14462 4528 14518 4584
rect 13726 3712 13782 3768
rect 13966 3834 14022 3836
rect 14046 3834 14102 3836
rect 14126 3834 14182 3836
rect 14206 3834 14262 3836
rect 13966 3782 14012 3834
rect 14012 3782 14022 3834
rect 14046 3782 14076 3834
rect 14076 3782 14088 3834
rect 14088 3782 14102 3834
rect 14126 3782 14140 3834
rect 14140 3782 14152 3834
rect 14152 3782 14182 3834
rect 14206 3782 14216 3834
rect 14216 3782 14262 3834
rect 13966 3780 14022 3782
rect 14046 3780 14102 3782
rect 14126 3780 14182 3782
rect 14206 3780 14262 3782
rect 13450 3188 13506 3224
rect 13450 3168 13452 3188
rect 13452 3168 13504 3188
rect 13504 3168 13506 3188
rect 13358 1944 13414 2000
rect 4666 570 4722 572
rect 4746 570 4802 572
rect 4826 570 4882 572
rect 4906 570 4962 572
rect 4666 518 4712 570
rect 4712 518 4722 570
rect 4746 518 4776 570
rect 4776 518 4788 570
rect 4788 518 4802 570
rect 4826 518 4840 570
rect 4840 518 4852 570
rect 4852 518 4882 570
rect 4906 518 4916 570
rect 4916 518 4962 570
rect 4666 516 4722 518
rect 4746 516 4802 518
rect 4826 516 4882 518
rect 4906 516 4962 518
rect 7766 570 7822 572
rect 7846 570 7902 572
rect 7926 570 7982 572
rect 8006 570 8062 572
rect 7766 518 7812 570
rect 7812 518 7822 570
rect 7846 518 7876 570
rect 7876 518 7888 570
rect 7888 518 7902 570
rect 7926 518 7940 570
rect 7940 518 7952 570
rect 7952 518 7982 570
rect 8006 518 8016 570
rect 8016 518 8062 570
rect 7766 516 7822 518
rect 7846 516 7902 518
rect 7926 516 7982 518
rect 8006 516 8062 518
rect 10866 570 10922 572
rect 10946 570 11002 572
rect 11026 570 11082 572
rect 11106 570 11162 572
rect 10866 518 10912 570
rect 10912 518 10922 570
rect 10946 518 10976 570
rect 10976 518 10988 570
rect 10988 518 11002 570
rect 11026 518 11040 570
rect 11040 518 11052 570
rect 11052 518 11082 570
rect 11106 518 11116 570
rect 11116 518 11162 570
rect 10866 516 10922 518
rect 10946 516 11002 518
rect 11026 516 11082 518
rect 11106 516 11162 518
rect 12416 1114 12472 1116
rect 12496 1114 12552 1116
rect 12576 1114 12632 1116
rect 12656 1114 12712 1116
rect 12416 1062 12462 1114
rect 12462 1062 12472 1114
rect 12496 1062 12526 1114
rect 12526 1062 12538 1114
rect 12538 1062 12552 1114
rect 12576 1062 12590 1114
rect 12590 1062 12602 1114
rect 12602 1062 12632 1114
rect 12656 1062 12666 1114
rect 12666 1062 12712 1114
rect 12416 1060 12472 1062
rect 12496 1060 12552 1062
rect 12576 1060 12632 1062
rect 12656 1060 12712 1062
rect 12806 756 12808 776
rect 12808 756 12860 776
rect 12860 756 12862 776
rect 12806 720 12862 756
rect 13818 3304 13874 3360
rect 14186 3168 14242 3224
rect 13966 2746 14022 2748
rect 14046 2746 14102 2748
rect 14126 2746 14182 2748
rect 14206 2746 14262 2748
rect 13966 2694 14012 2746
rect 14012 2694 14022 2746
rect 14046 2694 14076 2746
rect 14076 2694 14088 2746
rect 14088 2694 14102 2746
rect 14126 2694 14140 2746
rect 14140 2694 14152 2746
rect 14152 2694 14182 2746
rect 14206 2694 14216 2746
rect 14216 2694 14262 2746
rect 13966 2692 14022 2694
rect 14046 2692 14102 2694
rect 14126 2692 14182 2694
rect 14206 2692 14262 2694
rect 13910 2524 13912 2544
rect 13912 2524 13964 2544
rect 13964 2524 13966 2544
rect 13910 2488 13966 2524
rect 14186 2508 14242 2544
rect 14186 2488 14188 2508
rect 14188 2488 14240 2508
rect 14240 2488 14242 2508
rect 13266 992 13322 1048
rect 13966 1658 14022 1660
rect 14046 1658 14102 1660
rect 14126 1658 14182 1660
rect 14206 1658 14262 1660
rect 13966 1606 14012 1658
rect 14012 1606 14022 1658
rect 14046 1606 14076 1658
rect 14076 1606 14088 1658
rect 14088 1606 14102 1658
rect 14126 1606 14140 1658
rect 14140 1606 14152 1658
rect 14152 1606 14182 1658
rect 14206 1606 14216 1658
rect 14216 1606 14262 1658
rect 13966 1604 14022 1606
rect 14046 1604 14102 1606
rect 14126 1604 14182 1606
rect 14206 1604 14262 1606
rect 13266 876 13322 912
rect 13266 856 13268 876
rect 13268 856 13320 876
rect 13320 856 13322 876
rect 14094 1400 14150 1456
rect 14278 992 14334 1048
rect 14922 6740 14924 6760
rect 14924 6740 14976 6760
rect 14976 6740 14978 6760
rect 14922 6704 14978 6740
rect 15106 6160 15162 6216
rect 14922 5208 14978 5264
rect 14738 3304 14794 3360
rect 14738 1944 14794 2000
rect 15106 4800 15162 4856
rect 15014 4004 15070 4040
rect 15014 3984 15016 4004
rect 15016 3984 15068 4004
rect 15068 3984 15070 4004
rect 15516 10906 15572 10908
rect 15596 10906 15652 10908
rect 15676 10906 15732 10908
rect 15756 10906 15812 10908
rect 15516 10854 15562 10906
rect 15562 10854 15572 10906
rect 15596 10854 15626 10906
rect 15626 10854 15638 10906
rect 15638 10854 15652 10906
rect 15676 10854 15690 10906
rect 15690 10854 15702 10906
rect 15702 10854 15732 10906
rect 15756 10854 15766 10906
rect 15766 10854 15812 10906
rect 15516 10852 15572 10854
rect 15596 10852 15652 10854
rect 15676 10852 15732 10854
rect 15756 10852 15812 10854
rect 15516 9818 15572 9820
rect 15596 9818 15652 9820
rect 15676 9818 15732 9820
rect 15756 9818 15812 9820
rect 15516 9766 15562 9818
rect 15562 9766 15572 9818
rect 15596 9766 15626 9818
rect 15626 9766 15638 9818
rect 15638 9766 15652 9818
rect 15676 9766 15690 9818
rect 15690 9766 15702 9818
rect 15702 9766 15732 9818
rect 15756 9766 15766 9818
rect 15766 9766 15812 9818
rect 15516 9764 15572 9766
rect 15596 9764 15652 9766
rect 15676 9764 15732 9766
rect 15756 9764 15812 9766
rect 15516 8730 15572 8732
rect 15596 8730 15652 8732
rect 15676 8730 15732 8732
rect 15756 8730 15812 8732
rect 15516 8678 15562 8730
rect 15562 8678 15572 8730
rect 15596 8678 15626 8730
rect 15626 8678 15638 8730
rect 15638 8678 15652 8730
rect 15676 8678 15690 8730
rect 15690 8678 15702 8730
rect 15702 8678 15732 8730
rect 15756 8678 15766 8730
rect 15766 8678 15812 8730
rect 15516 8676 15572 8678
rect 15596 8676 15652 8678
rect 15676 8676 15732 8678
rect 15756 8676 15812 8678
rect 16302 10512 16358 10568
rect 15516 7642 15572 7644
rect 15596 7642 15652 7644
rect 15676 7642 15732 7644
rect 15756 7642 15812 7644
rect 15516 7590 15562 7642
rect 15562 7590 15572 7642
rect 15596 7590 15626 7642
rect 15626 7590 15638 7642
rect 15638 7590 15652 7642
rect 15676 7590 15690 7642
rect 15690 7590 15702 7642
rect 15702 7590 15732 7642
rect 15756 7590 15766 7642
rect 15766 7590 15812 7642
rect 15516 7588 15572 7590
rect 15596 7588 15652 7590
rect 15676 7588 15732 7590
rect 15756 7588 15812 7590
rect 15516 6554 15572 6556
rect 15596 6554 15652 6556
rect 15676 6554 15732 6556
rect 15756 6554 15812 6556
rect 15516 6502 15562 6554
rect 15562 6502 15572 6554
rect 15596 6502 15626 6554
rect 15626 6502 15638 6554
rect 15638 6502 15652 6554
rect 15676 6502 15690 6554
rect 15690 6502 15702 6554
rect 15702 6502 15732 6554
rect 15756 6502 15766 6554
rect 15766 6502 15812 6554
rect 15516 6500 15572 6502
rect 15596 6500 15652 6502
rect 15676 6500 15732 6502
rect 15756 6500 15812 6502
rect 15516 5466 15572 5468
rect 15596 5466 15652 5468
rect 15676 5466 15732 5468
rect 15756 5466 15812 5468
rect 15516 5414 15562 5466
rect 15562 5414 15572 5466
rect 15596 5414 15626 5466
rect 15626 5414 15638 5466
rect 15638 5414 15652 5466
rect 15676 5414 15690 5466
rect 15690 5414 15702 5466
rect 15702 5414 15732 5466
rect 15756 5414 15766 5466
rect 15766 5414 15812 5466
rect 15516 5412 15572 5414
rect 15596 5412 15652 5414
rect 15676 5412 15732 5414
rect 15756 5412 15812 5414
rect 15566 5208 15622 5264
rect 15934 6296 15990 6352
rect 15750 4700 15752 4720
rect 15752 4700 15804 4720
rect 15804 4700 15806 4720
rect 15750 4664 15806 4700
rect 15516 4378 15572 4380
rect 15596 4378 15652 4380
rect 15676 4378 15732 4380
rect 15756 4378 15812 4380
rect 15516 4326 15562 4378
rect 15562 4326 15572 4378
rect 15596 4326 15626 4378
rect 15626 4326 15638 4378
rect 15638 4326 15652 4378
rect 15676 4326 15690 4378
rect 15690 4326 15702 4378
rect 15702 4326 15732 4378
rect 15756 4326 15766 4378
rect 15766 4326 15812 4378
rect 15516 4324 15572 4326
rect 15596 4324 15652 4326
rect 15676 4324 15732 4326
rect 15756 4324 15812 4326
rect 16210 7384 16266 7440
rect 16026 5616 16082 5672
rect 14278 756 14280 776
rect 14280 756 14332 776
rect 14332 756 14334 776
rect 14278 720 14334 756
rect 15198 2352 15254 2408
rect 15014 1944 15070 2000
rect 13966 570 14022 572
rect 14046 570 14102 572
rect 14126 570 14182 572
rect 14206 570 14262 572
rect 13966 518 14012 570
rect 14012 518 14022 570
rect 14046 518 14076 570
rect 14076 518 14088 570
rect 14088 518 14102 570
rect 14126 518 14140 570
rect 14140 518 14152 570
rect 14152 518 14182 570
rect 14206 518 14216 570
rect 14216 518 14262 570
rect 13966 516 14022 518
rect 14046 516 14102 518
rect 14126 516 14182 518
rect 14206 516 14262 518
rect 15516 3290 15572 3292
rect 15596 3290 15652 3292
rect 15676 3290 15732 3292
rect 15756 3290 15812 3292
rect 15516 3238 15562 3290
rect 15562 3238 15572 3290
rect 15596 3238 15626 3290
rect 15626 3238 15638 3290
rect 15638 3238 15652 3290
rect 15676 3238 15690 3290
rect 15690 3238 15702 3290
rect 15702 3238 15732 3290
rect 15756 3238 15766 3290
rect 15766 3238 15812 3290
rect 15516 3236 15572 3238
rect 15596 3236 15652 3238
rect 15676 3236 15732 3238
rect 15756 3236 15812 3238
rect 15842 2488 15898 2544
rect 15516 2202 15572 2204
rect 15596 2202 15652 2204
rect 15676 2202 15732 2204
rect 15756 2202 15812 2204
rect 15516 2150 15562 2202
rect 15562 2150 15572 2202
rect 15596 2150 15626 2202
rect 15626 2150 15638 2202
rect 15638 2150 15652 2202
rect 15676 2150 15690 2202
rect 15690 2150 15702 2202
rect 15702 2150 15732 2202
rect 15756 2150 15766 2202
rect 15766 2150 15812 2202
rect 15516 2148 15572 2150
rect 15596 2148 15652 2150
rect 15676 2148 15732 2150
rect 15756 2148 15812 2150
rect 15474 1828 15530 1864
rect 15474 1808 15476 1828
rect 15476 1808 15528 1828
rect 15528 1808 15530 1828
rect 15658 1808 15714 1864
rect 15516 1114 15572 1116
rect 15596 1114 15652 1116
rect 15676 1114 15732 1116
rect 15756 1114 15812 1116
rect 15516 1062 15562 1114
rect 15562 1062 15572 1114
rect 15596 1062 15626 1114
rect 15626 1062 15638 1114
rect 15638 1062 15652 1114
rect 15676 1062 15690 1114
rect 15690 1062 15702 1114
rect 15702 1062 15732 1114
rect 15756 1062 15766 1114
rect 15766 1062 15812 1114
rect 15516 1060 15572 1062
rect 15596 1060 15652 1062
rect 15676 1060 15732 1062
rect 15756 1060 15812 1062
rect 15842 856 15898 912
rect 18418 11056 18474 11112
rect 17066 10362 17122 10364
rect 17146 10362 17202 10364
rect 17226 10362 17282 10364
rect 17306 10362 17362 10364
rect 17066 10310 17112 10362
rect 17112 10310 17122 10362
rect 17146 10310 17176 10362
rect 17176 10310 17188 10362
rect 17188 10310 17202 10362
rect 17226 10310 17240 10362
rect 17240 10310 17252 10362
rect 17252 10310 17282 10362
rect 17306 10310 17316 10362
rect 17316 10310 17362 10362
rect 17066 10308 17122 10310
rect 17146 10308 17202 10310
rect 17226 10308 17282 10310
rect 17306 10308 17362 10310
rect 17066 9274 17122 9276
rect 17146 9274 17202 9276
rect 17226 9274 17282 9276
rect 17306 9274 17362 9276
rect 17066 9222 17112 9274
rect 17112 9222 17122 9274
rect 17146 9222 17176 9274
rect 17176 9222 17188 9274
rect 17188 9222 17202 9274
rect 17226 9222 17240 9274
rect 17240 9222 17252 9274
rect 17252 9222 17282 9274
rect 17306 9222 17316 9274
rect 17316 9222 17362 9274
rect 17066 9220 17122 9222
rect 17146 9220 17202 9222
rect 17226 9220 17282 9222
rect 17306 9220 17362 9222
rect 16302 6296 16358 6352
rect 16394 6160 16450 6216
rect 16118 4800 16174 4856
rect 16762 6840 16818 6896
rect 17066 8186 17122 8188
rect 17146 8186 17202 8188
rect 17226 8186 17282 8188
rect 17306 8186 17362 8188
rect 17066 8134 17112 8186
rect 17112 8134 17122 8186
rect 17146 8134 17176 8186
rect 17176 8134 17188 8186
rect 17188 8134 17202 8186
rect 17226 8134 17240 8186
rect 17240 8134 17252 8186
rect 17252 8134 17282 8186
rect 17306 8134 17316 8186
rect 17316 8134 17362 8186
rect 17066 8132 17122 8134
rect 17146 8132 17202 8134
rect 17226 8132 17282 8134
rect 17306 8132 17362 8134
rect 17066 7098 17122 7100
rect 17146 7098 17202 7100
rect 17226 7098 17282 7100
rect 17306 7098 17362 7100
rect 17066 7046 17112 7098
rect 17112 7046 17122 7098
rect 17146 7046 17176 7098
rect 17176 7046 17188 7098
rect 17188 7046 17202 7098
rect 17226 7046 17240 7098
rect 17240 7046 17252 7098
rect 17252 7046 17282 7098
rect 17306 7046 17316 7098
rect 17316 7046 17362 7098
rect 17066 7044 17122 7046
rect 17146 7044 17202 7046
rect 17226 7044 17282 7046
rect 17306 7044 17362 7046
rect 16394 4392 16450 4448
rect 16394 4120 16450 4176
rect 16302 3304 16358 3360
rect 16670 5228 16726 5264
rect 16670 5208 16672 5228
rect 16672 5208 16724 5228
rect 16724 5208 16726 5228
rect 16670 4664 16726 4720
rect 16578 4004 16634 4040
rect 16578 3984 16580 4004
rect 16580 3984 16632 4004
rect 16632 3984 16634 4004
rect 16394 2352 16450 2408
rect 16302 2100 16358 2136
rect 16302 2080 16304 2100
rect 16304 2080 16356 2100
rect 16356 2080 16358 2100
rect 16302 1944 16358 2000
rect 16578 2624 16634 2680
rect 16762 2760 16818 2816
rect 17130 6704 17186 6760
rect 17066 6010 17122 6012
rect 17146 6010 17202 6012
rect 17226 6010 17282 6012
rect 17306 6010 17362 6012
rect 17066 5958 17112 6010
rect 17112 5958 17122 6010
rect 17146 5958 17176 6010
rect 17176 5958 17188 6010
rect 17188 5958 17202 6010
rect 17226 5958 17240 6010
rect 17240 5958 17252 6010
rect 17252 5958 17282 6010
rect 17306 5958 17316 6010
rect 17316 5958 17362 6010
rect 17066 5956 17122 5958
rect 17146 5956 17202 5958
rect 17226 5956 17282 5958
rect 17306 5956 17362 5958
rect 17130 5752 17186 5808
rect 17222 5208 17278 5264
rect 18418 10548 18420 10568
rect 18420 10548 18472 10568
rect 18472 10548 18474 10568
rect 18418 10512 18474 10548
rect 17958 5752 18014 5808
rect 17866 5208 17922 5264
rect 17066 4922 17122 4924
rect 17146 4922 17202 4924
rect 17226 4922 17282 4924
rect 17306 4922 17362 4924
rect 17066 4870 17112 4922
rect 17112 4870 17122 4922
rect 17146 4870 17176 4922
rect 17176 4870 17188 4922
rect 17188 4870 17202 4922
rect 17226 4870 17240 4922
rect 17240 4870 17252 4922
rect 17252 4870 17282 4922
rect 17306 4870 17316 4922
rect 17316 4870 17362 4922
rect 17066 4868 17122 4870
rect 17146 4868 17202 4870
rect 17226 4868 17282 4870
rect 17306 4868 17362 4870
rect 17130 4392 17186 4448
rect 17498 4528 17554 4584
rect 17314 4428 17316 4448
rect 17316 4428 17368 4448
rect 17368 4428 17370 4448
rect 17314 4392 17370 4428
rect 17066 3834 17122 3836
rect 17146 3834 17202 3836
rect 17226 3834 17282 3836
rect 17306 3834 17362 3836
rect 17066 3782 17112 3834
rect 17112 3782 17122 3834
rect 17146 3782 17176 3834
rect 17176 3782 17188 3834
rect 17188 3782 17202 3834
rect 17226 3782 17240 3834
rect 17240 3782 17252 3834
rect 17252 3782 17282 3834
rect 17306 3782 17316 3834
rect 17316 3782 17362 3834
rect 17066 3780 17122 3782
rect 17146 3780 17202 3782
rect 17226 3780 17282 3782
rect 17306 3780 17362 3782
rect 16946 3304 17002 3360
rect 16854 2352 16910 2408
rect 17314 3576 17370 3632
rect 17222 3032 17278 3088
rect 17498 3304 17554 3360
rect 17682 3304 17738 3360
rect 18050 5480 18106 5536
rect 18326 8472 18382 8528
rect 18616 10906 18672 10908
rect 18696 10906 18752 10908
rect 18776 10906 18832 10908
rect 18856 10906 18912 10908
rect 18616 10854 18662 10906
rect 18662 10854 18672 10906
rect 18696 10854 18726 10906
rect 18726 10854 18738 10906
rect 18738 10854 18752 10906
rect 18776 10854 18790 10906
rect 18790 10854 18802 10906
rect 18802 10854 18832 10906
rect 18856 10854 18866 10906
rect 18866 10854 18912 10906
rect 18616 10852 18672 10854
rect 18696 10852 18752 10854
rect 18776 10852 18832 10854
rect 18856 10852 18912 10854
rect 18616 9818 18672 9820
rect 18696 9818 18752 9820
rect 18776 9818 18832 9820
rect 18856 9818 18912 9820
rect 18616 9766 18662 9818
rect 18662 9766 18672 9818
rect 18696 9766 18726 9818
rect 18726 9766 18738 9818
rect 18738 9766 18752 9818
rect 18776 9766 18790 9818
rect 18790 9766 18802 9818
rect 18802 9766 18832 9818
rect 18856 9766 18866 9818
rect 18866 9766 18912 9818
rect 18616 9764 18672 9766
rect 18696 9764 18752 9766
rect 18776 9764 18832 9766
rect 18856 9764 18912 9766
rect 18616 8730 18672 8732
rect 18696 8730 18752 8732
rect 18776 8730 18832 8732
rect 18856 8730 18912 8732
rect 18616 8678 18662 8730
rect 18662 8678 18672 8730
rect 18696 8678 18726 8730
rect 18726 8678 18738 8730
rect 18738 8678 18752 8730
rect 18776 8678 18790 8730
rect 18790 8678 18802 8730
rect 18802 8678 18832 8730
rect 18856 8678 18866 8730
rect 18866 8678 18912 8730
rect 18616 8676 18672 8678
rect 18696 8676 18752 8678
rect 18776 8676 18832 8678
rect 18856 8676 18912 8678
rect 18970 8200 19026 8256
rect 18616 7642 18672 7644
rect 18696 7642 18752 7644
rect 18776 7642 18832 7644
rect 18856 7642 18912 7644
rect 18616 7590 18662 7642
rect 18662 7590 18672 7642
rect 18696 7590 18726 7642
rect 18726 7590 18738 7642
rect 18738 7590 18752 7642
rect 18776 7590 18790 7642
rect 18790 7590 18802 7642
rect 18802 7590 18832 7642
rect 18856 7590 18866 7642
rect 18866 7590 18912 7642
rect 18616 7588 18672 7590
rect 18696 7588 18752 7590
rect 18776 7588 18832 7590
rect 18856 7588 18912 7590
rect 18510 6704 18566 6760
rect 18616 6554 18672 6556
rect 18696 6554 18752 6556
rect 18776 6554 18832 6556
rect 18856 6554 18912 6556
rect 18616 6502 18662 6554
rect 18662 6502 18672 6554
rect 18696 6502 18726 6554
rect 18726 6502 18738 6554
rect 18738 6502 18752 6554
rect 18776 6502 18790 6554
rect 18790 6502 18802 6554
rect 18802 6502 18832 6554
rect 18856 6502 18866 6554
rect 18866 6502 18912 6554
rect 18616 6500 18672 6502
rect 18696 6500 18752 6502
rect 18776 6500 18832 6502
rect 18856 6500 18912 6502
rect 18510 5616 18566 5672
rect 18616 5466 18672 5468
rect 18696 5466 18752 5468
rect 18776 5466 18832 5468
rect 18856 5466 18912 5468
rect 18616 5414 18662 5466
rect 18662 5414 18672 5466
rect 18696 5414 18726 5466
rect 18726 5414 18738 5466
rect 18738 5414 18752 5466
rect 18776 5414 18790 5466
rect 18790 5414 18802 5466
rect 18802 5414 18832 5466
rect 18856 5414 18866 5466
rect 18866 5414 18912 5466
rect 18616 5412 18672 5414
rect 18696 5412 18752 5414
rect 18776 5412 18832 5414
rect 18856 5412 18912 5414
rect 18970 5208 19026 5264
rect 17066 2746 17122 2748
rect 17146 2746 17202 2748
rect 17226 2746 17282 2748
rect 17306 2746 17362 2748
rect 17066 2694 17112 2746
rect 17112 2694 17122 2746
rect 17146 2694 17176 2746
rect 17176 2694 17188 2746
rect 17188 2694 17202 2746
rect 17226 2694 17240 2746
rect 17240 2694 17252 2746
rect 17252 2694 17282 2746
rect 17306 2694 17316 2746
rect 17316 2694 17362 2746
rect 17066 2692 17122 2694
rect 17146 2692 17202 2694
rect 17226 2692 17282 2694
rect 17306 2692 17362 2694
rect 17066 1658 17122 1660
rect 17146 1658 17202 1660
rect 17226 1658 17282 1660
rect 17306 1658 17362 1660
rect 17066 1606 17112 1658
rect 17112 1606 17122 1658
rect 17146 1606 17176 1658
rect 17176 1606 17188 1658
rect 17188 1606 17202 1658
rect 17226 1606 17240 1658
rect 17240 1606 17252 1658
rect 17252 1606 17282 1658
rect 17306 1606 17316 1658
rect 17316 1606 17362 1658
rect 17066 1604 17122 1606
rect 17146 1604 17202 1606
rect 17226 1604 17282 1606
rect 17306 1604 17362 1606
rect 17406 1300 17408 1320
rect 17408 1300 17460 1320
rect 17460 1300 17462 1320
rect 17406 1264 17462 1300
rect 17682 3032 17738 3088
rect 17774 2352 17830 2408
rect 18050 2896 18106 2952
rect 17958 2080 18014 2136
rect 17866 1944 17922 2000
rect 18234 3440 18290 3496
rect 18050 1420 18106 1456
rect 18050 1400 18052 1420
rect 18052 1400 18104 1420
rect 18104 1400 18106 1420
rect 17866 756 17868 776
rect 17868 756 17920 776
rect 17920 756 17922 776
rect 17866 720 17922 756
rect 18616 4378 18672 4380
rect 18696 4378 18752 4380
rect 18776 4378 18832 4380
rect 18856 4378 18912 4380
rect 18616 4326 18662 4378
rect 18662 4326 18672 4378
rect 18696 4326 18726 4378
rect 18726 4326 18738 4378
rect 18738 4326 18752 4378
rect 18776 4326 18790 4378
rect 18790 4326 18802 4378
rect 18802 4326 18832 4378
rect 18856 4326 18866 4378
rect 18866 4326 18912 4378
rect 18616 4324 18672 4326
rect 18696 4324 18752 4326
rect 18776 4324 18832 4326
rect 18856 4324 18912 4326
rect 18970 4120 19026 4176
rect 18970 3712 19026 3768
rect 18616 3290 18672 3292
rect 18696 3290 18752 3292
rect 18776 3290 18832 3292
rect 18856 3290 18912 3292
rect 18616 3238 18662 3290
rect 18662 3238 18672 3290
rect 18696 3238 18726 3290
rect 18726 3238 18738 3290
rect 18738 3238 18752 3290
rect 18776 3238 18790 3290
rect 18790 3238 18802 3290
rect 18802 3238 18832 3290
rect 18856 3238 18866 3290
rect 18866 3238 18912 3290
rect 18616 3236 18672 3238
rect 18696 3236 18752 3238
rect 18776 3236 18832 3238
rect 18856 3236 18912 3238
rect 19062 2216 19118 2272
rect 18616 2202 18672 2204
rect 18696 2202 18752 2204
rect 18776 2202 18832 2204
rect 18856 2202 18912 2204
rect 18616 2150 18662 2202
rect 18662 2150 18672 2202
rect 18696 2150 18726 2202
rect 18726 2150 18738 2202
rect 18738 2150 18752 2202
rect 18776 2150 18790 2202
rect 18790 2150 18802 2202
rect 18802 2150 18832 2202
rect 18856 2150 18866 2202
rect 18866 2150 18912 2202
rect 18616 2148 18672 2150
rect 18696 2148 18752 2150
rect 18776 2148 18832 2150
rect 18856 2148 18912 2150
rect 18510 1944 18566 2000
rect 18616 1114 18672 1116
rect 18696 1114 18752 1116
rect 18776 1114 18832 1116
rect 18856 1114 18912 1116
rect 18616 1062 18662 1114
rect 18662 1062 18672 1114
rect 18696 1062 18726 1114
rect 18726 1062 18738 1114
rect 18738 1062 18752 1114
rect 18776 1062 18790 1114
rect 18790 1062 18802 1114
rect 18802 1062 18832 1114
rect 18856 1062 18866 1114
rect 18866 1062 18912 1114
rect 18616 1060 18672 1062
rect 18696 1060 18752 1062
rect 18776 1060 18832 1062
rect 18856 1060 18912 1062
rect 17066 570 17122 572
rect 17146 570 17202 572
rect 17226 570 17282 572
rect 17306 570 17362 572
rect 17066 518 17112 570
rect 17112 518 17122 570
rect 17146 518 17176 570
rect 17176 518 17188 570
rect 17188 518 17202 570
rect 17226 518 17240 570
rect 17240 518 17252 570
rect 17252 518 17282 570
rect 17306 518 17316 570
rect 17316 518 17362 570
rect 17066 516 17122 518
rect 17146 516 17202 518
rect 17226 516 17282 518
rect 17306 516 17362 518
<< metal3 >>
rect 19200 11250 20000 11280
rect 18462 11190 20000 11250
rect 18462 11117 18522 11190
rect 19200 11160 20000 11190
rect 18413 11112 18522 11117
rect 18413 11056 18418 11112
rect 18474 11056 18522 11112
rect 18413 11054 18522 11056
rect 18413 11051 18479 11054
rect 3106 10912 3422 10913
rect 3106 10848 3112 10912
rect 3176 10848 3192 10912
rect 3256 10848 3272 10912
rect 3336 10848 3352 10912
rect 3416 10848 3422 10912
rect 3106 10847 3422 10848
rect 6206 10912 6522 10913
rect 6206 10848 6212 10912
rect 6276 10848 6292 10912
rect 6356 10848 6372 10912
rect 6436 10848 6452 10912
rect 6516 10848 6522 10912
rect 6206 10847 6522 10848
rect 9306 10912 9622 10913
rect 9306 10848 9312 10912
rect 9376 10848 9392 10912
rect 9456 10848 9472 10912
rect 9536 10848 9552 10912
rect 9616 10848 9622 10912
rect 9306 10847 9622 10848
rect 12406 10912 12722 10913
rect 12406 10848 12412 10912
rect 12476 10848 12492 10912
rect 12556 10848 12572 10912
rect 12636 10848 12652 10912
rect 12716 10848 12722 10912
rect 12406 10847 12722 10848
rect 15506 10912 15822 10913
rect 15506 10848 15512 10912
rect 15576 10848 15592 10912
rect 15656 10848 15672 10912
rect 15736 10848 15752 10912
rect 15816 10848 15822 10912
rect 15506 10847 15822 10848
rect 18606 10912 18922 10913
rect 18606 10848 18612 10912
rect 18676 10848 18692 10912
rect 18756 10848 18772 10912
rect 18836 10848 18852 10912
rect 18916 10848 18922 10912
rect 18606 10847 18922 10848
rect 2497 10706 2563 10709
rect 9305 10706 9371 10709
rect 2497 10704 9371 10706
rect 2497 10648 2502 10704
rect 2558 10648 9310 10704
rect 9366 10648 9371 10704
rect 2497 10646 9371 10648
rect 2497 10643 2563 10646
rect 9305 10643 9371 10646
rect 4061 10570 4127 10573
rect 5533 10570 5599 10573
rect 4061 10568 5599 10570
rect 4061 10512 4066 10568
rect 4122 10512 5538 10568
rect 5594 10512 5599 10568
rect 4061 10510 5599 10512
rect 4061 10507 4127 10510
rect 5533 10507 5599 10510
rect 10133 10570 10199 10573
rect 15193 10570 15259 10573
rect 10133 10568 15259 10570
rect 10133 10512 10138 10568
rect 10194 10512 15198 10568
rect 15254 10512 15259 10568
rect 10133 10510 15259 10512
rect 10133 10507 10199 10510
rect 15193 10507 15259 10510
rect 16297 10570 16363 10573
rect 18413 10570 18479 10573
rect 16297 10568 18479 10570
rect 16297 10512 16302 10568
rect 16358 10512 18418 10568
rect 18474 10512 18479 10568
rect 16297 10510 18479 10512
rect 16297 10507 16363 10510
rect 18413 10507 18479 10510
rect 4656 10368 4972 10369
rect 4656 10304 4662 10368
rect 4726 10304 4742 10368
rect 4806 10304 4822 10368
rect 4886 10304 4902 10368
rect 4966 10304 4972 10368
rect 4656 10303 4972 10304
rect 7756 10368 8072 10369
rect 7756 10304 7762 10368
rect 7826 10304 7842 10368
rect 7906 10304 7922 10368
rect 7986 10304 8002 10368
rect 8066 10304 8072 10368
rect 7756 10303 8072 10304
rect 10856 10368 11172 10369
rect 10856 10304 10862 10368
rect 10926 10304 10942 10368
rect 11006 10304 11022 10368
rect 11086 10304 11102 10368
rect 11166 10304 11172 10368
rect 10856 10303 11172 10304
rect 13956 10368 14272 10369
rect 13956 10304 13962 10368
rect 14026 10304 14042 10368
rect 14106 10304 14122 10368
rect 14186 10304 14202 10368
rect 14266 10304 14272 10368
rect 13956 10303 14272 10304
rect 17056 10368 17372 10369
rect 17056 10304 17062 10368
rect 17126 10304 17142 10368
rect 17206 10304 17222 10368
rect 17286 10304 17302 10368
rect 17366 10304 17372 10368
rect 17056 10303 17372 10304
rect 1117 10162 1183 10165
rect 4429 10162 4495 10165
rect 1117 10160 4495 10162
rect 1117 10104 1122 10160
rect 1178 10104 4434 10160
rect 4490 10104 4495 10160
rect 1117 10102 4495 10104
rect 1117 10099 1183 10102
rect 4429 10099 4495 10102
rect 10133 10162 10199 10165
rect 11973 10162 12039 10165
rect 10133 10160 12039 10162
rect 10133 10104 10138 10160
rect 10194 10104 11978 10160
rect 12034 10104 12039 10160
rect 10133 10102 12039 10104
rect 10133 10099 10199 10102
rect 11973 10099 12039 10102
rect 3141 10026 3207 10029
rect 3509 10026 3575 10029
rect 4889 10026 4955 10029
rect 3141 10024 4955 10026
rect 3141 9968 3146 10024
rect 3202 9968 3514 10024
rect 3570 9968 4894 10024
rect 4950 9968 4955 10024
rect 3141 9966 4955 9968
rect 3141 9963 3207 9966
rect 3509 9963 3575 9966
rect 4889 9963 4955 9966
rect 9581 10026 9647 10029
rect 10409 10026 10475 10029
rect 9581 10024 10475 10026
rect 9581 9968 9586 10024
rect 9642 9968 10414 10024
rect 10470 9968 10475 10024
rect 9581 9966 10475 9968
rect 9581 9963 9647 9966
rect 10409 9963 10475 9966
rect 15193 10026 15259 10029
rect 15193 10024 19074 10026
rect 15193 9968 15198 10024
rect 15254 9968 19074 10024
rect 15193 9966 19074 9968
rect 15193 9963 15259 9966
rect 3106 9824 3422 9825
rect 3106 9760 3112 9824
rect 3176 9760 3192 9824
rect 3256 9760 3272 9824
rect 3336 9760 3352 9824
rect 3416 9760 3422 9824
rect 3106 9759 3422 9760
rect 6206 9824 6522 9825
rect 6206 9760 6212 9824
rect 6276 9760 6292 9824
rect 6356 9760 6372 9824
rect 6436 9760 6452 9824
rect 6516 9760 6522 9824
rect 6206 9759 6522 9760
rect 9306 9824 9622 9825
rect 9306 9760 9312 9824
rect 9376 9760 9392 9824
rect 9456 9760 9472 9824
rect 9536 9760 9552 9824
rect 9616 9760 9622 9824
rect 9306 9759 9622 9760
rect 12406 9824 12722 9825
rect 12406 9760 12412 9824
rect 12476 9760 12492 9824
rect 12556 9760 12572 9824
rect 12636 9760 12652 9824
rect 12716 9760 12722 9824
rect 12406 9759 12722 9760
rect 15506 9824 15822 9825
rect 15506 9760 15512 9824
rect 15576 9760 15592 9824
rect 15656 9760 15672 9824
rect 15736 9760 15752 9824
rect 15816 9760 15822 9824
rect 15506 9759 15822 9760
rect 18606 9824 18922 9825
rect 18606 9760 18612 9824
rect 18676 9760 18692 9824
rect 18756 9760 18772 9824
rect 18836 9760 18852 9824
rect 18916 9760 18922 9824
rect 18606 9759 18922 9760
rect 19014 9754 19074 9966
rect 19200 9754 20000 9784
rect 19014 9694 20000 9754
rect 19200 9664 20000 9694
rect 657 9482 723 9485
rect 1761 9482 1827 9485
rect 657 9480 1827 9482
rect 657 9424 662 9480
rect 718 9424 1766 9480
rect 1822 9424 1827 9480
rect 657 9422 1827 9424
rect 657 9419 723 9422
rect 1761 9419 1827 9422
rect 4656 9280 4972 9281
rect 4656 9216 4662 9280
rect 4726 9216 4742 9280
rect 4806 9216 4822 9280
rect 4886 9216 4902 9280
rect 4966 9216 4972 9280
rect 4656 9215 4972 9216
rect 7756 9280 8072 9281
rect 7756 9216 7762 9280
rect 7826 9216 7842 9280
rect 7906 9216 7922 9280
rect 7986 9216 8002 9280
rect 8066 9216 8072 9280
rect 7756 9215 8072 9216
rect 10856 9280 11172 9281
rect 10856 9216 10862 9280
rect 10926 9216 10942 9280
rect 11006 9216 11022 9280
rect 11086 9216 11102 9280
rect 11166 9216 11172 9280
rect 10856 9215 11172 9216
rect 13956 9280 14272 9281
rect 13956 9216 13962 9280
rect 14026 9216 14042 9280
rect 14106 9216 14122 9280
rect 14186 9216 14202 9280
rect 14266 9216 14272 9280
rect 13956 9215 14272 9216
rect 17056 9280 17372 9281
rect 17056 9216 17062 9280
rect 17126 9216 17142 9280
rect 17206 9216 17222 9280
rect 17286 9216 17302 9280
rect 17366 9216 17372 9280
rect 17056 9215 17372 9216
rect 3106 8736 3422 8737
rect 3106 8672 3112 8736
rect 3176 8672 3192 8736
rect 3256 8672 3272 8736
rect 3336 8672 3352 8736
rect 3416 8672 3422 8736
rect 3106 8671 3422 8672
rect 6206 8736 6522 8737
rect 6206 8672 6212 8736
rect 6276 8672 6292 8736
rect 6356 8672 6372 8736
rect 6436 8672 6452 8736
rect 6516 8672 6522 8736
rect 6206 8671 6522 8672
rect 9306 8736 9622 8737
rect 9306 8672 9312 8736
rect 9376 8672 9392 8736
rect 9456 8672 9472 8736
rect 9536 8672 9552 8736
rect 9616 8672 9622 8736
rect 9306 8671 9622 8672
rect 12406 8736 12722 8737
rect 12406 8672 12412 8736
rect 12476 8672 12492 8736
rect 12556 8672 12572 8736
rect 12636 8672 12652 8736
rect 12716 8672 12722 8736
rect 12406 8671 12722 8672
rect 15506 8736 15822 8737
rect 15506 8672 15512 8736
rect 15576 8672 15592 8736
rect 15656 8672 15672 8736
rect 15736 8672 15752 8736
rect 15816 8672 15822 8736
rect 15506 8671 15822 8672
rect 18606 8736 18922 8737
rect 18606 8672 18612 8736
rect 18676 8672 18692 8736
rect 18756 8672 18772 8736
rect 18836 8672 18852 8736
rect 18916 8672 18922 8736
rect 18606 8671 18922 8672
rect 16798 8468 16804 8532
rect 16868 8530 16874 8532
rect 18321 8530 18387 8533
rect 16868 8528 18387 8530
rect 16868 8472 18326 8528
rect 18382 8472 18387 8528
rect 16868 8470 18387 8472
rect 16868 8468 16874 8470
rect 18321 8467 18387 8470
rect 565 8394 631 8397
rect 1025 8394 1091 8397
rect 4981 8394 5047 8397
rect 565 8392 5047 8394
rect 565 8336 570 8392
rect 626 8336 1030 8392
rect 1086 8336 4986 8392
rect 5042 8336 5047 8392
rect 565 8334 5047 8336
rect 565 8331 631 8334
rect 1025 8331 1091 8334
rect 4981 8331 5047 8334
rect 10777 8394 10843 8397
rect 12341 8394 12407 8397
rect 10777 8392 12407 8394
rect 10777 8336 10782 8392
rect 10838 8336 12346 8392
rect 12402 8336 12407 8392
rect 10777 8334 12407 8336
rect 10777 8331 10843 8334
rect 12341 8331 12407 8334
rect 18965 8258 19031 8261
rect 19200 8258 20000 8288
rect 18965 8256 20000 8258
rect 18965 8200 18970 8256
rect 19026 8200 20000 8256
rect 18965 8198 20000 8200
rect 18965 8195 19031 8198
rect 4656 8192 4972 8193
rect 4656 8128 4662 8192
rect 4726 8128 4742 8192
rect 4806 8128 4822 8192
rect 4886 8128 4902 8192
rect 4966 8128 4972 8192
rect 4656 8127 4972 8128
rect 7756 8192 8072 8193
rect 7756 8128 7762 8192
rect 7826 8128 7842 8192
rect 7906 8128 7922 8192
rect 7986 8128 8002 8192
rect 8066 8128 8072 8192
rect 7756 8127 8072 8128
rect 10856 8192 11172 8193
rect 10856 8128 10862 8192
rect 10926 8128 10942 8192
rect 11006 8128 11022 8192
rect 11086 8128 11102 8192
rect 11166 8128 11172 8192
rect 10856 8127 11172 8128
rect 13956 8192 14272 8193
rect 13956 8128 13962 8192
rect 14026 8128 14042 8192
rect 14106 8128 14122 8192
rect 14186 8128 14202 8192
rect 14266 8128 14272 8192
rect 13956 8127 14272 8128
rect 17056 8192 17372 8193
rect 17056 8128 17062 8192
rect 17126 8128 17142 8192
rect 17206 8128 17222 8192
rect 17286 8128 17302 8192
rect 17366 8128 17372 8192
rect 19200 8168 20000 8198
rect 17056 8127 17372 8128
rect 657 7986 723 7989
rect 2313 7986 2379 7989
rect 657 7984 2379 7986
rect 657 7928 662 7984
rect 718 7928 2318 7984
rect 2374 7928 2379 7984
rect 657 7926 2379 7928
rect 657 7923 723 7926
rect 2313 7923 2379 7926
rect 11697 7986 11763 7989
rect 12157 7986 12223 7989
rect 11697 7984 12223 7986
rect 11697 7928 11702 7984
rect 11758 7928 12162 7984
rect 12218 7928 12223 7984
rect 11697 7926 12223 7928
rect 11697 7923 11763 7926
rect 12157 7923 12223 7926
rect 3106 7648 3422 7649
rect 3106 7584 3112 7648
rect 3176 7584 3192 7648
rect 3256 7584 3272 7648
rect 3336 7584 3352 7648
rect 3416 7584 3422 7648
rect 3106 7583 3422 7584
rect 6206 7648 6522 7649
rect 6206 7584 6212 7648
rect 6276 7584 6292 7648
rect 6356 7584 6372 7648
rect 6436 7584 6452 7648
rect 6516 7584 6522 7648
rect 6206 7583 6522 7584
rect 9306 7648 9622 7649
rect 9306 7584 9312 7648
rect 9376 7584 9392 7648
rect 9456 7584 9472 7648
rect 9536 7584 9552 7648
rect 9616 7584 9622 7648
rect 9306 7583 9622 7584
rect 12406 7648 12722 7649
rect 12406 7584 12412 7648
rect 12476 7584 12492 7648
rect 12556 7584 12572 7648
rect 12636 7584 12652 7648
rect 12716 7584 12722 7648
rect 12406 7583 12722 7584
rect 15506 7648 15822 7649
rect 15506 7584 15512 7648
rect 15576 7584 15592 7648
rect 15656 7584 15672 7648
rect 15736 7584 15752 7648
rect 15816 7584 15822 7648
rect 15506 7583 15822 7584
rect 18606 7648 18922 7649
rect 18606 7584 18612 7648
rect 18676 7584 18692 7648
rect 18756 7584 18772 7648
rect 18836 7584 18852 7648
rect 18916 7584 18922 7648
rect 18606 7583 18922 7584
rect 933 7442 999 7445
rect 3785 7442 3851 7445
rect 933 7440 3851 7442
rect 933 7384 938 7440
rect 994 7384 3790 7440
rect 3846 7384 3851 7440
rect 933 7382 3851 7384
rect 933 7379 999 7382
rect 3785 7379 3851 7382
rect 16062 7380 16068 7444
rect 16132 7442 16138 7444
rect 16205 7442 16271 7445
rect 16132 7440 16271 7442
rect 16132 7384 16210 7440
rect 16266 7384 16271 7440
rect 16132 7382 16271 7384
rect 16132 7380 16138 7382
rect 16205 7379 16271 7382
rect 565 7306 631 7309
rect 2497 7306 2563 7309
rect 4245 7306 4311 7309
rect 565 7304 4311 7306
rect 565 7248 570 7304
rect 626 7248 2502 7304
rect 2558 7248 4250 7304
rect 4306 7248 4311 7304
rect 565 7246 4311 7248
rect 565 7243 631 7246
rect 2497 7243 2563 7246
rect 4245 7243 4311 7246
rect 10409 7306 10475 7309
rect 16798 7306 16804 7308
rect 10409 7304 16804 7306
rect 10409 7248 10414 7304
rect 10470 7248 16804 7304
rect 10409 7246 16804 7248
rect 10409 7243 10475 7246
rect 16798 7244 16804 7246
rect 16868 7244 16874 7308
rect 1209 7170 1275 7173
rect 3049 7170 3115 7173
rect 1209 7168 3115 7170
rect 1209 7112 1214 7168
rect 1270 7112 3054 7168
rect 3110 7112 3115 7168
rect 1209 7110 3115 7112
rect 1209 7107 1275 7110
rect 3049 7107 3115 7110
rect 4656 7104 4972 7105
rect 4656 7040 4662 7104
rect 4726 7040 4742 7104
rect 4806 7040 4822 7104
rect 4886 7040 4902 7104
rect 4966 7040 4972 7104
rect 4656 7039 4972 7040
rect 7756 7104 8072 7105
rect 7756 7040 7762 7104
rect 7826 7040 7842 7104
rect 7906 7040 7922 7104
rect 7986 7040 8002 7104
rect 8066 7040 8072 7104
rect 7756 7039 8072 7040
rect 10856 7104 11172 7105
rect 10856 7040 10862 7104
rect 10926 7040 10942 7104
rect 11006 7040 11022 7104
rect 11086 7040 11102 7104
rect 11166 7040 11172 7104
rect 10856 7039 11172 7040
rect 13956 7104 14272 7105
rect 13956 7040 13962 7104
rect 14026 7040 14042 7104
rect 14106 7040 14122 7104
rect 14186 7040 14202 7104
rect 14266 7040 14272 7104
rect 13956 7039 14272 7040
rect 17056 7104 17372 7105
rect 17056 7040 17062 7104
rect 17126 7040 17142 7104
rect 17206 7040 17222 7104
rect 17286 7040 17302 7104
rect 17366 7040 17372 7104
rect 17056 7039 17372 7040
rect 841 7034 907 7037
rect 2405 7034 2471 7037
rect 841 7032 2471 7034
rect 841 6976 846 7032
rect 902 6976 2410 7032
rect 2466 6976 2471 7032
rect 841 6974 2471 6976
rect 841 6971 907 6974
rect 2405 6971 2471 6974
rect 2957 7034 3023 7037
rect 4153 7034 4219 7037
rect 2957 7032 4219 7034
rect 2957 6976 2962 7032
rect 3018 6976 4158 7032
rect 4214 6976 4219 7032
rect 2957 6974 4219 6976
rect 2957 6971 3023 6974
rect 4153 6971 4219 6974
rect 749 6898 815 6901
rect 5441 6898 5507 6901
rect 749 6896 5507 6898
rect 749 6840 754 6896
rect 810 6840 5446 6896
rect 5502 6840 5507 6896
rect 749 6838 5507 6840
rect 749 6835 815 6838
rect 5441 6835 5507 6838
rect 6085 6898 6151 6901
rect 7189 6898 7255 6901
rect 6085 6896 7255 6898
rect 6085 6840 6090 6896
rect 6146 6840 7194 6896
rect 7250 6840 7255 6896
rect 6085 6838 7255 6840
rect 6085 6835 6151 6838
rect 7189 6835 7255 6838
rect 10041 6898 10107 6901
rect 14641 6898 14707 6901
rect 16757 6898 16823 6901
rect 10041 6896 16823 6898
rect 10041 6840 10046 6896
rect 10102 6840 14646 6896
rect 14702 6840 16762 6896
rect 16818 6840 16823 6896
rect 10041 6838 16823 6840
rect 10041 6835 10107 6838
rect 14641 6835 14707 6838
rect 16757 6835 16823 6838
rect 1301 6762 1367 6765
rect 3417 6762 3483 6765
rect 1301 6760 3483 6762
rect 1301 6704 1306 6760
rect 1362 6704 3422 6760
rect 3478 6704 3483 6760
rect 1301 6702 3483 6704
rect 1301 6699 1367 6702
rect 3417 6699 3483 6702
rect 6729 6762 6795 6765
rect 7925 6762 7991 6765
rect 6729 6760 7991 6762
rect 6729 6704 6734 6760
rect 6790 6704 7930 6760
rect 7986 6704 7991 6760
rect 6729 6702 7991 6704
rect 6729 6699 6795 6702
rect 7925 6699 7991 6702
rect 14917 6762 14983 6765
rect 16430 6762 16436 6764
rect 14917 6760 16436 6762
rect 14917 6704 14922 6760
rect 14978 6704 16436 6760
rect 14917 6702 16436 6704
rect 14917 6699 14983 6702
rect 16430 6700 16436 6702
rect 16500 6762 16506 6764
rect 17125 6762 17191 6765
rect 16500 6760 17191 6762
rect 16500 6704 17130 6760
rect 17186 6704 17191 6760
rect 16500 6702 17191 6704
rect 16500 6700 16506 6702
rect 17125 6699 17191 6702
rect 18505 6762 18571 6765
rect 19200 6762 20000 6792
rect 18505 6760 20000 6762
rect 18505 6704 18510 6760
rect 18566 6704 20000 6760
rect 18505 6702 20000 6704
rect 18505 6699 18571 6702
rect 19200 6672 20000 6702
rect 3106 6560 3422 6561
rect 3106 6496 3112 6560
rect 3176 6496 3192 6560
rect 3256 6496 3272 6560
rect 3336 6496 3352 6560
rect 3416 6496 3422 6560
rect 3106 6495 3422 6496
rect 6206 6560 6522 6561
rect 6206 6496 6212 6560
rect 6276 6496 6292 6560
rect 6356 6496 6372 6560
rect 6436 6496 6452 6560
rect 6516 6496 6522 6560
rect 6206 6495 6522 6496
rect 9306 6560 9622 6561
rect 9306 6496 9312 6560
rect 9376 6496 9392 6560
rect 9456 6496 9472 6560
rect 9536 6496 9552 6560
rect 9616 6496 9622 6560
rect 9306 6495 9622 6496
rect 12406 6560 12722 6561
rect 12406 6496 12412 6560
rect 12476 6496 12492 6560
rect 12556 6496 12572 6560
rect 12636 6496 12652 6560
rect 12716 6496 12722 6560
rect 12406 6495 12722 6496
rect 15506 6560 15822 6561
rect 15506 6496 15512 6560
rect 15576 6496 15592 6560
rect 15656 6496 15672 6560
rect 15736 6496 15752 6560
rect 15816 6496 15822 6560
rect 15506 6495 15822 6496
rect 18606 6560 18922 6561
rect 18606 6496 18612 6560
rect 18676 6496 18692 6560
rect 18756 6496 18772 6560
rect 18836 6496 18852 6560
rect 18916 6496 18922 6560
rect 18606 6495 18922 6496
rect 2129 6354 2195 6357
rect 3233 6354 3299 6357
rect 2129 6352 3299 6354
rect 2129 6296 2134 6352
rect 2190 6296 3238 6352
rect 3294 6296 3299 6352
rect 2129 6294 3299 6296
rect 2129 6291 2195 6294
rect 3233 6291 3299 6294
rect 15929 6354 15995 6357
rect 16297 6354 16363 6357
rect 15929 6352 16363 6354
rect 15929 6296 15934 6352
rect 15990 6296 16302 6352
rect 16358 6296 16363 6352
rect 15929 6294 16363 6296
rect 15929 6291 15995 6294
rect 16297 6291 16363 6294
rect 841 6218 907 6221
rect 4245 6218 4311 6221
rect 841 6216 4311 6218
rect 841 6160 846 6216
rect 902 6160 4250 6216
rect 4306 6160 4311 6216
rect 841 6158 4311 6160
rect 841 6155 907 6158
rect 4245 6155 4311 6158
rect 11973 6218 12039 6221
rect 13537 6218 13603 6221
rect 11973 6216 13603 6218
rect 11973 6160 11978 6216
rect 12034 6160 13542 6216
rect 13598 6160 13603 6216
rect 11973 6158 13603 6160
rect 11973 6155 12039 6158
rect 13537 6155 13603 6158
rect 15101 6218 15167 6221
rect 16389 6218 16455 6221
rect 15101 6216 16455 6218
rect 15101 6160 15106 6216
rect 15162 6160 16394 6216
rect 16450 6160 16455 6216
rect 15101 6158 16455 6160
rect 15101 6155 15167 6158
rect 16389 6155 16455 6158
rect 4656 6016 4972 6017
rect 4656 5952 4662 6016
rect 4726 5952 4742 6016
rect 4806 5952 4822 6016
rect 4886 5952 4902 6016
rect 4966 5952 4972 6016
rect 4656 5951 4972 5952
rect 7756 6016 8072 6017
rect 7756 5952 7762 6016
rect 7826 5952 7842 6016
rect 7906 5952 7922 6016
rect 7986 5952 8002 6016
rect 8066 5952 8072 6016
rect 7756 5951 8072 5952
rect 10856 6016 11172 6017
rect 10856 5952 10862 6016
rect 10926 5952 10942 6016
rect 11006 5952 11022 6016
rect 11086 5952 11102 6016
rect 11166 5952 11172 6016
rect 10856 5951 11172 5952
rect 13956 6016 14272 6017
rect 13956 5952 13962 6016
rect 14026 5952 14042 6016
rect 14106 5952 14122 6016
rect 14186 5952 14202 6016
rect 14266 5952 14272 6016
rect 13956 5951 14272 5952
rect 17056 6016 17372 6017
rect 17056 5952 17062 6016
rect 17126 5952 17142 6016
rect 17206 5952 17222 6016
rect 17286 5952 17302 6016
rect 17366 5952 17372 6016
rect 17056 5951 17372 5952
rect 5901 5810 5967 5813
rect 7097 5810 7163 5813
rect 7925 5810 7991 5813
rect 5901 5808 7991 5810
rect 5901 5752 5906 5808
rect 5962 5752 7102 5808
rect 7158 5752 7930 5808
rect 7986 5752 7991 5808
rect 5901 5750 7991 5752
rect 5901 5747 5967 5750
rect 7097 5747 7163 5750
rect 7925 5747 7991 5750
rect 17125 5810 17191 5813
rect 17953 5810 18019 5813
rect 17125 5808 18019 5810
rect 17125 5752 17130 5808
rect 17186 5752 17958 5808
rect 18014 5752 18019 5808
rect 17125 5750 18019 5752
rect 17125 5747 17191 5750
rect 17953 5747 18019 5750
rect 5441 5674 5507 5677
rect 9397 5674 9463 5677
rect 5441 5672 9463 5674
rect 5441 5616 5446 5672
rect 5502 5616 9402 5672
rect 9458 5616 9463 5672
rect 5441 5614 9463 5616
rect 5441 5611 5507 5614
rect 9397 5611 9463 5614
rect 16021 5674 16087 5677
rect 18505 5674 18571 5677
rect 16021 5672 18571 5674
rect 16021 5616 16026 5672
rect 16082 5616 18510 5672
rect 18566 5616 18571 5672
rect 16021 5614 18571 5616
rect 16021 5611 16087 5614
rect 18505 5611 18571 5614
rect 17534 5476 17540 5540
rect 17604 5538 17610 5540
rect 18045 5538 18111 5541
rect 17604 5536 18111 5538
rect 17604 5480 18050 5536
rect 18106 5480 18111 5536
rect 17604 5478 18111 5480
rect 17604 5476 17610 5478
rect 18045 5475 18111 5478
rect 3106 5472 3422 5473
rect 3106 5408 3112 5472
rect 3176 5408 3192 5472
rect 3256 5408 3272 5472
rect 3336 5408 3352 5472
rect 3416 5408 3422 5472
rect 3106 5407 3422 5408
rect 6206 5472 6522 5473
rect 6206 5408 6212 5472
rect 6276 5408 6292 5472
rect 6356 5408 6372 5472
rect 6436 5408 6452 5472
rect 6516 5408 6522 5472
rect 6206 5407 6522 5408
rect 9306 5472 9622 5473
rect 9306 5408 9312 5472
rect 9376 5408 9392 5472
rect 9456 5408 9472 5472
rect 9536 5408 9552 5472
rect 9616 5408 9622 5472
rect 9306 5407 9622 5408
rect 12406 5472 12722 5473
rect 12406 5408 12412 5472
rect 12476 5408 12492 5472
rect 12556 5408 12572 5472
rect 12636 5408 12652 5472
rect 12716 5408 12722 5472
rect 12406 5407 12722 5408
rect 15506 5472 15822 5473
rect 15506 5408 15512 5472
rect 15576 5408 15592 5472
rect 15656 5408 15672 5472
rect 15736 5408 15752 5472
rect 15816 5408 15822 5472
rect 15506 5407 15822 5408
rect 18606 5472 18922 5473
rect 18606 5408 18612 5472
rect 18676 5408 18692 5472
rect 18756 5408 18772 5472
rect 18836 5408 18852 5472
rect 18916 5408 18922 5472
rect 18606 5407 18922 5408
rect 13537 5266 13603 5269
rect 14917 5266 14983 5269
rect 15561 5266 15627 5269
rect 16062 5266 16068 5268
rect 13537 5264 16068 5266
rect 13537 5208 13542 5264
rect 13598 5208 14922 5264
rect 14978 5208 15566 5264
rect 15622 5208 16068 5264
rect 13537 5206 16068 5208
rect 13537 5203 13603 5206
rect 14917 5203 14983 5206
rect 15561 5203 15627 5206
rect 16062 5204 16068 5206
rect 16132 5204 16138 5268
rect 16665 5266 16731 5269
rect 16798 5266 16804 5268
rect 16665 5264 16804 5266
rect 16665 5208 16670 5264
rect 16726 5208 16804 5264
rect 16665 5206 16804 5208
rect 16665 5203 16731 5206
rect 16798 5204 16804 5206
rect 16868 5204 16874 5268
rect 17217 5266 17283 5269
rect 17861 5266 17927 5269
rect 17217 5264 17927 5266
rect 17217 5208 17222 5264
rect 17278 5208 17866 5264
rect 17922 5208 17927 5264
rect 17217 5206 17927 5208
rect 17217 5203 17283 5206
rect 17861 5203 17927 5206
rect 18965 5266 19031 5269
rect 19200 5266 20000 5296
rect 18965 5264 20000 5266
rect 18965 5208 18970 5264
rect 19026 5208 20000 5264
rect 18965 5206 20000 5208
rect 18965 5203 19031 5206
rect 19200 5176 20000 5206
rect 4656 4928 4972 4929
rect 4656 4864 4662 4928
rect 4726 4864 4742 4928
rect 4806 4864 4822 4928
rect 4886 4864 4902 4928
rect 4966 4864 4972 4928
rect 4656 4863 4972 4864
rect 7756 4928 8072 4929
rect 7756 4864 7762 4928
rect 7826 4864 7842 4928
rect 7906 4864 7922 4928
rect 7986 4864 8002 4928
rect 8066 4864 8072 4928
rect 7756 4863 8072 4864
rect 10856 4928 11172 4929
rect 10856 4864 10862 4928
rect 10926 4864 10942 4928
rect 11006 4864 11022 4928
rect 11086 4864 11102 4928
rect 11166 4864 11172 4928
rect 10856 4863 11172 4864
rect 13956 4928 14272 4929
rect 13956 4864 13962 4928
rect 14026 4864 14042 4928
rect 14106 4864 14122 4928
rect 14186 4864 14202 4928
rect 14266 4864 14272 4928
rect 13956 4863 14272 4864
rect 17056 4928 17372 4929
rect 17056 4864 17062 4928
rect 17126 4864 17142 4928
rect 17206 4864 17222 4928
rect 17286 4864 17302 4928
rect 17366 4864 17372 4928
rect 17056 4863 17372 4864
rect 5901 4858 5967 4861
rect 6729 4858 6795 4861
rect 5901 4856 6795 4858
rect 5901 4800 5906 4856
rect 5962 4800 6734 4856
rect 6790 4800 6795 4856
rect 5901 4798 6795 4800
rect 5901 4795 5967 4798
rect 6729 4795 6795 4798
rect 15101 4858 15167 4861
rect 16113 4858 16179 4861
rect 15101 4856 16179 4858
rect 15101 4800 15106 4856
rect 15162 4800 16118 4856
rect 16174 4800 16179 4856
rect 15101 4798 16179 4800
rect 15101 4795 15167 4798
rect 16113 4795 16179 4798
rect 4337 4722 4403 4725
rect 6085 4722 6151 4725
rect 4337 4720 6151 4722
rect 4337 4664 4342 4720
rect 4398 4664 6090 4720
rect 6146 4664 6151 4720
rect 4337 4662 6151 4664
rect 4337 4659 4403 4662
rect 6085 4659 6151 4662
rect 15745 4722 15811 4725
rect 16665 4722 16731 4725
rect 15745 4720 16731 4722
rect 15745 4664 15750 4720
rect 15806 4664 16670 4720
rect 16726 4664 16731 4720
rect 15745 4662 16731 4664
rect 15745 4659 15811 4662
rect 16665 4659 16731 4662
rect 11329 4586 11395 4589
rect 12617 4586 12683 4589
rect 11329 4584 12683 4586
rect 11329 4528 11334 4584
rect 11390 4528 12622 4584
rect 12678 4528 12683 4584
rect 11329 4526 12683 4528
rect 11329 4523 11395 4526
rect 12617 4523 12683 4526
rect 14457 4586 14523 4589
rect 17493 4586 17559 4589
rect 14457 4584 17559 4586
rect 14457 4528 14462 4584
rect 14518 4528 17498 4584
rect 17554 4528 17559 4584
rect 14457 4526 17559 4528
rect 14457 4523 14523 4526
rect 17493 4523 17559 4526
rect 16246 4388 16252 4452
rect 16316 4450 16322 4452
rect 16389 4450 16455 4453
rect 17125 4450 17191 4453
rect 17309 4450 17375 4453
rect 16316 4448 17375 4450
rect 16316 4392 16394 4448
rect 16450 4392 17130 4448
rect 17186 4392 17314 4448
rect 17370 4392 17375 4448
rect 16316 4390 17375 4392
rect 16316 4388 16322 4390
rect 16389 4387 16455 4390
rect 17125 4387 17191 4390
rect 17309 4387 17375 4390
rect 3106 4384 3422 4385
rect 3106 4320 3112 4384
rect 3176 4320 3192 4384
rect 3256 4320 3272 4384
rect 3336 4320 3352 4384
rect 3416 4320 3422 4384
rect 3106 4319 3422 4320
rect 6206 4384 6522 4385
rect 6206 4320 6212 4384
rect 6276 4320 6292 4384
rect 6356 4320 6372 4384
rect 6436 4320 6452 4384
rect 6516 4320 6522 4384
rect 6206 4319 6522 4320
rect 9306 4384 9622 4385
rect 9306 4320 9312 4384
rect 9376 4320 9392 4384
rect 9456 4320 9472 4384
rect 9536 4320 9552 4384
rect 9616 4320 9622 4384
rect 9306 4319 9622 4320
rect 12406 4384 12722 4385
rect 12406 4320 12412 4384
rect 12476 4320 12492 4384
rect 12556 4320 12572 4384
rect 12636 4320 12652 4384
rect 12716 4320 12722 4384
rect 12406 4319 12722 4320
rect 15506 4384 15822 4385
rect 15506 4320 15512 4384
rect 15576 4320 15592 4384
rect 15656 4320 15672 4384
rect 15736 4320 15752 4384
rect 15816 4320 15822 4384
rect 15506 4319 15822 4320
rect 18606 4384 18922 4385
rect 18606 4320 18612 4384
rect 18676 4320 18692 4384
rect 18756 4320 18772 4384
rect 18836 4320 18852 4384
rect 18916 4320 18922 4384
rect 18606 4319 18922 4320
rect 6637 4314 6703 4317
rect 8201 4314 8267 4317
rect 6637 4312 8267 4314
rect 6637 4256 6642 4312
rect 6698 4256 8206 4312
rect 8262 4256 8267 4312
rect 6637 4254 8267 4256
rect 6637 4251 6703 4254
rect 8201 4251 8267 4254
rect 16389 4178 16455 4181
rect 18965 4178 19031 4181
rect 16389 4176 19031 4178
rect 16389 4120 16394 4176
rect 16450 4120 18970 4176
rect 19026 4120 19031 4176
rect 16389 4118 19031 4120
rect 16389 4115 16455 4118
rect 18965 4115 19031 4118
rect 6177 4042 6243 4045
rect 8017 4042 8083 4045
rect 15009 4042 15075 4045
rect 16573 4042 16639 4045
rect 6177 4040 8218 4042
rect 6177 3984 6182 4040
rect 6238 3984 8022 4040
rect 8078 3984 8218 4040
rect 6177 3982 8218 3984
rect 6177 3979 6243 3982
rect 8017 3979 8083 3982
rect 4656 3840 4972 3841
rect 4656 3776 4662 3840
rect 4726 3776 4742 3840
rect 4806 3776 4822 3840
rect 4886 3776 4902 3840
rect 4966 3776 4972 3840
rect 4656 3775 4972 3776
rect 7756 3840 8072 3841
rect 7756 3776 7762 3840
rect 7826 3776 7842 3840
rect 7906 3776 7922 3840
rect 7986 3776 8002 3840
rect 8066 3776 8072 3840
rect 7756 3775 8072 3776
rect 5901 3770 5967 3773
rect 7373 3770 7439 3773
rect 5901 3768 7439 3770
rect 5901 3712 5906 3768
rect 5962 3712 7378 3768
rect 7434 3712 7439 3768
rect 5901 3710 7439 3712
rect 5901 3707 5967 3710
rect 7373 3707 7439 3710
rect 8158 3637 8218 3982
rect 15009 4040 16639 4042
rect 15009 3984 15014 4040
rect 15070 3984 16578 4040
rect 16634 3984 16639 4040
rect 15009 3982 16639 3984
rect 15009 3979 15075 3982
rect 16573 3979 16639 3982
rect 10856 3840 11172 3841
rect 10856 3776 10862 3840
rect 10926 3776 10942 3840
rect 11006 3776 11022 3840
rect 11086 3776 11102 3840
rect 11166 3776 11172 3840
rect 10856 3775 11172 3776
rect 13956 3840 14272 3841
rect 13956 3776 13962 3840
rect 14026 3776 14042 3840
rect 14106 3776 14122 3840
rect 14186 3776 14202 3840
rect 14266 3776 14272 3840
rect 13956 3775 14272 3776
rect 17056 3840 17372 3841
rect 17056 3776 17062 3840
rect 17126 3776 17142 3840
rect 17206 3776 17222 3840
rect 17286 3776 17302 3840
rect 17366 3776 17372 3840
rect 17056 3775 17372 3776
rect 12801 3770 12867 3773
rect 13721 3770 13787 3773
rect 12801 3768 13787 3770
rect 12801 3712 12806 3768
rect 12862 3712 13726 3768
rect 13782 3712 13787 3768
rect 12801 3710 13787 3712
rect 12801 3707 12867 3710
rect 13721 3707 13787 3710
rect 18965 3770 19031 3773
rect 19200 3770 20000 3800
rect 18965 3768 20000 3770
rect 18965 3712 18970 3768
rect 19026 3712 20000 3768
rect 18965 3710 20000 3712
rect 18965 3707 19031 3710
rect 19200 3680 20000 3710
rect 5625 3634 5691 3637
rect 7833 3634 7899 3637
rect 5625 3632 7899 3634
rect 5625 3576 5630 3632
rect 5686 3576 7838 3632
rect 7894 3576 7899 3632
rect 5625 3574 7899 3576
rect 5625 3571 5691 3574
rect 7833 3571 7899 3574
rect 8109 3632 8218 3637
rect 8109 3576 8114 3632
rect 8170 3576 8218 3632
rect 8109 3574 8218 3576
rect 11881 3634 11947 3637
rect 17309 3634 17375 3637
rect 11881 3632 17375 3634
rect 11881 3576 11886 3632
rect 11942 3576 17314 3632
rect 17370 3576 17375 3632
rect 11881 3574 17375 3576
rect 8109 3571 8175 3574
rect 11881 3571 11947 3574
rect 17309 3571 17375 3574
rect 4797 3498 4863 3501
rect 8937 3498 9003 3501
rect 4797 3496 9003 3498
rect 4797 3440 4802 3496
rect 4858 3440 8942 3496
rect 8998 3440 9003 3496
rect 4797 3438 9003 3440
rect 4797 3435 4863 3438
rect 8937 3435 9003 3438
rect 13169 3498 13235 3501
rect 18229 3498 18295 3501
rect 13169 3496 18295 3498
rect 13169 3440 13174 3496
rect 13230 3440 18234 3496
rect 18290 3440 18295 3496
rect 13169 3438 18295 3440
rect 13169 3435 13235 3438
rect 18229 3435 18295 3438
rect 6821 3362 6887 3365
rect 7925 3362 7991 3365
rect 6821 3360 7991 3362
rect 6821 3304 6826 3360
rect 6882 3304 7930 3360
rect 7986 3304 7991 3360
rect 6821 3302 7991 3304
rect 6821 3299 6887 3302
rect 7925 3299 7991 3302
rect 13813 3362 13879 3365
rect 14733 3362 14799 3365
rect 13813 3360 14799 3362
rect 13813 3304 13818 3360
rect 13874 3304 14738 3360
rect 14794 3304 14799 3360
rect 13813 3302 14799 3304
rect 13813 3299 13879 3302
rect 14733 3299 14799 3302
rect 16297 3362 16363 3365
rect 16430 3362 16436 3364
rect 16297 3360 16436 3362
rect 16297 3304 16302 3360
rect 16358 3304 16436 3360
rect 16297 3302 16436 3304
rect 16297 3299 16363 3302
rect 16430 3300 16436 3302
rect 16500 3300 16506 3364
rect 16941 3362 17007 3365
rect 17493 3362 17559 3365
rect 16941 3360 17559 3362
rect 16941 3304 16946 3360
rect 17002 3304 17498 3360
rect 17554 3304 17559 3360
rect 16941 3302 17559 3304
rect 16941 3299 17007 3302
rect 17493 3299 17559 3302
rect 17677 3362 17743 3365
rect 17677 3360 17786 3362
rect 17677 3304 17682 3360
rect 17738 3304 17786 3360
rect 17677 3299 17786 3304
rect 3106 3296 3422 3297
rect 3106 3232 3112 3296
rect 3176 3232 3192 3296
rect 3256 3232 3272 3296
rect 3336 3232 3352 3296
rect 3416 3232 3422 3296
rect 3106 3231 3422 3232
rect 6206 3296 6522 3297
rect 6206 3232 6212 3296
rect 6276 3232 6292 3296
rect 6356 3232 6372 3296
rect 6436 3232 6452 3296
rect 6516 3232 6522 3296
rect 6206 3231 6522 3232
rect 9306 3296 9622 3297
rect 9306 3232 9312 3296
rect 9376 3232 9392 3296
rect 9456 3232 9472 3296
rect 9536 3232 9552 3296
rect 9616 3232 9622 3296
rect 9306 3231 9622 3232
rect 12406 3296 12722 3297
rect 12406 3232 12412 3296
rect 12476 3232 12492 3296
rect 12556 3232 12572 3296
rect 12636 3232 12652 3296
rect 12716 3232 12722 3296
rect 12406 3231 12722 3232
rect 15506 3296 15822 3297
rect 15506 3232 15512 3296
rect 15576 3232 15592 3296
rect 15656 3232 15672 3296
rect 15736 3232 15752 3296
rect 15816 3232 15822 3296
rect 15506 3231 15822 3232
rect 7373 3226 7439 3229
rect 8109 3226 8175 3229
rect 7373 3224 8175 3226
rect 7373 3168 7378 3224
rect 7434 3168 8114 3224
rect 8170 3168 8175 3224
rect 7373 3166 8175 3168
rect 7373 3163 7439 3166
rect 8109 3163 8175 3166
rect 13445 3226 13511 3229
rect 14181 3226 14247 3229
rect 13445 3224 14247 3226
rect 13445 3168 13450 3224
rect 13506 3168 14186 3224
rect 14242 3168 14247 3224
rect 13445 3166 14247 3168
rect 13445 3163 13511 3166
rect 14181 3163 14247 3166
rect 17726 3093 17786 3299
rect 18606 3296 18922 3297
rect 18606 3232 18612 3296
rect 18676 3232 18692 3296
rect 18756 3232 18772 3296
rect 18836 3232 18852 3296
rect 18916 3232 18922 3296
rect 18606 3231 18922 3232
rect 6177 3090 6243 3093
rect 8109 3090 8175 3093
rect 6177 3088 8175 3090
rect 6177 3032 6182 3088
rect 6238 3032 8114 3088
rect 8170 3032 8175 3088
rect 6177 3030 8175 3032
rect 6177 3027 6243 3030
rect 8109 3027 8175 3030
rect 8385 3090 8451 3093
rect 11237 3090 11303 3093
rect 8385 3088 11303 3090
rect 8385 3032 8390 3088
rect 8446 3032 11242 3088
rect 11298 3032 11303 3088
rect 8385 3030 11303 3032
rect 8385 3027 8451 3030
rect 11237 3027 11303 3030
rect 17217 3088 17283 3093
rect 17217 3032 17222 3088
rect 17278 3032 17283 3088
rect 17217 3027 17283 3032
rect 17677 3088 17786 3093
rect 17677 3032 17682 3088
rect 17738 3032 17786 3088
rect 17677 3030 17786 3032
rect 17677 3027 17743 3030
rect 6729 2954 6795 2957
rect 8845 2954 8911 2957
rect 6729 2952 8911 2954
rect 6729 2896 6734 2952
rect 6790 2896 8850 2952
rect 8906 2896 8911 2952
rect 6729 2894 8911 2896
rect 6729 2891 6795 2894
rect 8845 2891 8911 2894
rect 12709 2954 12775 2957
rect 13261 2954 13327 2957
rect 12709 2952 13327 2954
rect 12709 2896 12714 2952
rect 12770 2896 13266 2952
rect 13322 2896 13327 2952
rect 12709 2894 13327 2896
rect 17220 2954 17280 3027
rect 18045 2954 18111 2957
rect 17220 2952 18111 2954
rect 17220 2896 18050 2952
rect 18106 2896 18111 2952
rect 17220 2894 18111 2896
rect 12709 2891 12775 2894
rect 13261 2891 13327 2894
rect 18045 2891 18111 2894
rect 16614 2756 16620 2820
rect 16684 2818 16690 2820
rect 16757 2818 16823 2821
rect 16684 2816 16823 2818
rect 16684 2760 16762 2816
rect 16818 2760 16823 2816
rect 16684 2758 16823 2760
rect 16684 2756 16690 2758
rect 16757 2755 16823 2758
rect 4656 2752 4972 2753
rect 4656 2688 4662 2752
rect 4726 2688 4742 2752
rect 4806 2688 4822 2752
rect 4886 2688 4902 2752
rect 4966 2688 4972 2752
rect 4656 2687 4972 2688
rect 7756 2752 8072 2753
rect 7756 2688 7762 2752
rect 7826 2688 7842 2752
rect 7906 2688 7922 2752
rect 7986 2688 8002 2752
rect 8066 2688 8072 2752
rect 7756 2687 8072 2688
rect 10856 2752 11172 2753
rect 10856 2688 10862 2752
rect 10926 2688 10942 2752
rect 11006 2688 11022 2752
rect 11086 2688 11102 2752
rect 11166 2688 11172 2752
rect 10856 2687 11172 2688
rect 13956 2752 14272 2753
rect 13956 2688 13962 2752
rect 14026 2688 14042 2752
rect 14106 2688 14122 2752
rect 14186 2688 14202 2752
rect 14266 2688 14272 2752
rect 13956 2687 14272 2688
rect 17056 2752 17372 2753
rect 17056 2688 17062 2752
rect 17126 2688 17142 2752
rect 17206 2688 17222 2752
rect 17286 2688 17302 2752
rect 17366 2688 17372 2752
rect 17056 2687 17372 2688
rect 6821 2682 6887 2685
rect 7281 2682 7347 2685
rect 6821 2680 7347 2682
rect 6821 2624 6826 2680
rect 6882 2624 7286 2680
rect 7342 2624 7347 2680
rect 6821 2622 7347 2624
rect 6821 2619 6887 2622
rect 7281 2619 7347 2622
rect 8477 2682 8543 2685
rect 8937 2682 9003 2685
rect 16573 2684 16639 2685
rect 16573 2682 16620 2684
rect 8477 2680 9003 2682
rect 8477 2624 8482 2680
rect 8538 2624 8942 2680
rect 8998 2624 9003 2680
rect 8477 2622 9003 2624
rect 16528 2680 16620 2682
rect 16528 2624 16578 2680
rect 16528 2622 16620 2624
rect 8477 2619 8543 2622
rect 8937 2619 9003 2622
rect 16573 2620 16620 2622
rect 16684 2620 16690 2684
rect 16573 2619 16639 2620
rect 5349 2546 5415 2549
rect 8109 2546 8175 2549
rect 5349 2544 8175 2546
rect 5349 2488 5354 2544
rect 5410 2488 8114 2544
rect 8170 2488 8175 2544
rect 5349 2486 8175 2488
rect 5349 2483 5415 2486
rect 8109 2483 8175 2486
rect 11237 2546 11303 2549
rect 13905 2546 13971 2549
rect 11237 2544 13971 2546
rect 11237 2488 11242 2544
rect 11298 2488 13910 2544
rect 13966 2488 13971 2544
rect 11237 2486 13971 2488
rect 11237 2483 11303 2486
rect 13905 2483 13971 2486
rect 14181 2546 14247 2549
rect 14406 2546 14412 2548
rect 14181 2544 14412 2546
rect 14181 2488 14186 2544
rect 14242 2488 14412 2544
rect 14181 2486 14412 2488
rect 14181 2483 14247 2486
rect 14406 2484 14412 2486
rect 14476 2546 14482 2548
rect 15837 2546 15903 2549
rect 14476 2544 15903 2546
rect 14476 2488 15842 2544
rect 15898 2488 15903 2544
rect 14476 2486 15903 2488
rect 14476 2484 14482 2486
rect 15837 2483 15903 2486
rect 15193 2410 15259 2413
rect 16389 2410 16455 2413
rect 15193 2408 16455 2410
rect 15193 2352 15198 2408
rect 15254 2352 16394 2408
rect 16450 2352 16455 2408
rect 15193 2350 16455 2352
rect 15193 2347 15259 2350
rect 16389 2347 16455 2350
rect 16849 2410 16915 2413
rect 17769 2410 17835 2413
rect 16849 2408 17835 2410
rect 16849 2352 16854 2408
rect 16910 2352 17774 2408
rect 17830 2352 17835 2408
rect 16849 2350 17835 2352
rect 16849 2347 16915 2350
rect 17769 2347 17835 2350
rect 16852 2274 16912 2347
rect 15886 2214 16912 2274
rect 19057 2274 19123 2277
rect 19200 2274 20000 2304
rect 19057 2272 20000 2274
rect 19057 2216 19062 2272
rect 19118 2216 20000 2272
rect 19057 2214 20000 2216
rect 3106 2208 3422 2209
rect 3106 2144 3112 2208
rect 3176 2144 3192 2208
rect 3256 2144 3272 2208
rect 3336 2144 3352 2208
rect 3416 2144 3422 2208
rect 3106 2143 3422 2144
rect 6206 2208 6522 2209
rect 6206 2144 6212 2208
rect 6276 2144 6292 2208
rect 6356 2144 6372 2208
rect 6436 2144 6452 2208
rect 6516 2144 6522 2208
rect 6206 2143 6522 2144
rect 9306 2208 9622 2209
rect 9306 2144 9312 2208
rect 9376 2144 9392 2208
rect 9456 2144 9472 2208
rect 9536 2144 9552 2208
rect 9616 2144 9622 2208
rect 9306 2143 9622 2144
rect 12406 2208 12722 2209
rect 12406 2144 12412 2208
rect 12476 2144 12492 2208
rect 12556 2144 12572 2208
rect 12636 2144 12652 2208
rect 12716 2144 12722 2208
rect 12406 2143 12722 2144
rect 15506 2208 15822 2209
rect 15506 2144 15512 2208
rect 15576 2144 15592 2208
rect 15656 2144 15672 2208
rect 15736 2144 15752 2208
rect 15816 2144 15822 2208
rect 15506 2143 15822 2144
rect 8845 2002 8911 2005
rect 9581 2002 9647 2005
rect 8845 2000 9647 2002
rect 8845 1944 8850 2000
rect 8906 1944 9586 2000
rect 9642 1944 9647 2000
rect 8845 1942 9647 1944
rect 8845 1939 8911 1942
rect 9581 1939 9647 1942
rect 13353 2002 13419 2005
rect 14733 2002 14799 2005
rect 15009 2002 15075 2005
rect 15886 2002 15946 2214
rect 19057 2211 19123 2214
rect 18606 2208 18922 2209
rect 18606 2144 18612 2208
rect 18676 2144 18692 2208
rect 18756 2144 18772 2208
rect 18836 2144 18852 2208
rect 18916 2144 18922 2208
rect 19200 2184 20000 2214
rect 18606 2143 18922 2144
rect 16297 2138 16363 2141
rect 17953 2138 18019 2141
rect 16297 2136 18019 2138
rect 16297 2080 16302 2136
rect 16358 2080 17958 2136
rect 18014 2080 18019 2136
rect 16297 2078 18019 2080
rect 16297 2075 16363 2078
rect 17953 2075 18019 2078
rect 16297 2004 16363 2005
rect 16246 2002 16252 2004
rect 13353 2000 15946 2002
rect 13353 1944 13358 2000
rect 13414 1944 14738 2000
rect 14794 1944 15014 2000
rect 15070 1944 15946 2000
rect 13353 1942 15946 1944
rect 16206 1942 16252 2002
rect 16316 2000 16363 2004
rect 17861 2002 17927 2005
rect 18505 2002 18571 2005
rect 16358 1944 16363 2000
rect 13353 1939 13419 1942
rect 14733 1939 14799 1942
rect 15009 1939 15075 1942
rect 16246 1940 16252 1942
rect 16316 1940 16363 1944
rect 16297 1939 16363 1940
rect 16622 2000 18571 2002
rect 16622 1944 17866 2000
rect 17922 1944 18510 2000
rect 18566 1944 18571 2000
rect 16622 1942 18571 1944
rect 12065 1866 12131 1869
rect 15469 1866 15535 1869
rect 12065 1864 15535 1866
rect 12065 1808 12070 1864
rect 12126 1808 15474 1864
rect 15530 1808 15535 1864
rect 12065 1806 15535 1808
rect 12065 1803 12131 1806
rect 15469 1803 15535 1806
rect 15653 1866 15719 1869
rect 16622 1866 16682 1942
rect 17861 1939 17927 1942
rect 18505 1939 18571 1942
rect 15653 1864 16682 1866
rect 15653 1808 15658 1864
rect 15714 1808 16682 1864
rect 15653 1806 16682 1808
rect 15653 1803 15719 1806
rect 4656 1664 4972 1665
rect 4656 1600 4662 1664
rect 4726 1600 4742 1664
rect 4806 1600 4822 1664
rect 4886 1600 4902 1664
rect 4966 1600 4972 1664
rect 4656 1599 4972 1600
rect 7756 1664 8072 1665
rect 7756 1600 7762 1664
rect 7826 1600 7842 1664
rect 7906 1600 7922 1664
rect 7986 1600 8002 1664
rect 8066 1600 8072 1664
rect 7756 1599 8072 1600
rect 10856 1664 11172 1665
rect 10856 1600 10862 1664
rect 10926 1600 10942 1664
rect 11006 1600 11022 1664
rect 11086 1600 11102 1664
rect 11166 1600 11172 1664
rect 10856 1599 11172 1600
rect 13956 1664 14272 1665
rect 13956 1600 13962 1664
rect 14026 1600 14042 1664
rect 14106 1600 14122 1664
rect 14186 1600 14202 1664
rect 14266 1600 14272 1664
rect 13956 1599 14272 1600
rect 17056 1664 17372 1665
rect 17056 1600 17062 1664
rect 17126 1600 17142 1664
rect 17206 1600 17222 1664
rect 17286 1600 17302 1664
rect 17366 1600 17372 1664
rect 17056 1599 17372 1600
rect 14089 1458 14155 1461
rect 18045 1458 18111 1461
rect 14089 1456 18111 1458
rect 14089 1400 14094 1456
rect 14150 1400 18050 1456
rect 18106 1400 18111 1456
rect 14089 1398 18111 1400
rect 14089 1395 14155 1398
rect 18045 1395 18111 1398
rect 17401 1322 17467 1325
rect 17534 1322 17540 1324
rect 17401 1320 17540 1322
rect 17401 1264 17406 1320
rect 17462 1264 17540 1320
rect 17401 1262 17540 1264
rect 17401 1259 17467 1262
rect 17534 1260 17540 1262
rect 17604 1260 17610 1324
rect 3106 1120 3422 1121
rect 3106 1056 3112 1120
rect 3176 1056 3192 1120
rect 3256 1056 3272 1120
rect 3336 1056 3352 1120
rect 3416 1056 3422 1120
rect 3106 1055 3422 1056
rect 6206 1120 6522 1121
rect 6206 1056 6212 1120
rect 6276 1056 6292 1120
rect 6356 1056 6372 1120
rect 6436 1056 6452 1120
rect 6516 1056 6522 1120
rect 6206 1055 6522 1056
rect 9306 1120 9622 1121
rect 9306 1056 9312 1120
rect 9376 1056 9392 1120
rect 9456 1056 9472 1120
rect 9536 1056 9552 1120
rect 9616 1056 9622 1120
rect 9306 1055 9622 1056
rect 12406 1120 12722 1121
rect 12406 1056 12412 1120
rect 12476 1056 12492 1120
rect 12556 1056 12572 1120
rect 12636 1056 12652 1120
rect 12716 1056 12722 1120
rect 12406 1055 12722 1056
rect 15506 1120 15822 1121
rect 15506 1056 15512 1120
rect 15576 1056 15592 1120
rect 15656 1056 15672 1120
rect 15736 1056 15752 1120
rect 15816 1056 15822 1120
rect 15506 1055 15822 1056
rect 18606 1120 18922 1121
rect 18606 1056 18612 1120
rect 18676 1056 18692 1120
rect 18756 1056 18772 1120
rect 18836 1056 18852 1120
rect 18916 1056 18922 1120
rect 18606 1055 18922 1056
rect 13261 1050 13327 1053
rect 14273 1050 14339 1053
rect 14406 1050 14412 1052
rect 13261 1048 14412 1050
rect 13261 992 13266 1048
rect 13322 992 14278 1048
rect 14334 992 14412 1048
rect 13261 990 14412 992
rect 13261 987 13327 990
rect 14273 987 14339 990
rect 14406 988 14412 990
rect 14476 988 14482 1052
rect 13261 914 13327 917
rect 15837 914 15903 917
rect 13261 912 15903 914
rect 13261 856 13266 912
rect 13322 856 15842 912
rect 15898 856 15903 912
rect 13261 854 15903 856
rect 13261 851 13327 854
rect 15837 851 15903 854
rect 12801 778 12867 781
rect 14273 778 14339 781
rect 12801 776 14339 778
rect 12801 720 12806 776
rect 12862 720 14278 776
rect 14334 720 14339 776
rect 12801 718 14339 720
rect 12801 715 12867 718
rect 14273 715 14339 718
rect 17861 778 17927 781
rect 19200 778 20000 808
rect 17861 776 20000 778
rect 17861 720 17866 776
rect 17922 720 20000 776
rect 17861 718 20000 720
rect 17861 715 17927 718
rect 19200 688 20000 718
rect 4656 576 4972 577
rect 4656 512 4662 576
rect 4726 512 4742 576
rect 4806 512 4822 576
rect 4886 512 4902 576
rect 4966 512 4972 576
rect 4656 511 4972 512
rect 7756 576 8072 577
rect 7756 512 7762 576
rect 7826 512 7842 576
rect 7906 512 7922 576
rect 7986 512 8002 576
rect 8066 512 8072 576
rect 7756 511 8072 512
rect 10856 576 11172 577
rect 10856 512 10862 576
rect 10926 512 10942 576
rect 11006 512 11022 576
rect 11086 512 11102 576
rect 11166 512 11172 576
rect 10856 511 11172 512
rect 13956 576 14272 577
rect 13956 512 13962 576
rect 14026 512 14042 576
rect 14106 512 14122 576
rect 14186 512 14202 576
rect 14266 512 14272 576
rect 13956 511 14272 512
rect 17056 576 17372 577
rect 17056 512 17062 576
rect 17126 512 17142 576
rect 17206 512 17222 576
rect 17286 512 17302 576
rect 17366 512 17372 576
rect 17056 511 17372 512
<< via3 >>
rect 3112 10908 3176 10912
rect 3112 10852 3116 10908
rect 3116 10852 3172 10908
rect 3172 10852 3176 10908
rect 3112 10848 3176 10852
rect 3192 10908 3256 10912
rect 3192 10852 3196 10908
rect 3196 10852 3252 10908
rect 3252 10852 3256 10908
rect 3192 10848 3256 10852
rect 3272 10908 3336 10912
rect 3272 10852 3276 10908
rect 3276 10852 3332 10908
rect 3332 10852 3336 10908
rect 3272 10848 3336 10852
rect 3352 10908 3416 10912
rect 3352 10852 3356 10908
rect 3356 10852 3412 10908
rect 3412 10852 3416 10908
rect 3352 10848 3416 10852
rect 6212 10908 6276 10912
rect 6212 10852 6216 10908
rect 6216 10852 6272 10908
rect 6272 10852 6276 10908
rect 6212 10848 6276 10852
rect 6292 10908 6356 10912
rect 6292 10852 6296 10908
rect 6296 10852 6352 10908
rect 6352 10852 6356 10908
rect 6292 10848 6356 10852
rect 6372 10908 6436 10912
rect 6372 10852 6376 10908
rect 6376 10852 6432 10908
rect 6432 10852 6436 10908
rect 6372 10848 6436 10852
rect 6452 10908 6516 10912
rect 6452 10852 6456 10908
rect 6456 10852 6512 10908
rect 6512 10852 6516 10908
rect 6452 10848 6516 10852
rect 9312 10908 9376 10912
rect 9312 10852 9316 10908
rect 9316 10852 9372 10908
rect 9372 10852 9376 10908
rect 9312 10848 9376 10852
rect 9392 10908 9456 10912
rect 9392 10852 9396 10908
rect 9396 10852 9452 10908
rect 9452 10852 9456 10908
rect 9392 10848 9456 10852
rect 9472 10908 9536 10912
rect 9472 10852 9476 10908
rect 9476 10852 9532 10908
rect 9532 10852 9536 10908
rect 9472 10848 9536 10852
rect 9552 10908 9616 10912
rect 9552 10852 9556 10908
rect 9556 10852 9612 10908
rect 9612 10852 9616 10908
rect 9552 10848 9616 10852
rect 12412 10908 12476 10912
rect 12412 10852 12416 10908
rect 12416 10852 12472 10908
rect 12472 10852 12476 10908
rect 12412 10848 12476 10852
rect 12492 10908 12556 10912
rect 12492 10852 12496 10908
rect 12496 10852 12552 10908
rect 12552 10852 12556 10908
rect 12492 10848 12556 10852
rect 12572 10908 12636 10912
rect 12572 10852 12576 10908
rect 12576 10852 12632 10908
rect 12632 10852 12636 10908
rect 12572 10848 12636 10852
rect 12652 10908 12716 10912
rect 12652 10852 12656 10908
rect 12656 10852 12712 10908
rect 12712 10852 12716 10908
rect 12652 10848 12716 10852
rect 15512 10908 15576 10912
rect 15512 10852 15516 10908
rect 15516 10852 15572 10908
rect 15572 10852 15576 10908
rect 15512 10848 15576 10852
rect 15592 10908 15656 10912
rect 15592 10852 15596 10908
rect 15596 10852 15652 10908
rect 15652 10852 15656 10908
rect 15592 10848 15656 10852
rect 15672 10908 15736 10912
rect 15672 10852 15676 10908
rect 15676 10852 15732 10908
rect 15732 10852 15736 10908
rect 15672 10848 15736 10852
rect 15752 10908 15816 10912
rect 15752 10852 15756 10908
rect 15756 10852 15812 10908
rect 15812 10852 15816 10908
rect 15752 10848 15816 10852
rect 18612 10908 18676 10912
rect 18612 10852 18616 10908
rect 18616 10852 18672 10908
rect 18672 10852 18676 10908
rect 18612 10848 18676 10852
rect 18692 10908 18756 10912
rect 18692 10852 18696 10908
rect 18696 10852 18752 10908
rect 18752 10852 18756 10908
rect 18692 10848 18756 10852
rect 18772 10908 18836 10912
rect 18772 10852 18776 10908
rect 18776 10852 18832 10908
rect 18832 10852 18836 10908
rect 18772 10848 18836 10852
rect 18852 10908 18916 10912
rect 18852 10852 18856 10908
rect 18856 10852 18912 10908
rect 18912 10852 18916 10908
rect 18852 10848 18916 10852
rect 4662 10364 4726 10368
rect 4662 10308 4666 10364
rect 4666 10308 4722 10364
rect 4722 10308 4726 10364
rect 4662 10304 4726 10308
rect 4742 10364 4806 10368
rect 4742 10308 4746 10364
rect 4746 10308 4802 10364
rect 4802 10308 4806 10364
rect 4742 10304 4806 10308
rect 4822 10364 4886 10368
rect 4822 10308 4826 10364
rect 4826 10308 4882 10364
rect 4882 10308 4886 10364
rect 4822 10304 4886 10308
rect 4902 10364 4966 10368
rect 4902 10308 4906 10364
rect 4906 10308 4962 10364
rect 4962 10308 4966 10364
rect 4902 10304 4966 10308
rect 7762 10364 7826 10368
rect 7762 10308 7766 10364
rect 7766 10308 7822 10364
rect 7822 10308 7826 10364
rect 7762 10304 7826 10308
rect 7842 10364 7906 10368
rect 7842 10308 7846 10364
rect 7846 10308 7902 10364
rect 7902 10308 7906 10364
rect 7842 10304 7906 10308
rect 7922 10364 7986 10368
rect 7922 10308 7926 10364
rect 7926 10308 7982 10364
rect 7982 10308 7986 10364
rect 7922 10304 7986 10308
rect 8002 10364 8066 10368
rect 8002 10308 8006 10364
rect 8006 10308 8062 10364
rect 8062 10308 8066 10364
rect 8002 10304 8066 10308
rect 10862 10364 10926 10368
rect 10862 10308 10866 10364
rect 10866 10308 10922 10364
rect 10922 10308 10926 10364
rect 10862 10304 10926 10308
rect 10942 10364 11006 10368
rect 10942 10308 10946 10364
rect 10946 10308 11002 10364
rect 11002 10308 11006 10364
rect 10942 10304 11006 10308
rect 11022 10364 11086 10368
rect 11022 10308 11026 10364
rect 11026 10308 11082 10364
rect 11082 10308 11086 10364
rect 11022 10304 11086 10308
rect 11102 10364 11166 10368
rect 11102 10308 11106 10364
rect 11106 10308 11162 10364
rect 11162 10308 11166 10364
rect 11102 10304 11166 10308
rect 13962 10364 14026 10368
rect 13962 10308 13966 10364
rect 13966 10308 14022 10364
rect 14022 10308 14026 10364
rect 13962 10304 14026 10308
rect 14042 10364 14106 10368
rect 14042 10308 14046 10364
rect 14046 10308 14102 10364
rect 14102 10308 14106 10364
rect 14042 10304 14106 10308
rect 14122 10364 14186 10368
rect 14122 10308 14126 10364
rect 14126 10308 14182 10364
rect 14182 10308 14186 10364
rect 14122 10304 14186 10308
rect 14202 10364 14266 10368
rect 14202 10308 14206 10364
rect 14206 10308 14262 10364
rect 14262 10308 14266 10364
rect 14202 10304 14266 10308
rect 17062 10364 17126 10368
rect 17062 10308 17066 10364
rect 17066 10308 17122 10364
rect 17122 10308 17126 10364
rect 17062 10304 17126 10308
rect 17142 10364 17206 10368
rect 17142 10308 17146 10364
rect 17146 10308 17202 10364
rect 17202 10308 17206 10364
rect 17142 10304 17206 10308
rect 17222 10364 17286 10368
rect 17222 10308 17226 10364
rect 17226 10308 17282 10364
rect 17282 10308 17286 10364
rect 17222 10304 17286 10308
rect 17302 10364 17366 10368
rect 17302 10308 17306 10364
rect 17306 10308 17362 10364
rect 17362 10308 17366 10364
rect 17302 10304 17366 10308
rect 3112 9820 3176 9824
rect 3112 9764 3116 9820
rect 3116 9764 3172 9820
rect 3172 9764 3176 9820
rect 3112 9760 3176 9764
rect 3192 9820 3256 9824
rect 3192 9764 3196 9820
rect 3196 9764 3252 9820
rect 3252 9764 3256 9820
rect 3192 9760 3256 9764
rect 3272 9820 3336 9824
rect 3272 9764 3276 9820
rect 3276 9764 3332 9820
rect 3332 9764 3336 9820
rect 3272 9760 3336 9764
rect 3352 9820 3416 9824
rect 3352 9764 3356 9820
rect 3356 9764 3412 9820
rect 3412 9764 3416 9820
rect 3352 9760 3416 9764
rect 6212 9820 6276 9824
rect 6212 9764 6216 9820
rect 6216 9764 6272 9820
rect 6272 9764 6276 9820
rect 6212 9760 6276 9764
rect 6292 9820 6356 9824
rect 6292 9764 6296 9820
rect 6296 9764 6352 9820
rect 6352 9764 6356 9820
rect 6292 9760 6356 9764
rect 6372 9820 6436 9824
rect 6372 9764 6376 9820
rect 6376 9764 6432 9820
rect 6432 9764 6436 9820
rect 6372 9760 6436 9764
rect 6452 9820 6516 9824
rect 6452 9764 6456 9820
rect 6456 9764 6512 9820
rect 6512 9764 6516 9820
rect 6452 9760 6516 9764
rect 9312 9820 9376 9824
rect 9312 9764 9316 9820
rect 9316 9764 9372 9820
rect 9372 9764 9376 9820
rect 9312 9760 9376 9764
rect 9392 9820 9456 9824
rect 9392 9764 9396 9820
rect 9396 9764 9452 9820
rect 9452 9764 9456 9820
rect 9392 9760 9456 9764
rect 9472 9820 9536 9824
rect 9472 9764 9476 9820
rect 9476 9764 9532 9820
rect 9532 9764 9536 9820
rect 9472 9760 9536 9764
rect 9552 9820 9616 9824
rect 9552 9764 9556 9820
rect 9556 9764 9612 9820
rect 9612 9764 9616 9820
rect 9552 9760 9616 9764
rect 12412 9820 12476 9824
rect 12412 9764 12416 9820
rect 12416 9764 12472 9820
rect 12472 9764 12476 9820
rect 12412 9760 12476 9764
rect 12492 9820 12556 9824
rect 12492 9764 12496 9820
rect 12496 9764 12552 9820
rect 12552 9764 12556 9820
rect 12492 9760 12556 9764
rect 12572 9820 12636 9824
rect 12572 9764 12576 9820
rect 12576 9764 12632 9820
rect 12632 9764 12636 9820
rect 12572 9760 12636 9764
rect 12652 9820 12716 9824
rect 12652 9764 12656 9820
rect 12656 9764 12712 9820
rect 12712 9764 12716 9820
rect 12652 9760 12716 9764
rect 15512 9820 15576 9824
rect 15512 9764 15516 9820
rect 15516 9764 15572 9820
rect 15572 9764 15576 9820
rect 15512 9760 15576 9764
rect 15592 9820 15656 9824
rect 15592 9764 15596 9820
rect 15596 9764 15652 9820
rect 15652 9764 15656 9820
rect 15592 9760 15656 9764
rect 15672 9820 15736 9824
rect 15672 9764 15676 9820
rect 15676 9764 15732 9820
rect 15732 9764 15736 9820
rect 15672 9760 15736 9764
rect 15752 9820 15816 9824
rect 15752 9764 15756 9820
rect 15756 9764 15812 9820
rect 15812 9764 15816 9820
rect 15752 9760 15816 9764
rect 18612 9820 18676 9824
rect 18612 9764 18616 9820
rect 18616 9764 18672 9820
rect 18672 9764 18676 9820
rect 18612 9760 18676 9764
rect 18692 9820 18756 9824
rect 18692 9764 18696 9820
rect 18696 9764 18752 9820
rect 18752 9764 18756 9820
rect 18692 9760 18756 9764
rect 18772 9820 18836 9824
rect 18772 9764 18776 9820
rect 18776 9764 18832 9820
rect 18832 9764 18836 9820
rect 18772 9760 18836 9764
rect 18852 9820 18916 9824
rect 18852 9764 18856 9820
rect 18856 9764 18912 9820
rect 18912 9764 18916 9820
rect 18852 9760 18916 9764
rect 4662 9276 4726 9280
rect 4662 9220 4666 9276
rect 4666 9220 4722 9276
rect 4722 9220 4726 9276
rect 4662 9216 4726 9220
rect 4742 9276 4806 9280
rect 4742 9220 4746 9276
rect 4746 9220 4802 9276
rect 4802 9220 4806 9276
rect 4742 9216 4806 9220
rect 4822 9276 4886 9280
rect 4822 9220 4826 9276
rect 4826 9220 4882 9276
rect 4882 9220 4886 9276
rect 4822 9216 4886 9220
rect 4902 9276 4966 9280
rect 4902 9220 4906 9276
rect 4906 9220 4962 9276
rect 4962 9220 4966 9276
rect 4902 9216 4966 9220
rect 7762 9276 7826 9280
rect 7762 9220 7766 9276
rect 7766 9220 7822 9276
rect 7822 9220 7826 9276
rect 7762 9216 7826 9220
rect 7842 9276 7906 9280
rect 7842 9220 7846 9276
rect 7846 9220 7902 9276
rect 7902 9220 7906 9276
rect 7842 9216 7906 9220
rect 7922 9276 7986 9280
rect 7922 9220 7926 9276
rect 7926 9220 7982 9276
rect 7982 9220 7986 9276
rect 7922 9216 7986 9220
rect 8002 9276 8066 9280
rect 8002 9220 8006 9276
rect 8006 9220 8062 9276
rect 8062 9220 8066 9276
rect 8002 9216 8066 9220
rect 10862 9276 10926 9280
rect 10862 9220 10866 9276
rect 10866 9220 10922 9276
rect 10922 9220 10926 9276
rect 10862 9216 10926 9220
rect 10942 9276 11006 9280
rect 10942 9220 10946 9276
rect 10946 9220 11002 9276
rect 11002 9220 11006 9276
rect 10942 9216 11006 9220
rect 11022 9276 11086 9280
rect 11022 9220 11026 9276
rect 11026 9220 11082 9276
rect 11082 9220 11086 9276
rect 11022 9216 11086 9220
rect 11102 9276 11166 9280
rect 11102 9220 11106 9276
rect 11106 9220 11162 9276
rect 11162 9220 11166 9276
rect 11102 9216 11166 9220
rect 13962 9276 14026 9280
rect 13962 9220 13966 9276
rect 13966 9220 14022 9276
rect 14022 9220 14026 9276
rect 13962 9216 14026 9220
rect 14042 9276 14106 9280
rect 14042 9220 14046 9276
rect 14046 9220 14102 9276
rect 14102 9220 14106 9276
rect 14042 9216 14106 9220
rect 14122 9276 14186 9280
rect 14122 9220 14126 9276
rect 14126 9220 14182 9276
rect 14182 9220 14186 9276
rect 14122 9216 14186 9220
rect 14202 9276 14266 9280
rect 14202 9220 14206 9276
rect 14206 9220 14262 9276
rect 14262 9220 14266 9276
rect 14202 9216 14266 9220
rect 17062 9276 17126 9280
rect 17062 9220 17066 9276
rect 17066 9220 17122 9276
rect 17122 9220 17126 9276
rect 17062 9216 17126 9220
rect 17142 9276 17206 9280
rect 17142 9220 17146 9276
rect 17146 9220 17202 9276
rect 17202 9220 17206 9276
rect 17142 9216 17206 9220
rect 17222 9276 17286 9280
rect 17222 9220 17226 9276
rect 17226 9220 17282 9276
rect 17282 9220 17286 9276
rect 17222 9216 17286 9220
rect 17302 9276 17366 9280
rect 17302 9220 17306 9276
rect 17306 9220 17362 9276
rect 17362 9220 17366 9276
rect 17302 9216 17366 9220
rect 3112 8732 3176 8736
rect 3112 8676 3116 8732
rect 3116 8676 3172 8732
rect 3172 8676 3176 8732
rect 3112 8672 3176 8676
rect 3192 8732 3256 8736
rect 3192 8676 3196 8732
rect 3196 8676 3252 8732
rect 3252 8676 3256 8732
rect 3192 8672 3256 8676
rect 3272 8732 3336 8736
rect 3272 8676 3276 8732
rect 3276 8676 3332 8732
rect 3332 8676 3336 8732
rect 3272 8672 3336 8676
rect 3352 8732 3416 8736
rect 3352 8676 3356 8732
rect 3356 8676 3412 8732
rect 3412 8676 3416 8732
rect 3352 8672 3416 8676
rect 6212 8732 6276 8736
rect 6212 8676 6216 8732
rect 6216 8676 6272 8732
rect 6272 8676 6276 8732
rect 6212 8672 6276 8676
rect 6292 8732 6356 8736
rect 6292 8676 6296 8732
rect 6296 8676 6352 8732
rect 6352 8676 6356 8732
rect 6292 8672 6356 8676
rect 6372 8732 6436 8736
rect 6372 8676 6376 8732
rect 6376 8676 6432 8732
rect 6432 8676 6436 8732
rect 6372 8672 6436 8676
rect 6452 8732 6516 8736
rect 6452 8676 6456 8732
rect 6456 8676 6512 8732
rect 6512 8676 6516 8732
rect 6452 8672 6516 8676
rect 9312 8732 9376 8736
rect 9312 8676 9316 8732
rect 9316 8676 9372 8732
rect 9372 8676 9376 8732
rect 9312 8672 9376 8676
rect 9392 8732 9456 8736
rect 9392 8676 9396 8732
rect 9396 8676 9452 8732
rect 9452 8676 9456 8732
rect 9392 8672 9456 8676
rect 9472 8732 9536 8736
rect 9472 8676 9476 8732
rect 9476 8676 9532 8732
rect 9532 8676 9536 8732
rect 9472 8672 9536 8676
rect 9552 8732 9616 8736
rect 9552 8676 9556 8732
rect 9556 8676 9612 8732
rect 9612 8676 9616 8732
rect 9552 8672 9616 8676
rect 12412 8732 12476 8736
rect 12412 8676 12416 8732
rect 12416 8676 12472 8732
rect 12472 8676 12476 8732
rect 12412 8672 12476 8676
rect 12492 8732 12556 8736
rect 12492 8676 12496 8732
rect 12496 8676 12552 8732
rect 12552 8676 12556 8732
rect 12492 8672 12556 8676
rect 12572 8732 12636 8736
rect 12572 8676 12576 8732
rect 12576 8676 12632 8732
rect 12632 8676 12636 8732
rect 12572 8672 12636 8676
rect 12652 8732 12716 8736
rect 12652 8676 12656 8732
rect 12656 8676 12712 8732
rect 12712 8676 12716 8732
rect 12652 8672 12716 8676
rect 15512 8732 15576 8736
rect 15512 8676 15516 8732
rect 15516 8676 15572 8732
rect 15572 8676 15576 8732
rect 15512 8672 15576 8676
rect 15592 8732 15656 8736
rect 15592 8676 15596 8732
rect 15596 8676 15652 8732
rect 15652 8676 15656 8732
rect 15592 8672 15656 8676
rect 15672 8732 15736 8736
rect 15672 8676 15676 8732
rect 15676 8676 15732 8732
rect 15732 8676 15736 8732
rect 15672 8672 15736 8676
rect 15752 8732 15816 8736
rect 15752 8676 15756 8732
rect 15756 8676 15812 8732
rect 15812 8676 15816 8732
rect 15752 8672 15816 8676
rect 18612 8732 18676 8736
rect 18612 8676 18616 8732
rect 18616 8676 18672 8732
rect 18672 8676 18676 8732
rect 18612 8672 18676 8676
rect 18692 8732 18756 8736
rect 18692 8676 18696 8732
rect 18696 8676 18752 8732
rect 18752 8676 18756 8732
rect 18692 8672 18756 8676
rect 18772 8732 18836 8736
rect 18772 8676 18776 8732
rect 18776 8676 18832 8732
rect 18832 8676 18836 8732
rect 18772 8672 18836 8676
rect 18852 8732 18916 8736
rect 18852 8676 18856 8732
rect 18856 8676 18912 8732
rect 18912 8676 18916 8732
rect 18852 8672 18916 8676
rect 16804 8468 16868 8532
rect 4662 8188 4726 8192
rect 4662 8132 4666 8188
rect 4666 8132 4722 8188
rect 4722 8132 4726 8188
rect 4662 8128 4726 8132
rect 4742 8188 4806 8192
rect 4742 8132 4746 8188
rect 4746 8132 4802 8188
rect 4802 8132 4806 8188
rect 4742 8128 4806 8132
rect 4822 8188 4886 8192
rect 4822 8132 4826 8188
rect 4826 8132 4882 8188
rect 4882 8132 4886 8188
rect 4822 8128 4886 8132
rect 4902 8188 4966 8192
rect 4902 8132 4906 8188
rect 4906 8132 4962 8188
rect 4962 8132 4966 8188
rect 4902 8128 4966 8132
rect 7762 8188 7826 8192
rect 7762 8132 7766 8188
rect 7766 8132 7822 8188
rect 7822 8132 7826 8188
rect 7762 8128 7826 8132
rect 7842 8188 7906 8192
rect 7842 8132 7846 8188
rect 7846 8132 7902 8188
rect 7902 8132 7906 8188
rect 7842 8128 7906 8132
rect 7922 8188 7986 8192
rect 7922 8132 7926 8188
rect 7926 8132 7982 8188
rect 7982 8132 7986 8188
rect 7922 8128 7986 8132
rect 8002 8188 8066 8192
rect 8002 8132 8006 8188
rect 8006 8132 8062 8188
rect 8062 8132 8066 8188
rect 8002 8128 8066 8132
rect 10862 8188 10926 8192
rect 10862 8132 10866 8188
rect 10866 8132 10922 8188
rect 10922 8132 10926 8188
rect 10862 8128 10926 8132
rect 10942 8188 11006 8192
rect 10942 8132 10946 8188
rect 10946 8132 11002 8188
rect 11002 8132 11006 8188
rect 10942 8128 11006 8132
rect 11022 8188 11086 8192
rect 11022 8132 11026 8188
rect 11026 8132 11082 8188
rect 11082 8132 11086 8188
rect 11022 8128 11086 8132
rect 11102 8188 11166 8192
rect 11102 8132 11106 8188
rect 11106 8132 11162 8188
rect 11162 8132 11166 8188
rect 11102 8128 11166 8132
rect 13962 8188 14026 8192
rect 13962 8132 13966 8188
rect 13966 8132 14022 8188
rect 14022 8132 14026 8188
rect 13962 8128 14026 8132
rect 14042 8188 14106 8192
rect 14042 8132 14046 8188
rect 14046 8132 14102 8188
rect 14102 8132 14106 8188
rect 14042 8128 14106 8132
rect 14122 8188 14186 8192
rect 14122 8132 14126 8188
rect 14126 8132 14182 8188
rect 14182 8132 14186 8188
rect 14122 8128 14186 8132
rect 14202 8188 14266 8192
rect 14202 8132 14206 8188
rect 14206 8132 14262 8188
rect 14262 8132 14266 8188
rect 14202 8128 14266 8132
rect 17062 8188 17126 8192
rect 17062 8132 17066 8188
rect 17066 8132 17122 8188
rect 17122 8132 17126 8188
rect 17062 8128 17126 8132
rect 17142 8188 17206 8192
rect 17142 8132 17146 8188
rect 17146 8132 17202 8188
rect 17202 8132 17206 8188
rect 17142 8128 17206 8132
rect 17222 8188 17286 8192
rect 17222 8132 17226 8188
rect 17226 8132 17282 8188
rect 17282 8132 17286 8188
rect 17222 8128 17286 8132
rect 17302 8188 17366 8192
rect 17302 8132 17306 8188
rect 17306 8132 17362 8188
rect 17362 8132 17366 8188
rect 17302 8128 17366 8132
rect 3112 7644 3176 7648
rect 3112 7588 3116 7644
rect 3116 7588 3172 7644
rect 3172 7588 3176 7644
rect 3112 7584 3176 7588
rect 3192 7644 3256 7648
rect 3192 7588 3196 7644
rect 3196 7588 3252 7644
rect 3252 7588 3256 7644
rect 3192 7584 3256 7588
rect 3272 7644 3336 7648
rect 3272 7588 3276 7644
rect 3276 7588 3332 7644
rect 3332 7588 3336 7644
rect 3272 7584 3336 7588
rect 3352 7644 3416 7648
rect 3352 7588 3356 7644
rect 3356 7588 3412 7644
rect 3412 7588 3416 7644
rect 3352 7584 3416 7588
rect 6212 7644 6276 7648
rect 6212 7588 6216 7644
rect 6216 7588 6272 7644
rect 6272 7588 6276 7644
rect 6212 7584 6276 7588
rect 6292 7644 6356 7648
rect 6292 7588 6296 7644
rect 6296 7588 6352 7644
rect 6352 7588 6356 7644
rect 6292 7584 6356 7588
rect 6372 7644 6436 7648
rect 6372 7588 6376 7644
rect 6376 7588 6432 7644
rect 6432 7588 6436 7644
rect 6372 7584 6436 7588
rect 6452 7644 6516 7648
rect 6452 7588 6456 7644
rect 6456 7588 6512 7644
rect 6512 7588 6516 7644
rect 6452 7584 6516 7588
rect 9312 7644 9376 7648
rect 9312 7588 9316 7644
rect 9316 7588 9372 7644
rect 9372 7588 9376 7644
rect 9312 7584 9376 7588
rect 9392 7644 9456 7648
rect 9392 7588 9396 7644
rect 9396 7588 9452 7644
rect 9452 7588 9456 7644
rect 9392 7584 9456 7588
rect 9472 7644 9536 7648
rect 9472 7588 9476 7644
rect 9476 7588 9532 7644
rect 9532 7588 9536 7644
rect 9472 7584 9536 7588
rect 9552 7644 9616 7648
rect 9552 7588 9556 7644
rect 9556 7588 9612 7644
rect 9612 7588 9616 7644
rect 9552 7584 9616 7588
rect 12412 7644 12476 7648
rect 12412 7588 12416 7644
rect 12416 7588 12472 7644
rect 12472 7588 12476 7644
rect 12412 7584 12476 7588
rect 12492 7644 12556 7648
rect 12492 7588 12496 7644
rect 12496 7588 12552 7644
rect 12552 7588 12556 7644
rect 12492 7584 12556 7588
rect 12572 7644 12636 7648
rect 12572 7588 12576 7644
rect 12576 7588 12632 7644
rect 12632 7588 12636 7644
rect 12572 7584 12636 7588
rect 12652 7644 12716 7648
rect 12652 7588 12656 7644
rect 12656 7588 12712 7644
rect 12712 7588 12716 7644
rect 12652 7584 12716 7588
rect 15512 7644 15576 7648
rect 15512 7588 15516 7644
rect 15516 7588 15572 7644
rect 15572 7588 15576 7644
rect 15512 7584 15576 7588
rect 15592 7644 15656 7648
rect 15592 7588 15596 7644
rect 15596 7588 15652 7644
rect 15652 7588 15656 7644
rect 15592 7584 15656 7588
rect 15672 7644 15736 7648
rect 15672 7588 15676 7644
rect 15676 7588 15732 7644
rect 15732 7588 15736 7644
rect 15672 7584 15736 7588
rect 15752 7644 15816 7648
rect 15752 7588 15756 7644
rect 15756 7588 15812 7644
rect 15812 7588 15816 7644
rect 15752 7584 15816 7588
rect 18612 7644 18676 7648
rect 18612 7588 18616 7644
rect 18616 7588 18672 7644
rect 18672 7588 18676 7644
rect 18612 7584 18676 7588
rect 18692 7644 18756 7648
rect 18692 7588 18696 7644
rect 18696 7588 18752 7644
rect 18752 7588 18756 7644
rect 18692 7584 18756 7588
rect 18772 7644 18836 7648
rect 18772 7588 18776 7644
rect 18776 7588 18832 7644
rect 18832 7588 18836 7644
rect 18772 7584 18836 7588
rect 18852 7644 18916 7648
rect 18852 7588 18856 7644
rect 18856 7588 18912 7644
rect 18912 7588 18916 7644
rect 18852 7584 18916 7588
rect 16068 7380 16132 7444
rect 16804 7244 16868 7308
rect 4662 7100 4726 7104
rect 4662 7044 4666 7100
rect 4666 7044 4722 7100
rect 4722 7044 4726 7100
rect 4662 7040 4726 7044
rect 4742 7100 4806 7104
rect 4742 7044 4746 7100
rect 4746 7044 4802 7100
rect 4802 7044 4806 7100
rect 4742 7040 4806 7044
rect 4822 7100 4886 7104
rect 4822 7044 4826 7100
rect 4826 7044 4882 7100
rect 4882 7044 4886 7100
rect 4822 7040 4886 7044
rect 4902 7100 4966 7104
rect 4902 7044 4906 7100
rect 4906 7044 4962 7100
rect 4962 7044 4966 7100
rect 4902 7040 4966 7044
rect 7762 7100 7826 7104
rect 7762 7044 7766 7100
rect 7766 7044 7822 7100
rect 7822 7044 7826 7100
rect 7762 7040 7826 7044
rect 7842 7100 7906 7104
rect 7842 7044 7846 7100
rect 7846 7044 7902 7100
rect 7902 7044 7906 7100
rect 7842 7040 7906 7044
rect 7922 7100 7986 7104
rect 7922 7044 7926 7100
rect 7926 7044 7982 7100
rect 7982 7044 7986 7100
rect 7922 7040 7986 7044
rect 8002 7100 8066 7104
rect 8002 7044 8006 7100
rect 8006 7044 8062 7100
rect 8062 7044 8066 7100
rect 8002 7040 8066 7044
rect 10862 7100 10926 7104
rect 10862 7044 10866 7100
rect 10866 7044 10922 7100
rect 10922 7044 10926 7100
rect 10862 7040 10926 7044
rect 10942 7100 11006 7104
rect 10942 7044 10946 7100
rect 10946 7044 11002 7100
rect 11002 7044 11006 7100
rect 10942 7040 11006 7044
rect 11022 7100 11086 7104
rect 11022 7044 11026 7100
rect 11026 7044 11082 7100
rect 11082 7044 11086 7100
rect 11022 7040 11086 7044
rect 11102 7100 11166 7104
rect 11102 7044 11106 7100
rect 11106 7044 11162 7100
rect 11162 7044 11166 7100
rect 11102 7040 11166 7044
rect 13962 7100 14026 7104
rect 13962 7044 13966 7100
rect 13966 7044 14022 7100
rect 14022 7044 14026 7100
rect 13962 7040 14026 7044
rect 14042 7100 14106 7104
rect 14042 7044 14046 7100
rect 14046 7044 14102 7100
rect 14102 7044 14106 7100
rect 14042 7040 14106 7044
rect 14122 7100 14186 7104
rect 14122 7044 14126 7100
rect 14126 7044 14182 7100
rect 14182 7044 14186 7100
rect 14122 7040 14186 7044
rect 14202 7100 14266 7104
rect 14202 7044 14206 7100
rect 14206 7044 14262 7100
rect 14262 7044 14266 7100
rect 14202 7040 14266 7044
rect 17062 7100 17126 7104
rect 17062 7044 17066 7100
rect 17066 7044 17122 7100
rect 17122 7044 17126 7100
rect 17062 7040 17126 7044
rect 17142 7100 17206 7104
rect 17142 7044 17146 7100
rect 17146 7044 17202 7100
rect 17202 7044 17206 7100
rect 17142 7040 17206 7044
rect 17222 7100 17286 7104
rect 17222 7044 17226 7100
rect 17226 7044 17282 7100
rect 17282 7044 17286 7100
rect 17222 7040 17286 7044
rect 17302 7100 17366 7104
rect 17302 7044 17306 7100
rect 17306 7044 17362 7100
rect 17362 7044 17366 7100
rect 17302 7040 17366 7044
rect 16436 6700 16500 6764
rect 3112 6556 3176 6560
rect 3112 6500 3116 6556
rect 3116 6500 3172 6556
rect 3172 6500 3176 6556
rect 3112 6496 3176 6500
rect 3192 6556 3256 6560
rect 3192 6500 3196 6556
rect 3196 6500 3252 6556
rect 3252 6500 3256 6556
rect 3192 6496 3256 6500
rect 3272 6556 3336 6560
rect 3272 6500 3276 6556
rect 3276 6500 3332 6556
rect 3332 6500 3336 6556
rect 3272 6496 3336 6500
rect 3352 6556 3416 6560
rect 3352 6500 3356 6556
rect 3356 6500 3412 6556
rect 3412 6500 3416 6556
rect 3352 6496 3416 6500
rect 6212 6556 6276 6560
rect 6212 6500 6216 6556
rect 6216 6500 6272 6556
rect 6272 6500 6276 6556
rect 6212 6496 6276 6500
rect 6292 6556 6356 6560
rect 6292 6500 6296 6556
rect 6296 6500 6352 6556
rect 6352 6500 6356 6556
rect 6292 6496 6356 6500
rect 6372 6556 6436 6560
rect 6372 6500 6376 6556
rect 6376 6500 6432 6556
rect 6432 6500 6436 6556
rect 6372 6496 6436 6500
rect 6452 6556 6516 6560
rect 6452 6500 6456 6556
rect 6456 6500 6512 6556
rect 6512 6500 6516 6556
rect 6452 6496 6516 6500
rect 9312 6556 9376 6560
rect 9312 6500 9316 6556
rect 9316 6500 9372 6556
rect 9372 6500 9376 6556
rect 9312 6496 9376 6500
rect 9392 6556 9456 6560
rect 9392 6500 9396 6556
rect 9396 6500 9452 6556
rect 9452 6500 9456 6556
rect 9392 6496 9456 6500
rect 9472 6556 9536 6560
rect 9472 6500 9476 6556
rect 9476 6500 9532 6556
rect 9532 6500 9536 6556
rect 9472 6496 9536 6500
rect 9552 6556 9616 6560
rect 9552 6500 9556 6556
rect 9556 6500 9612 6556
rect 9612 6500 9616 6556
rect 9552 6496 9616 6500
rect 12412 6556 12476 6560
rect 12412 6500 12416 6556
rect 12416 6500 12472 6556
rect 12472 6500 12476 6556
rect 12412 6496 12476 6500
rect 12492 6556 12556 6560
rect 12492 6500 12496 6556
rect 12496 6500 12552 6556
rect 12552 6500 12556 6556
rect 12492 6496 12556 6500
rect 12572 6556 12636 6560
rect 12572 6500 12576 6556
rect 12576 6500 12632 6556
rect 12632 6500 12636 6556
rect 12572 6496 12636 6500
rect 12652 6556 12716 6560
rect 12652 6500 12656 6556
rect 12656 6500 12712 6556
rect 12712 6500 12716 6556
rect 12652 6496 12716 6500
rect 15512 6556 15576 6560
rect 15512 6500 15516 6556
rect 15516 6500 15572 6556
rect 15572 6500 15576 6556
rect 15512 6496 15576 6500
rect 15592 6556 15656 6560
rect 15592 6500 15596 6556
rect 15596 6500 15652 6556
rect 15652 6500 15656 6556
rect 15592 6496 15656 6500
rect 15672 6556 15736 6560
rect 15672 6500 15676 6556
rect 15676 6500 15732 6556
rect 15732 6500 15736 6556
rect 15672 6496 15736 6500
rect 15752 6556 15816 6560
rect 15752 6500 15756 6556
rect 15756 6500 15812 6556
rect 15812 6500 15816 6556
rect 15752 6496 15816 6500
rect 18612 6556 18676 6560
rect 18612 6500 18616 6556
rect 18616 6500 18672 6556
rect 18672 6500 18676 6556
rect 18612 6496 18676 6500
rect 18692 6556 18756 6560
rect 18692 6500 18696 6556
rect 18696 6500 18752 6556
rect 18752 6500 18756 6556
rect 18692 6496 18756 6500
rect 18772 6556 18836 6560
rect 18772 6500 18776 6556
rect 18776 6500 18832 6556
rect 18832 6500 18836 6556
rect 18772 6496 18836 6500
rect 18852 6556 18916 6560
rect 18852 6500 18856 6556
rect 18856 6500 18912 6556
rect 18912 6500 18916 6556
rect 18852 6496 18916 6500
rect 4662 6012 4726 6016
rect 4662 5956 4666 6012
rect 4666 5956 4722 6012
rect 4722 5956 4726 6012
rect 4662 5952 4726 5956
rect 4742 6012 4806 6016
rect 4742 5956 4746 6012
rect 4746 5956 4802 6012
rect 4802 5956 4806 6012
rect 4742 5952 4806 5956
rect 4822 6012 4886 6016
rect 4822 5956 4826 6012
rect 4826 5956 4882 6012
rect 4882 5956 4886 6012
rect 4822 5952 4886 5956
rect 4902 6012 4966 6016
rect 4902 5956 4906 6012
rect 4906 5956 4962 6012
rect 4962 5956 4966 6012
rect 4902 5952 4966 5956
rect 7762 6012 7826 6016
rect 7762 5956 7766 6012
rect 7766 5956 7822 6012
rect 7822 5956 7826 6012
rect 7762 5952 7826 5956
rect 7842 6012 7906 6016
rect 7842 5956 7846 6012
rect 7846 5956 7902 6012
rect 7902 5956 7906 6012
rect 7842 5952 7906 5956
rect 7922 6012 7986 6016
rect 7922 5956 7926 6012
rect 7926 5956 7982 6012
rect 7982 5956 7986 6012
rect 7922 5952 7986 5956
rect 8002 6012 8066 6016
rect 8002 5956 8006 6012
rect 8006 5956 8062 6012
rect 8062 5956 8066 6012
rect 8002 5952 8066 5956
rect 10862 6012 10926 6016
rect 10862 5956 10866 6012
rect 10866 5956 10922 6012
rect 10922 5956 10926 6012
rect 10862 5952 10926 5956
rect 10942 6012 11006 6016
rect 10942 5956 10946 6012
rect 10946 5956 11002 6012
rect 11002 5956 11006 6012
rect 10942 5952 11006 5956
rect 11022 6012 11086 6016
rect 11022 5956 11026 6012
rect 11026 5956 11082 6012
rect 11082 5956 11086 6012
rect 11022 5952 11086 5956
rect 11102 6012 11166 6016
rect 11102 5956 11106 6012
rect 11106 5956 11162 6012
rect 11162 5956 11166 6012
rect 11102 5952 11166 5956
rect 13962 6012 14026 6016
rect 13962 5956 13966 6012
rect 13966 5956 14022 6012
rect 14022 5956 14026 6012
rect 13962 5952 14026 5956
rect 14042 6012 14106 6016
rect 14042 5956 14046 6012
rect 14046 5956 14102 6012
rect 14102 5956 14106 6012
rect 14042 5952 14106 5956
rect 14122 6012 14186 6016
rect 14122 5956 14126 6012
rect 14126 5956 14182 6012
rect 14182 5956 14186 6012
rect 14122 5952 14186 5956
rect 14202 6012 14266 6016
rect 14202 5956 14206 6012
rect 14206 5956 14262 6012
rect 14262 5956 14266 6012
rect 14202 5952 14266 5956
rect 17062 6012 17126 6016
rect 17062 5956 17066 6012
rect 17066 5956 17122 6012
rect 17122 5956 17126 6012
rect 17062 5952 17126 5956
rect 17142 6012 17206 6016
rect 17142 5956 17146 6012
rect 17146 5956 17202 6012
rect 17202 5956 17206 6012
rect 17142 5952 17206 5956
rect 17222 6012 17286 6016
rect 17222 5956 17226 6012
rect 17226 5956 17282 6012
rect 17282 5956 17286 6012
rect 17222 5952 17286 5956
rect 17302 6012 17366 6016
rect 17302 5956 17306 6012
rect 17306 5956 17362 6012
rect 17362 5956 17366 6012
rect 17302 5952 17366 5956
rect 17540 5476 17604 5540
rect 3112 5468 3176 5472
rect 3112 5412 3116 5468
rect 3116 5412 3172 5468
rect 3172 5412 3176 5468
rect 3112 5408 3176 5412
rect 3192 5468 3256 5472
rect 3192 5412 3196 5468
rect 3196 5412 3252 5468
rect 3252 5412 3256 5468
rect 3192 5408 3256 5412
rect 3272 5468 3336 5472
rect 3272 5412 3276 5468
rect 3276 5412 3332 5468
rect 3332 5412 3336 5468
rect 3272 5408 3336 5412
rect 3352 5468 3416 5472
rect 3352 5412 3356 5468
rect 3356 5412 3412 5468
rect 3412 5412 3416 5468
rect 3352 5408 3416 5412
rect 6212 5468 6276 5472
rect 6212 5412 6216 5468
rect 6216 5412 6272 5468
rect 6272 5412 6276 5468
rect 6212 5408 6276 5412
rect 6292 5468 6356 5472
rect 6292 5412 6296 5468
rect 6296 5412 6352 5468
rect 6352 5412 6356 5468
rect 6292 5408 6356 5412
rect 6372 5468 6436 5472
rect 6372 5412 6376 5468
rect 6376 5412 6432 5468
rect 6432 5412 6436 5468
rect 6372 5408 6436 5412
rect 6452 5468 6516 5472
rect 6452 5412 6456 5468
rect 6456 5412 6512 5468
rect 6512 5412 6516 5468
rect 6452 5408 6516 5412
rect 9312 5468 9376 5472
rect 9312 5412 9316 5468
rect 9316 5412 9372 5468
rect 9372 5412 9376 5468
rect 9312 5408 9376 5412
rect 9392 5468 9456 5472
rect 9392 5412 9396 5468
rect 9396 5412 9452 5468
rect 9452 5412 9456 5468
rect 9392 5408 9456 5412
rect 9472 5468 9536 5472
rect 9472 5412 9476 5468
rect 9476 5412 9532 5468
rect 9532 5412 9536 5468
rect 9472 5408 9536 5412
rect 9552 5468 9616 5472
rect 9552 5412 9556 5468
rect 9556 5412 9612 5468
rect 9612 5412 9616 5468
rect 9552 5408 9616 5412
rect 12412 5468 12476 5472
rect 12412 5412 12416 5468
rect 12416 5412 12472 5468
rect 12472 5412 12476 5468
rect 12412 5408 12476 5412
rect 12492 5468 12556 5472
rect 12492 5412 12496 5468
rect 12496 5412 12552 5468
rect 12552 5412 12556 5468
rect 12492 5408 12556 5412
rect 12572 5468 12636 5472
rect 12572 5412 12576 5468
rect 12576 5412 12632 5468
rect 12632 5412 12636 5468
rect 12572 5408 12636 5412
rect 12652 5468 12716 5472
rect 12652 5412 12656 5468
rect 12656 5412 12712 5468
rect 12712 5412 12716 5468
rect 12652 5408 12716 5412
rect 15512 5468 15576 5472
rect 15512 5412 15516 5468
rect 15516 5412 15572 5468
rect 15572 5412 15576 5468
rect 15512 5408 15576 5412
rect 15592 5468 15656 5472
rect 15592 5412 15596 5468
rect 15596 5412 15652 5468
rect 15652 5412 15656 5468
rect 15592 5408 15656 5412
rect 15672 5468 15736 5472
rect 15672 5412 15676 5468
rect 15676 5412 15732 5468
rect 15732 5412 15736 5468
rect 15672 5408 15736 5412
rect 15752 5468 15816 5472
rect 15752 5412 15756 5468
rect 15756 5412 15812 5468
rect 15812 5412 15816 5468
rect 15752 5408 15816 5412
rect 18612 5468 18676 5472
rect 18612 5412 18616 5468
rect 18616 5412 18672 5468
rect 18672 5412 18676 5468
rect 18612 5408 18676 5412
rect 18692 5468 18756 5472
rect 18692 5412 18696 5468
rect 18696 5412 18752 5468
rect 18752 5412 18756 5468
rect 18692 5408 18756 5412
rect 18772 5468 18836 5472
rect 18772 5412 18776 5468
rect 18776 5412 18832 5468
rect 18832 5412 18836 5468
rect 18772 5408 18836 5412
rect 18852 5468 18916 5472
rect 18852 5412 18856 5468
rect 18856 5412 18912 5468
rect 18912 5412 18916 5468
rect 18852 5408 18916 5412
rect 16068 5204 16132 5268
rect 16804 5204 16868 5268
rect 4662 4924 4726 4928
rect 4662 4868 4666 4924
rect 4666 4868 4722 4924
rect 4722 4868 4726 4924
rect 4662 4864 4726 4868
rect 4742 4924 4806 4928
rect 4742 4868 4746 4924
rect 4746 4868 4802 4924
rect 4802 4868 4806 4924
rect 4742 4864 4806 4868
rect 4822 4924 4886 4928
rect 4822 4868 4826 4924
rect 4826 4868 4882 4924
rect 4882 4868 4886 4924
rect 4822 4864 4886 4868
rect 4902 4924 4966 4928
rect 4902 4868 4906 4924
rect 4906 4868 4962 4924
rect 4962 4868 4966 4924
rect 4902 4864 4966 4868
rect 7762 4924 7826 4928
rect 7762 4868 7766 4924
rect 7766 4868 7822 4924
rect 7822 4868 7826 4924
rect 7762 4864 7826 4868
rect 7842 4924 7906 4928
rect 7842 4868 7846 4924
rect 7846 4868 7902 4924
rect 7902 4868 7906 4924
rect 7842 4864 7906 4868
rect 7922 4924 7986 4928
rect 7922 4868 7926 4924
rect 7926 4868 7982 4924
rect 7982 4868 7986 4924
rect 7922 4864 7986 4868
rect 8002 4924 8066 4928
rect 8002 4868 8006 4924
rect 8006 4868 8062 4924
rect 8062 4868 8066 4924
rect 8002 4864 8066 4868
rect 10862 4924 10926 4928
rect 10862 4868 10866 4924
rect 10866 4868 10922 4924
rect 10922 4868 10926 4924
rect 10862 4864 10926 4868
rect 10942 4924 11006 4928
rect 10942 4868 10946 4924
rect 10946 4868 11002 4924
rect 11002 4868 11006 4924
rect 10942 4864 11006 4868
rect 11022 4924 11086 4928
rect 11022 4868 11026 4924
rect 11026 4868 11082 4924
rect 11082 4868 11086 4924
rect 11022 4864 11086 4868
rect 11102 4924 11166 4928
rect 11102 4868 11106 4924
rect 11106 4868 11162 4924
rect 11162 4868 11166 4924
rect 11102 4864 11166 4868
rect 13962 4924 14026 4928
rect 13962 4868 13966 4924
rect 13966 4868 14022 4924
rect 14022 4868 14026 4924
rect 13962 4864 14026 4868
rect 14042 4924 14106 4928
rect 14042 4868 14046 4924
rect 14046 4868 14102 4924
rect 14102 4868 14106 4924
rect 14042 4864 14106 4868
rect 14122 4924 14186 4928
rect 14122 4868 14126 4924
rect 14126 4868 14182 4924
rect 14182 4868 14186 4924
rect 14122 4864 14186 4868
rect 14202 4924 14266 4928
rect 14202 4868 14206 4924
rect 14206 4868 14262 4924
rect 14262 4868 14266 4924
rect 14202 4864 14266 4868
rect 17062 4924 17126 4928
rect 17062 4868 17066 4924
rect 17066 4868 17122 4924
rect 17122 4868 17126 4924
rect 17062 4864 17126 4868
rect 17142 4924 17206 4928
rect 17142 4868 17146 4924
rect 17146 4868 17202 4924
rect 17202 4868 17206 4924
rect 17142 4864 17206 4868
rect 17222 4924 17286 4928
rect 17222 4868 17226 4924
rect 17226 4868 17282 4924
rect 17282 4868 17286 4924
rect 17222 4864 17286 4868
rect 17302 4924 17366 4928
rect 17302 4868 17306 4924
rect 17306 4868 17362 4924
rect 17362 4868 17366 4924
rect 17302 4864 17366 4868
rect 16252 4388 16316 4452
rect 3112 4380 3176 4384
rect 3112 4324 3116 4380
rect 3116 4324 3172 4380
rect 3172 4324 3176 4380
rect 3112 4320 3176 4324
rect 3192 4380 3256 4384
rect 3192 4324 3196 4380
rect 3196 4324 3252 4380
rect 3252 4324 3256 4380
rect 3192 4320 3256 4324
rect 3272 4380 3336 4384
rect 3272 4324 3276 4380
rect 3276 4324 3332 4380
rect 3332 4324 3336 4380
rect 3272 4320 3336 4324
rect 3352 4380 3416 4384
rect 3352 4324 3356 4380
rect 3356 4324 3412 4380
rect 3412 4324 3416 4380
rect 3352 4320 3416 4324
rect 6212 4380 6276 4384
rect 6212 4324 6216 4380
rect 6216 4324 6272 4380
rect 6272 4324 6276 4380
rect 6212 4320 6276 4324
rect 6292 4380 6356 4384
rect 6292 4324 6296 4380
rect 6296 4324 6352 4380
rect 6352 4324 6356 4380
rect 6292 4320 6356 4324
rect 6372 4380 6436 4384
rect 6372 4324 6376 4380
rect 6376 4324 6432 4380
rect 6432 4324 6436 4380
rect 6372 4320 6436 4324
rect 6452 4380 6516 4384
rect 6452 4324 6456 4380
rect 6456 4324 6512 4380
rect 6512 4324 6516 4380
rect 6452 4320 6516 4324
rect 9312 4380 9376 4384
rect 9312 4324 9316 4380
rect 9316 4324 9372 4380
rect 9372 4324 9376 4380
rect 9312 4320 9376 4324
rect 9392 4380 9456 4384
rect 9392 4324 9396 4380
rect 9396 4324 9452 4380
rect 9452 4324 9456 4380
rect 9392 4320 9456 4324
rect 9472 4380 9536 4384
rect 9472 4324 9476 4380
rect 9476 4324 9532 4380
rect 9532 4324 9536 4380
rect 9472 4320 9536 4324
rect 9552 4380 9616 4384
rect 9552 4324 9556 4380
rect 9556 4324 9612 4380
rect 9612 4324 9616 4380
rect 9552 4320 9616 4324
rect 12412 4380 12476 4384
rect 12412 4324 12416 4380
rect 12416 4324 12472 4380
rect 12472 4324 12476 4380
rect 12412 4320 12476 4324
rect 12492 4380 12556 4384
rect 12492 4324 12496 4380
rect 12496 4324 12552 4380
rect 12552 4324 12556 4380
rect 12492 4320 12556 4324
rect 12572 4380 12636 4384
rect 12572 4324 12576 4380
rect 12576 4324 12632 4380
rect 12632 4324 12636 4380
rect 12572 4320 12636 4324
rect 12652 4380 12716 4384
rect 12652 4324 12656 4380
rect 12656 4324 12712 4380
rect 12712 4324 12716 4380
rect 12652 4320 12716 4324
rect 15512 4380 15576 4384
rect 15512 4324 15516 4380
rect 15516 4324 15572 4380
rect 15572 4324 15576 4380
rect 15512 4320 15576 4324
rect 15592 4380 15656 4384
rect 15592 4324 15596 4380
rect 15596 4324 15652 4380
rect 15652 4324 15656 4380
rect 15592 4320 15656 4324
rect 15672 4380 15736 4384
rect 15672 4324 15676 4380
rect 15676 4324 15732 4380
rect 15732 4324 15736 4380
rect 15672 4320 15736 4324
rect 15752 4380 15816 4384
rect 15752 4324 15756 4380
rect 15756 4324 15812 4380
rect 15812 4324 15816 4380
rect 15752 4320 15816 4324
rect 18612 4380 18676 4384
rect 18612 4324 18616 4380
rect 18616 4324 18672 4380
rect 18672 4324 18676 4380
rect 18612 4320 18676 4324
rect 18692 4380 18756 4384
rect 18692 4324 18696 4380
rect 18696 4324 18752 4380
rect 18752 4324 18756 4380
rect 18692 4320 18756 4324
rect 18772 4380 18836 4384
rect 18772 4324 18776 4380
rect 18776 4324 18832 4380
rect 18832 4324 18836 4380
rect 18772 4320 18836 4324
rect 18852 4380 18916 4384
rect 18852 4324 18856 4380
rect 18856 4324 18912 4380
rect 18912 4324 18916 4380
rect 18852 4320 18916 4324
rect 4662 3836 4726 3840
rect 4662 3780 4666 3836
rect 4666 3780 4722 3836
rect 4722 3780 4726 3836
rect 4662 3776 4726 3780
rect 4742 3836 4806 3840
rect 4742 3780 4746 3836
rect 4746 3780 4802 3836
rect 4802 3780 4806 3836
rect 4742 3776 4806 3780
rect 4822 3836 4886 3840
rect 4822 3780 4826 3836
rect 4826 3780 4882 3836
rect 4882 3780 4886 3836
rect 4822 3776 4886 3780
rect 4902 3836 4966 3840
rect 4902 3780 4906 3836
rect 4906 3780 4962 3836
rect 4962 3780 4966 3836
rect 4902 3776 4966 3780
rect 7762 3836 7826 3840
rect 7762 3780 7766 3836
rect 7766 3780 7822 3836
rect 7822 3780 7826 3836
rect 7762 3776 7826 3780
rect 7842 3836 7906 3840
rect 7842 3780 7846 3836
rect 7846 3780 7902 3836
rect 7902 3780 7906 3836
rect 7842 3776 7906 3780
rect 7922 3836 7986 3840
rect 7922 3780 7926 3836
rect 7926 3780 7982 3836
rect 7982 3780 7986 3836
rect 7922 3776 7986 3780
rect 8002 3836 8066 3840
rect 8002 3780 8006 3836
rect 8006 3780 8062 3836
rect 8062 3780 8066 3836
rect 8002 3776 8066 3780
rect 10862 3836 10926 3840
rect 10862 3780 10866 3836
rect 10866 3780 10922 3836
rect 10922 3780 10926 3836
rect 10862 3776 10926 3780
rect 10942 3836 11006 3840
rect 10942 3780 10946 3836
rect 10946 3780 11002 3836
rect 11002 3780 11006 3836
rect 10942 3776 11006 3780
rect 11022 3836 11086 3840
rect 11022 3780 11026 3836
rect 11026 3780 11082 3836
rect 11082 3780 11086 3836
rect 11022 3776 11086 3780
rect 11102 3836 11166 3840
rect 11102 3780 11106 3836
rect 11106 3780 11162 3836
rect 11162 3780 11166 3836
rect 11102 3776 11166 3780
rect 13962 3836 14026 3840
rect 13962 3780 13966 3836
rect 13966 3780 14022 3836
rect 14022 3780 14026 3836
rect 13962 3776 14026 3780
rect 14042 3836 14106 3840
rect 14042 3780 14046 3836
rect 14046 3780 14102 3836
rect 14102 3780 14106 3836
rect 14042 3776 14106 3780
rect 14122 3836 14186 3840
rect 14122 3780 14126 3836
rect 14126 3780 14182 3836
rect 14182 3780 14186 3836
rect 14122 3776 14186 3780
rect 14202 3836 14266 3840
rect 14202 3780 14206 3836
rect 14206 3780 14262 3836
rect 14262 3780 14266 3836
rect 14202 3776 14266 3780
rect 17062 3836 17126 3840
rect 17062 3780 17066 3836
rect 17066 3780 17122 3836
rect 17122 3780 17126 3836
rect 17062 3776 17126 3780
rect 17142 3836 17206 3840
rect 17142 3780 17146 3836
rect 17146 3780 17202 3836
rect 17202 3780 17206 3836
rect 17142 3776 17206 3780
rect 17222 3836 17286 3840
rect 17222 3780 17226 3836
rect 17226 3780 17282 3836
rect 17282 3780 17286 3836
rect 17222 3776 17286 3780
rect 17302 3836 17366 3840
rect 17302 3780 17306 3836
rect 17306 3780 17362 3836
rect 17362 3780 17366 3836
rect 17302 3776 17366 3780
rect 16436 3300 16500 3364
rect 3112 3292 3176 3296
rect 3112 3236 3116 3292
rect 3116 3236 3172 3292
rect 3172 3236 3176 3292
rect 3112 3232 3176 3236
rect 3192 3292 3256 3296
rect 3192 3236 3196 3292
rect 3196 3236 3252 3292
rect 3252 3236 3256 3292
rect 3192 3232 3256 3236
rect 3272 3292 3336 3296
rect 3272 3236 3276 3292
rect 3276 3236 3332 3292
rect 3332 3236 3336 3292
rect 3272 3232 3336 3236
rect 3352 3292 3416 3296
rect 3352 3236 3356 3292
rect 3356 3236 3412 3292
rect 3412 3236 3416 3292
rect 3352 3232 3416 3236
rect 6212 3292 6276 3296
rect 6212 3236 6216 3292
rect 6216 3236 6272 3292
rect 6272 3236 6276 3292
rect 6212 3232 6276 3236
rect 6292 3292 6356 3296
rect 6292 3236 6296 3292
rect 6296 3236 6352 3292
rect 6352 3236 6356 3292
rect 6292 3232 6356 3236
rect 6372 3292 6436 3296
rect 6372 3236 6376 3292
rect 6376 3236 6432 3292
rect 6432 3236 6436 3292
rect 6372 3232 6436 3236
rect 6452 3292 6516 3296
rect 6452 3236 6456 3292
rect 6456 3236 6512 3292
rect 6512 3236 6516 3292
rect 6452 3232 6516 3236
rect 9312 3292 9376 3296
rect 9312 3236 9316 3292
rect 9316 3236 9372 3292
rect 9372 3236 9376 3292
rect 9312 3232 9376 3236
rect 9392 3292 9456 3296
rect 9392 3236 9396 3292
rect 9396 3236 9452 3292
rect 9452 3236 9456 3292
rect 9392 3232 9456 3236
rect 9472 3292 9536 3296
rect 9472 3236 9476 3292
rect 9476 3236 9532 3292
rect 9532 3236 9536 3292
rect 9472 3232 9536 3236
rect 9552 3292 9616 3296
rect 9552 3236 9556 3292
rect 9556 3236 9612 3292
rect 9612 3236 9616 3292
rect 9552 3232 9616 3236
rect 12412 3292 12476 3296
rect 12412 3236 12416 3292
rect 12416 3236 12472 3292
rect 12472 3236 12476 3292
rect 12412 3232 12476 3236
rect 12492 3292 12556 3296
rect 12492 3236 12496 3292
rect 12496 3236 12552 3292
rect 12552 3236 12556 3292
rect 12492 3232 12556 3236
rect 12572 3292 12636 3296
rect 12572 3236 12576 3292
rect 12576 3236 12632 3292
rect 12632 3236 12636 3292
rect 12572 3232 12636 3236
rect 12652 3292 12716 3296
rect 12652 3236 12656 3292
rect 12656 3236 12712 3292
rect 12712 3236 12716 3292
rect 12652 3232 12716 3236
rect 15512 3292 15576 3296
rect 15512 3236 15516 3292
rect 15516 3236 15572 3292
rect 15572 3236 15576 3292
rect 15512 3232 15576 3236
rect 15592 3292 15656 3296
rect 15592 3236 15596 3292
rect 15596 3236 15652 3292
rect 15652 3236 15656 3292
rect 15592 3232 15656 3236
rect 15672 3292 15736 3296
rect 15672 3236 15676 3292
rect 15676 3236 15732 3292
rect 15732 3236 15736 3292
rect 15672 3232 15736 3236
rect 15752 3292 15816 3296
rect 15752 3236 15756 3292
rect 15756 3236 15812 3292
rect 15812 3236 15816 3292
rect 15752 3232 15816 3236
rect 18612 3292 18676 3296
rect 18612 3236 18616 3292
rect 18616 3236 18672 3292
rect 18672 3236 18676 3292
rect 18612 3232 18676 3236
rect 18692 3292 18756 3296
rect 18692 3236 18696 3292
rect 18696 3236 18752 3292
rect 18752 3236 18756 3292
rect 18692 3232 18756 3236
rect 18772 3292 18836 3296
rect 18772 3236 18776 3292
rect 18776 3236 18832 3292
rect 18832 3236 18836 3292
rect 18772 3232 18836 3236
rect 18852 3292 18916 3296
rect 18852 3236 18856 3292
rect 18856 3236 18912 3292
rect 18912 3236 18916 3292
rect 18852 3232 18916 3236
rect 16620 2756 16684 2820
rect 4662 2748 4726 2752
rect 4662 2692 4666 2748
rect 4666 2692 4722 2748
rect 4722 2692 4726 2748
rect 4662 2688 4726 2692
rect 4742 2748 4806 2752
rect 4742 2692 4746 2748
rect 4746 2692 4802 2748
rect 4802 2692 4806 2748
rect 4742 2688 4806 2692
rect 4822 2748 4886 2752
rect 4822 2692 4826 2748
rect 4826 2692 4882 2748
rect 4882 2692 4886 2748
rect 4822 2688 4886 2692
rect 4902 2748 4966 2752
rect 4902 2692 4906 2748
rect 4906 2692 4962 2748
rect 4962 2692 4966 2748
rect 4902 2688 4966 2692
rect 7762 2748 7826 2752
rect 7762 2692 7766 2748
rect 7766 2692 7822 2748
rect 7822 2692 7826 2748
rect 7762 2688 7826 2692
rect 7842 2748 7906 2752
rect 7842 2692 7846 2748
rect 7846 2692 7902 2748
rect 7902 2692 7906 2748
rect 7842 2688 7906 2692
rect 7922 2748 7986 2752
rect 7922 2692 7926 2748
rect 7926 2692 7982 2748
rect 7982 2692 7986 2748
rect 7922 2688 7986 2692
rect 8002 2748 8066 2752
rect 8002 2692 8006 2748
rect 8006 2692 8062 2748
rect 8062 2692 8066 2748
rect 8002 2688 8066 2692
rect 10862 2748 10926 2752
rect 10862 2692 10866 2748
rect 10866 2692 10922 2748
rect 10922 2692 10926 2748
rect 10862 2688 10926 2692
rect 10942 2748 11006 2752
rect 10942 2692 10946 2748
rect 10946 2692 11002 2748
rect 11002 2692 11006 2748
rect 10942 2688 11006 2692
rect 11022 2748 11086 2752
rect 11022 2692 11026 2748
rect 11026 2692 11082 2748
rect 11082 2692 11086 2748
rect 11022 2688 11086 2692
rect 11102 2748 11166 2752
rect 11102 2692 11106 2748
rect 11106 2692 11162 2748
rect 11162 2692 11166 2748
rect 11102 2688 11166 2692
rect 13962 2748 14026 2752
rect 13962 2692 13966 2748
rect 13966 2692 14022 2748
rect 14022 2692 14026 2748
rect 13962 2688 14026 2692
rect 14042 2748 14106 2752
rect 14042 2692 14046 2748
rect 14046 2692 14102 2748
rect 14102 2692 14106 2748
rect 14042 2688 14106 2692
rect 14122 2748 14186 2752
rect 14122 2692 14126 2748
rect 14126 2692 14182 2748
rect 14182 2692 14186 2748
rect 14122 2688 14186 2692
rect 14202 2748 14266 2752
rect 14202 2692 14206 2748
rect 14206 2692 14262 2748
rect 14262 2692 14266 2748
rect 14202 2688 14266 2692
rect 17062 2748 17126 2752
rect 17062 2692 17066 2748
rect 17066 2692 17122 2748
rect 17122 2692 17126 2748
rect 17062 2688 17126 2692
rect 17142 2748 17206 2752
rect 17142 2692 17146 2748
rect 17146 2692 17202 2748
rect 17202 2692 17206 2748
rect 17142 2688 17206 2692
rect 17222 2748 17286 2752
rect 17222 2692 17226 2748
rect 17226 2692 17282 2748
rect 17282 2692 17286 2748
rect 17222 2688 17286 2692
rect 17302 2748 17366 2752
rect 17302 2692 17306 2748
rect 17306 2692 17362 2748
rect 17362 2692 17366 2748
rect 17302 2688 17366 2692
rect 16620 2680 16684 2684
rect 16620 2624 16634 2680
rect 16634 2624 16684 2680
rect 16620 2620 16684 2624
rect 14412 2484 14476 2548
rect 3112 2204 3176 2208
rect 3112 2148 3116 2204
rect 3116 2148 3172 2204
rect 3172 2148 3176 2204
rect 3112 2144 3176 2148
rect 3192 2204 3256 2208
rect 3192 2148 3196 2204
rect 3196 2148 3252 2204
rect 3252 2148 3256 2204
rect 3192 2144 3256 2148
rect 3272 2204 3336 2208
rect 3272 2148 3276 2204
rect 3276 2148 3332 2204
rect 3332 2148 3336 2204
rect 3272 2144 3336 2148
rect 3352 2204 3416 2208
rect 3352 2148 3356 2204
rect 3356 2148 3412 2204
rect 3412 2148 3416 2204
rect 3352 2144 3416 2148
rect 6212 2204 6276 2208
rect 6212 2148 6216 2204
rect 6216 2148 6272 2204
rect 6272 2148 6276 2204
rect 6212 2144 6276 2148
rect 6292 2204 6356 2208
rect 6292 2148 6296 2204
rect 6296 2148 6352 2204
rect 6352 2148 6356 2204
rect 6292 2144 6356 2148
rect 6372 2204 6436 2208
rect 6372 2148 6376 2204
rect 6376 2148 6432 2204
rect 6432 2148 6436 2204
rect 6372 2144 6436 2148
rect 6452 2204 6516 2208
rect 6452 2148 6456 2204
rect 6456 2148 6512 2204
rect 6512 2148 6516 2204
rect 6452 2144 6516 2148
rect 9312 2204 9376 2208
rect 9312 2148 9316 2204
rect 9316 2148 9372 2204
rect 9372 2148 9376 2204
rect 9312 2144 9376 2148
rect 9392 2204 9456 2208
rect 9392 2148 9396 2204
rect 9396 2148 9452 2204
rect 9452 2148 9456 2204
rect 9392 2144 9456 2148
rect 9472 2204 9536 2208
rect 9472 2148 9476 2204
rect 9476 2148 9532 2204
rect 9532 2148 9536 2204
rect 9472 2144 9536 2148
rect 9552 2204 9616 2208
rect 9552 2148 9556 2204
rect 9556 2148 9612 2204
rect 9612 2148 9616 2204
rect 9552 2144 9616 2148
rect 12412 2204 12476 2208
rect 12412 2148 12416 2204
rect 12416 2148 12472 2204
rect 12472 2148 12476 2204
rect 12412 2144 12476 2148
rect 12492 2204 12556 2208
rect 12492 2148 12496 2204
rect 12496 2148 12552 2204
rect 12552 2148 12556 2204
rect 12492 2144 12556 2148
rect 12572 2204 12636 2208
rect 12572 2148 12576 2204
rect 12576 2148 12632 2204
rect 12632 2148 12636 2204
rect 12572 2144 12636 2148
rect 12652 2204 12716 2208
rect 12652 2148 12656 2204
rect 12656 2148 12712 2204
rect 12712 2148 12716 2204
rect 12652 2144 12716 2148
rect 15512 2204 15576 2208
rect 15512 2148 15516 2204
rect 15516 2148 15572 2204
rect 15572 2148 15576 2204
rect 15512 2144 15576 2148
rect 15592 2204 15656 2208
rect 15592 2148 15596 2204
rect 15596 2148 15652 2204
rect 15652 2148 15656 2204
rect 15592 2144 15656 2148
rect 15672 2204 15736 2208
rect 15672 2148 15676 2204
rect 15676 2148 15732 2204
rect 15732 2148 15736 2204
rect 15672 2144 15736 2148
rect 15752 2204 15816 2208
rect 15752 2148 15756 2204
rect 15756 2148 15812 2204
rect 15812 2148 15816 2204
rect 15752 2144 15816 2148
rect 18612 2204 18676 2208
rect 18612 2148 18616 2204
rect 18616 2148 18672 2204
rect 18672 2148 18676 2204
rect 18612 2144 18676 2148
rect 18692 2204 18756 2208
rect 18692 2148 18696 2204
rect 18696 2148 18752 2204
rect 18752 2148 18756 2204
rect 18692 2144 18756 2148
rect 18772 2204 18836 2208
rect 18772 2148 18776 2204
rect 18776 2148 18832 2204
rect 18832 2148 18836 2204
rect 18772 2144 18836 2148
rect 18852 2204 18916 2208
rect 18852 2148 18856 2204
rect 18856 2148 18912 2204
rect 18912 2148 18916 2204
rect 18852 2144 18916 2148
rect 16252 2000 16316 2004
rect 16252 1944 16302 2000
rect 16302 1944 16316 2000
rect 16252 1940 16316 1944
rect 4662 1660 4726 1664
rect 4662 1604 4666 1660
rect 4666 1604 4722 1660
rect 4722 1604 4726 1660
rect 4662 1600 4726 1604
rect 4742 1660 4806 1664
rect 4742 1604 4746 1660
rect 4746 1604 4802 1660
rect 4802 1604 4806 1660
rect 4742 1600 4806 1604
rect 4822 1660 4886 1664
rect 4822 1604 4826 1660
rect 4826 1604 4882 1660
rect 4882 1604 4886 1660
rect 4822 1600 4886 1604
rect 4902 1660 4966 1664
rect 4902 1604 4906 1660
rect 4906 1604 4962 1660
rect 4962 1604 4966 1660
rect 4902 1600 4966 1604
rect 7762 1660 7826 1664
rect 7762 1604 7766 1660
rect 7766 1604 7822 1660
rect 7822 1604 7826 1660
rect 7762 1600 7826 1604
rect 7842 1660 7906 1664
rect 7842 1604 7846 1660
rect 7846 1604 7902 1660
rect 7902 1604 7906 1660
rect 7842 1600 7906 1604
rect 7922 1660 7986 1664
rect 7922 1604 7926 1660
rect 7926 1604 7982 1660
rect 7982 1604 7986 1660
rect 7922 1600 7986 1604
rect 8002 1660 8066 1664
rect 8002 1604 8006 1660
rect 8006 1604 8062 1660
rect 8062 1604 8066 1660
rect 8002 1600 8066 1604
rect 10862 1660 10926 1664
rect 10862 1604 10866 1660
rect 10866 1604 10922 1660
rect 10922 1604 10926 1660
rect 10862 1600 10926 1604
rect 10942 1660 11006 1664
rect 10942 1604 10946 1660
rect 10946 1604 11002 1660
rect 11002 1604 11006 1660
rect 10942 1600 11006 1604
rect 11022 1660 11086 1664
rect 11022 1604 11026 1660
rect 11026 1604 11082 1660
rect 11082 1604 11086 1660
rect 11022 1600 11086 1604
rect 11102 1660 11166 1664
rect 11102 1604 11106 1660
rect 11106 1604 11162 1660
rect 11162 1604 11166 1660
rect 11102 1600 11166 1604
rect 13962 1660 14026 1664
rect 13962 1604 13966 1660
rect 13966 1604 14022 1660
rect 14022 1604 14026 1660
rect 13962 1600 14026 1604
rect 14042 1660 14106 1664
rect 14042 1604 14046 1660
rect 14046 1604 14102 1660
rect 14102 1604 14106 1660
rect 14042 1600 14106 1604
rect 14122 1660 14186 1664
rect 14122 1604 14126 1660
rect 14126 1604 14182 1660
rect 14182 1604 14186 1660
rect 14122 1600 14186 1604
rect 14202 1660 14266 1664
rect 14202 1604 14206 1660
rect 14206 1604 14262 1660
rect 14262 1604 14266 1660
rect 14202 1600 14266 1604
rect 17062 1660 17126 1664
rect 17062 1604 17066 1660
rect 17066 1604 17122 1660
rect 17122 1604 17126 1660
rect 17062 1600 17126 1604
rect 17142 1660 17206 1664
rect 17142 1604 17146 1660
rect 17146 1604 17202 1660
rect 17202 1604 17206 1660
rect 17142 1600 17206 1604
rect 17222 1660 17286 1664
rect 17222 1604 17226 1660
rect 17226 1604 17282 1660
rect 17282 1604 17286 1660
rect 17222 1600 17286 1604
rect 17302 1660 17366 1664
rect 17302 1604 17306 1660
rect 17306 1604 17362 1660
rect 17362 1604 17366 1660
rect 17302 1600 17366 1604
rect 17540 1260 17604 1324
rect 3112 1116 3176 1120
rect 3112 1060 3116 1116
rect 3116 1060 3172 1116
rect 3172 1060 3176 1116
rect 3112 1056 3176 1060
rect 3192 1116 3256 1120
rect 3192 1060 3196 1116
rect 3196 1060 3252 1116
rect 3252 1060 3256 1116
rect 3192 1056 3256 1060
rect 3272 1116 3336 1120
rect 3272 1060 3276 1116
rect 3276 1060 3332 1116
rect 3332 1060 3336 1116
rect 3272 1056 3336 1060
rect 3352 1116 3416 1120
rect 3352 1060 3356 1116
rect 3356 1060 3412 1116
rect 3412 1060 3416 1116
rect 3352 1056 3416 1060
rect 6212 1116 6276 1120
rect 6212 1060 6216 1116
rect 6216 1060 6272 1116
rect 6272 1060 6276 1116
rect 6212 1056 6276 1060
rect 6292 1116 6356 1120
rect 6292 1060 6296 1116
rect 6296 1060 6352 1116
rect 6352 1060 6356 1116
rect 6292 1056 6356 1060
rect 6372 1116 6436 1120
rect 6372 1060 6376 1116
rect 6376 1060 6432 1116
rect 6432 1060 6436 1116
rect 6372 1056 6436 1060
rect 6452 1116 6516 1120
rect 6452 1060 6456 1116
rect 6456 1060 6512 1116
rect 6512 1060 6516 1116
rect 6452 1056 6516 1060
rect 9312 1116 9376 1120
rect 9312 1060 9316 1116
rect 9316 1060 9372 1116
rect 9372 1060 9376 1116
rect 9312 1056 9376 1060
rect 9392 1116 9456 1120
rect 9392 1060 9396 1116
rect 9396 1060 9452 1116
rect 9452 1060 9456 1116
rect 9392 1056 9456 1060
rect 9472 1116 9536 1120
rect 9472 1060 9476 1116
rect 9476 1060 9532 1116
rect 9532 1060 9536 1116
rect 9472 1056 9536 1060
rect 9552 1116 9616 1120
rect 9552 1060 9556 1116
rect 9556 1060 9612 1116
rect 9612 1060 9616 1116
rect 9552 1056 9616 1060
rect 12412 1116 12476 1120
rect 12412 1060 12416 1116
rect 12416 1060 12472 1116
rect 12472 1060 12476 1116
rect 12412 1056 12476 1060
rect 12492 1116 12556 1120
rect 12492 1060 12496 1116
rect 12496 1060 12552 1116
rect 12552 1060 12556 1116
rect 12492 1056 12556 1060
rect 12572 1116 12636 1120
rect 12572 1060 12576 1116
rect 12576 1060 12632 1116
rect 12632 1060 12636 1116
rect 12572 1056 12636 1060
rect 12652 1116 12716 1120
rect 12652 1060 12656 1116
rect 12656 1060 12712 1116
rect 12712 1060 12716 1116
rect 12652 1056 12716 1060
rect 15512 1116 15576 1120
rect 15512 1060 15516 1116
rect 15516 1060 15572 1116
rect 15572 1060 15576 1116
rect 15512 1056 15576 1060
rect 15592 1116 15656 1120
rect 15592 1060 15596 1116
rect 15596 1060 15652 1116
rect 15652 1060 15656 1116
rect 15592 1056 15656 1060
rect 15672 1116 15736 1120
rect 15672 1060 15676 1116
rect 15676 1060 15732 1116
rect 15732 1060 15736 1116
rect 15672 1056 15736 1060
rect 15752 1116 15816 1120
rect 15752 1060 15756 1116
rect 15756 1060 15812 1116
rect 15812 1060 15816 1116
rect 15752 1056 15816 1060
rect 18612 1116 18676 1120
rect 18612 1060 18616 1116
rect 18616 1060 18672 1116
rect 18672 1060 18676 1116
rect 18612 1056 18676 1060
rect 18692 1116 18756 1120
rect 18692 1060 18696 1116
rect 18696 1060 18752 1116
rect 18752 1060 18756 1116
rect 18692 1056 18756 1060
rect 18772 1116 18836 1120
rect 18772 1060 18776 1116
rect 18776 1060 18832 1116
rect 18832 1060 18836 1116
rect 18772 1056 18836 1060
rect 18852 1116 18916 1120
rect 18852 1060 18856 1116
rect 18856 1060 18912 1116
rect 18912 1060 18916 1116
rect 18852 1056 18916 1060
rect 14412 988 14476 1052
rect 4662 572 4726 576
rect 4662 516 4666 572
rect 4666 516 4722 572
rect 4722 516 4726 572
rect 4662 512 4726 516
rect 4742 572 4806 576
rect 4742 516 4746 572
rect 4746 516 4802 572
rect 4802 516 4806 572
rect 4742 512 4806 516
rect 4822 572 4886 576
rect 4822 516 4826 572
rect 4826 516 4882 572
rect 4882 516 4886 572
rect 4822 512 4886 516
rect 4902 572 4966 576
rect 4902 516 4906 572
rect 4906 516 4962 572
rect 4962 516 4966 572
rect 4902 512 4966 516
rect 7762 572 7826 576
rect 7762 516 7766 572
rect 7766 516 7822 572
rect 7822 516 7826 572
rect 7762 512 7826 516
rect 7842 572 7906 576
rect 7842 516 7846 572
rect 7846 516 7902 572
rect 7902 516 7906 572
rect 7842 512 7906 516
rect 7922 572 7986 576
rect 7922 516 7926 572
rect 7926 516 7982 572
rect 7982 516 7986 572
rect 7922 512 7986 516
rect 8002 572 8066 576
rect 8002 516 8006 572
rect 8006 516 8062 572
rect 8062 516 8066 572
rect 8002 512 8066 516
rect 10862 572 10926 576
rect 10862 516 10866 572
rect 10866 516 10922 572
rect 10922 516 10926 572
rect 10862 512 10926 516
rect 10942 572 11006 576
rect 10942 516 10946 572
rect 10946 516 11002 572
rect 11002 516 11006 572
rect 10942 512 11006 516
rect 11022 572 11086 576
rect 11022 516 11026 572
rect 11026 516 11082 572
rect 11082 516 11086 572
rect 11022 512 11086 516
rect 11102 572 11166 576
rect 11102 516 11106 572
rect 11106 516 11162 572
rect 11162 516 11166 572
rect 11102 512 11166 516
rect 13962 572 14026 576
rect 13962 516 13966 572
rect 13966 516 14022 572
rect 14022 516 14026 572
rect 13962 512 14026 516
rect 14042 572 14106 576
rect 14042 516 14046 572
rect 14046 516 14102 572
rect 14102 516 14106 572
rect 14042 512 14106 516
rect 14122 572 14186 576
rect 14122 516 14126 572
rect 14126 516 14182 572
rect 14182 516 14186 572
rect 14122 512 14186 516
rect 14202 572 14266 576
rect 14202 516 14206 572
rect 14206 516 14262 572
rect 14262 516 14266 572
rect 14202 512 14266 516
rect 17062 572 17126 576
rect 17062 516 17066 572
rect 17066 516 17122 572
rect 17122 516 17126 572
rect 17062 512 17126 516
rect 17142 572 17206 576
rect 17142 516 17146 572
rect 17146 516 17202 572
rect 17202 516 17206 572
rect 17142 512 17206 516
rect 17222 572 17286 576
rect 17222 516 17226 572
rect 17226 516 17282 572
rect 17282 516 17286 572
rect 17222 512 17286 516
rect 17302 572 17366 576
rect 17302 516 17306 572
rect 17306 516 17362 572
rect 17362 516 17366 572
rect 17302 512 17366 516
<< metal4 >>
rect 3104 10912 3424 10928
rect 3104 10848 3112 10912
rect 3176 10848 3192 10912
rect 3256 10848 3272 10912
rect 3336 10848 3352 10912
rect 3416 10848 3424 10912
rect 3104 10160 3424 10848
rect 3104 9924 3146 10160
rect 3382 9924 3424 10160
rect 3104 9824 3424 9924
rect 3104 9760 3112 9824
rect 3176 9760 3192 9824
rect 3256 9760 3272 9824
rect 3336 9760 3352 9824
rect 3416 9760 3424 9824
rect 3104 8736 3424 9760
rect 3104 8672 3112 8736
rect 3176 8672 3192 8736
rect 3256 8672 3272 8736
rect 3336 8672 3352 8736
rect 3416 8672 3424 8736
rect 3104 7648 3424 8672
rect 3104 7584 3112 7648
rect 3176 7584 3192 7648
rect 3256 7584 3272 7648
rect 3336 7584 3352 7648
rect 3416 7584 3424 7648
rect 3104 6780 3424 7584
rect 3104 6560 3146 6780
rect 3382 6560 3424 6780
rect 3104 6496 3112 6560
rect 3176 6496 3192 6544
rect 3256 6496 3272 6544
rect 3336 6496 3352 6544
rect 3416 6496 3424 6560
rect 3104 5472 3424 6496
rect 3104 5408 3112 5472
rect 3176 5408 3192 5472
rect 3256 5408 3272 5472
rect 3336 5408 3352 5472
rect 3416 5408 3424 5472
rect 3104 4384 3424 5408
rect 3104 4320 3112 4384
rect 3176 4320 3192 4384
rect 3256 4320 3272 4384
rect 3336 4320 3352 4384
rect 3416 4320 3424 4384
rect 3104 3400 3424 4320
rect 3104 3296 3146 3400
rect 3382 3296 3424 3400
rect 3104 3232 3112 3296
rect 3416 3232 3424 3296
rect 3104 3164 3146 3232
rect 3382 3164 3424 3232
rect 3104 2208 3424 3164
rect 3104 2144 3112 2208
rect 3176 2144 3192 2208
rect 3256 2144 3272 2208
rect 3336 2144 3352 2208
rect 3416 2144 3424 2208
rect 3104 1120 3424 2144
rect 3104 1056 3112 1120
rect 3176 1056 3192 1120
rect 3256 1056 3272 1120
rect 3336 1056 3352 1120
rect 3416 1056 3424 1120
rect 3104 496 3424 1056
rect 4654 10368 4974 10928
rect 4654 10304 4662 10368
rect 4726 10304 4742 10368
rect 4806 10304 4822 10368
rect 4886 10304 4902 10368
rect 4966 10304 4974 10368
rect 4654 9280 4974 10304
rect 4654 9216 4662 9280
rect 4726 9216 4742 9280
rect 4806 9216 4822 9280
rect 4886 9216 4902 9280
rect 4966 9216 4974 9280
rect 4654 8470 4974 9216
rect 4654 8234 4696 8470
rect 4932 8234 4974 8470
rect 4654 8192 4974 8234
rect 4654 8128 4662 8192
rect 4726 8128 4742 8192
rect 4806 8128 4822 8192
rect 4886 8128 4902 8192
rect 4966 8128 4974 8192
rect 4654 7104 4974 8128
rect 4654 7040 4662 7104
rect 4726 7040 4742 7104
rect 4806 7040 4822 7104
rect 4886 7040 4902 7104
rect 4966 7040 4974 7104
rect 4654 6016 4974 7040
rect 4654 5952 4662 6016
rect 4726 5952 4742 6016
rect 4806 5952 4822 6016
rect 4886 5952 4902 6016
rect 4966 5952 4974 6016
rect 4654 5090 4974 5952
rect 4654 4928 4696 5090
rect 4932 4928 4974 5090
rect 4654 4864 4662 4928
rect 4966 4864 4974 4928
rect 4654 4854 4696 4864
rect 4932 4854 4974 4864
rect 4654 3840 4974 4854
rect 4654 3776 4662 3840
rect 4726 3776 4742 3840
rect 4806 3776 4822 3840
rect 4886 3776 4902 3840
rect 4966 3776 4974 3840
rect 4654 2752 4974 3776
rect 4654 2688 4662 2752
rect 4726 2688 4742 2752
rect 4806 2688 4822 2752
rect 4886 2688 4902 2752
rect 4966 2688 4974 2752
rect 4654 1664 4974 2688
rect 4654 1600 4662 1664
rect 4726 1600 4742 1664
rect 4806 1600 4822 1664
rect 4886 1600 4902 1664
rect 4966 1600 4974 1664
rect 4654 576 4974 1600
rect 4654 512 4662 576
rect 4726 512 4742 576
rect 4806 512 4822 576
rect 4886 512 4902 576
rect 4966 512 4974 576
rect 4654 496 4974 512
rect 6204 10912 6524 10928
rect 6204 10848 6212 10912
rect 6276 10848 6292 10912
rect 6356 10848 6372 10912
rect 6436 10848 6452 10912
rect 6516 10848 6524 10912
rect 6204 10160 6524 10848
rect 6204 9924 6246 10160
rect 6482 9924 6524 10160
rect 6204 9824 6524 9924
rect 6204 9760 6212 9824
rect 6276 9760 6292 9824
rect 6356 9760 6372 9824
rect 6436 9760 6452 9824
rect 6516 9760 6524 9824
rect 6204 8736 6524 9760
rect 6204 8672 6212 8736
rect 6276 8672 6292 8736
rect 6356 8672 6372 8736
rect 6436 8672 6452 8736
rect 6516 8672 6524 8736
rect 6204 7648 6524 8672
rect 6204 7584 6212 7648
rect 6276 7584 6292 7648
rect 6356 7584 6372 7648
rect 6436 7584 6452 7648
rect 6516 7584 6524 7648
rect 6204 6780 6524 7584
rect 6204 6560 6246 6780
rect 6482 6560 6524 6780
rect 6204 6496 6212 6560
rect 6276 6496 6292 6544
rect 6356 6496 6372 6544
rect 6436 6496 6452 6544
rect 6516 6496 6524 6560
rect 6204 5472 6524 6496
rect 6204 5408 6212 5472
rect 6276 5408 6292 5472
rect 6356 5408 6372 5472
rect 6436 5408 6452 5472
rect 6516 5408 6524 5472
rect 6204 4384 6524 5408
rect 6204 4320 6212 4384
rect 6276 4320 6292 4384
rect 6356 4320 6372 4384
rect 6436 4320 6452 4384
rect 6516 4320 6524 4384
rect 6204 3400 6524 4320
rect 6204 3296 6246 3400
rect 6482 3296 6524 3400
rect 6204 3232 6212 3296
rect 6516 3232 6524 3296
rect 6204 3164 6246 3232
rect 6482 3164 6524 3232
rect 6204 2208 6524 3164
rect 6204 2144 6212 2208
rect 6276 2144 6292 2208
rect 6356 2144 6372 2208
rect 6436 2144 6452 2208
rect 6516 2144 6524 2208
rect 6204 1120 6524 2144
rect 6204 1056 6212 1120
rect 6276 1056 6292 1120
rect 6356 1056 6372 1120
rect 6436 1056 6452 1120
rect 6516 1056 6524 1120
rect 6204 496 6524 1056
rect 7754 10368 8074 10928
rect 7754 10304 7762 10368
rect 7826 10304 7842 10368
rect 7906 10304 7922 10368
rect 7986 10304 8002 10368
rect 8066 10304 8074 10368
rect 7754 9280 8074 10304
rect 7754 9216 7762 9280
rect 7826 9216 7842 9280
rect 7906 9216 7922 9280
rect 7986 9216 8002 9280
rect 8066 9216 8074 9280
rect 7754 8470 8074 9216
rect 7754 8234 7796 8470
rect 8032 8234 8074 8470
rect 7754 8192 8074 8234
rect 7754 8128 7762 8192
rect 7826 8128 7842 8192
rect 7906 8128 7922 8192
rect 7986 8128 8002 8192
rect 8066 8128 8074 8192
rect 7754 7104 8074 8128
rect 7754 7040 7762 7104
rect 7826 7040 7842 7104
rect 7906 7040 7922 7104
rect 7986 7040 8002 7104
rect 8066 7040 8074 7104
rect 7754 6016 8074 7040
rect 7754 5952 7762 6016
rect 7826 5952 7842 6016
rect 7906 5952 7922 6016
rect 7986 5952 8002 6016
rect 8066 5952 8074 6016
rect 7754 5090 8074 5952
rect 7754 4928 7796 5090
rect 8032 4928 8074 5090
rect 7754 4864 7762 4928
rect 8066 4864 8074 4928
rect 7754 4854 7796 4864
rect 8032 4854 8074 4864
rect 7754 3840 8074 4854
rect 7754 3776 7762 3840
rect 7826 3776 7842 3840
rect 7906 3776 7922 3840
rect 7986 3776 8002 3840
rect 8066 3776 8074 3840
rect 7754 2752 8074 3776
rect 7754 2688 7762 2752
rect 7826 2688 7842 2752
rect 7906 2688 7922 2752
rect 7986 2688 8002 2752
rect 8066 2688 8074 2752
rect 7754 1664 8074 2688
rect 7754 1600 7762 1664
rect 7826 1600 7842 1664
rect 7906 1600 7922 1664
rect 7986 1600 8002 1664
rect 8066 1600 8074 1664
rect 7754 576 8074 1600
rect 7754 512 7762 576
rect 7826 512 7842 576
rect 7906 512 7922 576
rect 7986 512 8002 576
rect 8066 512 8074 576
rect 7754 496 8074 512
rect 9304 10912 9624 10928
rect 9304 10848 9312 10912
rect 9376 10848 9392 10912
rect 9456 10848 9472 10912
rect 9536 10848 9552 10912
rect 9616 10848 9624 10912
rect 9304 10160 9624 10848
rect 9304 9924 9346 10160
rect 9582 9924 9624 10160
rect 9304 9824 9624 9924
rect 9304 9760 9312 9824
rect 9376 9760 9392 9824
rect 9456 9760 9472 9824
rect 9536 9760 9552 9824
rect 9616 9760 9624 9824
rect 9304 8736 9624 9760
rect 9304 8672 9312 8736
rect 9376 8672 9392 8736
rect 9456 8672 9472 8736
rect 9536 8672 9552 8736
rect 9616 8672 9624 8736
rect 9304 7648 9624 8672
rect 9304 7584 9312 7648
rect 9376 7584 9392 7648
rect 9456 7584 9472 7648
rect 9536 7584 9552 7648
rect 9616 7584 9624 7648
rect 9304 6780 9624 7584
rect 9304 6560 9346 6780
rect 9582 6560 9624 6780
rect 9304 6496 9312 6560
rect 9376 6496 9392 6544
rect 9456 6496 9472 6544
rect 9536 6496 9552 6544
rect 9616 6496 9624 6560
rect 9304 5472 9624 6496
rect 9304 5408 9312 5472
rect 9376 5408 9392 5472
rect 9456 5408 9472 5472
rect 9536 5408 9552 5472
rect 9616 5408 9624 5472
rect 9304 4384 9624 5408
rect 9304 4320 9312 4384
rect 9376 4320 9392 4384
rect 9456 4320 9472 4384
rect 9536 4320 9552 4384
rect 9616 4320 9624 4384
rect 9304 3400 9624 4320
rect 9304 3296 9346 3400
rect 9582 3296 9624 3400
rect 9304 3232 9312 3296
rect 9616 3232 9624 3296
rect 9304 3164 9346 3232
rect 9582 3164 9624 3232
rect 9304 2208 9624 3164
rect 9304 2144 9312 2208
rect 9376 2144 9392 2208
rect 9456 2144 9472 2208
rect 9536 2144 9552 2208
rect 9616 2144 9624 2208
rect 9304 1120 9624 2144
rect 9304 1056 9312 1120
rect 9376 1056 9392 1120
rect 9456 1056 9472 1120
rect 9536 1056 9552 1120
rect 9616 1056 9624 1120
rect 9304 496 9624 1056
rect 10854 10368 11174 10928
rect 10854 10304 10862 10368
rect 10926 10304 10942 10368
rect 11006 10304 11022 10368
rect 11086 10304 11102 10368
rect 11166 10304 11174 10368
rect 10854 9280 11174 10304
rect 10854 9216 10862 9280
rect 10926 9216 10942 9280
rect 11006 9216 11022 9280
rect 11086 9216 11102 9280
rect 11166 9216 11174 9280
rect 10854 8470 11174 9216
rect 10854 8234 10896 8470
rect 11132 8234 11174 8470
rect 10854 8192 11174 8234
rect 10854 8128 10862 8192
rect 10926 8128 10942 8192
rect 11006 8128 11022 8192
rect 11086 8128 11102 8192
rect 11166 8128 11174 8192
rect 10854 7104 11174 8128
rect 10854 7040 10862 7104
rect 10926 7040 10942 7104
rect 11006 7040 11022 7104
rect 11086 7040 11102 7104
rect 11166 7040 11174 7104
rect 10854 6016 11174 7040
rect 10854 5952 10862 6016
rect 10926 5952 10942 6016
rect 11006 5952 11022 6016
rect 11086 5952 11102 6016
rect 11166 5952 11174 6016
rect 10854 5090 11174 5952
rect 10854 4928 10896 5090
rect 11132 4928 11174 5090
rect 10854 4864 10862 4928
rect 11166 4864 11174 4928
rect 10854 4854 10896 4864
rect 11132 4854 11174 4864
rect 10854 3840 11174 4854
rect 10854 3776 10862 3840
rect 10926 3776 10942 3840
rect 11006 3776 11022 3840
rect 11086 3776 11102 3840
rect 11166 3776 11174 3840
rect 10854 2752 11174 3776
rect 10854 2688 10862 2752
rect 10926 2688 10942 2752
rect 11006 2688 11022 2752
rect 11086 2688 11102 2752
rect 11166 2688 11174 2752
rect 10854 1664 11174 2688
rect 10854 1600 10862 1664
rect 10926 1600 10942 1664
rect 11006 1600 11022 1664
rect 11086 1600 11102 1664
rect 11166 1600 11174 1664
rect 10854 576 11174 1600
rect 10854 512 10862 576
rect 10926 512 10942 576
rect 11006 512 11022 576
rect 11086 512 11102 576
rect 11166 512 11174 576
rect 10854 496 11174 512
rect 12404 10912 12724 10928
rect 12404 10848 12412 10912
rect 12476 10848 12492 10912
rect 12556 10848 12572 10912
rect 12636 10848 12652 10912
rect 12716 10848 12724 10912
rect 12404 10160 12724 10848
rect 12404 9924 12446 10160
rect 12682 9924 12724 10160
rect 12404 9824 12724 9924
rect 12404 9760 12412 9824
rect 12476 9760 12492 9824
rect 12556 9760 12572 9824
rect 12636 9760 12652 9824
rect 12716 9760 12724 9824
rect 12404 8736 12724 9760
rect 12404 8672 12412 8736
rect 12476 8672 12492 8736
rect 12556 8672 12572 8736
rect 12636 8672 12652 8736
rect 12716 8672 12724 8736
rect 12404 7648 12724 8672
rect 12404 7584 12412 7648
rect 12476 7584 12492 7648
rect 12556 7584 12572 7648
rect 12636 7584 12652 7648
rect 12716 7584 12724 7648
rect 12404 6780 12724 7584
rect 12404 6560 12446 6780
rect 12682 6560 12724 6780
rect 12404 6496 12412 6560
rect 12476 6496 12492 6544
rect 12556 6496 12572 6544
rect 12636 6496 12652 6544
rect 12716 6496 12724 6560
rect 12404 5472 12724 6496
rect 12404 5408 12412 5472
rect 12476 5408 12492 5472
rect 12556 5408 12572 5472
rect 12636 5408 12652 5472
rect 12716 5408 12724 5472
rect 12404 4384 12724 5408
rect 12404 4320 12412 4384
rect 12476 4320 12492 4384
rect 12556 4320 12572 4384
rect 12636 4320 12652 4384
rect 12716 4320 12724 4384
rect 12404 3400 12724 4320
rect 12404 3296 12446 3400
rect 12682 3296 12724 3400
rect 12404 3232 12412 3296
rect 12716 3232 12724 3296
rect 12404 3164 12446 3232
rect 12682 3164 12724 3232
rect 12404 2208 12724 3164
rect 12404 2144 12412 2208
rect 12476 2144 12492 2208
rect 12556 2144 12572 2208
rect 12636 2144 12652 2208
rect 12716 2144 12724 2208
rect 12404 1120 12724 2144
rect 12404 1056 12412 1120
rect 12476 1056 12492 1120
rect 12556 1056 12572 1120
rect 12636 1056 12652 1120
rect 12716 1056 12724 1120
rect 12404 496 12724 1056
rect 13954 10368 14274 10928
rect 13954 10304 13962 10368
rect 14026 10304 14042 10368
rect 14106 10304 14122 10368
rect 14186 10304 14202 10368
rect 14266 10304 14274 10368
rect 13954 9280 14274 10304
rect 13954 9216 13962 9280
rect 14026 9216 14042 9280
rect 14106 9216 14122 9280
rect 14186 9216 14202 9280
rect 14266 9216 14274 9280
rect 13954 8470 14274 9216
rect 13954 8234 13996 8470
rect 14232 8234 14274 8470
rect 13954 8192 14274 8234
rect 13954 8128 13962 8192
rect 14026 8128 14042 8192
rect 14106 8128 14122 8192
rect 14186 8128 14202 8192
rect 14266 8128 14274 8192
rect 13954 7104 14274 8128
rect 13954 7040 13962 7104
rect 14026 7040 14042 7104
rect 14106 7040 14122 7104
rect 14186 7040 14202 7104
rect 14266 7040 14274 7104
rect 13954 6016 14274 7040
rect 13954 5952 13962 6016
rect 14026 5952 14042 6016
rect 14106 5952 14122 6016
rect 14186 5952 14202 6016
rect 14266 5952 14274 6016
rect 13954 5090 14274 5952
rect 13954 4928 13996 5090
rect 14232 4928 14274 5090
rect 13954 4864 13962 4928
rect 14266 4864 14274 4928
rect 13954 4854 13996 4864
rect 14232 4854 14274 4864
rect 13954 3840 14274 4854
rect 13954 3776 13962 3840
rect 14026 3776 14042 3840
rect 14106 3776 14122 3840
rect 14186 3776 14202 3840
rect 14266 3776 14274 3840
rect 13954 2752 14274 3776
rect 13954 2688 13962 2752
rect 14026 2688 14042 2752
rect 14106 2688 14122 2752
rect 14186 2688 14202 2752
rect 14266 2688 14274 2752
rect 13954 1664 14274 2688
rect 15504 10912 15824 10928
rect 15504 10848 15512 10912
rect 15576 10848 15592 10912
rect 15656 10848 15672 10912
rect 15736 10848 15752 10912
rect 15816 10848 15824 10912
rect 15504 10160 15824 10848
rect 15504 9924 15546 10160
rect 15782 9924 15824 10160
rect 15504 9824 15824 9924
rect 15504 9760 15512 9824
rect 15576 9760 15592 9824
rect 15656 9760 15672 9824
rect 15736 9760 15752 9824
rect 15816 9760 15824 9824
rect 15504 8736 15824 9760
rect 15504 8672 15512 8736
rect 15576 8672 15592 8736
rect 15656 8672 15672 8736
rect 15736 8672 15752 8736
rect 15816 8672 15824 8736
rect 15504 7648 15824 8672
rect 17054 10368 17374 10928
rect 17054 10304 17062 10368
rect 17126 10304 17142 10368
rect 17206 10304 17222 10368
rect 17286 10304 17302 10368
rect 17366 10304 17374 10368
rect 17054 9280 17374 10304
rect 17054 9216 17062 9280
rect 17126 9216 17142 9280
rect 17206 9216 17222 9280
rect 17286 9216 17302 9280
rect 17366 9216 17374 9280
rect 16803 8532 16869 8533
rect 16803 8468 16804 8532
rect 16868 8468 16869 8532
rect 16803 8467 16869 8468
rect 17054 8470 17374 9216
rect 15504 7584 15512 7648
rect 15576 7584 15592 7648
rect 15656 7584 15672 7648
rect 15736 7584 15752 7648
rect 15816 7584 15824 7648
rect 15504 6780 15824 7584
rect 16067 7444 16133 7445
rect 16067 7380 16068 7444
rect 16132 7380 16133 7444
rect 16067 7379 16133 7380
rect 15504 6560 15546 6780
rect 15782 6560 15824 6780
rect 15504 6496 15512 6560
rect 15576 6496 15592 6544
rect 15656 6496 15672 6544
rect 15736 6496 15752 6544
rect 15816 6496 15824 6560
rect 15504 5472 15824 6496
rect 15504 5408 15512 5472
rect 15576 5408 15592 5472
rect 15656 5408 15672 5472
rect 15736 5408 15752 5472
rect 15816 5408 15824 5472
rect 15504 4384 15824 5408
rect 16070 5269 16130 7379
rect 16806 7309 16866 8467
rect 17054 8234 17096 8470
rect 17332 8234 17374 8470
rect 17054 8192 17374 8234
rect 17054 8128 17062 8192
rect 17126 8128 17142 8192
rect 17206 8128 17222 8192
rect 17286 8128 17302 8192
rect 17366 8128 17374 8192
rect 16803 7308 16869 7309
rect 16803 7244 16804 7308
rect 16868 7244 16869 7308
rect 16803 7243 16869 7244
rect 16435 6764 16501 6765
rect 16435 6700 16436 6764
rect 16500 6700 16501 6764
rect 16435 6699 16501 6700
rect 16067 5268 16133 5269
rect 16067 5204 16068 5268
rect 16132 5204 16133 5268
rect 16067 5203 16133 5204
rect 16251 4452 16317 4453
rect 16251 4388 16252 4452
rect 16316 4388 16317 4452
rect 16251 4387 16317 4388
rect 15504 4320 15512 4384
rect 15576 4320 15592 4384
rect 15656 4320 15672 4384
rect 15736 4320 15752 4384
rect 15816 4320 15824 4384
rect 15504 3400 15824 4320
rect 15504 3296 15546 3400
rect 15782 3296 15824 3400
rect 15504 3232 15512 3296
rect 15816 3232 15824 3296
rect 15504 3164 15546 3232
rect 15782 3164 15824 3232
rect 14411 2548 14477 2549
rect 14411 2484 14412 2548
rect 14476 2484 14477 2548
rect 14411 2483 14477 2484
rect 13954 1600 13962 1664
rect 14026 1600 14042 1664
rect 14106 1600 14122 1664
rect 14186 1600 14202 1664
rect 14266 1600 14274 1664
rect 13954 576 14274 1600
rect 14414 1053 14474 2483
rect 15504 2208 15824 3164
rect 15504 2144 15512 2208
rect 15576 2144 15592 2208
rect 15656 2144 15672 2208
rect 15736 2144 15752 2208
rect 15816 2144 15824 2208
rect 15504 1120 15824 2144
rect 16254 2005 16314 4387
rect 16438 3365 16498 6699
rect 16806 5269 16866 7243
rect 17054 7104 17374 8128
rect 17054 7040 17062 7104
rect 17126 7040 17142 7104
rect 17206 7040 17222 7104
rect 17286 7040 17302 7104
rect 17366 7040 17374 7104
rect 17054 6016 17374 7040
rect 17054 5952 17062 6016
rect 17126 5952 17142 6016
rect 17206 5952 17222 6016
rect 17286 5952 17302 6016
rect 17366 5952 17374 6016
rect 16803 5268 16869 5269
rect 16803 5204 16804 5268
rect 16868 5204 16869 5268
rect 16803 5203 16869 5204
rect 17054 5090 17374 5952
rect 18604 10912 18924 10928
rect 18604 10848 18612 10912
rect 18676 10848 18692 10912
rect 18756 10848 18772 10912
rect 18836 10848 18852 10912
rect 18916 10848 18924 10912
rect 18604 10160 18924 10848
rect 18604 9924 18646 10160
rect 18882 9924 18924 10160
rect 18604 9824 18924 9924
rect 18604 9760 18612 9824
rect 18676 9760 18692 9824
rect 18756 9760 18772 9824
rect 18836 9760 18852 9824
rect 18916 9760 18924 9824
rect 18604 8736 18924 9760
rect 18604 8672 18612 8736
rect 18676 8672 18692 8736
rect 18756 8672 18772 8736
rect 18836 8672 18852 8736
rect 18916 8672 18924 8736
rect 18604 7648 18924 8672
rect 18604 7584 18612 7648
rect 18676 7584 18692 7648
rect 18756 7584 18772 7648
rect 18836 7584 18852 7648
rect 18916 7584 18924 7648
rect 18604 6780 18924 7584
rect 18604 6560 18646 6780
rect 18882 6560 18924 6780
rect 18604 6496 18612 6560
rect 18676 6496 18692 6544
rect 18756 6496 18772 6544
rect 18836 6496 18852 6544
rect 18916 6496 18924 6560
rect 17539 5540 17605 5541
rect 17539 5476 17540 5540
rect 17604 5476 17605 5540
rect 17539 5475 17605 5476
rect 17054 4928 17096 5090
rect 17332 4928 17374 5090
rect 17054 4864 17062 4928
rect 17366 4864 17374 4928
rect 17054 4854 17096 4864
rect 17332 4854 17374 4864
rect 17054 3840 17374 4854
rect 17054 3776 17062 3840
rect 17126 3776 17142 3840
rect 17206 3776 17222 3840
rect 17286 3776 17302 3840
rect 17366 3776 17374 3840
rect 16435 3364 16501 3365
rect 16435 3300 16436 3364
rect 16500 3300 16501 3364
rect 16435 3299 16501 3300
rect 16619 2820 16685 2821
rect 16619 2756 16620 2820
rect 16684 2756 16685 2820
rect 16619 2755 16685 2756
rect 16622 2685 16682 2755
rect 17054 2752 17374 3776
rect 17054 2688 17062 2752
rect 17126 2688 17142 2752
rect 17206 2688 17222 2752
rect 17286 2688 17302 2752
rect 17366 2688 17374 2752
rect 16619 2684 16685 2685
rect 16619 2620 16620 2684
rect 16684 2620 16685 2684
rect 16619 2619 16685 2620
rect 16251 2004 16317 2005
rect 16251 1940 16252 2004
rect 16316 1940 16317 2004
rect 16251 1939 16317 1940
rect 15504 1056 15512 1120
rect 15576 1056 15592 1120
rect 15656 1056 15672 1120
rect 15736 1056 15752 1120
rect 15816 1056 15824 1120
rect 14411 1052 14477 1053
rect 14411 988 14412 1052
rect 14476 988 14477 1052
rect 14411 987 14477 988
rect 13954 512 13962 576
rect 14026 512 14042 576
rect 14106 512 14122 576
rect 14186 512 14202 576
rect 14266 512 14274 576
rect 13954 496 14274 512
rect 15504 496 15824 1056
rect 17054 1664 17374 2688
rect 17054 1600 17062 1664
rect 17126 1600 17142 1664
rect 17206 1600 17222 1664
rect 17286 1600 17302 1664
rect 17366 1600 17374 1664
rect 17054 576 17374 1600
rect 17542 1325 17602 5475
rect 18604 5472 18924 6496
rect 18604 5408 18612 5472
rect 18676 5408 18692 5472
rect 18756 5408 18772 5472
rect 18836 5408 18852 5472
rect 18916 5408 18924 5472
rect 18604 4384 18924 5408
rect 18604 4320 18612 4384
rect 18676 4320 18692 4384
rect 18756 4320 18772 4384
rect 18836 4320 18852 4384
rect 18916 4320 18924 4384
rect 18604 3400 18924 4320
rect 18604 3296 18646 3400
rect 18882 3296 18924 3400
rect 18604 3232 18612 3296
rect 18916 3232 18924 3296
rect 18604 3164 18646 3232
rect 18882 3164 18924 3232
rect 18604 2208 18924 3164
rect 18604 2144 18612 2208
rect 18676 2144 18692 2208
rect 18756 2144 18772 2208
rect 18836 2144 18852 2208
rect 18916 2144 18924 2208
rect 17539 1324 17605 1325
rect 17539 1260 17540 1324
rect 17604 1260 17605 1324
rect 17539 1259 17605 1260
rect 17054 512 17062 576
rect 17126 512 17142 576
rect 17206 512 17222 576
rect 17286 512 17302 576
rect 17366 512 17374 576
rect 17054 496 17374 512
rect 18604 1120 18924 2144
rect 18604 1056 18612 1120
rect 18676 1056 18692 1120
rect 18756 1056 18772 1120
rect 18836 1056 18852 1120
rect 18916 1056 18924 1120
rect 18604 496 18924 1056
<< via4 >>
rect 3146 9924 3382 10160
rect 3146 6560 3382 6780
rect 3146 6544 3176 6560
rect 3176 6544 3192 6560
rect 3192 6544 3256 6560
rect 3256 6544 3272 6560
rect 3272 6544 3336 6560
rect 3336 6544 3352 6560
rect 3352 6544 3382 6560
rect 3146 3296 3382 3400
rect 3146 3232 3176 3296
rect 3176 3232 3192 3296
rect 3192 3232 3256 3296
rect 3256 3232 3272 3296
rect 3272 3232 3336 3296
rect 3336 3232 3352 3296
rect 3352 3232 3382 3296
rect 3146 3164 3382 3232
rect 4696 8234 4932 8470
rect 4696 4928 4932 5090
rect 4696 4864 4726 4928
rect 4726 4864 4742 4928
rect 4742 4864 4806 4928
rect 4806 4864 4822 4928
rect 4822 4864 4886 4928
rect 4886 4864 4902 4928
rect 4902 4864 4932 4928
rect 4696 4854 4932 4864
rect 6246 9924 6482 10160
rect 6246 6560 6482 6780
rect 6246 6544 6276 6560
rect 6276 6544 6292 6560
rect 6292 6544 6356 6560
rect 6356 6544 6372 6560
rect 6372 6544 6436 6560
rect 6436 6544 6452 6560
rect 6452 6544 6482 6560
rect 6246 3296 6482 3400
rect 6246 3232 6276 3296
rect 6276 3232 6292 3296
rect 6292 3232 6356 3296
rect 6356 3232 6372 3296
rect 6372 3232 6436 3296
rect 6436 3232 6452 3296
rect 6452 3232 6482 3296
rect 6246 3164 6482 3232
rect 7796 8234 8032 8470
rect 7796 4928 8032 5090
rect 7796 4864 7826 4928
rect 7826 4864 7842 4928
rect 7842 4864 7906 4928
rect 7906 4864 7922 4928
rect 7922 4864 7986 4928
rect 7986 4864 8002 4928
rect 8002 4864 8032 4928
rect 7796 4854 8032 4864
rect 9346 9924 9582 10160
rect 9346 6560 9582 6780
rect 9346 6544 9376 6560
rect 9376 6544 9392 6560
rect 9392 6544 9456 6560
rect 9456 6544 9472 6560
rect 9472 6544 9536 6560
rect 9536 6544 9552 6560
rect 9552 6544 9582 6560
rect 9346 3296 9582 3400
rect 9346 3232 9376 3296
rect 9376 3232 9392 3296
rect 9392 3232 9456 3296
rect 9456 3232 9472 3296
rect 9472 3232 9536 3296
rect 9536 3232 9552 3296
rect 9552 3232 9582 3296
rect 9346 3164 9582 3232
rect 10896 8234 11132 8470
rect 10896 4928 11132 5090
rect 10896 4864 10926 4928
rect 10926 4864 10942 4928
rect 10942 4864 11006 4928
rect 11006 4864 11022 4928
rect 11022 4864 11086 4928
rect 11086 4864 11102 4928
rect 11102 4864 11132 4928
rect 10896 4854 11132 4864
rect 12446 9924 12682 10160
rect 12446 6560 12682 6780
rect 12446 6544 12476 6560
rect 12476 6544 12492 6560
rect 12492 6544 12556 6560
rect 12556 6544 12572 6560
rect 12572 6544 12636 6560
rect 12636 6544 12652 6560
rect 12652 6544 12682 6560
rect 12446 3296 12682 3400
rect 12446 3232 12476 3296
rect 12476 3232 12492 3296
rect 12492 3232 12556 3296
rect 12556 3232 12572 3296
rect 12572 3232 12636 3296
rect 12636 3232 12652 3296
rect 12652 3232 12682 3296
rect 12446 3164 12682 3232
rect 13996 8234 14232 8470
rect 13996 4928 14232 5090
rect 13996 4864 14026 4928
rect 14026 4864 14042 4928
rect 14042 4864 14106 4928
rect 14106 4864 14122 4928
rect 14122 4864 14186 4928
rect 14186 4864 14202 4928
rect 14202 4864 14232 4928
rect 13996 4854 14232 4864
rect 15546 9924 15782 10160
rect 15546 6560 15782 6780
rect 15546 6544 15576 6560
rect 15576 6544 15592 6560
rect 15592 6544 15656 6560
rect 15656 6544 15672 6560
rect 15672 6544 15736 6560
rect 15736 6544 15752 6560
rect 15752 6544 15782 6560
rect 17096 8234 17332 8470
rect 15546 3296 15782 3400
rect 15546 3232 15576 3296
rect 15576 3232 15592 3296
rect 15592 3232 15656 3296
rect 15656 3232 15672 3296
rect 15672 3232 15736 3296
rect 15736 3232 15752 3296
rect 15752 3232 15782 3296
rect 15546 3164 15782 3232
rect 18646 9924 18882 10160
rect 18646 6560 18882 6780
rect 18646 6544 18676 6560
rect 18676 6544 18692 6560
rect 18692 6544 18756 6560
rect 18756 6544 18772 6560
rect 18772 6544 18836 6560
rect 18836 6544 18852 6560
rect 18852 6544 18882 6560
rect 17096 4928 17332 5090
rect 17096 4864 17126 4928
rect 17126 4864 17142 4928
rect 17142 4864 17206 4928
rect 17206 4864 17222 4928
rect 17222 4864 17286 4928
rect 17286 4864 17302 4928
rect 17302 4864 17332 4928
rect 17096 4854 17332 4864
rect 18646 3296 18882 3400
rect 18646 3232 18676 3296
rect 18676 3232 18692 3296
rect 18692 3232 18756 3296
rect 18756 3232 18772 3296
rect 18772 3232 18836 3296
rect 18836 3232 18852 3296
rect 18852 3232 18882 3296
rect 18646 3164 18882 3232
<< metal5 >>
rect 136 10160 18924 10202
rect 136 9924 3146 10160
rect 3382 9924 6246 10160
rect 6482 9924 9346 10160
rect 9582 9924 12446 10160
rect 12682 9924 15546 10160
rect 15782 9924 18646 10160
rect 18882 9924 18924 10160
rect 136 9882 18924 9924
rect 136 8470 18908 8512
rect 136 8234 4696 8470
rect 4932 8234 7796 8470
rect 8032 8234 10896 8470
rect 11132 8234 13996 8470
rect 14232 8234 17096 8470
rect 17332 8234 18908 8470
rect 136 8192 18908 8234
rect 136 6780 18924 6822
rect 136 6544 3146 6780
rect 3382 6544 6246 6780
rect 6482 6544 9346 6780
rect 9582 6544 12446 6780
rect 12682 6544 15546 6780
rect 15782 6544 18646 6780
rect 18882 6544 18924 6780
rect 136 6502 18924 6544
rect 136 5090 18908 5132
rect 136 4854 4696 5090
rect 4932 4854 7796 5090
rect 8032 4854 10896 5090
rect 11132 4854 13996 5090
rect 14232 4854 17096 5090
rect 17332 4854 18908 5090
rect 136 4812 18908 4854
rect 136 3400 18924 3442
rect 136 3164 3146 3400
rect 3382 3164 6246 3400
rect 6482 3164 9346 3400
rect 9582 3164 12446 3400
rect 12682 3164 15546 3400
rect 15782 3164 18646 3400
rect 18882 3164 18924 3400
rect 136 3122 18924 3164
use sky130_fd_sc_hd__diode_2  ANTENNA__233__A1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 5336 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__A1
timestamp 1665323087
transform -1 0 4140 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__S
timestamp 1665323087
transform 1 0 5152 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__A1
timestamp 1665323087
transform 1 0 4508 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__A1
timestamp 1665323087
transform 1 0 3496 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__S
timestamp 1665323087
transform -1 0 644 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__A1
timestamp 1665323087
transform 1 0 3864 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__238__A1
timestamp 1665323087
transform 1 0 3312 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__S
timestamp 1665323087
transform 1 0 12236 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__A1
timestamp 1665323087
transform 1 0 7176 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__242__A1
timestamp 1665323087
transform 1 0 4600 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__242__S
timestamp 1665323087
transform 1 0 4784 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A1
timestamp 1665323087
transform 1 0 7452 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__A1
timestamp 1665323087
transform 1 0 5152 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__A0
timestamp 1665323087
transform -1 0 13892 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__A0
timestamp 1665323087
transform -1 0 17204 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__A
timestamp 1665323087
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__B
timestamp 1665323087
transform 1 0 14628 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__A1
timestamp 1665323087
transform -1 0 18584 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__B1
timestamp 1665323087
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__277__A1
timestamp 1665323087
transform 1 0 7176 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__277__A2
timestamp 1665323087
transform 1 0 6440 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__277__B1
timestamp 1665323087
transform 1 0 6256 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__A1
timestamp 1665323087
transform 1 0 8372 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__A2
timestamp 1665323087
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__B1
timestamp 1665323087
transform -1 0 9752 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__A2
timestamp 1665323087
transform -1 0 17848 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__A1
timestamp 1665323087
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__306__B
timestamp 1665323087
transform 1 0 460 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__313__A_N
timestamp 1665323087
transform 1 0 11960 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__316__A2
timestamp 1665323087
transform -1 0 13708 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__333__A
timestamp 1665323087
transform 1 0 4140 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__333__B
timestamp 1665323087
transform 1 0 3956 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__A
timestamp 1665323087
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__B
timestamp 1665323087
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__C
timestamp 1665323087
transform 1 0 5060 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__336__A1
timestamp 1665323087
transform 1 0 2392 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__336__A2
timestamp 1665323087
transform -1 0 828 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__336__B1
timestamp 1665323087
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__351__B1
timestamp 1665323087
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__381__A1
timestamp 1665323087
transform 1 0 12696 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__387__A_N
timestamp 1665323087
transform 1 0 16744 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__388__A
timestamp 1665323087
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__390__A1
timestamp 1665323087
transform -1 0 14536 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__390__A2
timestamp 1665323087
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__397__A1
timestamp 1665323087
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__397__A2
timestamp 1665323087
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__398__A1
timestamp 1665323087
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__398__A3
timestamp 1665323087
transform 1 0 6072 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__399__A1
timestamp 1665323087
transform -1 0 8924 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__399__A2
timestamp 1665323087
transform 1 0 7176 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__400__A1
timestamp 1665323087
transform 1 0 3588 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__400__A3
timestamp 1665323087
transform 1 0 2944 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__401__A2
timestamp 1665323087
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__402__A1
timestamp 1665323087
transform 1 0 5060 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__402__A3
timestamp 1665323087
transform 1 0 4784 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__408__A
timestamp 1665323087
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__409__A1
timestamp 1665323087
transform -1 0 16928 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__417__SET_B
timestamp 1665323087
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__421__RESET_B
timestamp 1665323087
transform 1 0 8648 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__SET_B
timestamp 1665323087
transform 1 0 12236 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__437__SET_B
timestamp 1665323087
transform 1 0 13340 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__438__RESET_B
timestamp 1665323087
transform -1 0 14352 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__450__D
timestamp 1665323087
transform 1 0 17020 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__452__SET_B
timestamp 1665323087
transform -1 0 14904 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__453__RESET_B
timestamp 1665323087
transform 1 0 13156 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__457__SET_B
timestamp 1665323087
transform 1 0 9568 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__461__RESET_B
timestamp 1665323087
transform 1 0 12236 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__463__RESET_B
timestamp 1665323087
transform 1 0 11040 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__465__SET_B
timestamp 1665323087
transform 1 0 5060 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__466__RESET_B
timestamp 1665323087
transform -1 0 18124 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__467__RESET_B
timestamp 1665323087
transform -1 0 16652 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__468__RESET_B
timestamp 1665323087
transform 1 0 16468 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__469__SET_B
timestamp 1665323087
transform -1 0 13616 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__470__RESET_B
timestamp 1665323087
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__471__RESET_B
timestamp 1665323087
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__472__SET_B
timestamp 1665323087
transform -1 0 14812 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__473__RESET_B
timestamp 1665323087
transform 1 0 14260 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_ext_clk_A
timestamp 1665323087
transform -1 0 4324 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_pll_clk90_A
timestamp 1665323087
transform -1 0 13340 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_pll_clk_A
timestamp 1665323087
transform 1 0 10764 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout21_A
timestamp 1665323087
transform 1 0 3680 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout27_A
timestamp 1665323087
transform 1 0 9660 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout28_A
timestamp 1665323087
transform -1 0 920 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1665323087
transform -1 0 12420 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1665323087
transform -1 0 11960 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1665323087
transform -1 0 2852 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1665323087
transform -1 0 12696 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1665323087
transform -1 0 15548 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1665323087
transform -1 0 15732 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1665323087
transform -1 0 12144 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1665323087
transform -1 0 12604 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1665323087
transform -1 0 12788 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 460 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1196 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1472 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27
timestamp 1665323087
transform 1 0 2668 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40
timestamp 1665323087
transform 1 0 3864 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53
timestamp 1665323087
transform 1 0 5060 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 6256 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 6624 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_88 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 8280 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_96
timestamp 1665323087
transform 1 0 9016 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 10304 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116
timestamp 1665323087
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_118
timestamp 1665323087
transform 1 0 11040 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_126
timestamp 1665323087
transform 1 0 11776 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_144
timestamp 1665323087
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_179
timestamp 1665323087
transform 1 0 16652 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_185
timestamp 1665323087
transform 1 0 17204 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_196
timestamp 1665323087
transform 1 0 18216 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1665323087
transform 1 0 460 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_15
timestamp 1665323087
transform 1 0 1564 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_23
timestamp 1665323087
transform 1 0 2300 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_27
timestamp 1665323087
transform 1 0 2668 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_50
timestamp 1665323087
transform 1 0 4784 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_56
timestamp 1665323087
transform 1 0 5336 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_69
timestamp 1665323087
transform 1 0 6532 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_77
timestamp 1665323087
transform 1 0 7268 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_83
timestamp 1665323087
transform 1 0 7820 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_95
timestamp 1665323087
transform 1 0 8924 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_99
timestamp 1665323087
transform 1 0 9292 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_124
timestamp 1665323087
transform 1 0 11592 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_135
timestamp 1665323087
transform 1 0 12604 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_157
timestamp 1665323087
transform 1 0 14628 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_185
timestamp 1665323087
transform 1 0 17204 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp 1665323087
transform 1 0 460 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_11
timestamp 1665323087
transform 1 0 1196 0 1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_14
timestamp 1665323087
transform 1 0 1472 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_26
timestamp 1665323087
transform 1 0 2576 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_35
timestamp 1665323087
transform 1 0 3404 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_40
timestamp 1665323087
transform 1 0 3864 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_90
timestamp 1665323087
transform 1 0 8464 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_92
timestamp 1665323087
transform 1 0 8648 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_133
timestamp 1665323087
transform 1 0 12420 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_196
timestamp 1665323087
transform 1 0 18216 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1665323087
transform 1 0 460 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_15
timestamp 1665323087
transform 1 0 1564 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_24
timestamp 1665323087
transform 1 0 2392 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_27
timestamp 1665323087
transform 1 0 2668 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_45
timestamp 1665323087
transform 1 0 4324 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_56
timestamp 1665323087
transform 1 0 5336 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_103
timestamp 1665323087
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_125
timestamp 1665323087
transform 1 0 11684 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_155
timestamp 1665323087
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_159
timestamp 1665323087
transform 1 0 14812 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_199
timestamp 1665323087
transform 1 0 18492 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_3
timestamp 1665323087
transform 1 0 460 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_11
timestamp 1665323087
transform 1 0 1196 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_14
timestamp 1665323087
transform 1 0 1472 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_92
timestamp 1665323087
transform 1 0 8648 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_120
timestamp 1665323087
transform 1 0 11224 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_142
timestamp 1665323087
transform 1 0 13248 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_196
timestamp 1665323087
transform 1 0 18216 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1665323087
transform 1 0 460 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_15
timestamp 1665323087
transform 1 0 1564 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_53
timestamp 1665323087
transform 1 0 5060 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_88
timestamp 1665323087
transform 1 0 8280 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_175
timestamp 1665323087
transform 1 0 16284 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1665323087
transform 1 0 460 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_11
timestamp 1665323087
transform 1 0 1196 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_14
timestamp 1665323087
transform 1 0 1472 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_18
timestamp 1665323087
transform 1 0 1840 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_40
timestamp 1665323087
transform 1 0 3864 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_116
timestamp 1665323087
transform 1 0 10856 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_121
timestamp 1665323087
transform 1 0 11316 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1665323087
transform 1 0 460 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_15
timestamp 1665323087
transform 1 0 1564 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_23
timestamp 1665323087
transform 1 0 2300 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_27
timestamp 1665323087
transform 1 0 2668 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_181
timestamp 1665323087
transform 1 0 16836 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_183
timestamp 1665323087
transform 1 0 17020 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_3
timestamp 1665323087
transform 1 0 460 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_11
timestamp 1665323087
transform 1 0 1196 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_34
timestamp 1665323087
transform 1 0 3312 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_64
timestamp 1665323087
transform 1 0 6072 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_66
timestamp 1665323087
transform 1 0 6256 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_168
timestamp 1665323087
transform 1 0 15640 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3
timestamp 1665323087
transform 1 0 460 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_29
timestamp 1665323087
transform 1 0 2852 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_47
timestamp 1665323087
transform 1 0 4508 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_79
timestamp 1665323087
transform 1 0 7452 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_103
timestamp 1665323087
transform 1 0 9660 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_155
timestamp 1665323087
transform 1 0 14444 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_199
timestamp 1665323087
transform 1 0 18492 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_35
timestamp 1665323087
transform 1 0 3404 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_55
timestamp 1665323087
transform 1 0 5244 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_70
timestamp 1665323087
transform 1 0 6624 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_148
timestamp 1665323087
transform 1 0 13800 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_199
timestamp 1665323087
transform 1 0 18492 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1665323087
transform 1 0 460 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_49
timestamp 1665323087
transform 1 0 4692 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_75
timestamp 1665323087
transform 1 0 7084 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_79
timestamp 1665323087
transform 1 0 7452 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_129
timestamp 1665323087
transform 1 0 12052 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_199
timestamp 1665323087
transform 1 0 18492 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_54
timestamp 1665323087
transform 1 0 5152 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_138
timestamp 1665323087
transform 1 0 12880 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_196
timestamp 1665323087
transform 1 0 18216 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_79
timestamp 1665323087
transform 1 0 7452 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_103
timestamp 1665323087
transform 1 0 9660 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_125
timestamp 1665323087
transform 1 0 11684 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_195
timestamp 1665323087
transform 1 0 18124 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_199
timestamp 1665323087
transform 1 0 18492 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_142
timestamp 1665323087
transform 1 0 13248 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1665323087
transform 1 0 460 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_75
timestamp 1665323087
transform 1 0 7084 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_199
timestamp 1665323087
transform 1 0 18492 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_44
timestamp 1665323087
transform 1 0 4232 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_120
timestamp 1665323087
transform 1 0 11224 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_142
timestamp 1665323087
transform 1 0 13248 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_53
timestamp 1665323087
transform 1 0 5060 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_199
timestamp 1665323087
transform 1 0 18492 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_40
timestamp 1665323087
transform 1 0 3864 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_53
timestamp 1665323087
transform 1 0 5060 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_88
timestamp 1665323087
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_92
timestamp 1665323087
transform 1 0 8648 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_116
timestamp 1665323087
transform 1 0 10856 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_155
timestamp 1665323087
transform 1 0 14444 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_168
timestamp 1665323087
transform 1 0 15640 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_199
timestamp 1665323087
transform 1 0 18492 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1665323087
transform 1 0 184 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1665323087
transform -1 0 18860 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1665323087
transform 1 0 184 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1665323087
transform -1 0 18860 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1665323087
transform 1 0 184 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1665323087
transform -1 0 18860 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1665323087
transform 1 0 184 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1665323087
transform -1 0 18860 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1665323087
transform 1 0 184 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1665323087
transform -1 0 18860 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1665323087
transform 1 0 184 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1665323087
transform -1 0 18860 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1665323087
transform 1 0 184 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1665323087
transform -1 0 18860 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1665323087
transform 1 0 184 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1665323087
transform -1 0 18860 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1665323087
transform 1 0 184 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1665323087
transform -1 0 18860 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1665323087
transform 1 0 184 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1665323087
transform -1 0 18860 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1665323087
transform 1 0 184 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1665323087
transform -1 0 18860 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1665323087
transform 1 0 184 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1665323087
transform -1 0 18860 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1665323087
transform 1 0 184 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1665323087
transform -1 0 18860 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1665323087
transform 1 0 184 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1665323087
transform -1 0 18860 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1665323087
transform 1 0 184 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1665323087
transform -1 0 18860 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1665323087
transform 1 0 184 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1665323087
transform -1 0 18860 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1665323087
transform 1 0 184 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1665323087
transform -1 0 18860 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1665323087
transform 1 0 184 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1665323087
transform -1 0 18860 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1665323087
transform 1 0 184 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1665323087
transform -1 0 18860 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1380 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1665323087
transform 1 0 2576 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1665323087
transform 1 0 3772 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1665323087
transform 1 0 4968 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1665323087
transform 1 0 6164 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1665323087
transform 1 0 7360 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1665323087
transform 1 0 8556 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1665323087
transform 1 0 9752 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1665323087
transform 1 0 10948 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1665323087
transform 1 0 12144 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1665323087
transform 1 0 13340 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1665323087
transform 1 0 14536 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1665323087
transform 1 0 15732 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1665323087
transform 1 0 16928 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1665323087
transform 1 0 18124 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1665323087
transform 1 0 2576 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1665323087
transform 1 0 4968 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1665323087
transform 1 0 7360 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1665323087
transform 1 0 9752 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1665323087
transform 1 0 12144 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1665323087
transform 1 0 14536 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1665323087
transform 1 0 16928 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1665323087
transform 1 0 1380 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1665323087
transform 1 0 3772 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1665323087
transform 1 0 6164 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1665323087
transform 1 0 8556 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1665323087
transform 1 0 10948 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1665323087
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1665323087
transform 1 0 15732 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1665323087
transform 1 0 18124 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1665323087
transform 1 0 2576 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1665323087
transform 1 0 4968 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1665323087
transform 1 0 7360 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1665323087
transform 1 0 9752 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1665323087
transform 1 0 12144 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1665323087
transform 1 0 14536 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1665323087
transform 1 0 16928 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1665323087
transform 1 0 1380 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1665323087
transform 1 0 3772 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1665323087
transform 1 0 6164 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1665323087
transform 1 0 8556 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1665323087
transform 1 0 10948 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1665323087
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1665323087
transform 1 0 15732 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1665323087
transform 1 0 18124 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1665323087
transform 1 0 2576 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1665323087
transform 1 0 4968 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1665323087
transform 1 0 7360 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1665323087
transform 1 0 9752 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1665323087
transform 1 0 12144 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1665323087
transform 1 0 14536 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1665323087
transform 1 0 16928 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1665323087
transform 1 0 1380 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1665323087
transform 1 0 3772 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1665323087
transform 1 0 6164 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1665323087
transform 1 0 8556 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1665323087
transform 1 0 10948 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1665323087
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1665323087
transform 1 0 15732 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1665323087
transform 1 0 18124 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1665323087
transform 1 0 2576 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1665323087
transform 1 0 4968 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1665323087
transform 1 0 7360 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1665323087
transform 1 0 9752 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1665323087
transform 1 0 12144 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1665323087
transform 1 0 14536 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1665323087
transform 1 0 16928 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1665323087
transform 1 0 1380 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1665323087
transform 1 0 3772 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1665323087
transform 1 0 6164 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1665323087
transform 1 0 8556 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1665323087
transform 1 0 10948 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1665323087
transform 1 0 13340 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1665323087
transform 1 0 15732 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1665323087
transform 1 0 18124 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1665323087
transform 1 0 2576 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1665323087
transform 1 0 4968 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1665323087
transform 1 0 7360 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1665323087
transform 1 0 9752 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1665323087
transform 1 0 12144 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1665323087
transform 1 0 14536 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1665323087
transform 1 0 16928 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1665323087
transform 1 0 1380 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1665323087
transform 1 0 3772 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1665323087
transform 1 0 6164 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1665323087
transform 1 0 8556 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1665323087
transform 1 0 10948 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1665323087
transform 1 0 13340 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1665323087
transform 1 0 15732 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1665323087
transform 1 0 18124 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1665323087
transform 1 0 2576 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1665323087
transform 1 0 4968 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1665323087
transform 1 0 7360 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1665323087
transform 1 0 9752 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1665323087
transform 1 0 12144 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1665323087
transform 1 0 14536 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1665323087
transform 1 0 16928 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1665323087
transform 1 0 1380 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1665323087
transform 1 0 3772 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1665323087
transform 1 0 6164 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1665323087
transform 1 0 8556 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1665323087
transform 1 0 10948 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1665323087
transform 1 0 13340 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1665323087
transform 1 0 15732 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1665323087
transform 1 0 18124 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1665323087
transform 1 0 2576 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1665323087
transform 1 0 4968 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1665323087
transform 1 0 7360 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1665323087
transform 1 0 9752 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1665323087
transform 1 0 12144 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1665323087
transform 1 0 14536 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1665323087
transform 1 0 16928 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1665323087
transform 1 0 1380 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1665323087
transform 1 0 3772 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1665323087
transform 1 0 6164 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1665323087
transform 1 0 8556 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1665323087
transform 1 0 10948 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1665323087
transform 1 0 13340 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1665323087
transform 1 0 15732 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1665323087
transform 1 0 18124 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1665323087
transform 1 0 2576 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1665323087
transform 1 0 4968 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1665323087
transform 1 0 7360 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1665323087
transform 1 0 9752 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1665323087
transform 1 0 12144 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1665323087
transform 1 0 14536 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1665323087
transform 1 0 16928 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1665323087
transform 1 0 1380 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1665323087
transform 1 0 3772 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1665323087
transform 1 0 6164 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1665323087
transform 1 0 8556 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1665323087
transform 1 0 10948 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1665323087
transform 1 0 13340 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1665323087
transform 1 0 15732 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1665323087
transform 1 0 18124 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1665323087
transform 1 0 2576 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1665323087
transform 1 0 4968 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1665323087
transform 1 0 7360 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1665323087
transform 1 0 9752 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1665323087
transform 1 0 12144 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1665323087
transform 1 0 14536 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1665323087
transform 1 0 16928 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1665323087
transform 1 0 1380 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1665323087
transform 1 0 2576 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1665323087
transform 1 0 3772 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1665323087
transform 1 0 4968 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1665323087
transform 1 0 6164 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1665323087
transform 1 0 7360 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1665323087
transform 1 0 8556 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1665323087
transform 1 0 9752 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1665323087
transform 1 0 10948 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1665323087
transform 1 0 12144 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1665323087
transform 1 0 13340 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1665323087
transform 1 0 14536 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1665323087
transform 1 0 15732 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1665323087
transform 1 0 16928 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1665323087
transform 1 0 18124 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _206_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 6256 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _207_
timestamp 1665323087
transform 1 0 1748 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _208_
timestamp 1665323087
transform 1 0 8924 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _209_
timestamp 1665323087
transform -1 0 2576 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _210_
timestamp 1665323087
transform 1 0 10028 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _211_
timestamp 1665323087
transform -1 0 14444 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _212_
timestamp 1665323087
transform -1 0 11868 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _213_
timestamp 1665323087
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _214_
timestamp 1665323087
transform 1 0 4692 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _215_
timestamp 1665323087
transform 1 0 4324 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _216_
timestamp 1665323087
transform 1 0 7912 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _217_
timestamp 1665323087
transform -1 0 8188 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _218_
timestamp 1665323087
transform 1 0 7452 0 1 544
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _219_
timestamp 1665323087
transform 1 0 5704 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _220_
timestamp 1665323087
transform 1 0 11040 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _221_
timestamp 1665323087
transform -1 0 10672 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _222_
timestamp 1665323087
transform -1 0 14168 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _223_
timestamp 1665323087
transform 1 0 13432 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _224_
timestamp 1665323087
transform -1 0 16652 0 1 544
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _225_
timestamp 1665323087
transform 1 0 15824 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _226_
timestamp 1665323087
transform 1 0 17020 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _227_
timestamp 1665323087
transform -1 0 17848 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _228_
timestamp 1665323087
transform -1 0 7084 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _229_
timestamp 1665323087
transform 1 0 7360 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _230_
timestamp 1665323087
transform 1 0 3680 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _231_
timestamp 1665323087
transform 1 0 4416 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _232_
timestamp 1665323087
transform 1 0 3864 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _233_
timestamp 1665323087
transform 1 0 6532 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _234_
timestamp 1665323087
transform 1 0 5336 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _235_
timestamp 1665323087
transform 1 0 4140 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _236_
timestamp 1665323087
transform -1 0 3772 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _237_
timestamp 1665323087
transform 1 0 2668 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _238_
timestamp 1665323087
transform 1 0 1748 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _239_
timestamp 1665323087
transform -1 0 10120 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _240_
timestamp 1665323087
transform -1 0 10948 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _241_
timestamp 1665323087
transform 1 0 8188 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _242_
timestamp 1665323087
transform -1 0 7360 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _243_
timestamp 1665323087
transform 1 0 8188 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _244_
timestamp 1665323087
transform 1 0 7452 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _245_
timestamp 1665323087
transform -1 0 15640 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _246_
timestamp 1665323087
transform 1 0 17020 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_4  _247_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 1748 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _248_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 10948 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 1665323087
transform 1 0 3864 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_4  _250_
timestamp 1665323087
transform 1 0 5152 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  _251_
timestamp 1665323087
transform -1 0 10304 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1665323087
transform -1 0 5336 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _253_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 8556 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1665323087
transform 1 0 5152 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_4  _255_
timestamp 1665323087
transform 1 0 5520 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _256_
timestamp 1665323087
transform -1 0 9016 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  _257_
timestamp 1665323087
transform -1 0 13340 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _258_
timestamp 1665323087
transform -1 0 16192 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  _259_
timestamp 1665323087
transform -1 0 3680 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp 1665323087
transform 1 0 3496 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _261_
timestamp 1665323087
transform 1 0 6992 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  _262_
timestamp 1665323087
transform -1 0 9292 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _263_
timestamp 1665323087
transform 1 0 18308 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1665323087
transform -1 0 10856 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1665323087
transform 1 0 16652 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  _266__7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 13340 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _267_
timestamp 1665323087
transform 1 0 8188 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  _268__4
timestamp 1665323087
transform -1 0 3404 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _269_
timestamp 1665323087
transform 1 0 10672 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1665323087
transform -1 0 828 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  _271__1
timestamp 1665323087
transform 1 0 3312 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _272_
timestamp 1665323087
transform -1 0 1748 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _273_
timestamp 1665323087
transform -1 0 2208 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _274_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 3772 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _275_
timestamp 1665323087
transform 1 0 14260 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _276_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 18124 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__o2111ai_4  _277_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 5060 0 -1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  _278_
timestamp 1665323087
transform -1 0 736 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_2  _279_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 5244 0 1 7072
box -38 -48 958 592
use sky130_fd_sc_hd__o2111a_1  _280_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 9568 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__a41oi_1  _281_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 12880 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _282_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 9844 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_2  _283_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 4968 0 1 7072
box -38 -48 958 592
use sky130_fd_sc_hd__nand3b_1  _284_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 552 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _285_
timestamp 1665323087
transform -1 0 4232 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _286_
timestamp 1665323087
transform 1 0 2852 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _287_
timestamp 1665323087
transform -1 0 5336 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _288_
timestamp 1665323087
transform -1 0 13156 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _289_
timestamp 1665323087
transform 1 0 12236 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__o2111ai_4  _290_
timestamp 1665323087
transform 1 0 5428 0 -1 2720
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  _291_
timestamp 1665323087
transform 1 0 9384 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_2  _292_
timestamp 1665323087
transform 1 0 9844 0 -1 1632
box -38 -48 958 592
use sky130_fd_sc_hd__o2111a_1  _293_
timestamp 1665323087
transform -1 0 9200 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__a41oi_1  _294_
timestamp 1665323087
transform -1 0 9384 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _295_
timestamp 1665323087
transform -1 0 9660 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_2  _296_
timestamp 1665323087
transform 1 0 6256 0 1 1632
box -38 -48 958 592
use sky130_fd_sc_hd__nand3b_1  _297_
timestamp 1665323087
transform -1 0 4600 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _298_
timestamp 1665323087
transform -1 0 6164 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _299_
timestamp 1665323087
transform -1 0 7360 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _300_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 8004 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _301_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 4968 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _302_
timestamp 1665323087
transform -1 0 14444 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _303_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 15364 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _304_
timestamp 1665323087
transform -1 0 18492 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _305_
timestamp 1665323087
transform -1 0 18124 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _306_
timestamp 1665323087
transform 1 0 460 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _307_
timestamp 1665323087
transform -1 0 13248 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _308_
timestamp 1665323087
transform 1 0 9016 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_2  _309_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 8280 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _310_
timestamp 1665323087
transform -1 0 11316 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _311_
timestamp 1665323087
transform -1 0 12696 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_2  _312_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 10948 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_2  _313_
timestamp 1665323087
transform -1 0 17664 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _314_
timestamp 1665323087
transform 1 0 15272 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _315_
timestamp 1665323087
transform 1 0 14076 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_2  _316_
timestamp 1665323087
transform 1 0 15824 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _317_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 7728 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _318_
timestamp 1665323087
transform 1 0 3680 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _319_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 7452 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _320_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 7360 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _321_
timestamp 1665323087
transform 1 0 8004 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _322_
timestamp 1665323087
transform -1 0 4968 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _323_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 4600 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _324_
timestamp 1665323087
transform 1 0 6716 0 1 544
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _325_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 9844 0 1 544
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _326_
timestamp 1665323087
transform 1 0 9384 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _327_
timestamp 1665323087
transform 1 0 11316 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _328_
timestamp 1665323087
transform -1 0 18492 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _329_
timestamp 1665323087
transform -1 0 13340 0 -1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _330_
timestamp 1665323087
transform 1 0 16652 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _331_
timestamp 1665323087
transform -1 0 18124 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _332_
timestamp 1665323087
transform 1 0 5428 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _333_
timestamp 1665323087
transform -1 0 6348 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _334_
timestamp 1665323087
transform 1 0 1932 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _335_
timestamp 1665323087
transform 1 0 6256 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _336_
timestamp 1665323087
transform -1 0 1380 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _337_
timestamp 1665323087
transform 1 0 5796 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _338_
timestamp 1665323087
transform 1 0 828 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _339_
timestamp 1665323087
transform 1 0 828 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _340_
timestamp 1665323087
transform 1 0 736 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _341_
timestamp 1665323087
transform 1 0 3312 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _342_
timestamp 1665323087
transform -1 0 4968 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _343_
timestamp 1665323087
transform -1 0 4968 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _344_
timestamp 1665323087
transform -1 0 9660 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _345_
timestamp 1665323087
transform -1 0 10948 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _346_
timestamp 1665323087
transform -1 0 8556 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _347_
timestamp 1665323087
transform 1 0 7544 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _348_
timestamp 1665323087
transform -1 0 17940 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _349_
timestamp 1665323087
transform 1 0 11868 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o2111ai_1  _350_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 16652 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _351_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 11776 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _352_
timestamp 1665323087
transform -1 0 12144 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _353_
timestamp 1665323087
transform 1 0 8648 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nand4b_1  _354_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 7636 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _355_
timestamp 1665323087
transform 1 0 8648 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _356_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 17664 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _357_
timestamp 1665323087
transform 1 0 16468 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _358_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 18584 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _359_
timestamp 1665323087
transform -1 0 18584 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _360_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 17664 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _361_
timestamp 1665323087
transform -1 0 18584 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _362_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 18308 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _363_
timestamp 1665323087
transform 1 0 6256 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _364_
timestamp 1665323087
transform -1 0 7820 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _365_
timestamp 1665323087
transform 1 0 8740 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _366_
timestamp 1665323087
transform -1 0 9660 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _367_
timestamp 1665323087
transform -1 0 2576 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _368_
timestamp 1665323087
transform 1 0 3864 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _369_
timestamp 1665323087
transform 1 0 12236 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_1  _370_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 11868 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_1  _371_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 13340 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _372_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 14536 0 1 544
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _373_
timestamp 1665323087
transform 1 0 17848 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _374_
timestamp 1665323087
transform 1 0 17664 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _375_
timestamp 1665323087
transform 1 0 6348 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _376_
timestamp 1665323087
transform 1 0 5336 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_1  _377_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 10304 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _378_
timestamp 1665323087
transform -1 0 8188 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _379_
timestamp 1665323087
transform 1 0 11684 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _380_
timestamp 1665323087
transform -1 0 2576 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _381_
timestamp 1665323087
transform -1 0 18584 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nand4b_1  _382_
timestamp 1665323087
transform -1 0 18492 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _383_
timestamp 1665323087
transform -1 0 16928 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _384_
timestamp 1665323087
transform -1 0 15088 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _385_
timestamp 1665323087
transform 1 0 15272 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _386_
timestamp 1665323087
transform -1 0 16284 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _387_
timestamp 1665323087
transform 1 0 14628 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _388_
timestamp 1665323087
transform 1 0 15272 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _389_
timestamp 1665323087
transform 1 0 12972 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _390_
timestamp 1665323087
transform 1 0 13524 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _391_
timestamp 1665323087
transform -1 0 1380 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _392_
timestamp 1665323087
transform 1 0 460 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _393_
timestamp 1665323087
transform -1 0 1932 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _394_
timestamp 1665323087
transform 1 0 460 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _395_
timestamp 1665323087
transform 1 0 2668 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _396_
timestamp 1665323087
transform -1 0 1748 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _397_
timestamp 1665323087
transform -1 0 12052 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_1  _398_
timestamp 1665323087
transform 1 0 8004 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_1  _399_
timestamp 1665323087
transform 1 0 7452 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _400_
timestamp 1665323087
transform -1 0 5704 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _401_
timestamp 1665323087
transform 1 0 7452 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _402_
timestamp 1665323087
transform -1 0 8188 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o2111ai_1  _403_
timestamp 1665323087
transform 1 0 17020 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _404_
timestamp 1665323087
transform -1 0 14536 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _405_
timestamp 1665323087
transform 1 0 13432 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _406_
timestamp 1665323087
transform 1 0 17020 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _407_
timestamp 1665323087
transform 1 0 15824 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_1  _408_
timestamp 1665323087
transform -1 0 18124 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _409_
timestamp 1665323087
transform 1 0 17848 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _410_
timestamp 1665323087
transform -1 0 18124 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _411__8
timestamp 1665323087
transform -1 0 7912 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _412__9
timestamp 1665323087
transform 1 0 6256 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _413__5
timestamp 1665323087
transform -1 0 10304 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _414__6
timestamp 1665323087
transform -1 0 2392 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _415__2
timestamp 1665323087
transform -1 0 14536 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _416__3
timestamp 1665323087
transform 1 0 920 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__dfstp_1  _417_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 10212 0 -1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _418_
timestamp 1665323087
transform 1 0 7452 0 -1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _419__30 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 6256 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _419_
timestamp 1665323087
transform 1 0 6624 0 1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _420_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 11684 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _421_
timestamp 1665323087
transform 1 0 8832 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _422_
timestamp 1665323087
transform 1 0 11040 0 1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _423_
timestamp 1665323087
transform -1 0 6164 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _424_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 14904 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _425_
timestamp 1665323087
transform 1 0 14904 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _426_
timestamp 1665323087
transform 1 0 14260 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_1  _427_
timestamp 1665323087
transform 1 0 9016 0 1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _428_
timestamp 1665323087
transform 1 0 15824 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtn_1  _429_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 7452 0 -1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _430_
timestamp 1665323087
transform 1 0 2852 0 -1 1632
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtn_1  _431_
timestamp 1665323087
transform -1 0 11684 0 -1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _432_
timestamp 1665323087
transform 1 0 8648 0 1 3808
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtn_1  _433_
timestamp 1665323087
transform 1 0 1932 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_2  _434_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1840 0 1 2720
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtn_1  _435_
timestamp 1665323087
transform 1 0 2668 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _436_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 12236 0 -1 2720
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _437_
timestamp 1665323087
transform 1 0 13800 0 1 2720
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _438_
timestamp 1665323087
transform 1 0 15824 0 1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_2  _439_
timestamp 1665323087
transform 1 0 3864 0 1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _440_
timestamp 1665323087
transform 1 0 3128 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _441_
timestamp 1665323087
transform -1 0 8556 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _442_
timestamp 1665323087
transform 1 0 12420 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _443_
timestamp 1665323087
transform 1 0 11408 0 1 3808
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _444_
timestamp 1665323087
transform 1 0 10304 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _445_
timestamp 1665323087
transform 1 0 13432 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _446_
timestamp 1665323087
transform 1 0 13432 0 1 3808
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _447_
timestamp 1665323087
transform 1 0 12696 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _448_
timestamp 1665323087
transform 1 0 3496 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _449_
timestamp 1665323087
transform -1 0 16100 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _450_
timestamp 1665323087
transform 1 0 17020 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _451_
timestamp 1665323087
transform -1 0 16284 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_1  _452_
timestamp 1665323087
transform 1 0 16192 0 1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _453_
timestamp 1665323087
transform -1 0 14260 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtn_1  _454_
timestamp 1665323087
transform 1 0 1472 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _455_
timestamp 1665323087
transform -1 0 4600 0 -1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtn_1  _456_
timestamp 1665323087
transform 1 0 1472 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _457_
timestamp 1665323087
transform 1 0 9844 0 -1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtn_1  _458_
timestamp 1665323087
transform -1 0 3312 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_2  _459_
timestamp 1665323087
transform 1 0 1472 0 1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtn_1  _460_
timestamp 1665323087
transform 1 0 1472 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _461_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 11040 0 1 5984
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_1  _462_
timestamp 1665323087
transform 1 0 6256 0 1 7072
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _463_
timestamp 1665323087
transform 1 0 9844 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _464_
timestamp 1665323087
transform -1 0 13248 0 1 2720
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _465_
timestamp 1665323087
transform 1 0 14812 0 -1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _466_
timestamp 1665323087
transform 1 0 15824 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _467_
timestamp 1665323087
transform 1 0 16284 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _468_
timestamp 1665323087
transform -1 0 16928 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _469_
timestamp 1665323087
transform 1 0 11316 0 1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _470_
timestamp 1665323087
transform -1 0 16468 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _471_
timestamp 1665323087
transform 1 0 15088 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _472_
timestamp 1665323087
transform 1 0 12604 0 -1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _473_
timestamp 1665323087
transform 1 0 13892 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__037_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 12236 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_divider.out
timestamp 1665323087
transform 1 0 13432 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_divider2.out
timestamp 1665323087
transform -1 0 16468 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_ext_clk
timestamp 1665323087
transform 1 0 4324 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_net10
timestamp 1665323087
transform -1 0 9752 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_pll_clk90
timestamp 1665323087
transform -1 0 11684 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_pll_clk
timestamp 1665323087
transform -1 0 10764 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__037_
timestamp 1665323087
transform -1 0 7360 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_divider.out
timestamp 1665323087
transform -1 0 12880 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_divider2.out
timestamp 1665323087
transform -1 0 12880 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_ext_clk
timestamp 1665323087
transform -1 0 4508 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_net10
timestamp 1665323087
transform -1 0 7084 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_pll_clk90
timestamp 1665323087
transform -1 0 7084 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_pll_clk
timestamp 1665323087
transform -1 0 7084 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__037_
timestamp 1665323087
transform 1 0 13432 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_divider.out
timestamp 1665323087
transform -1 0 9660 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_divider2.out
timestamp 1665323087
transform 1 0 15824 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_ext_clk
timestamp 1665323087
transform 1 0 8648 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_net10
timestamp 1665323087
transform 1 0 6716 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_pll_clk90
timestamp 1665323087
transform 1 0 12236 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_pll_clk
timestamp 1665323087
transform 1 0 10304 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout13 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 16376 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout14
timestamp 1665323087
transform -1 0 16928 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout15
timestamp 1665323087
transform -1 0 17848 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 18584 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout17
timestamp 1665323087
transform -1 0 16928 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout18
timestamp 1665323087
transform 1 0 17112 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout19
timestamp 1665323087
transform -1 0 8556 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout20
timestamp 1665323087
transform 1 0 15364 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout21
timestamp 1665323087
transform 1 0 3864 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout22
timestamp 1665323087
transform 1 0 16284 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout23
timestamp 1665323087
transform -1 0 11316 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout24
timestamp 1665323087
transform -1 0 17848 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout25 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 644 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 828 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout27
timestamp 1665323087
transform 1 0 9200 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout28
timestamp 1665323087
transform 1 0 828 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout29
timestamp 1665323087
transform 1 0 1196 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 18124 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1665323087
transform 1 0 18216 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1665323087
transform 1 0 2668 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1665323087
transform 1 0 18308 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1665323087
transform 1 0 18216 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1665323087
transform -1 0 15732 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1665323087
transform 1 0 18308 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1665323087
transform 1 0 18308 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1665323087
transform 1 0 18308 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  output11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 17020 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  user_clk_out_buffer
timestamp 1665323087
transform 1 0 13432 0 1 9248
box -38 -48 1878 592
<< labels >>
flabel metal4 s 4654 496 4974 10928 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 7754 496 8074 10928 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 10854 496 11174 10928 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 13954 496 14274 10928 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17054 496 17374 10928 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 136 4812 18908 5132 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 136 8192 18908 8512 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 3104 496 3424 10928 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 6204 496 6524 10928 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 9304 496 9624 10928 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12404 496 12724 10928 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 15504 496 15824 10928 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 18604 496 18924 10928 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 136 3122 18924 3442 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 136 6502 18924 6822 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 136 9882 18924 10202 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 7102 11200 7158 12000 0 FreeSans 224 90 0 0 core_clk
port 2 nsew signal tristate
flabel metal2 s 4250 11200 4306 12000 0 FreeSans 224 90 0 0 ext_clk
port 3 nsew signal input
flabel metal3 s 19200 688 20000 808 0 FreeSans 480 0 0 0 ext_clk_sel
port 4 nsew signal input
flabel metal3 s 19200 11160 20000 11280 0 FreeSans 480 0 0 0 ext_reset
port 5 nsew signal input
flabel metal2 s 15658 11200 15714 12000 0 FreeSans 224 90 0 0 pll_clk
port 6 nsew signal input
flabel metal2 s 18510 11200 18566 12000 0 FreeSans 224 90 0 0 pll_clk90
port 7 nsew signal input
flabel metal2 s 1398 11200 1454 12000 0 FreeSans 224 90 0 0 resetb
port 8 nsew signal input
flabel metal2 s 12806 11200 12862 12000 0 FreeSans 224 90 0 0 resetb_sync
port 9 nsew signal tristate
flabel metal3 s 19200 6672 20000 6792 0 FreeSans 480 0 0 0 sel2[0]
port 10 nsew signal input
flabel metal3 s 19200 8168 20000 8288 0 FreeSans 480 0 0 0 sel2[1]
port 11 nsew signal input
flabel metal3 s 19200 9664 20000 9784 0 FreeSans 480 0 0 0 sel2[2]
port 12 nsew signal input
flabel metal3 s 19200 2184 20000 2304 0 FreeSans 480 0 0 0 sel[0]
port 13 nsew signal input
flabel metal3 s 19200 3680 20000 3800 0 FreeSans 480 0 0 0 sel[1]
port 14 nsew signal input
flabel metal3 s 19200 5176 20000 5296 0 FreeSans 480 0 0 0 sel[2]
port 15 nsew signal input
flabel metal2 s 9954 11200 10010 12000 0 FreeSans 224 90 0 0 user_clk
port 16 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 20000 12000
<< end >>
