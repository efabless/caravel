magic
tech sky130A
magscale 1 2
timestamp 1637281321
<< locali >>
rect 3709 10455 3743 10761
rect 5089 9435 5123 9537
rect 765 5559 799 9401
rect 5273 5015 5307 5321
rect 2697 2295 2731 4641
rect 2789 2363 2823 4913
rect 2881 2839 2915 4709
rect 9965 3519 9999 7293
rect 9907 3485 9999 3519
rect 2973 2839 3007 3009
rect 2965 2805 3007 2839
rect 2965 2771 2999 2805
rect 2881 2737 2999 2771
rect 2881 1887 2915 2737
rect 5549 2363 5583 2465
rect 2881 1547 2915 1853
rect 9965 1479 9999 2465
<< viali >>
rect 1501 11305 1535 11339
rect 1777 11305 1811 11339
rect 2605 11305 2639 11339
rect 2881 11305 2915 11339
rect 3157 11305 3191 11339
rect 6469 11305 6503 11339
rect 6929 11305 6963 11339
rect 7665 11305 7699 11339
rect 7941 11305 7975 11339
rect 8493 11305 8527 11339
rect 8769 11305 8803 11339
rect 1869 11237 1903 11271
rect 3985 11237 4019 11271
rect 4353 11237 4387 11271
rect 4445 11237 4479 11271
rect 4997 11237 5031 11271
rect 5457 11237 5491 11271
rect 6193 11237 6227 11271
rect 7389 11237 7423 11271
rect 1317 11101 1351 11135
rect 1593 11101 1627 11135
rect 2053 11101 2087 11135
rect 2145 11101 2179 11135
rect 2421 11101 2455 11135
rect 2697 11101 2731 11135
rect 2973 11101 3007 11135
rect 3433 11101 3467 11135
rect 3801 11101 3835 11135
rect 4169 11101 4203 11135
rect 4629 11101 4663 11135
rect 4813 11101 4847 11135
rect 5273 11101 5307 11135
rect 5641 11101 5675 11135
rect 5733 11101 5767 11135
rect 6653 11101 6687 11135
rect 7113 11101 7147 11135
rect 7573 11101 7607 11135
rect 8125 11101 8159 11135
rect 8309 11101 8343 11135
rect 8953 11101 8987 11135
rect 9321 11101 9355 11135
rect 3617 11033 3651 11067
rect 2329 10965 2363 10999
rect 3249 10965 3283 10999
rect 5089 10965 5123 10999
rect 5917 10965 5951 10999
rect 9137 10965 9171 10999
rect 9505 10965 9539 10999
rect 1501 10761 1535 10795
rect 2329 10761 2363 10795
rect 3065 10761 3099 10795
rect 3709 10761 3743 10795
rect 5457 10761 5491 10795
rect 8953 10761 8987 10795
rect 1317 10625 1351 10659
rect 1593 10625 1627 10659
rect 1869 10625 1903 10659
rect 2145 10625 2179 10659
rect 2421 10625 2455 10659
rect 3617 10625 3651 10659
rect 1777 10489 1811 10523
rect 3157 10489 3191 10523
rect 5641 10693 5675 10727
rect 5825 10693 5859 10727
rect 9045 10693 9079 10727
rect 4261 10625 4295 10659
rect 4353 10625 4387 10659
rect 4537 10625 4571 10659
rect 4813 10625 4847 10659
rect 5273 10625 5307 10659
rect 6009 10625 6043 10659
rect 8033 10625 8067 10659
rect 8585 10625 8619 10659
rect 8769 10625 8803 10659
rect 9229 10625 9263 10659
rect 3801 10557 3835 10591
rect 6193 10557 6227 10591
rect 6561 10557 6595 10591
rect 9413 10557 9447 10591
rect 8493 10489 8527 10523
rect 2053 10421 2087 10455
rect 3525 10421 3559 10455
rect 3709 10421 3743 10455
rect 3985 10421 4019 10455
rect 4721 10421 4755 10455
rect 4997 10421 5031 10455
rect 5181 10421 5215 10455
rect 3175 10217 3209 10251
rect 6101 10217 6135 10251
rect 7941 10217 7975 10251
rect 8125 10217 8159 10251
rect 8585 10149 8619 10183
rect 9137 10149 9171 10183
rect 9413 10149 9447 10183
rect 3709 10081 3743 10115
rect 1409 10013 1443 10047
rect 3433 10013 3467 10047
rect 4077 10013 4111 10047
rect 5549 10013 5583 10047
rect 7849 10013 7883 10047
rect 8401 10013 8435 10047
rect 9229 10013 9263 10047
rect 7573 9945 7607 9979
rect 8769 9945 8803 9979
rect 8953 9945 8987 9979
rect 1593 9877 1627 9911
rect 1685 9877 1719 9911
rect 6009 9877 6043 9911
rect 1501 9673 1535 9707
rect 2513 9673 2547 9707
rect 4997 9673 5031 9707
rect 6837 9673 6871 9707
rect 5181 9605 5215 9639
rect 1317 9537 1351 9571
rect 1409 9537 1443 9571
rect 1685 9537 1719 9571
rect 2605 9537 2639 9571
rect 4537 9537 4571 9571
rect 5089 9537 5123 9571
rect 5365 9537 5399 9571
rect 5549 9537 5583 9571
rect 5641 9537 5675 9571
rect 5825 9537 5859 9571
rect 6193 9537 6227 9571
rect 7113 9537 7147 9571
rect 7665 9537 7699 9571
rect 9505 9537 9539 9571
rect 2697 9469 2731 9503
rect 3065 9469 3099 9503
rect 9137 9469 9171 9503
rect 765 9401 799 9435
rect 5089 9401 5123 9435
rect 7021 9401 7055 9435
rect 2329 9333 2363 9367
rect 6009 9333 6043 9367
rect 7205 9333 7239 9367
rect 1501 9129 1535 9163
rect 2329 9129 2363 9163
rect 3433 9129 3467 9163
rect 3709 9129 3743 9163
rect 9413 9129 9447 9163
rect 2053 9061 2087 9095
rect 2881 9061 2915 9095
rect 3157 9061 3191 9095
rect 4813 9061 4847 9095
rect 5365 8993 5399 9027
rect 1317 8925 1351 8959
rect 1593 8925 1627 8959
rect 1869 8925 1903 8959
rect 2145 8925 2179 8959
rect 2605 8925 2639 8959
rect 2697 8925 2731 8959
rect 2973 8925 3007 8959
rect 3249 8925 3283 8959
rect 4077 8925 4111 8959
rect 4169 8925 4203 8959
rect 7389 8925 7423 8959
rect 8769 8925 8803 8959
rect 4905 8857 4939 8891
rect 5089 8857 5123 8891
rect 5273 8857 5307 8891
rect 5641 8857 5675 8891
rect 8125 8857 8159 8891
rect 1777 8789 1811 8823
rect 2421 8789 2455 8823
rect 3893 8789 3927 8823
rect 7113 8789 7147 8823
rect 2605 8517 2639 8551
rect 1317 8449 1351 8483
rect 2237 8449 2271 8483
rect 6193 8449 6227 8483
rect 6929 8449 6963 8483
rect 7665 8449 7699 8483
rect 9505 8449 9539 8483
rect 2329 8381 2363 8415
rect 4169 8381 4203 8415
rect 4445 8381 4479 8415
rect 5917 8381 5951 8415
rect 9137 8381 9171 8415
rect 7205 8313 7239 8347
rect 1501 8245 1535 8279
rect 1593 8245 1627 8279
rect 4077 8245 4111 8279
rect 6837 8245 6871 8279
rect 7113 8245 7147 8279
rect 1317 8041 1351 8075
rect 1501 8041 1535 8075
rect 3175 8041 3209 8075
rect 4353 8041 4387 8075
rect 4537 8041 4571 8075
rect 8217 8041 8251 8075
rect 8585 7973 8619 8007
rect 5181 7905 5215 7939
rect 5549 7905 5583 7939
rect 1409 7837 1443 7871
rect 3433 7837 3467 7871
rect 3617 7837 3651 7871
rect 4813 7837 4847 7871
rect 4905 7837 4939 7871
rect 7021 7837 7055 7871
rect 7573 7837 7607 7871
rect 8769 7837 8803 7871
rect 4261 7769 4295 7803
rect 8401 7769 8435 7803
rect 1685 7701 1719 7735
rect 5089 7701 5123 7735
rect 7481 7701 7515 7735
rect 9413 7701 9447 7735
rect 1409 7429 1443 7463
rect 6193 7429 6227 7463
rect 7941 7429 7975 7463
rect 1685 7361 1719 7395
rect 2329 7361 2363 7395
rect 2973 7361 3007 7395
rect 4445 7361 4479 7395
rect 4997 7361 5031 7395
rect 5733 7361 5767 7395
rect 8033 7361 8067 7395
rect 9045 7361 9079 7395
rect 2605 7293 2639 7327
rect 9137 7293 9171 7327
rect 9229 7293 9263 7327
rect 9965 7293 9999 7327
rect 2421 7225 2455 7259
rect 5641 7225 5675 7259
rect 5917 7225 5951 7259
rect 8677 7225 8711 7259
rect 1501 7157 1535 7191
rect 4905 7157 4939 7191
rect 8125 7157 8159 7191
rect 8493 7157 8527 7191
rect 1225 6953 1259 6987
rect 6101 6953 6135 6987
rect 6824 6953 6858 6987
rect 8309 6953 8343 6987
rect 6469 6885 6503 6919
rect 8401 6885 8435 6919
rect 5917 6817 5951 6851
rect 9321 6817 9355 6851
rect 1409 6749 1443 6783
rect 1685 6749 1719 6783
rect 3617 6749 3651 6783
rect 3985 6749 4019 6783
rect 5457 6749 5491 6783
rect 6009 6749 6043 6783
rect 6561 6749 6595 6783
rect 8585 6749 8619 6783
rect 1961 6681 1995 6715
rect 9137 6681 9171 6715
rect 1593 6613 1627 6647
rect 3433 6613 3467 6647
rect 8769 6613 8803 6647
rect 9229 6613 9263 6647
rect 1317 6409 1351 6443
rect 1593 6409 1627 6443
rect 2237 6409 2271 6443
rect 9321 6409 9355 6443
rect 2697 6341 2731 6375
rect 1501 6273 1535 6307
rect 1777 6273 1811 6307
rect 1869 6273 1903 6307
rect 2145 6273 2179 6307
rect 4261 6273 4295 6307
rect 4905 6273 4939 6307
rect 5641 6273 5675 6307
rect 6009 6273 6043 6307
rect 6837 6273 6871 6307
rect 8769 6273 8803 6307
rect 9505 6273 9539 6307
rect 2421 6205 2455 6239
rect 6929 6205 6963 6239
rect 7297 6205 7331 6239
rect 5825 6137 5859 6171
rect 2053 6069 2087 6103
rect 4169 6069 4203 6103
rect 4997 6069 5031 6103
rect 6193 6069 6227 6103
rect 9229 6069 9263 6103
rect 1409 5865 1443 5899
rect 1961 5865 1995 5899
rect 2237 5865 2271 5899
rect 2513 5865 2547 5899
rect 3801 5865 3835 5899
rect 6285 5865 6319 5899
rect 6653 5865 6687 5899
rect 8769 5865 8803 5899
rect 6837 5797 6871 5831
rect 4537 5729 4571 5763
rect 8585 5729 8619 5763
rect 1225 5661 1259 5695
rect 1501 5661 1535 5695
rect 1777 5661 1811 5695
rect 2053 5661 2087 5695
rect 2329 5661 2363 5695
rect 2789 5661 2823 5695
rect 2973 5661 3007 5695
rect 3249 5661 3283 5695
rect 3433 5661 3467 5695
rect 4077 5661 4111 5695
rect 4261 5661 4295 5695
rect 6193 5661 6227 5695
rect 9413 5661 9447 5695
rect 8309 5593 8343 5627
rect 765 5525 799 5559
rect 1685 5525 1719 5559
rect 2605 5525 2639 5559
rect 3065 5525 3099 5559
rect 3617 5525 3651 5559
rect 6009 5525 6043 5559
rect 5089 5321 5123 5355
rect 5273 5321 5307 5355
rect 9413 5321 9447 5355
rect 3617 5253 3651 5287
rect 3341 5185 3375 5219
rect 5365 5185 5399 5219
rect 5549 5185 5583 5219
rect 5733 5185 5767 5219
rect 7665 5185 7699 5219
rect 8309 5185 8343 5219
rect 5825 5117 5859 5151
rect 6193 5117 6227 5151
rect 8125 5117 8159 5151
rect 8677 5117 8711 5151
rect 8861 5117 8895 5151
rect 8493 5049 8527 5083
rect 5273 4981 5307 5015
rect 9321 4981 9355 5015
rect 2789 4913 2823 4947
rect 2697 4641 2731 4675
rect 3801 4777 3835 4811
rect 4445 4777 4479 4811
rect 9505 4777 9539 4811
rect 2881 4709 2915 4743
rect 6285 4641 6319 4675
rect 6561 4641 6595 4675
rect 3433 4573 3467 4607
rect 3709 4573 3743 4607
rect 4353 4573 4387 4607
rect 5549 4573 5583 4607
rect 8125 4573 8159 4607
rect 8769 4573 8803 4607
rect 8861 4573 8895 4607
rect 4905 4505 4939 4539
rect 5733 4505 5767 4539
rect 5917 4505 5951 4539
rect 3617 4437 3651 4471
rect 4169 4437 4203 4471
rect 4813 4437 4847 4471
rect 6101 4437 6135 4471
rect 8033 4437 8067 4471
rect 3525 4233 3559 4267
rect 9045 4165 9079 4199
rect 3341 4097 3375 4131
rect 3617 4097 3651 4131
rect 3985 4097 4019 4131
rect 5457 4097 5491 4131
rect 6101 4097 6135 4131
rect 6837 4097 6871 4131
rect 8125 4097 8159 4131
rect 8585 4097 8619 4131
rect 7573 4029 7607 4063
rect 7665 4029 7699 4063
rect 8861 4029 8895 4063
rect 8953 4029 8987 4063
rect 8401 3961 8435 3995
rect 5917 3893 5951 3927
rect 6745 3893 6779 3927
rect 7481 3893 7515 3927
rect 9413 3893 9447 3927
rect 4077 3689 4111 3723
rect 4537 3689 4571 3723
rect 5181 3689 5215 3723
rect 5365 3689 5399 3723
rect 6285 3689 6319 3723
rect 8861 3689 8895 3723
rect 9229 3689 9263 3723
rect 3525 3621 3559 3655
rect 3893 3621 3927 3655
rect 6929 3553 6963 3587
rect 3341 3485 3375 3519
rect 3617 3485 3651 3519
rect 4261 3485 4295 3519
rect 4353 3485 4387 3519
rect 4721 3485 4755 3519
rect 4997 3485 5031 3519
rect 5549 3485 5583 3519
rect 5733 3485 5767 3519
rect 6009 3485 6043 3519
rect 6561 3485 6595 3519
rect 8401 3485 8435 3519
rect 8953 3485 8987 3519
rect 9873 3485 9907 3519
rect 3801 3349 3835 3383
rect 4905 3349 4939 3383
rect 5917 3349 5951 3383
rect 6469 3349 6503 3383
rect 8585 3349 8619 3383
rect 9413 3349 9447 3383
rect 3801 3145 3835 3179
rect 4077 3145 4111 3179
rect 4261 3145 4295 3179
rect 6837 3145 6871 3179
rect 8677 3145 8711 3179
rect 9045 3145 9079 3179
rect 7573 3077 7607 3111
rect 7757 3077 7791 3111
rect 9137 3077 9171 3111
rect 2973 3009 3007 3043
rect 3341 3009 3375 3043
rect 3617 3009 3651 3043
rect 3893 3009 3927 3043
rect 4353 3009 4387 3043
rect 4721 3009 4755 3043
rect 6193 3009 6227 3043
rect 7481 3009 7515 3043
rect 8309 3009 8343 3043
rect 9229 2941 9263 2975
rect 3525 2873 3559 2907
rect 8493 2873 8527 2907
rect 2881 2805 2915 2839
rect 6653 2805 6687 2839
rect 7941 2805 7975 2839
rect 2789 2329 2823 2363
rect 2697 2261 2731 2295
rect 3525 2601 3559 2635
rect 4169 2601 4203 2635
rect 5457 2601 5491 2635
rect 6469 2601 6503 2635
rect 6929 2601 6963 2635
rect 7113 2601 7147 2635
rect 8125 2601 8159 2635
rect 9045 2601 9079 2635
rect 3617 2533 3651 2567
rect 4077 2533 4111 2567
rect 5089 2533 5123 2567
rect 5733 2533 5767 2567
rect 7481 2533 7515 2567
rect 8585 2533 8619 2567
rect 5549 2465 5583 2499
rect 7573 2465 7607 2499
rect 9965 2465 9999 2499
rect 3341 2397 3375 2431
rect 3801 2397 3835 2431
rect 3893 2397 3927 2431
rect 4353 2397 4387 2431
rect 4813 2397 4847 2431
rect 4905 2397 4939 2431
rect 5273 2397 5307 2431
rect 5917 2397 5951 2431
rect 6009 2397 6043 2431
rect 6285 2397 6319 2431
rect 6745 2397 6779 2431
rect 7205 2397 7239 2431
rect 7297 2397 7331 2431
rect 7757 2397 7791 2431
rect 7941 2397 7975 2431
rect 8309 2397 8343 2431
rect 8401 2397 8435 2431
rect 8769 2397 8803 2431
rect 9505 2397 9539 2431
rect 5549 2329 5583 2363
rect 4537 2261 4571 2295
rect 4629 2261 4663 2295
rect 6193 2261 6227 2295
rect 9229 2261 9263 2295
rect 9321 2261 9355 2295
rect 3617 2057 3651 2091
rect 5273 2057 5307 2091
rect 7573 2057 7607 2091
rect 7849 2057 7883 2091
rect 8125 2057 8159 2091
rect 8585 2057 8619 2091
rect 8861 2057 8895 2091
rect 9413 2057 9447 2091
rect 4629 1989 4663 2023
rect 4905 1989 4939 2023
rect 3341 1921 3375 1955
rect 3801 1921 3835 1955
rect 3893 1921 3927 1955
rect 4169 1921 4203 1955
rect 7665 1921 7699 1955
rect 7941 1921 7975 1955
rect 8401 1921 8435 1955
rect 8677 1921 8711 1955
rect 9137 1921 9171 1955
rect 9229 1921 9263 1955
rect 2881 1853 2915 1887
rect 4445 1853 4479 1887
rect 5365 1853 5399 1887
rect 4077 1785 4111 1819
rect 4353 1785 4387 1819
rect 3525 1717 3559 1751
rect 5089 1717 5123 1751
rect 8953 1717 8987 1751
rect 2881 1513 2915 1547
rect 3985 1513 4019 1547
rect 4169 1513 4203 1547
rect 8401 1513 8435 1547
rect 3617 1445 3651 1479
rect 9965 1445 9999 1479
rect 4353 1377 4387 1411
rect 9137 1377 9171 1411
rect 3341 1309 3375 1343
rect 8585 1309 8619 1343
rect 8677 1309 8711 1343
rect 9505 1309 9539 1343
rect 3525 1173 3559 1207
rect 3801 1173 3835 1207
rect 4537 1173 4571 1207
rect 8861 1173 8895 1207
rect 8953 1173 8987 1207
rect 9321 1173 9355 1207
<< metal1 >>
rect 1946 12112 1952 12164
rect 2004 12152 2010 12164
rect 2314 12152 2320 12164
rect 2004 12124 2320 12152
rect 2004 12112 2010 12124
rect 2314 12112 2320 12124
rect 2372 12112 2378 12164
rect 5994 12112 6000 12164
rect 6052 12152 6058 12164
rect 6362 12152 6368 12164
rect 6052 12124 6368 12152
rect 6052 12112 6058 12124
rect 6362 12112 6368 12124
rect 6420 12112 6426 12164
rect 4154 12044 4160 12096
rect 4212 12084 4218 12096
rect 5350 12084 5356 12096
rect 4212 12056 5356 12084
rect 4212 12044 4218 12056
rect 5350 12044 5356 12056
rect 5408 12044 5414 12096
rect 6086 12044 6092 12096
rect 6144 12084 6150 12096
rect 6454 12084 6460 12096
rect 6144 12056 6460 12084
rect 6144 12044 6150 12056
rect 6454 12044 6460 12056
rect 6512 12044 6518 12096
rect 2314 11976 2320 12028
rect 2372 12016 2378 12028
rect 7834 12016 7840 12028
rect 2372 11988 7840 12016
rect 2372 11976 2378 11988
rect 7834 11976 7840 11988
rect 7892 11976 7898 12028
rect 8570 11948 8576 11960
rect 2746 11920 8576 11948
rect 2406 11840 2412 11892
rect 2464 11880 2470 11892
rect 2746 11880 2774 11920
rect 8570 11908 8576 11920
rect 8628 11908 8634 11960
rect 2464 11852 2774 11880
rect 2464 11840 2470 11852
rect 2958 11840 2964 11892
rect 3016 11880 3022 11892
rect 8386 11880 8392 11892
rect 3016 11852 8392 11880
rect 3016 11840 3022 11852
rect 8386 11840 8392 11852
rect 8444 11840 8450 11892
rect 4338 11772 4344 11824
rect 4396 11812 4402 11824
rect 6086 11812 6092 11824
rect 4396 11784 6092 11812
rect 4396 11772 4402 11784
rect 6086 11772 6092 11784
rect 6144 11772 6150 11824
rect 6822 11772 6828 11824
rect 6880 11812 6886 11824
rect 8202 11812 8208 11824
rect 6880 11784 8208 11812
rect 6880 11772 6886 11784
rect 8202 11772 8208 11784
rect 8260 11772 8266 11824
rect 1486 11704 1492 11756
rect 1544 11744 1550 11756
rect 6914 11744 6920 11756
rect 1544 11716 6920 11744
rect 1544 11704 1550 11716
rect 6914 11704 6920 11716
rect 6972 11704 6978 11756
rect 2222 11636 2228 11688
rect 2280 11676 2286 11688
rect 4706 11676 4712 11688
rect 2280 11648 4712 11676
rect 2280 11636 2286 11648
rect 4706 11636 4712 11648
rect 4764 11636 4770 11688
rect 1302 11568 1308 11620
rect 1360 11608 1366 11620
rect 6178 11608 6184 11620
rect 1360 11580 6184 11608
rect 1360 11568 1366 11580
rect 6178 11568 6184 11580
rect 6236 11568 6242 11620
rect 7098 11568 7104 11620
rect 7156 11608 7162 11620
rect 9674 11608 9680 11620
rect 7156 11580 9680 11608
rect 7156 11568 7162 11580
rect 9674 11568 9680 11580
rect 9732 11568 9738 11620
rect 5258 11500 5264 11552
rect 5316 11540 5322 11552
rect 8294 11540 8300 11552
rect 5316 11512 8300 11540
rect 5316 11500 5322 11512
rect 8294 11500 8300 11512
rect 8352 11500 8358 11552
rect 8478 11500 8484 11552
rect 8536 11540 8542 11552
rect 10410 11540 10416 11552
rect 8536 11512 10416 11540
rect 8536 11500 8542 11512
rect 10410 11500 10416 11512
rect 10468 11500 10474 11552
rect 920 11450 9844 11472
rect 920 11398 2566 11450
rect 2618 11398 2630 11450
rect 2682 11398 2694 11450
rect 2746 11398 2758 11450
rect 2810 11398 2822 11450
rect 2874 11398 5666 11450
rect 5718 11398 5730 11450
rect 5782 11398 5794 11450
rect 5846 11398 5858 11450
rect 5910 11398 5922 11450
rect 5974 11398 8766 11450
rect 8818 11398 8830 11450
rect 8882 11398 8894 11450
rect 8946 11398 8958 11450
rect 9010 11398 9022 11450
rect 9074 11398 9844 11450
rect 920 11376 9844 11398
rect 1486 11336 1492 11348
rect 1447 11308 1492 11336
rect 1486 11296 1492 11308
rect 1544 11296 1550 11348
rect 1765 11339 1823 11345
rect 1765 11305 1777 11339
rect 1811 11336 1823 11339
rect 2222 11336 2228 11348
rect 1811 11308 2228 11336
rect 1811 11305 1823 11308
rect 1765 11299 1823 11305
rect 2222 11296 2228 11308
rect 2280 11296 2286 11348
rect 2314 11296 2320 11348
rect 2372 11336 2378 11348
rect 2593 11339 2651 11345
rect 2593 11336 2605 11339
rect 2372 11308 2605 11336
rect 2372 11296 2378 11308
rect 2593 11305 2605 11308
rect 2639 11305 2651 11339
rect 2593 11299 2651 11305
rect 2869 11339 2927 11345
rect 2869 11305 2881 11339
rect 2915 11336 2927 11339
rect 2958 11336 2964 11348
rect 2915 11308 2964 11336
rect 2915 11305 2927 11308
rect 2869 11299 2927 11305
rect 2958 11296 2964 11308
rect 3016 11296 3022 11348
rect 3145 11339 3203 11345
rect 3145 11305 3157 11339
rect 3191 11336 3203 11339
rect 6454 11336 6460 11348
rect 3191 11308 6316 11336
rect 6415 11308 6460 11336
rect 3191 11305 3203 11308
rect 3145 11299 3203 11305
rect 1857 11271 1915 11277
rect 1857 11237 1869 11271
rect 1903 11237 1915 11271
rect 1857 11231 1915 11237
rect 1302 11132 1308 11144
rect 1263 11104 1308 11132
rect 1302 11092 1308 11104
rect 1360 11092 1366 11144
rect 1581 11135 1639 11141
rect 1581 11101 1593 11135
rect 1627 11132 1639 11135
rect 1872 11132 1900 11231
rect 1946 11228 1952 11280
rect 2004 11268 2010 11280
rect 3973 11271 4031 11277
rect 3973 11268 3985 11271
rect 2004 11240 3985 11268
rect 2004 11228 2010 11240
rect 3973 11237 3985 11240
rect 4019 11237 4031 11271
rect 4338 11268 4344 11280
rect 4299 11240 4344 11268
rect 3973 11231 4031 11237
rect 4338 11228 4344 11240
rect 4396 11228 4402 11280
rect 4433 11271 4491 11277
rect 4433 11237 4445 11271
rect 4479 11268 4491 11271
rect 4798 11268 4804 11280
rect 4479 11240 4804 11268
rect 4479 11237 4491 11240
rect 4433 11231 4491 11237
rect 4798 11228 4804 11240
rect 4856 11228 4862 11280
rect 4985 11271 5043 11277
rect 4985 11237 4997 11271
rect 5031 11268 5043 11271
rect 5258 11268 5264 11280
rect 5031 11240 5264 11268
rect 5031 11237 5043 11240
rect 4985 11231 5043 11237
rect 5258 11228 5264 11240
rect 5316 11228 5322 11280
rect 5442 11268 5448 11280
rect 5403 11240 5448 11268
rect 5442 11228 5448 11240
rect 5500 11228 5506 11280
rect 6178 11268 6184 11280
rect 6139 11240 6184 11268
rect 6178 11228 6184 11240
rect 6236 11228 6242 11280
rect 6288 11268 6316 11308
rect 6454 11296 6460 11308
rect 6512 11296 6518 11348
rect 6917 11339 6975 11345
rect 6917 11305 6929 11339
rect 6963 11336 6975 11339
rect 7098 11336 7104 11348
rect 6963 11308 7104 11336
rect 6963 11305 6975 11308
rect 6917 11299 6975 11305
rect 7098 11296 7104 11308
rect 7156 11296 7162 11348
rect 7190 11296 7196 11348
rect 7248 11336 7254 11348
rect 7653 11339 7711 11345
rect 7653 11336 7665 11339
rect 7248 11308 7665 11336
rect 7248 11296 7254 11308
rect 7653 11305 7665 11308
rect 7699 11305 7711 11339
rect 7926 11336 7932 11348
rect 7887 11308 7932 11336
rect 7653 11299 7711 11305
rect 7926 11296 7932 11308
rect 7984 11296 7990 11348
rect 8478 11336 8484 11348
rect 8439 11308 8484 11336
rect 8478 11296 8484 11308
rect 8536 11296 8542 11348
rect 8662 11296 8668 11348
rect 8720 11336 8726 11348
rect 8757 11339 8815 11345
rect 8757 11336 8769 11339
rect 8720 11308 8769 11336
rect 8720 11296 8726 11308
rect 8757 11305 8769 11308
rect 8803 11305 8815 11339
rect 8757 11299 8815 11305
rect 6638 11268 6644 11280
rect 6288 11240 6644 11268
rect 6638 11228 6644 11240
rect 6696 11228 6702 11280
rect 7377 11271 7435 11277
rect 7377 11237 7389 11271
rect 7423 11237 7435 11271
rect 7377 11231 7435 11237
rect 7282 11200 7288 11212
rect 3436 11172 5304 11200
rect 3436 11144 3464 11172
rect 2038 11132 2044 11144
rect 1627 11104 1900 11132
rect 1999 11104 2044 11132
rect 1627 11101 1639 11104
rect 1581 11095 1639 11101
rect 2038 11092 2044 11104
rect 2096 11092 2102 11144
rect 2133 11135 2191 11141
rect 2133 11101 2145 11135
rect 2179 11132 2191 11135
rect 2222 11132 2228 11144
rect 2179 11104 2228 11132
rect 2179 11101 2191 11104
rect 2133 11095 2191 11101
rect 2222 11092 2228 11104
rect 2280 11092 2286 11144
rect 2406 11132 2412 11144
rect 2367 11104 2412 11132
rect 2406 11092 2412 11104
rect 2464 11092 2470 11144
rect 2682 11132 2688 11144
rect 2643 11104 2688 11132
rect 2682 11092 2688 11104
rect 2740 11092 2746 11144
rect 2958 11132 2964 11144
rect 2919 11104 2964 11132
rect 2958 11092 2964 11104
rect 3016 11092 3022 11144
rect 3418 11132 3424 11144
rect 3331 11104 3424 11132
rect 3418 11092 3424 11104
rect 3476 11092 3482 11144
rect 3510 11092 3516 11144
rect 3568 11132 3574 11144
rect 3789 11135 3847 11141
rect 3789 11132 3801 11135
rect 3568 11104 3801 11132
rect 3568 11092 3574 11104
rect 3789 11101 3801 11104
rect 3835 11101 3847 11135
rect 3789 11095 3847 11101
rect 3878 11092 3884 11144
rect 3936 11132 3942 11144
rect 4157 11135 4215 11141
rect 4157 11132 4169 11135
rect 3936 11104 4169 11132
rect 3936 11092 3942 11104
rect 4157 11101 4169 11104
rect 4203 11101 4215 11135
rect 4157 11095 4215 11101
rect 4522 11092 4528 11144
rect 4580 11132 4586 11144
rect 4617 11135 4675 11141
rect 4617 11132 4629 11135
rect 4580 11104 4629 11132
rect 4580 11092 4586 11104
rect 4617 11101 4629 11104
rect 4663 11101 4675 11135
rect 4617 11095 4675 11101
rect 4801 11135 4859 11141
rect 4801 11101 4813 11135
rect 4847 11134 4859 11135
rect 4847 11132 4936 11134
rect 5074 11132 5080 11144
rect 4847 11106 5080 11132
rect 4847 11101 4859 11106
rect 4908 11104 5080 11106
rect 4801 11095 4859 11101
rect 5074 11092 5080 11104
rect 5132 11092 5138 11144
rect 5276 11141 5304 11172
rect 5644 11172 7288 11200
rect 5644 11141 5672 11172
rect 7282 11160 7288 11172
rect 7340 11160 7346 11212
rect 7392 11200 7420 11231
rect 9858 11200 9864 11212
rect 7392 11172 9864 11200
rect 9858 11160 9864 11172
rect 9916 11160 9922 11212
rect 5261 11135 5319 11141
rect 5261 11101 5273 11135
rect 5307 11101 5319 11135
rect 5261 11095 5319 11101
rect 5629 11135 5687 11141
rect 5629 11101 5641 11135
rect 5675 11101 5687 11135
rect 5629 11095 5687 11101
rect 5721 11135 5779 11141
rect 5721 11101 5733 11135
rect 5767 11101 5779 11135
rect 5721 11095 5779 11101
rect 3602 11024 3608 11076
rect 3660 11064 3666 11076
rect 3660 11036 3705 11064
rect 3660 11024 3666 11036
rect 3970 11024 3976 11076
rect 4028 11064 4034 11076
rect 5736 11064 5764 11095
rect 5810 11092 5816 11144
rect 5868 11132 5874 11144
rect 6641 11135 6699 11141
rect 6641 11132 6653 11135
rect 5868 11104 6653 11132
rect 5868 11092 5874 11104
rect 6641 11101 6653 11104
rect 6687 11132 6699 11135
rect 6730 11132 6736 11144
rect 6687 11104 6736 11132
rect 6687 11101 6699 11104
rect 6641 11095 6699 11101
rect 6730 11092 6736 11104
rect 6788 11092 6794 11144
rect 7098 11132 7104 11144
rect 7059 11104 7104 11132
rect 7098 11092 7104 11104
rect 7156 11092 7162 11144
rect 7561 11135 7619 11141
rect 7561 11101 7573 11135
rect 7607 11132 7619 11135
rect 7650 11132 7656 11144
rect 7607 11104 7656 11132
rect 7607 11101 7619 11104
rect 7561 11095 7619 11101
rect 7650 11092 7656 11104
rect 7708 11092 7714 11144
rect 8110 11132 8116 11144
rect 8071 11104 8116 11132
rect 8110 11092 8116 11104
rect 8168 11092 8174 11144
rect 8202 11092 8208 11144
rect 8260 11132 8266 11144
rect 8297 11135 8355 11141
rect 8297 11132 8309 11135
rect 8260 11104 8309 11132
rect 8260 11092 8266 11104
rect 8297 11101 8309 11104
rect 8343 11101 8355 11135
rect 8297 11095 8355 11101
rect 8941 11135 8999 11141
rect 8941 11101 8953 11135
rect 8987 11132 8999 11135
rect 9122 11132 9128 11144
rect 8987 11104 9128 11132
rect 8987 11101 8999 11104
rect 8941 11095 8999 11101
rect 9122 11092 9128 11104
rect 9180 11092 9186 11144
rect 9309 11135 9367 11141
rect 9309 11101 9321 11135
rect 9355 11132 9367 11135
rect 9355 11104 9536 11132
rect 9355 11101 9367 11104
rect 9309 11095 9367 11101
rect 4028 11036 4752 11064
rect 4028 11024 4034 11036
rect 1854 10956 1860 11008
rect 1912 10996 1918 11008
rect 2130 10996 2136 11008
rect 1912 10968 2136 10996
rect 1912 10956 1918 10968
rect 2130 10956 2136 10968
rect 2188 10956 2194 11008
rect 2317 10999 2375 11005
rect 2317 10965 2329 10999
rect 2363 10996 2375 10999
rect 2406 10996 2412 11008
rect 2363 10968 2412 10996
rect 2363 10965 2375 10968
rect 2317 10959 2375 10965
rect 2406 10956 2412 10968
rect 2464 10956 2470 11008
rect 2958 10956 2964 11008
rect 3016 10996 3022 11008
rect 3237 10999 3295 11005
rect 3237 10996 3249 10999
rect 3016 10968 3249 10996
rect 3016 10956 3022 10968
rect 3237 10965 3249 10968
rect 3283 10965 3295 10999
rect 4724 10996 4752 11036
rect 4908 11036 5764 11064
rect 4908 10996 4936 11036
rect 6454 11024 6460 11076
rect 6512 11064 6518 11076
rect 7926 11064 7932 11076
rect 6512 11036 7932 11064
rect 6512 11024 6518 11036
rect 7926 11024 7932 11036
rect 7984 11024 7990 11076
rect 5074 10996 5080 11008
rect 4724 10968 4936 10996
rect 5035 10968 5080 10996
rect 3237 10959 3295 10965
rect 5074 10956 5080 10968
rect 5132 10956 5138 11008
rect 5902 10996 5908 11008
rect 5863 10968 5908 10996
rect 5902 10956 5908 10968
rect 5960 10956 5966 11008
rect 6270 10956 6276 11008
rect 6328 10996 6334 11008
rect 9508 11005 9536 11104
rect 9125 10999 9183 11005
rect 9125 10996 9137 10999
rect 6328 10968 9137 10996
rect 6328 10956 6334 10968
rect 9125 10965 9137 10968
rect 9171 10965 9183 10999
rect 9125 10959 9183 10965
rect 9493 10999 9551 11005
rect 9493 10965 9505 10999
rect 9539 10996 9551 10999
rect 9582 10996 9588 11008
rect 9539 10968 9588 10996
rect 9539 10965 9551 10968
rect 9493 10959 9551 10965
rect 9582 10956 9588 10968
rect 9640 10956 9646 11008
rect 920 10906 9844 10928
rect 920 10854 4116 10906
rect 4168 10854 4180 10906
rect 4232 10854 4244 10906
rect 4296 10854 4308 10906
rect 4360 10854 4372 10906
rect 4424 10854 7216 10906
rect 7268 10854 7280 10906
rect 7332 10854 7344 10906
rect 7396 10854 7408 10906
rect 7460 10854 7472 10906
rect 7524 10854 9844 10906
rect 920 10832 9844 10854
rect 1486 10792 1492 10804
rect 1447 10764 1492 10792
rect 1486 10752 1492 10764
rect 1544 10752 1550 10804
rect 2222 10752 2228 10804
rect 2280 10792 2286 10804
rect 2317 10795 2375 10801
rect 2317 10792 2329 10795
rect 2280 10764 2329 10792
rect 2280 10752 2286 10764
rect 2317 10761 2329 10764
rect 2363 10761 2375 10795
rect 3050 10792 3056 10804
rect 3011 10764 3056 10792
rect 2317 10755 2375 10761
rect 3050 10752 3056 10764
rect 3108 10752 3114 10804
rect 3326 10752 3332 10804
rect 3384 10792 3390 10804
rect 3510 10792 3516 10804
rect 3384 10764 3516 10792
rect 3384 10752 3390 10764
rect 3510 10752 3516 10764
rect 3568 10792 3574 10804
rect 3697 10795 3755 10801
rect 3697 10792 3709 10795
rect 3568 10764 3709 10792
rect 3568 10752 3574 10764
rect 3697 10761 3709 10764
rect 3743 10761 3755 10795
rect 5445 10795 5503 10801
rect 3697 10755 3755 10761
rect 4126 10764 5396 10792
rect 4126 10724 4154 10764
rect 1320 10696 4154 10724
rect 5368 10724 5396 10764
rect 5445 10761 5457 10795
rect 5491 10792 5503 10795
rect 7006 10792 7012 10804
rect 5491 10764 7012 10792
rect 5491 10761 5503 10764
rect 5445 10755 5503 10761
rect 7006 10752 7012 10764
rect 7064 10752 7070 10804
rect 8478 10752 8484 10804
rect 8536 10752 8542 10804
rect 8570 10752 8576 10804
rect 8628 10792 8634 10804
rect 8941 10795 8999 10801
rect 8941 10792 8953 10795
rect 8628 10764 8953 10792
rect 8628 10752 8634 10764
rect 8941 10761 8953 10764
rect 8987 10761 8999 10795
rect 8941 10755 8999 10761
rect 5629 10727 5687 10733
rect 5629 10724 5641 10727
rect 5368 10696 5641 10724
rect 1320 10665 1348 10696
rect 5629 10693 5641 10696
rect 5675 10693 5687 10727
rect 5810 10724 5816 10736
rect 5771 10696 5816 10724
rect 5629 10687 5687 10693
rect 5810 10684 5816 10696
rect 5868 10684 5874 10736
rect 6914 10684 6920 10736
rect 6972 10684 6978 10736
rect 8496 10724 8524 10752
rect 9033 10727 9091 10733
rect 9033 10724 9045 10727
rect 8496 10696 9045 10724
rect 9033 10693 9045 10696
rect 9079 10693 9091 10727
rect 9033 10687 9091 10693
rect 1305 10659 1363 10665
rect 1305 10625 1317 10659
rect 1351 10625 1363 10659
rect 1578 10656 1584 10668
rect 1539 10628 1584 10656
rect 1305 10619 1363 10625
rect 1578 10616 1584 10628
rect 1636 10616 1642 10668
rect 1857 10659 1915 10665
rect 1857 10625 1869 10659
rect 1903 10625 1915 10659
rect 1857 10619 1915 10625
rect 1872 10588 1900 10619
rect 1946 10616 1952 10668
rect 2004 10656 2010 10668
rect 2133 10659 2191 10665
rect 2133 10656 2145 10659
rect 2004 10628 2145 10656
rect 2004 10616 2010 10628
rect 2133 10625 2145 10628
rect 2179 10625 2191 10659
rect 2133 10619 2191 10625
rect 2222 10616 2228 10668
rect 2280 10656 2286 10668
rect 2409 10659 2467 10665
rect 2409 10656 2421 10659
rect 2280 10628 2421 10656
rect 2280 10616 2286 10628
rect 2409 10625 2421 10628
rect 2455 10625 2467 10659
rect 2409 10619 2467 10625
rect 2866 10616 2872 10668
rect 2924 10656 2930 10668
rect 3510 10656 3516 10668
rect 2924 10628 3516 10656
rect 2924 10616 2930 10628
rect 3510 10616 3516 10628
rect 3568 10616 3574 10668
rect 3602 10616 3608 10668
rect 3660 10656 3666 10668
rect 4246 10656 4252 10668
rect 3660 10628 3705 10656
rect 4207 10628 4252 10656
rect 3660 10616 3666 10628
rect 4246 10616 4252 10628
rect 4304 10656 4310 10668
rect 4341 10659 4399 10665
rect 4341 10656 4353 10659
rect 4304 10628 4353 10656
rect 4304 10616 4310 10628
rect 4341 10625 4353 10628
rect 4387 10625 4399 10659
rect 4341 10619 4399 10625
rect 4525 10659 4583 10665
rect 4525 10625 4537 10659
rect 4571 10625 4583 10659
rect 4525 10619 4583 10625
rect 4801 10659 4859 10665
rect 4801 10625 4813 10659
rect 4847 10656 4859 10659
rect 4890 10656 4896 10668
rect 4847 10628 4896 10656
rect 4847 10625 4859 10628
rect 4801 10619 4859 10625
rect 3789 10591 3847 10597
rect 3789 10588 3801 10591
rect 1872 10560 3801 10588
rect 3789 10557 3801 10560
rect 3835 10557 3847 10591
rect 3970 10588 3976 10600
rect 3789 10551 3847 10557
rect 3896 10560 3976 10588
rect 1765 10523 1823 10529
rect 1765 10489 1777 10523
rect 1811 10520 1823 10523
rect 2866 10520 2872 10532
rect 1811 10492 2872 10520
rect 1811 10489 1823 10492
rect 1765 10483 1823 10489
rect 2866 10480 2872 10492
rect 2924 10480 2930 10532
rect 2958 10480 2964 10532
rect 3016 10520 3022 10532
rect 3145 10523 3203 10529
rect 3145 10520 3157 10523
rect 3016 10492 3157 10520
rect 3016 10480 3022 10492
rect 3145 10489 3157 10492
rect 3191 10489 3203 10523
rect 3896 10520 3924 10560
rect 3970 10548 3976 10560
rect 4028 10548 4034 10600
rect 4540 10588 4568 10619
rect 4890 10616 4896 10628
rect 4948 10616 4954 10668
rect 4982 10616 4988 10668
rect 5040 10656 5046 10668
rect 5261 10659 5319 10665
rect 5261 10656 5273 10659
rect 5040 10628 5273 10656
rect 5040 10616 5046 10628
rect 5261 10625 5273 10628
rect 5307 10625 5319 10659
rect 5261 10619 5319 10625
rect 5997 10659 6055 10665
rect 5997 10625 6009 10659
rect 6043 10656 6055 10659
rect 6454 10656 6460 10668
rect 6043 10628 6460 10656
rect 6043 10625 6055 10628
rect 5997 10619 6055 10625
rect 6454 10616 6460 10628
rect 6512 10616 6518 10668
rect 8018 10656 8024 10668
rect 7979 10628 8024 10656
rect 8018 10616 8024 10628
rect 8076 10616 8082 10668
rect 8110 10616 8116 10668
rect 8168 10656 8174 10668
rect 8573 10662 8631 10665
rect 8496 10659 8631 10662
rect 8496 10656 8585 10659
rect 8168 10634 8585 10656
rect 8168 10628 8524 10634
rect 8168 10616 8174 10628
rect 8573 10625 8585 10634
rect 8619 10625 8631 10659
rect 8573 10619 8631 10625
rect 8757 10659 8815 10665
rect 8757 10625 8769 10659
rect 8803 10625 8815 10659
rect 8757 10619 8815 10625
rect 9217 10659 9275 10665
rect 9217 10625 9229 10659
rect 9263 10656 9275 10659
rect 9306 10656 9312 10668
rect 9263 10628 9312 10656
rect 9263 10625 9275 10628
rect 9217 10619 9275 10625
rect 4264 10560 4568 10588
rect 4264 10520 4292 10560
rect 4706 10548 4712 10600
rect 4764 10588 4770 10600
rect 6181 10591 6239 10597
rect 6181 10588 6193 10591
rect 4764 10560 6193 10588
rect 4764 10548 4770 10560
rect 6181 10557 6193 10560
rect 6227 10557 6239 10591
rect 6546 10588 6552 10600
rect 6507 10560 6552 10588
rect 6181 10551 6239 10557
rect 6546 10548 6552 10560
rect 6604 10548 6610 10600
rect 8772 10588 8800 10619
rect 9306 10616 9312 10628
rect 9364 10616 9370 10668
rect 8266 10560 8800 10588
rect 9401 10591 9459 10597
rect 3145 10483 3203 10489
rect 3252 10492 3924 10520
rect 4126 10492 4292 10520
rect 2041 10455 2099 10461
rect 2041 10421 2053 10455
rect 2087 10452 2099 10455
rect 3252 10452 3280 10492
rect 2087 10424 3280 10452
rect 3513 10455 3571 10461
rect 2087 10421 2099 10424
rect 2041 10415 2099 10421
rect 3513 10421 3525 10455
rect 3559 10452 3571 10455
rect 3697 10455 3755 10461
rect 3697 10452 3709 10455
rect 3559 10424 3709 10452
rect 3559 10421 3571 10424
rect 3513 10415 3571 10421
rect 3697 10421 3709 10424
rect 3743 10452 3755 10455
rect 3973 10455 4031 10461
rect 3973 10452 3985 10455
rect 3743 10424 3985 10452
rect 3743 10421 3755 10424
rect 3697 10415 3755 10421
rect 3973 10421 3985 10424
rect 4019 10452 4031 10455
rect 4126 10452 4154 10492
rect 4338 10480 4344 10532
rect 4396 10520 4402 10532
rect 4396 10492 4752 10520
rect 4396 10480 4402 10492
rect 4724 10461 4752 10492
rect 8018 10480 8024 10532
rect 8076 10520 8082 10532
rect 8266 10520 8294 10560
rect 9401 10557 9413 10591
rect 9447 10588 9459 10591
rect 9582 10588 9588 10600
rect 9447 10560 9588 10588
rect 9447 10557 9459 10560
rect 9401 10551 9459 10557
rect 9582 10548 9588 10560
rect 9640 10548 9646 10600
rect 8076 10492 8294 10520
rect 8481 10523 8539 10529
rect 8076 10480 8082 10492
rect 8481 10489 8493 10523
rect 8527 10520 8539 10523
rect 9214 10520 9220 10532
rect 8527 10492 9220 10520
rect 8527 10489 8539 10492
rect 8481 10483 8539 10489
rect 9214 10480 9220 10492
rect 9272 10480 9278 10532
rect 4019 10424 4154 10452
rect 4709 10455 4767 10461
rect 4019 10421 4031 10424
rect 3973 10415 4031 10421
rect 4709 10421 4721 10455
rect 4755 10421 4767 10455
rect 4982 10452 4988 10464
rect 4943 10424 4988 10452
rect 4709 10415 4767 10421
rect 4982 10412 4988 10424
rect 5040 10412 5046 10464
rect 5169 10455 5227 10461
rect 5169 10421 5181 10455
rect 5215 10452 5227 10455
rect 7006 10452 7012 10464
rect 5215 10424 7012 10452
rect 5215 10421 5227 10424
rect 5169 10415 5227 10421
rect 7006 10412 7012 10424
rect 7064 10412 7070 10464
rect 15194 10412 15200 10464
rect 15252 10452 15258 10464
rect 16574 10452 16580 10464
rect 15252 10424 16580 10452
rect 15252 10412 15258 10424
rect 16574 10412 16580 10424
rect 16632 10412 16638 10464
rect 920 10362 9844 10384
rect 920 10310 2566 10362
rect 2618 10310 2630 10362
rect 2682 10310 2694 10362
rect 2746 10310 2758 10362
rect 2810 10310 2822 10362
rect 2874 10310 5666 10362
rect 5718 10310 5730 10362
rect 5782 10310 5794 10362
rect 5846 10310 5858 10362
rect 5910 10310 5922 10362
rect 5974 10310 8766 10362
rect 8818 10310 8830 10362
rect 8882 10310 8894 10362
rect 8946 10310 8958 10362
rect 9010 10310 9022 10362
rect 9074 10310 9844 10362
rect 920 10288 9844 10310
rect 3163 10251 3221 10257
rect 3163 10217 3175 10251
rect 3209 10248 3221 10251
rect 6089 10251 6147 10257
rect 6089 10248 6101 10251
rect 3209 10220 6101 10248
rect 3209 10217 3221 10220
rect 3163 10211 3221 10217
rect 6089 10217 6101 10220
rect 6135 10248 6147 10251
rect 6178 10248 6184 10260
rect 6135 10220 6184 10248
rect 6135 10217 6147 10220
rect 6089 10211 6147 10217
rect 6178 10208 6184 10220
rect 6236 10208 6242 10260
rect 7558 10208 7564 10260
rect 7616 10248 7622 10260
rect 7929 10251 7987 10257
rect 7929 10248 7941 10251
rect 7616 10220 7941 10248
rect 7616 10208 7622 10220
rect 7929 10217 7941 10220
rect 7975 10217 7987 10251
rect 7929 10211 7987 10217
rect 8018 10208 8024 10260
rect 8076 10248 8082 10260
rect 8113 10251 8171 10257
rect 8113 10248 8125 10251
rect 8076 10220 8125 10248
rect 8076 10208 8082 10220
rect 8113 10217 8125 10220
rect 8159 10248 8171 10251
rect 8159 10220 8984 10248
rect 8159 10217 8171 10220
rect 8113 10211 8171 10217
rect 8956 10192 8984 10220
rect 5074 10140 5080 10192
rect 5132 10180 5138 10192
rect 5626 10180 5632 10192
rect 5132 10152 5632 10180
rect 5132 10140 5138 10152
rect 5626 10140 5632 10152
rect 5684 10140 5690 10192
rect 6454 10180 6460 10192
rect 6380 10152 6460 10180
rect 2406 10072 2412 10124
rect 2464 10112 2470 10124
rect 3697 10115 3755 10121
rect 3697 10112 3709 10115
rect 2464 10084 3709 10112
rect 2464 10072 2470 10084
rect 3697 10081 3709 10084
rect 3743 10081 3755 10115
rect 3697 10075 3755 10081
rect 1394 10044 1400 10056
rect 1355 10016 1400 10044
rect 1394 10004 1400 10016
rect 1452 10004 1458 10056
rect 3421 10047 3479 10053
rect 3421 10013 3433 10047
rect 3467 10013 3479 10047
rect 3421 10007 3479 10013
rect 2682 9936 2688 9988
rect 2740 9936 2746 9988
rect 3436 9976 3464 10007
rect 3602 10004 3608 10056
rect 3660 10044 3666 10056
rect 3878 10044 3884 10056
rect 3660 10016 3884 10044
rect 3660 10004 3666 10016
rect 3878 10004 3884 10016
rect 3936 10004 3942 10056
rect 3970 10004 3976 10056
rect 4028 10044 4034 10056
rect 4065 10047 4123 10053
rect 4065 10044 4077 10047
rect 4028 10016 4077 10044
rect 4028 10004 4034 10016
rect 4065 10013 4077 10016
rect 4111 10013 4123 10047
rect 4065 10007 4123 10013
rect 5537 10047 5595 10053
rect 5537 10013 5549 10047
rect 5583 10013 5595 10047
rect 5537 10007 5595 10013
rect 3344 9948 3464 9976
rect 3344 9920 3372 9948
rect 4430 9936 4436 9988
rect 4488 9936 4494 9988
rect 1578 9908 1584 9920
rect 1539 9880 1584 9908
rect 1578 9868 1584 9880
rect 1636 9868 1642 9920
rect 1673 9911 1731 9917
rect 1673 9877 1685 9911
rect 1719 9908 1731 9911
rect 1854 9908 1860 9920
rect 1719 9880 1860 9908
rect 1719 9877 1731 9880
rect 1673 9871 1731 9877
rect 1854 9868 1860 9880
rect 1912 9868 1918 9920
rect 3326 9868 3332 9920
rect 3384 9868 3390 9920
rect 3510 9868 3516 9920
rect 3568 9908 3574 9920
rect 5552 9908 5580 10007
rect 5810 9936 5816 9988
rect 5868 9976 5874 9988
rect 6380 9976 6408 10152
rect 6454 10140 6460 10152
rect 6512 10140 6518 10192
rect 8570 10180 8576 10192
rect 8531 10152 8576 10180
rect 8570 10140 8576 10152
rect 8628 10140 8634 10192
rect 8938 10140 8944 10192
rect 8996 10140 9002 10192
rect 9122 10180 9128 10192
rect 9083 10152 9128 10180
rect 9122 10140 9128 10152
rect 9180 10140 9186 10192
rect 9401 10183 9459 10189
rect 9401 10149 9413 10183
rect 9447 10149 9459 10183
rect 9401 10143 9459 10149
rect 7558 10072 7564 10124
rect 7616 10112 7622 10124
rect 9416 10112 9444 10143
rect 7616 10084 9444 10112
rect 7616 10072 7622 10084
rect 7837 10047 7895 10053
rect 7837 10013 7849 10047
rect 7883 10044 7895 10047
rect 8018 10044 8024 10056
rect 7883 10016 8024 10044
rect 7883 10013 7895 10016
rect 7837 10007 7895 10013
rect 8018 10004 8024 10016
rect 8076 10004 8082 10056
rect 8110 10004 8116 10056
rect 8168 10044 8174 10056
rect 8389 10047 8447 10053
rect 8389 10046 8401 10047
rect 8266 10044 8401 10046
rect 8168 10018 8401 10044
rect 8168 10016 8294 10018
rect 8168 10004 8174 10016
rect 8389 10013 8401 10018
rect 8435 10013 8447 10047
rect 8389 10007 8447 10013
rect 8846 10004 8852 10056
rect 8904 10044 8910 10056
rect 9217 10047 9275 10053
rect 9217 10044 9229 10047
rect 8904 10016 9229 10044
rect 8904 10004 8910 10016
rect 9217 10013 9229 10016
rect 9263 10013 9275 10047
rect 9217 10007 9275 10013
rect 5868 9962 6408 9976
rect 7561 9979 7619 9985
rect 5868 9948 6394 9962
rect 5868 9936 5874 9948
rect 7561 9945 7573 9979
rect 7607 9976 7619 9979
rect 7926 9976 7932 9988
rect 7607 9948 7932 9976
rect 7607 9945 7619 9948
rect 7561 9939 7619 9945
rect 7926 9936 7932 9948
rect 7984 9936 7990 9988
rect 8757 9979 8815 9985
rect 8757 9945 8769 9979
rect 8803 9945 8815 9979
rect 8938 9976 8944 9988
rect 8899 9948 8944 9976
rect 8757 9939 8815 9945
rect 3568 9880 5580 9908
rect 5997 9911 6055 9917
rect 3568 9868 3574 9880
rect 5997 9877 6009 9911
rect 6043 9908 6055 9911
rect 6638 9908 6644 9920
rect 6043 9880 6644 9908
rect 6043 9877 6055 9880
rect 5997 9871 6055 9877
rect 6638 9868 6644 9880
rect 6696 9868 6702 9920
rect 8018 9868 8024 9920
rect 8076 9908 8082 9920
rect 8772 9908 8800 9939
rect 8938 9936 8944 9948
rect 8996 9936 9002 9988
rect 8076 9880 8800 9908
rect 8076 9868 8082 9880
rect 920 9818 9844 9840
rect 920 9766 4116 9818
rect 4168 9766 4180 9818
rect 4232 9766 4244 9818
rect 4296 9766 4308 9818
rect 4360 9766 4372 9818
rect 4424 9766 7216 9818
rect 7268 9766 7280 9818
rect 7332 9766 7344 9818
rect 7396 9766 7408 9818
rect 7460 9766 7472 9818
rect 7524 9766 9844 9818
rect 920 9744 9844 9766
rect 1489 9707 1547 9713
rect 1489 9673 1501 9707
rect 1535 9704 1547 9707
rect 1946 9704 1952 9716
rect 1535 9676 1952 9704
rect 1535 9673 1547 9676
rect 1489 9667 1547 9673
rect 1946 9664 1952 9676
rect 2004 9664 2010 9716
rect 2038 9664 2044 9716
rect 2096 9704 2102 9716
rect 2501 9707 2559 9713
rect 2501 9704 2513 9707
rect 2096 9676 2513 9704
rect 2096 9664 2102 9676
rect 2501 9673 2513 9676
rect 2547 9673 2559 9707
rect 2501 9667 2559 9673
rect 2590 9664 2596 9716
rect 2648 9704 2654 9716
rect 3602 9704 3608 9716
rect 2648 9676 3608 9704
rect 2648 9664 2654 9676
rect 3602 9664 3608 9676
rect 3660 9664 3666 9716
rect 3786 9664 3792 9716
rect 3844 9704 3850 9716
rect 4985 9707 5043 9713
rect 3844 9676 4752 9704
rect 3844 9664 3850 9676
rect 1412 9608 2636 9636
rect 1302 9568 1308 9580
rect 1215 9540 1308 9568
rect 1302 9528 1308 9540
rect 1360 9568 1366 9580
rect 1412 9577 1440 9608
rect 1397 9571 1455 9577
rect 1397 9568 1409 9571
rect 1360 9540 1409 9568
rect 1360 9528 1366 9540
rect 1397 9537 1409 9540
rect 1443 9537 1455 9571
rect 1397 9531 1455 9537
rect 1673 9571 1731 9577
rect 1673 9537 1685 9571
rect 1719 9568 1731 9571
rect 1854 9568 1860 9580
rect 1719 9540 1860 9568
rect 1719 9537 1731 9540
rect 1673 9531 1731 9537
rect 1854 9528 1860 9540
rect 1912 9528 1918 9580
rect 2608 9577 2636 9608
rect 3510 9596 3516 9648
rect 3568 9596 3574 9648
rect 4724 9636 4752 9676
rect 4985 9673 4997 9707
rect 5031 9704 5043 9707
rect 5031 9676 6500 9704
rect 5031 9673 5043 9676
rect 4985 9667 5043 9673
rect 5169 9639 5227 9645
rect 5169 9636 5181 9639
rect 4724 9608 5181 9636
rect 5169 9605 5181 9608
rect 5215 9605 5227 9639
rect 5169 9599 5227 9605
rect 2593 9571 2651 9577
rect 2593 9537 2605 9571
rect 2639 9568 2651 9571
rect 2639 9540 3188 9568
rect 2639 9537 2651 9540
rect 2593 9531 2651 9537
rect 2314 9460 2320 9512
rect 2372 9500 2378 9512
rect 2685 9503 2743 9509
rect 2685 9500 2697 9503
rect 2372 9472 2697 9500
rect 2372 9460 2378 9472
rect 2685 9469 2697 9472
rect 2731 9469 2743 9503
rect 3050 9500 3056 9512
rect 3011 9472 3056 9500
rect 2685 9463 2743 9469
rect 3050 9460 3056 9472
rect 3108 9460 3114 9512
rect 3160 9500 3188 9540
rect 4062 9528 4068 9580
rect 4120 9568 4126 9580
rect 4525 9571 4583 9577
rect 4525 9568 4537 9571
rect 4120 9540 4537 9568
rect 4120 9528 4126 9540
rect 4525 9537 4537 9540
rect 4571 9537 4583 9571
rect 4525 9531 4583 9537
rect 5077 9571 5135 9577
rect 5077 9537 5089 9571
rect 5123 9568 5135 9571
rect 5353 9571 5411 9577
rect 5353 9568 5365 9571
rect 5123 9540 5365 9568
rect 5123 9537 5135 9540
rect 5077 9531 5135 9537
rect 5353 9537 5365 9540
rect 5399 9537 5411 9571
rect 5353 9531 5411 9537
rect 5537 9571 5595 9577
rect 5537 9537 5549 9571
rect 5583 9537 5595 9571
rect 5537 9531 5595 9537
rect 3694 9500 3700 9512
rect 3160 9472 3700 9500
rect 3694 9460 3700 9472
rect 3752 9460 3758 9512
rect 4890 9460 4896 9512
rect 4948 9500 4954 9512
rect 5552 9500 5580 9531
rect 5626 9528 5632 9580
rect 5684 9568 5690 9580
rect 5684 9540 5729 9568
rect 5684 9528 5690 9540
rect 5810 9528 5816 9580
rect 5868 9568 5874 9580
rect 6178 9568 6184 9580
rect 5868 9540 5961 9568
rect 6139 9540 6184 9568
rect 5868 9528 5874 9540
rect 6178 9528 6184 9540
rect 6236 9528 6242 9580
rect 5718 9500 5724 9512
rect 4948 9472 5724 9500
rect 4948 9460 4954 9472
rect 5718 9460 5724 9472
rect 5776 9460 5782 9512
rect 753 9435 811 9441
rect 753 9401 765 9435
rect 799 9432 811 9435
rect 2590 9432 2596 9444
rect 799 9404 2596 9432
rect 799 9401 811 9404
rect 753 9395 811 9401
rect 2590 9392 2596 9404
rect 2648 9392 2654 9444
rect 5077 9435 5135 9441
rect 5077 9401 5089 9435
rect 5123 9432 5135 9435
rect 5166 9432 5172 9444
rect 5123 9404 5172 9432
rect 5123 9401 5135 9404
rect 5077 9395 5135 9401
rect 5166 9392 5172 9404
rect 5224 9432 5230 9444
rect 5828 9432 5856 9528
rect 6472 9500 6500 9676
rect 6546 9664 6552 9716
rect 6604 9704 6610 9716
rect 6825 9707 6883 9713
rect 6825 9704 6837 9707
rect 6604 9676 6837 9704
rect 6604 9664 6610 9676
rect 6825 9673 6837 9676
rect 6871 9673 6883 9707
rect 8570 9704 8576 9716
rect 6825 9667 6883 9673
rect 7944 9676 8576 9704
rect 7944 9636 7972 9676
rect 8570 9664 8576 9676
rect 8628 9664 8634 9716
rect 7116 9608 7972 9636
rect 7116 9580 7144 9608
rect 8386 9596 8392 9648
rect 8444 9596 8450 9648
rect 7098 9528 7104 9580
rect 7156 9568 7162 9580
rect 7653 9571 7711 9577
rect 7156 9540 7249 9568
rect 7156 9528 7162 9540
rect 7653 9537 7665 9571
rect 7699 9568 7711 9571
rect 7834 9568 7840 9580
rect 7699 9540 7840 9568
rect 7699 9537 7711 9540
rect 7653 9531 7711 9537
rect 7834 9528 7840 9540
rect 7892 9528 7898 9580
rect 9490 9568 9496 9580
rect 9451 9540 9496 9568
rect 9490 9528 9496 9540
rect 9548 9528 9554 9580
rect 9125 9503 9183 9509
rect 6472 9472 7328 9500
rect 7009 9435 7067 9441
rect 7009 9432 7021 9435
rect 5224 9404 5856 9432
rect 5920 9404 7021 9432
rect 5224 9392 5230 9404
rect 2222 9324 2228 9376
rect 2280 9364 2286 9376
rect 2317 9367 2375 9373
rect 2317 9364 2329 9367
rect 2280 9336 2329 9364
rect 2280 9324 2286 9336
rect 2317 9333 2329 9336
rect 2363 9333 2375 9367
rect 2317 9327 2375 9333
rect 3050 9324 3056 9376
rect 3108 9364 3114 9376
rect 4062 9364 4068 9376
rect 3108 9336 4068 9364
rect 3108 9324 3114 9336
rect 4062 9324 4068 9336
rect 4120 9324 4126 9376
rect 4614 9324 4620 9376
rect 4672 9364 4678 9376
rect 5442 9364 5448 9376
rect 4672 9336 5448 9364
rect 4672 9324 4678 9336
rect 5442 9324 5448 9336
rect 5500 9324 5506 9376
rect 5534 9324 5540 9376
rect 5592 9364 5598 9376
rect 5920 9364 5948 9404
rect 7009 9401 7021 9404
rect 7055 9401 7067 9435
rect 7009 9395 7067 9401
rect 5592 9336 5948 9364
rect 5997 9367 6055 9373
rect 5592 9324 5598 9336
rect 5997 9333 6009 9367
rect 6043 9364 6055 9367
rect 6914 9364 6920 9376
rect 6043 9336 6920 9364
rect 6043 9333 6055 9336
rect 5997 9327 6055 9333
rect 6914 9324 6920 9336
rect 6972 9324 6978 9376
rect 7190 9364 7196 9376
rect 7151 9336 7196 9364
rect 7190 9324 7196 9336
rect 7248 9324 7254 9376
rect 7300 9364 7328 9472
rect 9125 9469 9137 9503
rect 9171 9500 9183 9503
rect 9398 9500 9404 9512
rect 9171 9472 9404 9500
rect 9171 9469 9183 9472
rect 9125 9463 9183 9469
rect 9398 9460 9404 9472
rect 9456 9460 9462 9512
rect 9582 9364 9588 9376
rect 7300 9336 9588 9364
rect 9582 9324 9588 9336
rect 9640 9324 9646 9376
rect 920 9274 9844 9296
rect 920 9222 2566 9274
rect 2618 9222 2630 9274
rect 2682 9222 2694 9274
rect 2746 9222 2758 9274
rect 2810 9222 2822 9274
rect 2874 9222 5666 9274
rect 5718 9222 5730 9274
rect 5782 9222 5794 9274
rect 5846 9222 5858 9274
rect 5910 9222 5922 9274
rect 5974 9222 8766 9274
rect 8818 9222 8830 9274
rect 8882 9222 8894 9274
rect 8946 9222 8958 9274
rect 9010 9222 9022 9274
rect 9074 9222 9844 9274
rect 920 9200 9844 9222
rect 1486 9160 1492 9172
rect 1447 9132 1492 9160
rect 1486 9120 1492 9132
rect 1544 9120 1550 9172
rect 2314 9160 2320 9172
rect 2275 9132 2320 9160
rect 2314 9120 2320 9132
rect 2372 9120 2378 9172
rect 3234 9160 3240 9172
rect 2700 9132 3240 9160
rect 2041 9095 2099 9101
rect 2041 9061 2053 9095
rect 2087 9092 2099 9095
rect 2700 9092 2728 9132
rect 3234 9120 3240 9132
rect 3292 9120 3298 9172
rect 3418 9160 3424 9172
rect 3379 9132 3424 9160
rect 3418 9120 3424 9132
rect 3476 9120 3482 9172
rect 3694 9160 3700 9172
rect 3607 9132 3700 9160
rect 3694 9120 3700 9132
rect 3752 9160 3758 9172
rect 7098 9160 7104 9172
rect 3752 9132 7104 9160
rect 3752 9120 3758 9132
rect 7098 9120 7104 9132
rect 7156 9120 7162 9172
rect 9398 9160 9404 9172
rect 9359 9132 9404 9160
rect 9398 9120 9404 9132
rect 9456 9120 9462 9172
rect 2087 9064 2728 9092
rect 2869 9095 2927 9101
rect 2087 9061 2099 9064
rect 2041 9055 2099 9061
rect 2869 9061 2881 9095
rect 2915 9092 2927 9095
rect 3050 9092 3056 9104
rect 2915 9064 3056 9092
rect 2915 9061 2927 9064
rect 2869 9055 2927 9061
rect 3050 9052 3056 9064
rect 3108 9052 3114 9104
rect 3145 9095 3203 9101
rect 3145 9061 3157 9095
rect 3191 9092 3203 9095
rect 3510 9092 3516 9104
rect 3191 9064 3516 9092
rect 3191 9061 3203 9064
rect 3145 9055 3203 9061
rect 3510 9052 3516 9064
rect 3568 9052 3574 9104
rect 3970 9052 3976 9104
rect 4028 9092 4034 9104
rect 4801 9095 4859 9101
rect 4801 9092 4813 9095
rect 4028 9064 4813 9092
rect 4028 9052 4034 9064
rect 4801 9061 4813 9064
rect 4847 9061 4859 9095
rect 4801 9055 4859 9061
rect 5074 9024 5080 9036
rect 1596 8996 5080 9024
rect 1210 8916 1216 8968
rect 1268 8956 1274 8968
rect 1596 8965 1624 8996
rect 5074 8984 5080 8996
rect 5132 8984 5138 9036
rect 5166 8984 5172 9036
rect 5224 9024 5230 9036
rect 5353 9027 5411 9033
rect 5224 8996 5304 9024
rect 5224 8984 5230 8996
rect 1305 8959 1363 8965
rect 1305 8956 1317 8959
rect 1268 8928 1317 8956
rect 1268 8916 1274 8928
rect 1305 8925 1317 8928
rect 1351 8925 1363 8959
rect 1305 8919 1363 8925
rect 1581 8959 1639 8965
rect 1581 8925 1593 8959
rect 1627 8925 1639 8959
rect 1581 8919 1639 8925
rect 1857 8959 1915 8965
rect 1857 8925 1869 8959
rect 1903 8956 1915 8959
rect 2038 8956 2044 8968
rect 1903 8928 2044 8956
rect 1903 8925 1915 8928
rect 1857 8919 1915 8925
rect 2038 8916 2044 8928
rect 2096 8916 2102 8968
rect 2133 8959 2191 8965
rect 2133 8925 2145 8959
rect 2179 8956 2191 8959
rect 2593 8959 2651 8965
rect 2179 8928 2452 8956
rect 2179 8925 2191 8928
rect 2133 8919 2191 8925
rect 1670 8848 1676 8900
rect 1728 8888 1734 8900
rect 2314 8888 2320 8900
rect 1728 8860 2320 8888
rect 1728 8848 1734 8860
rect 2314 8848 2320 8860
rect 2372 8848 2378 8900
rect 1762 8820 1768 8832
rect 1723 8792 1768 8820
rect 1762 8780 1768 8792
rect 1820 8780 1826 8832
rect 2424 8829 2452 8928
rect 2593 8925 2605 8959
rect 2639 8925 2651 8959
rect 2593 8919 2651 8925
rect 2498 8848 2504 8900
rect 2556 8888 2562 8900
rect 2608 8888 2636 8919
rect 2682 8916 2688 8968
rect 2740 8956 2746 8968
rect 2958 8956 2964 8968
rect 2740 8928 2785 8956
rect 2919 8928 2964 8956
rect 2740 8916 2746 8928
rect 2958 8916 2964 8928
rect 3016 8916 3022 8968
rect 3050 8916 3056 8968
rect 3108 8956 3114 8968
rect 3237 8959 3295 8965
rect 3237 8956 3249 8959
rect 3108 8928 3249 8956
rect 3108 8916 3114 8928
rect 3237 8925 3249 8928
rect 3283 8925 3295 8959
rect 3237 8919 3295 8925
rect 4065 8959 4123 8965
rect 4065 8925 4077 8959
rect 4111 8925 4123 8959
rect 4065 8919 4123 8925
rect 3418 8888 3424 8900
rect 2556 8860 3424 8888
rect 2556 8848 2562 8860
rect 3418 8848 3424 8860
rect 3476 8848 3482 8900
rect 2409 8823 2467 8829
rect 2409 8789 2421 8823
rect 2455 8789 2467 8823
rect 3878 8820 3884 8832
rect 3839 8792 3884 8820
rect 2409 8783 2467 8789
rect 3878 8780 3884 8792
rect 3936 8780 3942 8832
rect 4080 8820 4108 8919
rect 4154 8916 4160 8968
rect 4212 8956 4218 8968
rect 4212 8928 4257 8956
rect 4212 8916 4218 8928
rect 4614 8916 4620 8968
rect 4672 8956 4678 8968
rect 5276 8956 5304 8996
rect 5353 8993 5365 9027
rect 5399 9024 5411 9027
rect 8294 9024 8300 9036
rect 5399 8996 8300 9024
rect 5399 8993 5411 8996
rect 5353 8987 5411 8993
rect 8294 8984 8300 8996
rect 8352 9024 8358 9036
rect 8570 9024 8576 9036
rect 8352 8996 8576 9024
rect 8352 8984 8358 8996
rect 8570 8984 8576 8996
rect 8628 8984 8634 9036
rect 4672 8928 5212 8956
rect 5276 8928 5396 8956
rect 4672 8916 4678 8928
rect 4893 8891 4951 8897
rect 4893 8857 4905 8891
rect 4939 8857 4951 8891
rect 5074 8888 5080 8900
rect 5035 8860 5080 8888
rect 4893 8851 4951 8857
rect 4614 8820 4620 8832
rect 4080 8792 4620 8820
rect 4614 8780 4620 8792
rect 4672 8780 4678 8832
rect 4908 8820 4936 8851
rect 5074 8848 5080 8860
rect 5132 8848 5138 8900
rect 5184 8888 5212 8928
rect 5261 8891 5319 8897
rect 5261 8888 5273 8891
rect 5184 8860 5273 8888
rect 5261 8857 5273 8860
rect 5307 8857 5319 8891
rect 5261 8851 5319 8857
rect 5166 8820 5172 8832
rect 4908 8792 5172 8820
rect 5166 8780 5172 8792
rect 5224 8780 5230 8832
rect 5368 8820 5396 8928
rect 7006 8916 7012 8968
rect 7064 8956 7070 8968
rect 7377 8959 7435 8965
rect 7377 8956 7389 8959
rect 7064 8928 7389 8956
rect 7064 8916 7070 8928
rect 7377 8925 7389 8928
rect 7423 8956 7435 8959
rect 7423 8928 8248 8956
rect 7423 8925 7435 8928
rect 7377 8919 7435 8925
rect 5629 8891 5687 8897
rect 5629 8857 5641 8891
rect 5675 8888 5687 8891
rect 5902 8888 5908 8900
rect 5675 8860 5908 8888
rect 5675 8857 5687 8860
rect 5629 8851 5687 8857
rect 5902 8848 5908 8860
rect 5960 8848 5966 8900
rect 8113 8891 8171 8897
rect 8113 8888 8125 8891
rect 6854 8874 8125 8888
rect 6104 8820 6132 8874
rect 6840 8860 8125 8874
rect 6840 8820 6868 8860
rect 8113 8857 8125 8860
rect 8159 8857 8171 8891
rect 8220 8888 8248 8928
rect 8386 8916 8392 8968
rect 8444 8956 8450 8968
rect 8757 8959 8815 8965
rect 8757 8956 8769 8959
rect 8444 8928 8769 8956
rect 8444 8916 8450 8928
rect 8757 8925 8769 8928
rect 8803 8925 8815 8959
rect 8757 8919 8815 8925
rect 9398 8888 9404 8900
rect 8220 8860 9404 8888
rect 8113 8851 8171 8857
rect 9398 8848 9404 8860
rect 9456 8848 9462 8900
rect 5368 8792 6868 8820
rect 7006 8780 7012 8832
rect 7064 8820 7070 8832
rect 7101 8823 7159 8829
rect 7101 8820 7113 8823
rect 7064 8792 7113 8820
rect 7064 8780 7070 8792
rect 7101 8789 7113 8792
rect 7147 8789 7159 8823
rect 7101 8783 7159 8789
rect 8294 8780 8300 8832
rect 8352 8820 8358 8832
rect 9122 8820 9128 8832
rect 8352 8792 9128 8820
rect 8352 8780 8358 8792
rect 9122 8780 9128 8792
rect 9180 8780 9186 8832
rect 920 8730 9844 8752
rect 920 8678 4116 8730
rect 4168 8678 4180 8730
rect 4232 8678 4244 8730
rect 4296 8678 4308 8730
rect 4360 8678 4372 8730
rect 4424 8678 7216 8730
rect 7268 8678 7280 8730
rect 7332 8678 7344 8730
rect 7396 8678 7408 8730
rect 7460 8678 7472 8730
rect 7524 8678 9844 8730
rect 920 8656 9844 8678
rect 1762 8576 1768 8628
rect 1820 8616 1826 8628
rect 1820 8588 9536 8616
rect 1820 8576 1826 8588
rect 1854 8508 1860 8560
rect 1912 8548 1918 8560
rect 2593 8551 2651 8557
rect 2593 8548 2605 8551
rect 1912 8520 2605 8548
rect 1912 8508 1918 8520
rect 2593 8517 2605 8520
rect 2639 8517 2651 8551
rect 4430 8548 4436 8560
rect 3818 8520 4436 8548
rect 2593 8511 2651 8517
rect 4430 8508 4436 8520
rect 4488 8548 4494 8560
rect 5074 8554 5080 8560
rect 4908 8548 5080 8554
rect 4488 8526 5080 8548
rect 4488 8520 4922 8526
rect 4488 8508 4494 8520
rect 5074 8508 5080 8526
rect 5132 8508 5138 8560
rect 6086 8508 6092 8560
rect 6144 8548 6150 8560
rect 6144 8520 7696 8548
rect 6144 8508 6150 8520
rect 1305 8483 1363 8489
rect 1305 8449 1317 8483
rect 1351 8480 1363 8483
rect 1578 8480 1584 8492
rect 1351 8452 1584 8480
rect 1351 8449 1363 8452
rect 1305 8443 1363 8449
rect 1578 8440 1584 8452
rect 1636 8440 1642 8492
rect 2222 8480 2228 8492
rect 2183 8452 2228 8480
rect 2222 8440 2228 8452
rect 2280 8440 2286 8492
rect 6181 8483 6239 8489
rect 6181 8480 6193 8483
rect 5920 8452 6193 8480
rect 5920 8424 5948 8452
rect 6181 8449 6193 8452
rect 6227 8449 6239 8483
rect 6181 8443 6239 8449
rect 6546 8440 6552 8492
rect 6604 8480 6610 8492
rect 6730 8480 6736 8492
rect 6604 8452 6736 8480
rect 6604 8440 6610 8452
rect 6730 8440 6736 8452
rect 6788 8440 6794 8492
rect 6914 8480 6920 8492
rect 6875 8452 6920 8480
rect 6914 8440 6920 8452
rect 6972 8440 6978 8492
rect 7668 8489 7696 8520
rect 8202 8508 8208 8560
rect 8260 8508 8266 8560
rect 9508 8489 9536 8588
rect 7653 8483 7711 8489
rect 7653 8449 7665 8483
rect 7699 8449 7711 8483
rect 7653 8443 7711 8449
rect 9493 8483 9551 8489
rect 9493 8449 9505 8483
rect 9539 8449 9551 8483
rect 9493 8443 9551 8449
rect 2317 8415 2375 8421
rect 2317 8381 2329 8415
rect 2363 8381 2375 8415
rect 4157 8415 4215 8421
rect 4157 8412 4169 8415
rect 2317 8375 2375 8381
rect 3620 8384 4169 8412
rect 1486 8276 1492 8288
rect 1447 8248 1492 8276
rect 1486 8236 1492 8248
rect 1544 8236 1550 8288
rect 1581 8279 1639 8285
rect 1581 8245 1593 8279
rect 1627 8276 1639 8279
rect 1762 8276 1768 8288
rect 1627 8248 1768 8276
rect 1627 8245 1639 8248
rect 1581 8239 1639 8245
rect 1762 8236 1768 8248
rect 1820 8236 1826 8288
rect 2332 8276 2360 8375
rect 3326 8276 3332 8288
rect 2332 8248 3332 8276
rect 3326 8236 3332 8248
rect 3384 8276 3390 8288
rect 3620 8276 3648 8384
rect 4157 8381 4169 8384
rect 4203 8381 4215 8415
rect 4157 8375 4215 8381
rect 4433 8415 4491 8421
rect 4433 8381 4445 8415
rect 4479 8412 4491 8415
rect 5074 8412 5080 8424
rect 4479 8384 5080 8412
rect 4479 8381 4491 8384
rect 4433 8375 4491 8381
rect 5074 8372 5080 8384
rect 5132 8372 5138 8424
rect 5902 8412 5908 8424
rect 5863 8384 5908 8412
rect 5902 8372 5908 8384
rect 5960 8372 5966 8424
rect 9122 8412 9128 8424
rect 9083 8384 9128 8412
rect 9122 8372 9128 8384
rect 9180 8372 9186 8424
rect 7193 8347 7251 8353
rect 7193 8313 7205 8347
rect 7239 8344 7251 8347
rect 7650 8344 7656 8356
rect 7239 8316 7656 8344
rect 7239 8313 7251 8316
rect 7193 8307 7251 8313
rect 7650 8304 7656 8316
rect 7708 8304 7714 8356
rect 3384 8248 3648 8276
rect 3384 8236 3390 8248
rect 3970 8236 3976 8288
rect 4028 8276 4034 8288
rect 4065 8279 4123 8285
rect 4065 8276 4077 8279
rect 4028 8248 4077 8276
rect 4028 8236 4034 8248
rect 4065 8245 4077 8248
rect 4111 8245 4123 8279
rect 4065 8239 4123 8245
rect 4522 8236 4528 8288
rect 4580 8276 4586 8288
rect 5442 8276 5448 8288
rect 4580 8248 5448 8276
rect 4580 8236 4586 8248
rect 5442 8236 5448 8248
rect 5500 8236 5506 8288
rect 5994 8236 6000 8288
rect 6052 8276 6058 8288
rect 6825 8279 6883 8285
rect 6825 8276 6837 8279
rect 6052 8248 6837 8276
rect 6052 8236 6058 8248
rect 6825 8245 6837 8248
rect 6871 8245 6883 8279
rect 6825 8239 6883 8245
rect 7006 8236 7012 8288
rect 7064 8276 7070 8288
rect 7101 8279 7159 8285
rect 7101 8276 7113 8279
rect 7064 8248 7113 8276
rect 7064 8236 7070 8248
rect 7101 8245 7113 8248
rect 7147 8245 7159 8279
rect 7101 8239 7159 8245
rect 920 8186 9844 8208
rect 920 8134 2566 8186
rect 2618 8134 2630 8186
rect 2682 8134 2694 8186
rect 2746 8134 2758 8186
rect 2810 8134 2822 8186
rect 2874 8134 5666 8186
rect 5718 8134 5730 8186
rect 5782 8134 5794 8186
rect 5846 8134 5858 8186
rect 5910 8134 5922 8186
rect 5974 8134 8766 8186
rect 8818 8134 8830 8186
rect 8882 8134 8894 8186
rect 8946 8134 8958 8186
rect 9010 8134 9022 8186
rect 9074 8134 9844 8186
rect 920 8112 9844 8134
rect 1302 8072 1308 8084
rect 1263 8044 1308 8072
rect 1302 8032 1308 8044
rect 1360 8032 1366 8084
rect 1489 8075 1547 8081
rect 1489 8041 1501 8075
rect 1535 8072 1547 8075
rect 3050 8072 3056 8084
rect 1535 8044 3056 8072
rect 1535 8041 1547 8044
rect 1489 8035 1547 8041
rect 3050 8032 3056 8044
rect 3108 8032 3114 8084
rect 3163 8075 3221 8081
rect 3163 8041 3175 8075
rect 3209 8072 3221 8075
rect 3970 8072 3976 8084
rect 3209 8044 3976 8072
rect 3209 8041 3221 8044
rect 3163 8035 3221 8041
rect 3970 8032 3976 8044
rect 4028 8032 4034 8084
rect 4062 8032 4068 8084
rect 4120 8072 4126 8084
rect 4341 8075 4399 8081
rect 4341 8072 4353 8075
rect 4120 8044 4353 8072
rect 4120 8032 4126 8044
rect 4341 8041 4353 8044
rect 4387 8041 4399 8075
rect 4522 8072 4528 8084
rect 4483 8044 4528 8072
rect 4341 8035 4399 8041
rect 4522 8032 4528 8044
rect 4580 8032 4586 8084
rect 8205 8075 8263 8081
rect 8205 8041 8217 8075
rect 8251 8072 8263 8075
rect 8386 8072 8392 8084
rect 8251 8044 8392 8072
rect 8251 8041 8263 8044
rect 8205 8035 8263 8041
rect 8386 8032 8392 8044
rect 8444 8032 8450 8084
rect 8570 8004 8576 8016
rect 8531 7976 8576 8004
rect 8570 7964 8576 7976
rect 8628 7964 8634 8016
rect 1670 7896 1676 7948
rect 1728 7936 1734 7948
rect 5169 7939 5227 7945
rect 5169 7936 5181 7939
rect 1728 7908 5181 7936
rect 1728 7896 1734 7908
rect 5169 7905 5181 7908
rect 5215 7905 5227 7939
rect 5169 7899 5227 7905
rect 5537 7939 5595 7945
rect 5537 7905 5549 7939
rect 5583 7936 5595 7939
rect 5994 7936 6000 7948
rect 5583 7908 6000 7936
rect 5583 7905 5595 7908
rect 5537 7899 5595 7905
rect 5994 7896 6000 7908
rect 6052 7896 6058 7948
rect 1302 7828 1308 7880
rect 1360 7868 1366 7880
rect 1397 7871 1455 7877
rect 1397 7868 1409 7871
rect 1360 7840 1409 7868
rect 1360 7828 1366 7840
rect 1397 7837 1409 7840
rect 1443 7837 1455 7871
rect 1397 7831 1455 7837
rect 3418 7828 3424 7880
rect 3476 7868 3482 7880
rect 3605 7871 3663 7877
rect 3476 7840 3521 7868
rect 3476 7828 3482 7840
rect 3605 7837 3617 7871
rect 3651 7837 3663 7871
rect 4338 7868 4344 7880
rect 3605 7831 3663 7837
rect 4126 7840 4344 7868
rect 2682 7760 2688 7812
rect 2740 7760 2746 7812
rect 3510 7760 3516 7812
rect 3568 7800 3574 7812
rect 3620 7800 3648 7831
rect 3568 7772 3648 7800
rect 3568 7760 3574 7772
rect 1673 7735 1731 7741
rect 1673 7701 1685 7735
rect 1719 7732 1731 7735
rect 2222 7732 2228 7744
rect 1719 7704 2228 7732
rect 1719 7701 1731 7704
rect 1673 7695 1731 7701
rect 2222 7692 2228 7704
rect 2280 7692 2286 7744
rect 3418 7692 3424 7744
rect 3476 7732 3482 7744
rect 4126 7732 4154 7840
rect 4338 7828 4344 7840
rect 4396 7828 4402 7880
rect 4801 7871 4859 7877
rect 4801 7837 4813 7871
rect 4847 7837 4859 7871
rect 4801 7831 4859 7837
rect 4249 7803 4307 7809
rect 4249 7769 4261 7803
rect 4295 7800 4307 7803
rect 4614 7800 4620 7812
rect 4295 7772 4620 7800
rect 4295 7769 4307 7772
rect 4249 7763 4307 7769
rect 4614 7760 4620 7772
rect 4672 7760 4678 7812
rect 4816 7800 4844 7831
rect 4890 7828 4896 7880
rect 4948 7868 4954 7880
rect 7006 7868 7012 7880
rect 4948 7840 4993 7868
rect 6967 7840 7012 7868
rect 4948 7828 4954 7840
rect 7006 7828 7012 7840
rect 7064 7828 7070 7880
rect 7561 7871 7619 7877
rect 7561 7837 7573 7871
rect 7607 7837 7619 7871
rect 7561 7831 7619 7837
rect 4816 7772 5212 7800
rect 5184 7744 5212 7772
rect 3476 7704 4154 7732
rect 3476 7692 3482 7704
rect 4522 7692 4528 7744
rect 4580 7732 4586 7744
rect 5077 7735 5135 7741
rect 5077 7732 5089 7735
rect 4580 7704 5089 7732
rect 4580 7692 4586 7704
rect 5077 7701 5089 7704
rect 5123 7701 5135 7735
rect 5077 7695 5135 7701
rect 5166 7692 5172 7744
rect 5224 7692 5230 7744
rect 6656 7732 6684 7786
rect 6914 7760 6920 7812
rect 6972 7800 6978 7812
rect 7576 7800 7604 7831
rect 8294 7828 8300 7880
rect 8352 7868 8358 7880
rect 8757 7871 8815 7877
rect 8757 7868 8769 7871
rect 8352 7840 8769 7868
rect 8352 7828 8358 7840
rect 8757 7837 8769 7840
rect 8803 7837 8815 7871
rect 8757 7831 8815 7837
rect 8386 7800 8392 7812
rect 6972 7772 7604 7800
rect 8347 7772 8392 7800
rect 6972 7760 6978 7772
rect 8386 7760 8392 7772
rect 8444 7760 8450 7812
rect 7006 7732 7012 7744
rect 6656 7704 7012 7732
rect 7006 7692 7012 7704
rect 7064 7692 7070 7744
rect 7469 7735 7527 7741
rect 7469 7701 7481 7735
rect 7515 7732 7527 7735
rect 8110 7732 8116 7744
rect 7515 7704 8116 7732
rect 7515 7701 7527 7704
rect 7469 7695 7527 7701
rect 8110 7692 8116 7704
rect 8168 7692 8174 7744
rect 9398 7732 9404 7744
rect 9359 7704 9404 7732
rect 9398 7692 9404 7704
rect 9456 7692 9462 7744
rect 920 7642 9844 7664
rect 920 7590 4116 7642
rect 4168 7590 4180 7642
rect 4232 7590 4244 7642
rect 4296 7590 4308 7642
rect 4360 7590 4372 7642
rect 4424 7590 7216 7642
rect 7268 7590 7280 7642
rect 7332 7590 7344 7642
rect 7396 7590 7408 7642
rect 7460 7590 7472 7642
rect 7524 7590 9844 7642
rect 920 7568 9844 7590
rect 8386 7528 8392 7540
rect 1412 7500 8392 7528
rect 1412 7469 1440 7500
rect 1397 7463 1455 7469
rect 1397 7429 1409 7463
rect 1443 7429 1455 7463
rect 1397 7423 1455 7429
rect 3234 7420 3240 7472
rect 3292 7460 3298 7472
rect 3292 7432 3358 7460
rect 3292 7420 3298 7432
rect 4706 7420 4712 7472
rect 4764 7460 4770 7472
rect 5166 7460 5172 7472
rect 4764 7432 5172 7460
rect 4764 7420 4770 7432
rect 5166 7420 5172 7432
rect 5224 7420 5230 7472
rect 6196 7469 6224 7500
rect 8386 7488 8392 7500
rect 8444 7488 8450 7540
rect 6181 7463 6239 7469
rect 6181 7429 6193 7463
rect 6227 7429 6239 7463
rect 7926 7460 7932 7472
rect 7887 7432 7932 7460
rect 6181 7423 6239 7429
rect 7926 7420 7932 7432
rect 7984 7420 7990 7472
rect 1673 7395 1731 7401
rect 1673 7361 1685 7395
rect 1719 7392 1731 7395
rect 1762 7392 1768 7404
rect 1719 7364 1768 7392
rect 1719 7361 1731 7364
rect 1673 7355 1731 7361
rect 1762 7352 1768 7364
rect 1820 7352 1826 7404
rect 2317 7395 2375 7401
rect 2317 7361 2329 7395
rect 2363 7392 2375 7395
rect 2961 7395 3019 7401
rect 2961 7392 2973 7395
rect 2363 7364 2973 7392
rect 2363 7361 2375 7364
rect 2317 7355 2375 7361
rect 2961 7361 2973 7364
rect 3007 7361 3019 7395
rect 2961 7355 3019 7361
rect 4433 7395 4491 7401
rect 4433 7361 4445 7395
rect 4479 7392 4491 7395
rect 4798 7392 4804 7404
rect 4479 7364 4804 7392
rect 4479 7361 4491 7364
rect 4433 7355 4491 7361
rect 4798 7352 4804 7364
rect 4856 7352 4862 7404
rect 4985 7395 5043 7401
rect 4985 7361 4997 7395
rect 5031 7361 5043 7395
rect 4985 7355 5043 7361
rect 5721 7395 5779 7401
rect 5721 7361 5733 7395
rect 5767 7392 5779 7395
rect 6086 7392 6092 7404
rect 5767 7364 6092 7392
rect 5767 7361 5779 7364
rect 5721 7355 5779 7361
rect 1486 7284 1492 7336
rect 1544 7324 1550 7336
rect 2593 7327 2651 7333
rect 2593 7324 2605 7327
rect 1544 7296 2605 7324
rect 1544 7284 1550 7296
rect 2593 7293 2605 7296
rect 2639 7293 2651 7327
rect 2593 7287 2651 7293
rect 4706 7284 4712 7336
rect 4764 7324 4770 7336
rect 5000 7324 5028 7355
rect 6086 7352 6092 7364
rect 6144 7352 6150 7404
rect 6822 7352 6828 7404
rect 6880 7352 6886 7404
rect 7742 7352 7748 7404
rect 7800 7392 7806 7404
rect 8021 7395 8079 7401
rect 8021 7392 8033 7395
rect 7800 7364 8033 7392
rect 7800 7352 7806 7364
rect 8021 7361 8033 7364
rect 8067 7361 8079 7395
rect 8021 7355 8079 7361
rect 9033 7395 9091 7401
rect 9033 7361 9045 7395
rect 9079 7392 9091 7395
rect 9306 7392 9312 7404
rect 9079 7364 9312 7392
rect 9079 7361 9091 7364
rect 9033 7355 9091 7361
rect 9306 7352 9312 7364
rect 9364 7352 9370 7404
rect 6840 7324 6868 7352
rect 4764 7296 5028 7324
rect 5460 7296 6868 7324
rect 4764 7284 4770 7296
rect 1302 7216 1308 7268
rect 1360 7256 1366 7268
rect 2130 7256 2136 7268
rect 1360 7228 2136 7256
rect 1360 7216 1366 7228
rect 2130 7216 2136 7228
rect 2188 7256 2194 7268
rect 2409 7259 2467 7265
rect 2409 7256 2421 7259
rect 2188 7228 2421 7256
rect 2188 7216 2194 7228
rect 2409 7225 2421 7228
rect 2455 7225 2467 7259
rect 5460 7256 5488 7296
rect 8386 7284 8392 7336
rect 8444 7324 8450 7336
rect 9125 7327 9183 7333
rect 9125 7324 9137 7327
rect 8444 7296 9137 7324
rect 8444 7284 8450 7296
rect 9125 7293 9137 7296
rect 9171 7293 9183 7327
rect 9125 7287 9183 7293
rect 9214 7284 9220 7336
rect 9272 7324 9278 7336
rect 9272 7296 9317 7324
rect 9272 7284 9278 7296
rect 9582 7284 9588 7336
rect 9640 7324 9646 7336
rect 9953 7327 10011 7333
rect 9953 7324 9965 7327
rect 9640 7296 9965 7324
rect 9640 7284 9646 7296
rect 9953 7293 9965 7296
rect 9999 7293 10011 7327
rect 9953 7287 10011 7293
rect 2409 7219 2467 7225
rect 4908 7228 5488 7256
rect 5629 7259 5687 7265
rect 1489 7191 1547 7197
rect 1489 7157 1501 7191
rect 1535 7188 1547 7191
rect 1670 7188 1676 7200
rect 1535 7160 1676 7188
rect 1535 7157 1547 7160
rect 1489 7151 1547 7157
rect 1670 7148 1676 7160
rect 1728 7148 1734 7200
rect 4338 7148 4344 7200
rect 4396 7188 4402 7200
rect 4908 7197 4936 7228
rect 5629 7225 5641 7259
rect 5675 7256 5687 7259
rect 5810 7256 5816 7268
rect 5675 7228 5816 7256
rect 5675 7225 5687 7228
rect 5629 7219 5687 7225
rect 5810 7216 5816 7228
rect 5868 7216 5874 7268
rect 5905 7259 5963 7265
rect 5905 7225 5917 7259
rect 5951 7256 5963 7259
rect 6822 7256 6828 7268
rect 5951 7228 6828 7256
rect 5951 7225 5963 7228
rect 5905 7219 5963 7225
rect 6822 7216 6828 7228
rect 6880 7216 6886 7268
rect 7098 7216 7104 7268
rect 7156 7256 7162 7268
rect 8665 7259 8723 7265
rect 8665 7256 8677 7259
rect 7156 7228 8677 7256
rect 7156 7216 7162 7228
rect 8665 7225 8677 7228
rect 8711 7225 8723 7259
rect 8665 7219 8723 7225
rect 4893 7191 4951 7197
rect 4893 7188 4905 7191
rect 4396 7160 4905 7188
rect 4396 7148 4402 7160
rect 4893 7157 4905 7160
rect 4939 7157 4951 7191
rect 4893 7151 4951 7157
rect 7282 7148 7288 7200
rect 7340 7188 7346 7200
rect 8113 7191 8171 7197
rect 8113 7188 8125 7191
rect 7340 7160 8125 7188
rect 7340 7148 7346 7160
rect 8113 7157 8125 7160
rect 8159 7157 8171 7191
rect 8113 7151 8171 7157
rect 8481 7191 8539 7197
rect 8481 7157 8493 7191
rect 8527 7188 8539 7191
rect 9582 7188 9588 7200
rect 8527 7160 9588 7188
rect 8527 7157 8539 7160
rect 8481 7151 8539 7157
rect 9582 7148 9588 7160
rect 9640 7148 9646 7200
rect 920 7098 9844 7120
rect 920 7046 2566 7098
rect 2618 7046 2630 7098
rect 2682 7046 2694 7098
rect 2746 7046 2758 7098
rect 2810 7046 2822 7098
rect 2874 7046 5666 7098
rect 5718 7046 5730 7098
rect 5782 7046 5794 7098
rect 5846 7046 5858 7098
rect 5910 7046 5922 7098
rect 5974 7046 8766 7098
rect 8818 7046 8830 7098
rect 8882 7046 8894 7098
rect 8946 7046 8958 7098
rect 9010 7046 9022 7098
rect 9074 7046 9844 7098
rect 920 7024 9844 7046
rect 934 6944 940 6996
rect 992 6984 998 6996
rect 1213 6987 1271 6993
rect 1213 6984 1225 6987
rect 992 6956 1225 6984
rect 992 6944 998 6956
rect 1213 6953 1225 6956
rect 1259 6953 1271 6987
rect 1762 6984 1768 6996
rect 1213 6947 1271 6953
rect 1412 6956 1768 6984
rect 1412 6789 1440 6956
rect 1762 6944 1768 6956
rect 1820 6984 1826 6996
rect 2406 6984 2412 6996
rect 1820 6956 2412 6984
rect 1820 6944 1826 6956
rect 2406 6944 2412 6956
rect 2464 6944 2470 6996
rect 4338 6944 4344 6996
rect 4396 6984 4402 6996
rect 6089 6987 6147 6993
rect 4396 6956 5672 6984
rect 4396 6944 4402 6956
rect 5644 6928 5672 6956
rect 6089 6953 6101 6987
rect 6135 6953 6147 6987
rect 6089 6947 6147 6953
rect 5626 6876 5632 6928
rect 5684 6876 5690 6928
rect 5810 6876 5816 6928
rect 5868 6916 5874 6928
rect 6104 6916 6132 6947
rect 6178 6944 6184 6996
rect 6236 6944 6242 6996
rect 6812 6987 6870 6993
rect 6812 6953 6824 6987
rect 6858 6984 6870 6987
rect 6914 6984 6920 6996
rect 6858 6956 6920 6984
rect 6858 6953 6870 6956
rect 6812 6947 6870 6953
rect 6914 6944 6920 6956
rect 6972 6944 6978 6996
rect 7006 6944 7012 6996
rect 7064 6984 7070 6996
rect 8294 6984 8300 6996
rect 7064 6956 7880 6984
rect 8255 6956 8300 6984
rect 7064 6944 7070 6956
rect 5868 6888 6132 6916
rect 5868 6876 5874 6888
rect 1946 6808 1952 6860
rect 2004 6848 2010 6860
rect 4522 6848 4528 6860
rect 2004 6820 4528 6848
rect 2004 6808 2010 6820
rect 4522 6808 4528 6820
rect 4580 6808 4586 6860
rect 5905 6851 5963 6857
rect 5905 6817 5917 6851
rect 5951 6848 5963 6851
rect 6086 6848 6092 6860
rect 5951 6820 6092 6848
rect 5951 6817 5963 6820
rect 5905 6811 5963 6817
rect 6086 6808 6092 6820
rect 6144 6808 6150 6860
rect 1397 6783 1455 6789
rect 1397 6749 1409 6783
rect 1443 6749 1455 6783
rect 1670 6780 1676 6792
rect 1631 6752 1676 6780
rect 1397 6743 1455 6749
rect 1670 6740 1676 6752
rect 1728 6740 1734 6792
rect 3050 6740 3056 6792
rect 3108 6740 3114 6792
rect 3602 6780 3608 6792
rect 3563 6752 3608 6780
rect 3602 6740 3608 6752
rect 3660 6740 3666 6792
rect 3970 6780 3976 6792
rect 3931 6752 3976 6780
rect 3970 6740 3976 6752
rect 4028 6740 4034 6792
rect 4982 6740 4988 6792
rect 5040 6780 5046 6792
rect 5445 6783 5503 6789
rect 5445 6780 5457 6783
rect 5040 6752 5457 6780
rect 5040 6740 5046 6752
rect 5445 6749 5457 6752
rect 5491 6749 5503 6783
rect 5445 6743 5503 6749
rect 5997 6783 6055 6789
rect 5997 6749 6009 6783
rect 6043 6780 6055 6783
rect 6043 6752 6132 6780
rect 6043 6749 6055 6752
rect 5997 6743 6055 6749
rect 6104 6724 6132 6752
rect 1949 6715 2007 6721
rect 1949 6681 1961 6715
rect 1995 6712 2007 6715
rect 2222 6712 2228 6724
rect 1995 6684 2228 6712
rect 1995 6681 2007 6684
rect 1949 6675 2007 6681
rect 2222 6672 2228 6684
rect 2280 6672 2286 6724
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6644 1639 6647
rect 2038 6644 2044 6656
rect 1627 6616 2044 6644
rect 1627 6613 1639 6616
rect 1581 6607 1639 6613
rect 2038 6604 2044 6616
rect 2096 6604 2102 6656
rect 2682 6604 2688 6656
rect 2740 6644 2746 6656
rect 3421 6647 3479 6653
rect 3421 6644 3433 6647
rect 2740 6616 3433 6644
rect 2740 6604 2746 6616
rect 3421 6613 3433 6616
rect 3467 6644 3479 6647
rect 3510 6644 3516 6656
rect 3467 6616 3516 6644
rect 3467 6613 3479 6616
rect 3421 6607 3479 6613
rect 3510 6604 3516 6616
rect 3568 6604 3574 6656
rect 3786 6604 3792 6656
rect 3844 6644 3850 6656
rect 4356 6644 4384 6698
rect 6086 6672 6092 6724
rect 6144 6672 6150 6724
rect 3844 6616 4384 6644
rect 3844 6604 3850 6616
rect 4982 6604 4988 6656
rect 5040 6644 5046 6656
rect 6196 6644 6224 6944
rect 6457 6919 6515 6925
rect 6457 6885 6469 6919
rect 6503 6916 6515 6919
rect 7852 6916 7880 6956
rect 8294 6944 8300 6956
rect 8352 6944 8358 6996
rect 8389 6919 8447 6925
rect 8389 6916 8401 6919
rect 6503 6888 6684 6916
rect 7852 6888 8401 6916
rect 6503 6885 6515 6888
rect 6457 6879 6515 6885
rect 6656 6848 6684 6888
rect 8389 6885 8401 6888
rect 8435 6885 8447 6919
rect 8389 6879 8447 6885
rect 8478 6876 8484 6928
rect 8536 6916 8542 6928
rect 15194 6916 15200 6928
rect 8536 6888 8708 6916
rect 8536 6876 8542 6888
rect 6656 6820 8616 6848
rect 8588 6789 8616 6820
rect 8680 6792 8708 6888
rect 13832 6888 15200 6916
rect 9214 6808 9220 6860
rect 9272 6848 9278 6860
rect 9309 6851 9367 6857
rect 9309 6848 9321 6851
rect 9272 6820 9321 6848
rect 9272 6808 9278 6820
rect 9309 6817 9321 6820
rect 9355 6817 9367 6851
rect 9309 6811 9367 6817
rect 9950 6808 9956 6860
rect 10008 6848 10014 6860
rect 13832 6848 13860 6888
rect 15194 6876 15200 6888
rect 15252 6876 15258 6928
rect 10008 6820 13860 6848
rect 10008 6808 10014 6820
rect 6549 6783 6607 6789
rect 6549 6749 6561 6783
rect 6595 6749 6607 6783
rect 6549 6743 6607 6749
rect 8573 6783 8631 6789
rect 8573 6749 8585 6783
rect 8619 6749 8631 6783
rect 8573 6743 8631 6749
rect 5040 6616 6224 6644
rect 5040 6604 5046 6616
rect 6270 6604 6276 6656
rect 6328 6644 6334 6656
rect 6564 6644 6592 6743
rect 8662 6740 8668 6792
rect 8720 6740 8726 6792
rect 6914 6672 6920 6724
rect 6972 6712 6978 6724
rect 7282 6712 7288 6724
rect 6972 6684 7288 6712
rect 6972 6672 6978 6684
rect 7282 6672 7288 6684
rect 7340 6672 7346 6724
rect 8202 6672 8208 6724
rect 8260 6712 8266 6724
rect 9125 6715 9183 6721
rect 9125 6712 9137 6715
rect 8260 6684 9137 6712
rect 8260 6672 8266 6684
rect 9125 6681 9137 6684
rect 9171 6681 9183 6715
rect 9125 6675 9183 6681
rect 6328 6616 6592 6644
rect 6328 6604 6334 6616
rect 6730 6604 6736 6656
rect 6788 6644 6794 6656
rect 8757 6647 8815 6653
rect 8757 6644 8769 6647
rect 6788 6616 8769 6644
rect 6788 6604 6794 6616
rect 8757 6613 8769 6616
rect 8803 6613 8815 6647
rect 8757 6607 8815 6613
rect 9214 6604 9220 6656
rect 9272 6644 9278 6656
rect 9272 6616 9317 6644
rect 9272 6604 9278 6616
rect 920 6554 9844 6576
rect 920 6502 4116 6554
rect 4168 6502 4180 6554
rect 4232 6502 4244 6554
rect 4296 6502 4308 6554
rect 4360 6502 4372 6554
rect 4424 6502 7216 6554
rect 7268 6502 7280 6554
rect 7332 6502 7344 6554
rect 7396 6502 7408 6554
rect 7460 6502 7472 6554
rect 7524 6502 9844 6554
rect 920 6480 9844 6502
rect 1305 6443 1363 6449
rect 1305 6409 1317 6443
rect 1351 6440 1363 6443
rect 1394 6440 1400 6452
rect 1351 6412 1400 6440
rect 1351 6409 1363 6412
rect 1305 6403 1363 6409
rect 1394 6400 1400 6412
rect 1452 6400 1458 6452
rect 1578 6440 1584 6452
rect 1539 6412 1584 6440
rect 1578 6400 1584 6412
rect 1636 6400 1642 6452
rect 2225 6443 2283 6449
rect 2225 6409 2237 6443
rect 2271 6440 2283 6443
rect 4890 6440 4896 6452
rect 2271 6412 4896 6440
rect 2271 6409 2283 6412
rect 2225 6403 2283 6409
rect 4890 6400 4896 6412
rect 4948 6400 4954 6452
rect 7098 6440 7104 6452
rect 6012 6412 7104 6440
rect 2682 6372 2688 6384
rect 2643 6344 2688 6372
rect 2682 6332 2688 6344
rect 2740 6332 2746 6384
rect 2958 6332 2964 6384
rect 3016 6372 3022 6384
rect 3016 6344 3174 6372
rect 3016 6332 3022 6344
rect 3970 6332 3976 6384
rect 4028 6372 4034 6384
rect 4028 6344 4936 6372
rect 4028 6332 4034 6344
rect 1489 6307 1547 6313
rect 1489 6273 1501 6307
rect 1535 6273 1547 6307
rect 1762 6304 1768 6316
rect 1723 6276 1768 6304
rect 1489 6267 1547 6273
rect 1504 6168 1532 6267
rect 1762 6264 1768 6276
rect 1820 6264 1826 6316
rect 1857 6307 1915 6313
rect 1857 6273 1869 6307
rect 1903 6304 1915 6307
rect 1946 6304 1952 6316
rect 1903 6276 1952 6304
rect 1903 6273 1915 6276
rect 1857 6267 1915 6273
rect 1946 6264 1952 6276
rect 2004 6264 2010 6316
rect 2130 6304 2136 6316
rect 2091 6276 2136 6304
rect 2130 6264 2136 6276
rect 2188 6264 2194 6316
rect 4249 6307 4307 6313
rect 4249 6273 4261 6307
rect 4295 6304 4307 6307
rect 4614 6304 4620 6316
rect 4295 6276 4620 6304
rect 4295 6273 4307 6276
rect 4249 6267 4307 6273
rect 4614 6264 4620 6276
rect 4672 6264 4678 6316
rect 4908 6313 4936 6344
rect 4893 6307 4951 6313
rect 4893 6273 4905 6307
rect 4939 6273 4951 6307
rect 4893 6267 4951 6273
rect 5629 6307 5687 6313
rect 5629 6273 5641 6307
rect 5675 6304 5687 6307
rect 5902 6304 5908 6316
rect 5675 6276 5908 6304
rect 5675 6273 5687 6276
rect 5629 6267 5687 6273
rect 5902 6264 5908 6276
rect 5960 6264 5966 6316
rect 6012 6313 6040 6412
rect 7098 6400 7104 6412
rect 7156 6400 7162 6452
rect 7834 6400 7840 6452
rect 7892 6440 7898 6452
rect 8202 6440 8208 6452
rect 7892 6412 8208 6440
rect 7892 6400 7898 6412
rect 8202 6400 8208 6412
rect 8260 6400 8266 6452
rect 9309 6443 9367 6449
rect 9309 6409 9321 6443
rect 9355 6409 9367 6443
rect 9309 6403 9367 6409
rect 9324 6372 9352 6403
rect 8418 6344 9352 6372
rect 5997 6307 6055 6313
rect 5997 6273 6009 6307
rect 6043 6273 6055 6307
rect 5997 6267 6055 6273
rect 6730 6264 6736 6316
rect 6788 6304 6794 6316
rect 6825 6307 6883 6313
rect 6825 6304 6837 6307
rect 6788 6276 6837 6304
rect 6788 6264 6794 6276
rect 6825 6273 6837 6276
rect 6871 6273 6883 6307
rect 8754 6304 8760 6316
rect 8715 6276 8760 6304
rect 6825 6267 6883 6273
rect 8754 6264 8760 6276
rect 8812 6264 8818 6316
rect 9493 6307 9551 6313
rect 9493 6273 9505 6307
rect 9539 6273 9551 6307
rect 9493 6267 9551 6273
rect 1670 6196 1676 6248
rect 1728 6236 1734 6248
rect 2406 6236 2412 6248
rect 1728 6208 2412 6236
rect 1728 6196 1734 6208
rect 2406 6196 2412 6208
rect 2464 6196 2470 6248
rect 3050 6196 3056 6248
rect 3108 6236 3114 6248
rect 6917 6239 6975 6245
rect 6917 6236 6929 6239
rect 3108 6208 6929 6236
rect 3108 6196 3114 6208
rect 6917 6205 6929 6208
rect 6963 6205 6975 6239
rect 7285 6239 7343 6245
rect 7285 6236 7297 6239
rect 6917 6199 6975 6205
rect 7024 6208 7297 6236
rect 5534 6168 5540 6180
rect 1504 6140 2544 6168
rect 2041 6103 2099 6109
rect 2041 6069 2053 6103
rect 2087 6100 2099 6103
rect 2130 6100 2136 6112
rect 2087 6072 2136 6100
rect 2087 6069 2099 6072
rect 2041 6063 2099 6069
rect 2130 6060 2136 6072
rect 2188 6060 2194 6112
rect 2516 6100 2544 6140
rect 3712 6140 5540 6168
rect 3712 6100 3740 6140
rect 5534 6128 5540 6140
rect 5592 6128 5598 6180
rect 5813 6171 5871 6177
rect 5813 6137 5825 6171
rect 5859 6168 5871 6171
rect 6546 6168 6552 6180
rect 5859 6140 6552 6168
rect 5859 6137 5871 6140
rect 5813 6131 5871 6137
rect 6546 6128 6552 6140
rect 6604 6128 6610 6180
rect 2516 6072 3740 6100
rect 4157 6103 4215 6109
rect 4157 6069 4169 6103
rect 4203 6100 4215 6103
rect 4706 6100 4712 6112
rect 4203 6072 4712 6100
rect 4203 6069 4215 6072
rect 4157 6063 4215 6069
rect 4706 6060 4712 6072
rect 4764 6060 4770 6112
rect 4982 6100 4988 6112
rect 4943 6072 4988 6100
rect 4982 6060 4988 6072
rect 5040 6060 5046 6112
rect 6086 6060 6092 6112
rect 6144 6100 6150 6112
rect 6181 6103 6239 6109
rect 6181 6100 6193 6103
rect 6144 6072 6193 6100
rect 6144 6060 6150 6072
rect 6181 6069 6193 6072
rect 6227 6069 6239 6103
rect 7024 6100 7052 6208
rect 7285 6205 7297 6208
rect 7331 6205 7343 6239
rect 7285 6199 7343 6205
rect 8202 6128 8208 6180
rect 8260 6168 8266 6180
rect 9508 6168 9536 6267
rect 8260 6140 9536 6168
rect 8260 6128 8266 6140
rect 8478 6100 8484 6112
rect 7024 6072 8484 6100
rect 6181 6063 6239 6069
rect 8478 6060 8484 6072
rect 8536 6060 8542 6112
rect 9217 6103 9275 6109
rect 9217 6069 9229 6103
rect 9263 6100 9275 6103
rect 9306 6100 9312 6112
rect 9263 6072 9312 6100
rect 9263 6069 9275 6072
rect 9217 6063 9275 6069
rect 9306 6060 9312 6072
rect 9364 6060 9370 6112
rect 920 6010 9844 6032
rect 920 5958 2566 6010
rect 2618 5958 2630 6010
rect 2682 5958 2694 6010
rect 2746 5958 2758 6010
rect 2810 5958 2822 6010
rect 2874 5958 5666 6010
rect 5718 5958 5730 6010
rect 5782 5958 5794 6010
rect 5846 5958 5858 6010
rect 5910 5958 5922 6010
rect 5974 5958 8766 6010
rect 8818 5958 8830 6010
rect 8882 5958 8894 6010
rect 8946 5958 8958 6010
rect 9010 5958 9022 6010
rect 9074 5958 9844 6010
rect 920 5936 9844 5958
rect 1397 5899 1455 5905
rect 1397 5865 1409 5899
rect 1443 5896 1455 5899
rect 1486 5896 1492 5908
rect 1443 5868 1492 5896
rect 1443 5865 1455 5868
rect 1397 5859 1455 5865
rect 1486 5856 1492 5868
rect 1544 5856 1550 5908
rect 1946 5896 1952 5908
rect 1907 5868 1952 5896
rect 1946 5856 1952 5868
rect 2004 5856 2010 5908
rect 2222 5896 2228 5908
rect 2183 5868 2228 5896
rect 2222 5856 2228 5868
rect 2280 5856 2286 5908
rect 2501 5899 2559 5905
rect 2501 5865 2513 5899
rect 2547 5896 2559 5899
rect 3050 5896 3056 5908
rect 2547 5868 3056 5896
rect 2547 5865 2559 5868
rect 2501 5859 2559 5865
rect 3050 5856 3056 5868
rect 3108 5856 3114 5908
rect 3786 5896 3792 5908
rect 3160 5868 3792 5896
rect 1118 5788 1124 5840
rect 1176 5828 1182 5840
rect 1762 5828 1768 5840
rect 1176 5800 1768 5828
rect 1176 5788 1182 5800
rect 1762 5788 1768 5800
rect 1820 5788 1826 5840
rect 2958 5788 2964 5840
rect 3016 5828 3022 5840
rect 3160 5828 3188 5868
rect 3786 5856 3792 5868
rect 3844 5856 3850 5908
rect 3970 5856 3976 5908
rect 4028 5896 4034 5908
rect 4982 5896 4988 5908
rect 4028 5868 4988 5896
rect 4028 5856 4034 5868
rect 4982 5856 4988 5868
rect 5040 5856 5046 5908
rect 5534 5856 5540 5908
rect 5592 5896 5598 5908
rect 6273 5899 6331 5905
rect 6273 5896 6285 5899
rect 5592 5868 6285 5896
rect 5592 5856 5598 5868
rect 6273 5865 6285 5868
rect 6319 5865 6331 5899
rect 6273 5859 6331 5865
rect 6641 5899 6699 5905
rect 6641 5865 6653 5899
rect 6687 5896 6699 5899
rect 8202 5896 8208 5908
rect 6687 5868 8208 5896
rect 6687 5865 6699 5868
rect 6641 5859 6699 5865
rect 8202 5856 8208 5868
rect 8260 5856 8266 5908
rect 8757 5899 8815 5905
rect 8757 5865 8769 5899
rect 8803 5896 8815 5899
rect 9122 5896 9128 5908
rect 8803 5868 9128 5896
rect 8803 5865 8815 5868
rect 8757 5859 8815 5865
rect 9122 5856 9128 5868
rect 9180 5856 9186 5908
rect 3016 5800 3280 5828
rect 3016 5788 3022 5800
rect 2976 5760 3004 5788
rect 1504 5732 3004 5760
rect 934 5652 940 5704
rect 992 5692 998 5704
rect 1504 5701 1532 5732
rect 1213 5695 1271 5701
rect 1213 5692 1225 5695
rect 992 5664 1225 5692
rect 992 5652 998 5664
rect 1213 5661 1225 5664
rect 1259 5661 1271 5695
rect 1213 5655 1271 5661
rect 1489 5695 1547 5701
rect 1489 5661 1501 5695
rect 1535 5661 1547 5695
rect 1489 5655 1547 5661
rect 1670 5652 1676 5704
rect 1728 5692 1734 5704
rect 1765 5695 1823 5701
rect 1765 5692 1777 5695
rect 1728 5664 1777 5692
rect 1728 5652 1734 5664
rect 1765 5661 1777 5664
rect 1811 5661 1823 5695
rect 2038 5692 2044 5704
rect 1999 5664 2044 5692
rect 1765 5655 1823 5661
rect 2038 5652 2044 5664
rect 2096 5652 2102 5704
rect 2130 5652 2136 5704
rect 2188 5692 2194 5704
rect 2792 5701 2820 5732
rect 3252 5701 3280 5800
rect 4154 5788 4160 5840
rect 4212 5788 4218 5840
rect 6822 5828 6828 5840
rect 6196 5800 6828 5828
rect 4172 5760 4200 5788
rect 3528 5732 4200 5760
rect 4525 5763 4583 5769
rect 2317 5695 2375 5701
rect 2317 5692 2329 5695
rect 2188 5664 2329 5692
rect 2188 5652 2194 5664
rect 2317 5661 2329 5664
rect 2363 5661 2375 5695
rect 2317 5655 2375 5661
rect 2777 5695 2835 5701
rect 2777 5661 2789 5695
rect 2823 5661 2835 5695
rect 2777 5655 2835 5661
rect 2866 5648 2872 5700
rect 2924 5692 2930 5700
rect 2961 5695 3019 5701
rect 2961 5692 2973 5695
rect 2924 5664 2973 5692
rect 2924 5648 2930 5664
rect 2961 5661 2973 5664
rect 3007 5661 3019 5695
rect 2961 5655 3019 5661
rect 3237 5695 3295 5701
rect 3237 5661 3249 5695
rect 3283 5661 3295 5695
rect 3237 5655 3295 5661
rect 3421 5695 3479 5701
rect 3421 5661 3433 5695
rect 3467 5692 3479 5695
rect 3528 5692 3556 5732
rect 4525 5729 4537 5763
rect 4571 5760 4583 5763
rect 6196 5760 6224 5800
rect 6822 5788 6828 5800
rect 6880 5788 6886 5840
rect 4571 5732 6224 5760
rect 4571 5729 4583 5732
rect 4525 5723 4583 5729
rect 6270 5720 6276 5772
rect 6328 5760 6334 5772
rect 8570 5760 8576 5772
rect 6328 5732 8576 5760
rect 6328 5720 6334 5732
rect 8570 5720 8576 5732
rect 8628 5720 8634 5772
rect 3467 5664 3556 5692
rect 3467 5661 3479 5664
rect 3421 5655 3479 5661
rect 3602 5652 3608 5704
rect 3660 5692 3666 5704
rect 4065 5695 4123 5701
rect 4065 5692 4077 5695
rect 3660 5664 4077 5692
rect 3660 5652 3666 5664
rect 4065 5661 4077 5664
rect 4111 5661 4123 5695
rect 4246 5692 4252 5704
rect 4207 5664 4252 5692
rect 4065 5655 4123 5661
rect 4246 5652 4252 5664
rect 4304 5652 4310 5704
rect 5902 5652 5908 5704
rect 5960 5692 5966 5704
rect 6181 5695 6239 5701
rect 6181 5692 6193 5695
rect 5960 5664 6193 5692
rect 5960 5652 5966 5664
rect 6181 5661 6193 5664
rect 6227 5692 6239 5695
rect 9398 5692 9404 5704
rect 6227 5664 6684 5692
rect 9359 5664 9404 5692
rect 6227 5661 6239 5664
rect 6181 5655 6239 5661
rect 5534 5584 5540 5636
rect 5592 5584 5598 5636
rect 5810 5584 5816 5636
rect 5868 5624 5874 5636
rect 6086 5624 6092 5636
rect 5868 5596 6092 5624
rect 5868 5584 5874 5596
rect 6086 5584 6092 5596
rect 6144 5584 6150 5636
rect 753 5559 811 5565
rect 753 5525 765 5559
rect 799 5556 811 5559
rect 1673 5559 1731 5565
rect 1673 5556 1685 5559
rect 799 5528 1685 5556
rect 799 5525 811 5528
rect 753 5519 811 5525
rect 1673 5525 1685 5528
rect 1719 5525 1731 5559
rect 1673 5519 1731 5525
rect 1762 5516 1768 5568
rect 1820 5556 1826 5568
rect 2593 5559 2651 5565
rect 2593 5556 2605 5559
rect 1820 5528 2605 5556
rect 1820 5516 1826 5528
rect 2593 5525 2605 5528
rect 2639 5525 2651 5559
rect 2593 5519 2651 5525
rect 2866 5516 2872 5568
rect 2924 5556 2930 5568
rect 3053 5559 3111 5565
rect 3053 5556 3065 5559
rect 2924 5528 3065 5556
rect 2924 5516 2930 5528
rect 3053 5525 3065 5528
rect 3099 5525 3111 5559
rect 3053 5519 3111 5525
rect 3142 5516 3148 5568
rect 3200 5556 3206 5568
rect 3605 5559 3663 5565
rect 3605 5556 3617 5559
rect 3200 5528 3617 5556
rect 3200 5516 3206 5528
rect 3605 5525 3617 5528
rect 3651 5525 3663 5559
rect 3605 5519 3663 5525
rect 5997 5559 6055 5565
rect 5997 5525 6009 5559
rect 6043 5556 6055 5559
rect 6546 5556 6552 5568
rect 6043 5528 6552 5556
rect 6043 5525 6055 5528
rect 5997 5519 6055 5525
rect 6546 5516 6552 5528
rect 6604 5516 6610 5568
rect 6656 5556 6684 5664
rect 9398 5652 9404 5664
rect 9456 5652 9462 5704
rect 7006 5584 7012 5636
rect 7064 5624 7070 5636
rect 8294 5624 8300 5636
rect 7064 5596 7130 5624
rect 8255 5596 8300 5624
rect 7064 5584 7070 5596
rect 8294 5584 8300 5596
rect 8352 5584 8358 5636
rect 8018 5556 8024 5568
rect 6656 5528 8024 5556
rect 8018 5516 8024 5528
rect 8076 5516 8082 5568
rect 920 5466 9844 5488
rect 920 5414 4116 5466
rect 4168 5414 4180 5466
rect 4232 5414 4244 5466
rect 4296 5414 4308 5466
rect 4360 5414 4372 5466
rect 4424 5414 7216 5466
rect 7268 5414 7280 5466
rect 7332 5414 7344 5466
rect 7396 5414 7408 5466
rect 7460 5414 7472 5466
rect 7524 5414 9844 5466
rect 920 5392 9844 5414
rect 1854 5312 1860 5364
rect 1912 5352 1918 5364
rect 2590 5352 2596 5364
rect 1912 5324 2596 5352
rect 1912 5312 1918 5324
rect 2590 5312 2596 5324
rect 2648 5312 2654 5364
rect 4614 5352 4620 5364
rect 3620 5324 4620 5352
rect 1210 5244 1216 5296
rect 1268 5284 1274 5296
rect 2406 5284 2412 5296
rect 1268 5256 2412 5284
rect 1268 5244 1274 5256
rect 2406 5244 2412 5256
rect 2464 5244 2470 5296
rect 3620 5293 3648 5324
rect 4614 5312 4620 5324
rect 4672 5312 4678 5364
rect 5074 5352 5080 5364
rect 5035 5324 5080 5352
rect 5074 5312 5080 5324
rect 5132 5312 5138 5364
rect 5261 5355 5319 5361
rect 5261 5321 5273 5355
rect 5307 5352 5319 5355
rect 7742 5352 7748 5364
rect 5307 5324 7748 5352
rect 5307 5321 5319 5324
rect 5261 5315 5319 5321
rect 7742 5312 7748 5324
rect 7800 5312 7806 5364
rect 7926 5312 7932 5364
rect 7984 5352 7990 5364
rect 9401 5355 9459 5361
rect 9401 5352 9413 5355
rect 7984 5324 9413 5352
rect 7984 5312 7990 5324
rect 9401 5321 9413 5324
rect 9447 5321 9459 5355
rect 9401 5315 9459 5321
rect 3605 5287 3663 5293
rect 3605 5253 3617 5287
rect 3651 5253 3663 5287
rect 8018 5284 8024 5296
rect 4830 5256 5488 5284
rect 7314 5256 8024 5284
rect 3605 5247 3663 5253
rect 3326 5216 3332 5228
rect 3287 5188 3332 5216
rect 3326 5176 3332 5188
rect 3384 5176 3390 5228
rect 5353 5219 5411 5225
rect 5353 5185 5365 5219
rect 5399 5185 5411 5219
rect 5353 5179 5411 5185
rect 5460 5216 5488 5256
rect 8018 5244 8024 5256
rect 8076 5244 8082 5296
rect 9122 5244 9128 5296
rect 9180 5284 9186 5296
rect 9306 5284 9312 5296
rect 9180 5256 9312 5284
rect 9180 5244 9186 5256
rect 9306 5244 9312 5256
rect 9364 5244 9370 5296
rect 5534 5216 5540 5228
rect 5460 5188 5540 5216
rect 2958 5108 2964 5160
rect 3016 5148 3022 5160
rect 3602 5148 3608 5160
rect 3016 5120 3608 5148
rect 3016 5108 3022 5120
rect 3602 5108 3608 5120
rect 3660 5108 3666 5160
rect 4062 5108 4068 5160
rect 4120 5148 4126 5160
rect 5368 5148 5396 5179
rect 4120 5120 5396 5148
rect 4120 5108 4126 5120
rect 3326 4972 3332 5024
rect 3384 5012 3390 5024
rect 5261 5015 5319 5021
rect 5261 5012 5273 5015
rect 3384 4984 5273 5012
rect 3384 4972 3390 4984
rect 5261 4981 5273 4984
rect 5307 4981 5319 5015
rect 5460 5012 5488 5188
rect 5534 5176 5540 5188
rect 5592 5216 5598 5228
rect 5721 5219 5779 5225
rect 5592 5188 5685 5216
rect 5592 5176 5598 5188
rect 5721 5185 5733 5219
rect 5767 5216 5779 5219
rect 5994 5216 6000 5228
rect 5767 5188 6000 5216
rect 5767 5185 5779 5188
rect 5721 5179 5779 5185
rect 5994 5176 6000 5188
rect 6052 5176 6058 5228
rect 7653 5219 7711 5225
rect 7653 5185 7665 5219
rect 7699 5216 7711 5219
rect 7742 5216 7748 5228
rect 7699 5188 7748 5216
rect 7699 5185 7711 5188
rect 7653 5179 7711 5185
rect 7742 5176 7748 5188
rect 7800 5176 7806 5228
rect 8297 5219 8355 5225
rect 8297 5216 8309 5219
rect 8128 5188 8309 5216
rect 5813 5151 5871 5157
rect 5813 5148 5825 5151
rect 5552 5120 5825 5148
rect 5552 5092 5580 5120
rect 5813 5117 5825 5120
rect 5859 5117 5871 5151
rect 5813 5111 5871 5117
rect 5902 5108 5908 5160
rect 5960 5148 5966 5160
rect 8128 5157 8156 5188
rect 8297 5185 8309 5188
rect 8343 5216 8355 5219
rect 9398 5216 9404 5228
rect 8343 5188 9404 5216
rect 8343 5185 8355 5188
rect 8297 5179 8355 5185
rect 9398 5176 9404 5188
rect 9456 5176 9462 5228
rect 6181 5151 6239 5157
rect 6181 5148 6193 5151
rect 5960 5120 6193 5148
rect 5960 5108 5966 5120
rect 6181 5117 6193 5120
rect 6227 5117 6239 5151
rect 6181 5111 6239 5117
rect 8113 5151 8171 5157
rect 8113 5117 8125 5151
rect 8159 5117 8171 5151
rect 8662 5148 8668 5160
rect 8623 5120 8668 5148
rect 8113 5111 8171 5117
rect 8662 5108 8668 5120
rect 8720 5108 8726 5160
rect 8849 5151 8907 5157
rect 8849 5117 8861 5151
rect 8895 5148 8907 5151
rect 9582 5148 9588 5160
rect 8895 5120 9588 5148
rect 8895 5117 8907 5120
rect 8849 5111 8907 5117
rect 9582 5108 9588 5120
rect 9640 5108 9646 5160
rect 5534 5040 5540 5092
rect 5592 5040 5598 5092
rect 8481 5083 8539 5089
rect 8481 5049 8493 5083
rect 8527 5080 8539 5083
rect 16574 5080 16580 5092
rect 8527 5052 16580 5080
rect 8527 5049 8539 5052
rect 8481 5043 8539 5049
rect 16574 5040 16580 5052
rect 16632 5040 16638 5092
rect 7098 5012 7104 5024
rect 5460 4984 7104 5012
rect 5261 4975 5319 4981
rect 7098 4972 7104 4984
rect 7156 4972 7162 5024
rect 9306 5012 9312 5024
rect 9267 4984 9312 5012
rect 9306 4972 9312 4984
rect 9364 4972 9370 5024
rect 2774 4944 2780 4956
rect 2735 4916 2780 4944
rect 2774 4904 2780 4916
rect 2832 4904 2838 4956
rect 3036 4922 9844 4944
rect 3036 4870 5666 4922
rect 5718 4870 5730 4922
rect 5782 4870 5794 4922
rect 5846 4870 5858 4922
rect 5910 4870 5922 4922
rect 5974 4870 8766 4922
rect 8818 4870 8830 4922
rect 8882 4870 8894 4922
rect 8946 4870 8958 4922
rect 9010 4870 9022 4922
rect 9074 4870 9844 4922
rect 3036 4848 9844 4870
rect 2774 4768 2780 4820
rect 2832 4808 2838 4820
rect 3418 4808 3424 4820
rect 2832 4780 3424 4808
rect 2832 4768 2838 4780
rect 3418 4768 3424 4780
rect 3476 4768 3482 4820
rect 3786 4808 3792 4820
rect 3747 4780 3792 4808
rect 3786 4768 3792 4780
rect 3844 4808 3850 4820
rect 4430 4808 4436 4820
rect 3844 4780 4436 4808
rect 3844 4768 3850 4780
rect 4430 4768 4436 4780
rect 4488 4768 4494 4820
rect 4540 4780 7604 4808
rect 2869 4743 2927 4749
rect 2869 4709 2881 4743
rect 2915 4740 2927 4743
rect 4540 4740 4568 4780
rect 2915 4712 4568 4740
rect 7576 4740 7604 4780
rect 8478 4768 8484 4820
rect 8536 4808 8542 4820
rect 9493 4811 9551 4817
rect 9493 4808 9505 4811
rect 8536 4780 9505 4808
rect 8536 4768 8542 4780
rect 9493 4777 9505 4780
rect 9539 4777 9551 4811
rect 9493 4771 9551 4777
rect 11054 4740 11060 4752
rect 7576 4712 11060 4740
rect 2915 4709 2927 4712
rect 2869 4703 2927 4709
rect 11054 4700 11060 4712
rect 11112 4700 11118 4752
rect 17770 4700 17776 4752
rect 17828 4740 17834 4752
rect 20622 4740 20628 4752
rect 17828 4712 20628 4740
rect 17828 4700 17834 4712
rect 20622 4700 20628 4712
rect 20680 4700 20686 4752
rect 2682 4672 2688 4684
rect 2643 4644 2688 4672
rect 2682 4632 2688 4644
rect 2740 4632 2746 4684
rect 4430 4632 4436 4684
rect 4488 4672 4494 4684
rect 6270 4672 6276 4684
rect 4488 4644 5948 4672
rect 6231 4644 6276 4672
rect 4488 4632 4494 4644
rect 3418 4604 3424 4616
rect 3379 4576 3424 4604
rect 3418 4564 3424 4576
rect 3476 4564 3482 4616
rect 3697 4607 3755 4613
rect 3697 4573 3709 4607
rect 3743 4604 3755 4607
rect 4062 4604 4068 4616
rect 3743 4576 4068 4604
rect 3743 4573 3755 4576
rect 3697 4567 3755 4573
rect 1026 4496 1032 4548
rect 1084 4536 1090 4548
rect 2682 4536 2688 4548
rect 1084 4508 2688 4536
rect 1084 4496 1090 4508
rect 2682 4496 2688 4508
rect 2740 4496 2746 4548
rect 3142 4496 3148 4548
rect 3200 4536 3206 4548
rect 3712 4536 3740 4567
rect 4062 4564 4068 4576
rect 4120 4564 4126 4616
rect 4341 4607 4399 4613
rect 4341 4573 4353 4607
rect 4387 4604 4399 4607
rect 4387 4576 5028 4604
rect 4387 4573 4399 4576
rect 4341 4567 4399 4573
rect 5000 4548 5028 4576
rect 5074 4564 5080 4616
rect 5132 4604 5138 4616
rect 5537 4607 5595 4613
rect 5537 4604 5549 4607
rect 5132 4576 5549 4604
rect 5132 4564 5138 4576
rect 5537 4573 5549 4576
rect 5583 4573 5595 4607
rect 5537 4567 5595 4573
rect 3200 4508 3740 4536
rect 3200 4496 3206 4508
rect 4706 4496 4712 4548
rect 4764 4536 4770 4548
rect 4893 4539 4951 4545
rect 4893 4536 4905 4539
rect 4764 4508 4905 4536
rect 4764 4496 4770 4508
rect 4893 4505 4905 4508
rect 4939 4505 4951 4539
rect 4893 4499 4951 4505
rect 4982 4496 4988 4548
rect 5040 4536 5046 4548
rect 5920 4545 5948 4644
rect 6270 4632 6276 4644
rect 6328 4632 6334 4684
rect 6546 4672 6552 4684
rect 6507 4644 6552 4672
rect 6546 4632 6552 4644
rect 6604 4632 6610 4684
rect 8113 4607 8171 4613
rect 8113 4604 8125 4607
rect 8036 4576 8125 4604
rect 5721 4539 5779 4545
rect 5721 4536 5733 4539
rect 5040 4508 5733 4536
rect 5040 4496 5046 4508
rect 5721 4505 5733 4508
rect 5767 4505 5779 4539
rect 5721 4499 5779 4505
rect 5905 4539 5963 4545
rect 5905 4505 5917 4539
rect 5951 4536 5963 4539
rect 6270 4536 6276 4548
rect 5951 4508 6276 4536
rect 5951 4505 5963 4508
rect 5905 4499 5963 4505
rect 6270 4496 6276 4508
rect 6328 4496 6334 4548
rect 7098 4496 7104 4548
rect 7156 4496 7162 4548
rect 3602 4468 3608 4480
rect 3563 4440 3608 4468
rect 3602 4428 3608 4440
rect 3660 4428 3666 4480
rect 3786 4428 3792 4480
rect 3844 4468 3850 4480
rect 4157 4471 4215 4477
rect 4157 4468 4169 4471
rect 3844 4440 4169 4468
rect 3844 4428 3850 4440
rect 4157 4437 4169 4440
rect 4203 4437 4215 4471
rect 4798 4468 4804 4480
rect 4759 4440 4804 4468
rect 4157 4431 4215 4437
rect 4798 4428 4804 4440
rect 4856 4428 4862 4480
rect 6086 4468 6092 4480
rect 6047 4440 6092 4468
rect 6086 4428 6092 4440
rect 6144 4428 6150 4480
rect 7834 4428 7840 4480
rect 7892 4468 7898 4480
rect 8036 4477 8064 4576
rect 8113 4573 8125 4576
rect 8159 4573 8171 4607
rect 8113 4567 8171 4573
rect 8757 4607 8815 4613
rect 8757 4573 8769 4607
rect 8803 4604 8815 4607
rect 8849 4607 8907 4613
rect 8849 4604 8861 4607
rect 8803 4576 8861 4604
rect 8803 4573 8815 4576
rect 8757 4567 8815 4573
rect 8849 4573 8861 4576
rect 8895 4573 8907 4607
rect 8849 4567 8907 4573
rect 8021 4471 8079 4477
rect 8021 4468 8033 4471
rect 7892 4440 8033 4468
rect 7892 4428 7898 4440
rect 8021 4437 8033 4440
rect 8067 4437 8079 4471
rect 8021 4431 8079 4437
rect 3036 4378 9844 4400
rect 3036 4326 4116 4378
rect 4168 4326 4180 4378
rect 4232 4326 4244 4378
rect 4296 4326 4308 4378
rect 4360 4326 4372 4378
rect 4424 4326 7216 4378
rect 7268 4326 7280 4378
rect 7332 4326 7344 4378
rect 7396 4326 7408 4378
rect 7460 4326 7472 4378
rect 7524 4326 9844 4378
rect 3036 4304 9844 4326
rect 3513 4267 3571 4273
rect 3513 4233 3525 4267
rect 3559 4264 3571 4267
rect 4982 4264 4988 4276
rect 3559 4236 4988 4264
rect 3559 4233 3571 4236
rect 3513 4227 3571 4233
rect 4982 4224 4988 4236
rect 5040 4224 5046 4276
rect 9490 4224 9496 4276
rect 9548 4224 9554 4276
rect 4338 4156 4344 4208
rect 4396 4156 4402 4208
rect 8202 4156 8208 4208
rect 8260 4196 8266 4208
rect 9033 4199 9091 4205
rect 9033 4196 9045 4199
rect 8260 4168 9045 4196
rect 8260 4156 8266 4168
rect 9033 4165 9045 4168
rect 9079 4165 9091 4199
rect 9033 4159 9091 4165
rect 3329 4131 3387 4137
rect 3329 4097 3341 4131
rect 3375 4097 3387 4131
rect 3602 4128 3608 4140
rect 3563 4100 3608 4128
rect 3329 4091 3387 4097
rect 3344 4060 3372 4091
rect 3602 4088 3608 4100
rect 3660 4088 3666 4140
rect 3970 4128 3976 4140
rect 3931 4100 3976 4128
rect 3970 4088 3976 4100
rect 4028 4088 4034 4140
rect 4982 4088 4988 4140
rect 5040 4128 5046 4140
rect 5445 4131 5503 4137
rect 5445 4128 5457 4131
rect 5040 4100 5457 4128
rect 5040 4088 5046 4100
rect 5445 4097 5457 4100
rect 5491 4097 5503 4131
rect 5445 4091 5503 4097
rect 6089 4131 6147 4137
rect 6089 4097 6101 4131
rect 6135 4128 6147 4131
rect 6546 4128 6552 4140
rect 6135 4100 6552 4128
rect 6135 4097 6147 4100
rect 6089 4091 6147 4097
rect 6546 4088 6552 4100
rect 6604 4088 6610 4140
rect 6822 4128 6828 4140
rect 6783 4100 6828 4128
rect 6822 4088 6828 4100
rect 6880 4088 6886 4140
rect 6914 4088 6920 4140
rect 6972 4128 6978 4140
rect 8113 4131 8171 4137
rect 8113 4128 8125 4131
rect 6972 4100 8125 4128
rect 6972 4088 6978 4100
rect 8113 4097 8125 4100
rect 8159 4097 8171 4131
rect 8570 4128 8576 4140
rect 8531 4100 8576 4128
rect 8113 4091 8171 4097
rect 8570 4088 8576 4100
rect 8628 4088 8634 4140
rect 9508 4128 9536 4224
rect 8864 4100 9536 4128
rect 3694 4060 3700 4072
rect 3344 4032 3700 4060
rect 3694 4020 3700 4032
rect 3752 4020 3758 4072
rect 5994 4060 6000 4072
rect 5828 4032 6000 4060
rect 3602 3884 3608 3936
rect 3660 3924 3666 3936
rect 5828 3924 5856 4032
rect 5994 4020 6000 4032
rect 6052 4020 6058 4072
rect 7098 4020 7104 4072
rect 7156 4060 7162 4072
rect 7561 4063 7619 4069
rect 7561 4060 7573 4063
rect 7156 4032 7573 4060
rect 7156 4020 7162 4032
rect 7561 4029 7573 4032
rect 7607 4029 7619 4063
rect 7561 4023 7619 4029
rect 7650 4020 7656 4072
rect 7708 4060 7714 4072
rect 7708 4032 7753 4060
rect 7708 4020 7714 4032
rect 8294 4020 8300 4072
rect 8352 4060 8358 4072
rect 8864 4069 8892 4100
rect 8849 4063 8907 4069
rect 8849 4060 8861 4063
rect 8352 4032 8861 4060
rect 8352 4020 8358 4032
rect 8849 4029 8861 4032
rect 8895 4029 8907 4063
rect 8849 4023 8907 4029
rect 8941 4063 8999 4069
rect 8941 4029 8953 4063
rect 8987 4060 8999 4063
rect 9398 4060 9404 4072
rect 8987 4032 9404 4060
rect 8987 4029 8999 4032
rect 8941 4023 8999 4029
rect 9398 4020 9404 4032
rect 9456 4020 9462 4072
rect 6270 3952 6276 4004
rect 6328 3992 6334 4004
rect 7190 3992 7196 4004
rect 6328 3964 7196 3992
rect 6328 3952 6334 3964
rect 7190 3952 7196 3964
rect 7248 3992 7254 4004
rect 8389 3995 8447 4001
rect 7248 3964 7696 3992
rect 7248 3952 7254 3964
rect 7668 3936 7696 3964
rect 8389 3961 8401 3995
rect 8435 3992 8447 3995
rect 8435 3964 16574 3992
rect 8435 3961 8447 3964
rect 8389 3955 8447 3961
rect 3660 3896 5856 3924
rect 5905 3927 5963 3933
rect 3660 3884 3666 3896
rect 5905 3893 5917 3927
rect 5951 3924 5963 3927
rect 6546 3924 6552 3936
rect 5951 3896 6552 3924
rect 5951 3893 5963 3896
rect 5905 3887 5963 3893
rect 6546 3884 6552 3896
rect 6604 3884 6610 3936
rect 6730 3924 6736 3936
rect 6691 3896 6736 3924
rect 6730 3884 6736 3896
rect 6788 3884 6794 3936
rect 6914 3884 6920 3936
rect 6972 3924 6978 3936
rect 7469 3927 7527 3933
rect 7469 3924 7481 3927
rect 6972 3896 7481 3924
rect 6972 3884 6978 3896
rect 7469 3893 7481 3896
rect 7515 3893 7527 3927
rect 7469 3887 7527 3893
rect 7650 3884 7656 3936
rect 7708 3884 7714 3936
rect 9214 3884 9220 3936
rect 9272 3924 9278 3936
rect 9401 3927 9459 3933
rect 9401 3924 9413 3927
rect 9272 3896 9413 3924
rect 9272 3884 9278 3896
rect 9401 3893 9413 3896
rect 9447 3893 9459 3927
rect 9401 3887 9459 3893
rect 3036 3834 9844 3856
rect 3036 3782 5666 3834
rect 5718 3782 5730 3834
rect 5782 3782 5794 3834
rect 5846 3782 5858 3834
rect 5910 3782 5922 3834
rect 5974 3782 8766 3834
rect 8818 3782 8830 3834
rect 8882 3782 8894 3834
rect 8946 3782 8958 3834
rect 9010 3782 9022 3834
rect 9074 3782 9844 3834
rect 3036 3760 9844 3782
rect 16546 3732 16574 3964
rect 3418 3680 3424 3732
rect 3476 3720 3482 3732
rect 4065 3723 4123 3729
rect 4065 3720 4077 3723
rect 3476 3692 4077 3720
rect 3476 3680 3482 3692
rect 4065 3689 4077 3692
rect 4111 3689 4123 3723
rect 4065 3683 4123 3689
rect 4338 3680 4344 3732
rect 4396 3720 4402 3732
rect 4525 3723 4583 3729
rect 4525 3720 4537 3723
rect 4396 3692 4537 3720
rect 4396 3680 4402 3692
rect 4525 3689 4537 3692
rect 4571 3689 4583 3723
rect 5166 3720 5172 3732
rect 5127 3692 5172 3720
rect 4525 3683 4583 3689
rect 5166 3680 5172 3692
rect 5224 3680 5230 3732
rect 5353 3723 5411 3729
rect 5353 3689 5365 3723
rect 5399 3720 5411 3723
rect 6270 3720 6276 3732
rect 5399 3692 6132 3720
rect 6231 3692 6276 3720
rect 5399 3689 5411 3692
rect 5353 3683 5411 3689
rect 3513 3655 3571 3661
rect 3513 3621 3525 3655
rect 3559 3652 3571 3655
rect 3602 3652 3608 3664
rect 3559 3624 3608 3652
rect 3559 3621 3571 3624
rect 3513 3615 3571 3621
rect 3602 3612 3608 3624
rect 3660 3612 3666 3664
rect 3694 3612 3700 3664
rect 3752 3652 3758 3664
rect 3881 3655 3939 3661
rect 3881 3652 3893 3655
rect 3752 3624 3893 3652
rect 3752 3612 3758 3624
rect 3881 3621 3893 3624
rect 3927 3621 3939 3655
rect 5994 3652 6000 3664
rect 3881 3615 3939 3621
rect 5092 3624 6000 3652
rect 3786 3544 3792 3596
rect 3844 3584 3850 3596
rect 4522 3584 4528 3596
rect 3844 3556 4200 3584
rect 3844 3544 3850 3556
rect 3329 3519 3387 3525
rect 3329 3485 3341 3519
rect 3375 3516 3387 3519
rect 3418 3516 3424 3528
rect 3375 3488 3424 3516
rect 3375 3485 3387 3488
rect 3329 3479 3387 3485
rect 3418 3476 3424 3488
rect 3476 3476 3482 3528
rect 3605 3519 3663 3525
rect 3605 3485 3617 3519
rect 3651 3516 3663 3519
rect 3970 3516 3976 3528
rect 3651 3488 3976 3516
rect 3651 3485 3663 3488
rect 3605 3479 3663 3485
rect 3970 3476 3976 3488
rect 4028 3476 4034 3528
rect 4172 3448 4200 3556
rect 4264 3556 4528 3584
rect 4264 3525 4292 3556
rect 4522 3544 4528 3556
rect 4580 3544 4586 3596
rect 5092 3584 5120 3624
rect 5994 3612 6000 3624
rect 6052 3612 6058 3664
rect 6104 3652 6132 3692
rect 6270 3680 6276 3692
rect 6328 3680 6334 3732
rect 6546 3680 6552 3732
rect 6604 3720 6610 3732
rect 8294 3720 8300 3732
rect 6604 3692 8300 3720
rect 6604 3680 6610 3692
rect 8294 3680 8300 3692
rect 8352 3680 8358 3732
rect 8570 3680 8576 3732
rect 8628 3720 8634 3732
rect 8849 3723 8907 3729
rect 8849 3720 8861 3723
rect 8628 3692 8861 3720
rect 8628 3680 8634 3692
rect 8849 3689 8861 3692
rect 8895 3689 8907 3723
rect 9214 3720 9220 3732
rect 9175 3692 9220 3720
rect 8849 3683 8907 3689
rect 9214 3680 9220 3692
rect 9272 3680 9278 3732
rect 16546 3692 16580 3732
rect 16574 3680 16580 3692
rect 16632 3680 16638 3732
rect 6104 3624 6684 3652
rect 6086 3584 6092 3596
rect 4724 3556 5120 3584
rect 5736 3556 6092 3584
rect 4724 3525 4752 3556
rect 4249 3519 4307 3525
rect 4249 3485 4261 3519
rect 4295 3485 4307 3519
rect 4249 3479 4307 3485
rect 4341 3519 4399 3525
rect 4341 3485 4353 3519
rect 4387 3485 4399 3519
rect 4341 3479 4399 3485
rect 4709 3519 4767 3525
rect 4709 3485 4721 3519
rect 4755 3485 4767 3519
rect 4709 3479 4767 3485
rect 4356 3448 4384 3479
rect 4798 3476 4804 3528
rect 4856 3516 4862 3528
rect 4985 3519 5043 3525
rect 4985 3516 4997 3519
rect 4856 3488 4997 3516
rect 4856 3476 4862 3488
rect 4985 3485 4997 3488
rect 5031 3485 5043 3519
rect 4985 3479 5043 3485
rect 5537 3519 5595 3525
rect 5537 3485 5549 3519
rect 5583 3516 5595 3519
rect 5626 3516 5632 3528
rect 5583 3488 5632 3516
rect 5583 3485 5595 3488
rect 5537 3479 5595 3485
rect 5626 3476 5632 3488
rect 5684 3476 5690 3528
rect 5736 3525 5764 3556
rect 6086 3544 6092 3556
rect 6144 3544 6150 3596
rect 5721 3519 5779 3525
rect 5721 3485 5733 3519
rect 5767 3485 5779 3519
rect 5721 3479 5779 3485
rect 5997 3519 6055 3525
rect 5997 3485 6009 3519
rect 6043 3516 6055 3519
rect 6270 3516 6276 3528
rect 6043 3488 6276 3516
rect 6043 3485 6055 3488
rect 5997 3479 6055 3485
rect 6270 3476 6276 3488
rect 6328 3476 6334 3528
rect 6546 3516 6552 3528
rect 6507 3488 6552 3516
rect 6546 3476 6552 3488
rect 6604 3476 6610 3528
rect 6656 3516 6684 3624
rect 8386 3612 8392 3664
rect 8444 3652 8450 3664
rect 9398 3652 9404 3664
rect 8444 3624 8524 3652
rect 8444 3612 8450 3624
rect 6914 3584 6920 3596
rect 6875 3556 6920 3584
rect 6914 3544 6920 3556
rect 6972 3544 6978 3596
rect 7374 3584 7380 3596
rect 7024 3556 7380 3584
rect 7024 3516 7052 3556
rect 7374 3544 7380 3556
rect 7432 3544 7438 3596
rect 8386 3516 8392 3528
rect 6656 3488 7052 3516
rect 8347 3488 8392 3516
rect 8386 3476 8392 3488
rect 8444 3476 8450 3528
rect 8496 3516 8524 3624
rect 8588 3624 9404 3652
rect 8588 3596 8616 3624
rect 9398 3612 9404 3624
rect 9456 3612 9462 3664
rect 8570 3544 8576 3596
rect 8628 3544 8634 3596
rect 8846 3544 8852 3596
rect 8904 3584 8910 3596
rect 9950 3584 9956 3596
rect 8904 3556 9956 3584
rect 8904 3544 8910 3556
rect 9950 3544 9956 3556
rect 10008 3544 10014 3596
rect 8754 3516 8760 3528
rect 8496 3488 8760 3516
rect 8754 3476 8760 3488
rect 8812 3476 8818 3528
rect 8941 3519 8999 3525
rect 8941 3485 8953 3519
rect 8987 3516 8999 3519
rect 9861 3519 9919 3525
rect 9861 3516 9873 3519
rect 8987 3488 9873 3516
rect 8987 3485 8999 3488
rect 8941 3479 8999 3485
rect 9861 3485 9873 3488
rect 9907 3485 9919 3519
rect 9861 3479 9919 3485
rect 4172 3420 4384 3448
rect 4614 3408 4620 3460
rect 4672 3408 4678 3460
rect 13814 3448 13820 3460
rect 8496 3442 13820 3448
rect 3510 3340 3516 3392
rect 3568 3380 3574 3392
rect 3694 3380 3700 3392
rect 3568 3352 3700 3380
rect 3568 3340 3574 3352
rect 3694 3340 3700 3352
rect 3752 3340 3758 3392
rect 3789 3383 3847 3389
rect 3789 3349 3801 3383
rect 3835 3380 3847 3383
rect 4632 3380 4660 3408
rect 3835 3352 4660 3380
rect 4893 3383 4951 3389
rect 3835 3349 3847 3352
rect 3789 3343 3847 3349
rect 4893 3349 4905 3383
rect 4939 3380 4951 3383
rect 4982 3380 4988 3392
rect 4939 3352 4988 3380
rect 4939 3349 4951 3352
rect 4893 3343 4951 3349
rect 4982 3340 4988 3352
rect 5040 3340 5046 3392
rect 5905 3383 5963 3389
rect 5905 3349 5917 3383
rect 5951 3380 5963 3383
rect 5994 3380 6000 3392
rect 5951 3352 6000 3380
rect 5951 3349 5963 3352
rect 5905 3343 5963 3349
rect 5994 3340 6000 3352
rect 6052 3340 6058 3392
rect 6457 3383 6515 3389
rect 6457 3349 6469 3383
rect 6503 3380 6515 3383
rect 6730 3380 6736 3392
rect 6503 3352 6736 3380
rect 6503 3349 6515 3352
rect 6457 3343 6515 3349
rect 6730 3340 6736 3352
rect 6788 3340 6794 3392
rect 6914 3340 6920 3392
rect 6972 3380 6978 3392
rect 7300 3380 7328 3434
rect 8404 3420 13820 3442
rect 8404 3414 8524 3420
rect 6972 3352 7328 3380
rect 6972 3340 6978 3352
rect 7926 3340 7932 3392
rect 7984 3380 7990 3392
rect 8404 3380 8432 3414
rect 13814 3408 13820 3420
rect 13872 3408 13878 3460
rect 7984 3352 8432 3380
rect 8573 3383 8631 3389
rect 7984 3340 7990 3352
rect 8573 3349 8585 3383
rect 8619 3380 8631 3383
rect 9030 3380 9036 3392
rect 8619 3352 9036 3380
rect 8619 3349 8631 3352
rect 8573 3343 8631 3349
rect 9030 3340 9036 3352
rect 9088 3340 9094 3392
rect 9401 3383 9459 3389
rect 9401 3349 9413 3383
rect 9447 3380 9459 3383
rect 9490 3380 9496 3392
rect 9447 3352 9496 3380
rect 9447 3349 9459 3352
rect 9401 3343 9459 3349
rect 9490 3340 9496 3352
rect 9548 3340 9554 3392
rect 3036 3290 9844 3312
rect 3036 3238 4116 3290
rect 4168 3238 4180 3290
rect 4232 3238 4244 3290
rect 4296 3238 4308 3290
rect 4360 3238 4372 3290
rect 4424 3238 7216 3290
rect 7268 3238 7280 3290
rect 7332 3238 7344 3290
rect 7396 3238 7408 3290
rect 7460 3238 7472 3290
rect 7524 3238 9844 3290
rect 3036 3216 9844 3238
rect 3326 3136 3332 3188
rect 3384 3176 3390 3188
rect 3789 3179 3847 3185
rect 3789 3176 3801 3179
rect 3384 3148 3801 3176
rect 3384 3136 3390 3148
rect 3789 3145 3801 3148
rect 3835 3145 3847 3179
rect 3789 3139 3847 3145
rect 3878 3136 3884 3188
rect 3936 3176 3942 3188
rect 4065 3179 4123 3185
rect 4065 3176 4077 3179
rect 3936 3148 4077 3176
rect 3936 3136 3942 3148
rect 4065 3145 4077 3148
rect 4111 3145 4123 3179
rect 4065 3139 4123 3145
rect 4249 3179 4307 3185
rect 4249 3145 4261 3179
rect 4295 3176 4307 3179
rect 4614 3176 4620 3188
rect 4295 3148 4620 3176
rect 4295 3145 4307 3148
rect 4249 3139 4307 3145
rect 3418 3068 3424 3120
rect 3476 3108 3482 3120
rect 4264 3108 4292 3139
rect 4614 3136 4620 3148
rect 4672 3136 4678 3188
rect 6822 3176 6828 3188
rect 6783 3148 6828 3176
rect 6822 3136 6828 3148
rect 6880 3136 6886 3188
rect 8202 3136 8208 3188
rect 8260 3136 8266 3188
rect 8570 3136 8576 3188
rect 8628 3176 8634 3188
rect 8665 3179 8723 3185
rect 8665 3176 8677 3179
rect 8628 3148 8677 3176
rect 8628 3136 8634 3148
rect 8665 3145 8677 3148
rect 8711 3145 8723 3179
rect 9030 3176 9036 3188
rect 8991 3148 9036 3176
rect 8665 3139 8723 3145
rect 9030 3136 9036 3148
rect 9088 3136 9094 3188
rect 3476 3080 4292 3108
rect 3476 3068 3482 3080
rect 5166 3068 5172 3120
rect 5224 3068 5230 3120
rect 6086 3068 6092 3120
rect 6144 3108 6150 3120
rect 6270 3108 6276 3120
rect 6144 3080 6276 3108
rect 6144 3068 6150 3080
rect 6270 3068 6276 3080
rect 6328 3108 6334 3120
rect 7561 3111 7619 3117
rect 7561 3108 7573 3111
rect 6328 3080 7573 3108
rect 6328 3068 6334 3080
rect 7561 3077 7573 3080
rect 7607 3077 7619 3111
rect 7561 3071 7619 3077
rect 7650 3068 7656 3120
rect 7708 3108 7714 3120
rect 7745 3111 7803 3117
rect 7745 3108 7757 3111
rect 7708 3080 7757 3108
rect 7708 3068 7714 3080
rect 7745 3077 7757 3080
rect 7791 3077 7803 3111
rect 8220 3108 8248 3136
rect 9125 3111 9183 3117
rect 9125 3108 9137 3111
rect 8220 3080 9137 3108
rect 7745 3071 7803 3077
rect 9125 3077 9137 3080
rect 9171 3077 9183 3111
rect 9125 3071 9183 3077
rect 9214 3068 9220 3120
rect 9272 3108 9278 3120
rect 9272 3080 9674 3108
rect 9272 3068 9278 3080
rect 9646 3052 9674 3080
rect 2961 3043 3019 3049
rect 2961 3009 2973 3043
rect 3007 3040 3019 3043
rect 3329 3043 3387 3049
rect 3329 3040 3341 3043
rect 3007 3012 3341 3040
rect 3007 3009 3019 3012
rect 2961 3003 3019 3009
rect 3329 3009 3341 3012
rect 3375 3009 3387 3043
rect 3329 3003 3387 3009
rect 3605 3043 3663 3049
rect 3605 3009 3617 3043
rect 3651 3009 3663 3043
rect 3605 3003 3663 3009
rect 3881 3043 3939 3049
rect 3881 3009 3893 3043
rect 3927 3009 3939 3043
rect 3881 3003 3939 3009
rect 4341 3043 4399 3049
rect 4341 3009 4353 3043
rect 4387 3040 4399 3043
rect 4522 3040 4528 3052
rect 4387 3012 4528 3040
rect 4387 3009 4399 3012
rect 4341 3003 4399 3009
rect 2774 2864 2780 2916
rect 2832 2904 2838 2916
rect 3513 2907 3571 2913
rect 3513 2904 3525 2907
rect 2832 2876 3525 2904
rect 2832 2864 2838 2876
rect 3513 2873 3525 2876
rect 3559 2873 3571 2907
rect 3513 2867 3571 2873
rect 2869 2839 2927 2845
rect 2869 2805 2881 2839
rect 2915 2836 2927 2839
rect 3620 2836 3648 3003
rect 3896 2972 3924 3003
rect 4522 3000 4528 3012
rect 4580 3000 4586 3052
rect 4706 3040 4712 3052
rect 4667 3012 4712 3040
rect 4706 3000 4712 3012
rect 4764 3000 4770 3052
rect 5994 3000 6000 3052
rect 6052 3040 6058 3052
rect 6181 3043 6239 3049
rect 6181 3040 6193 3043
rect 6052 3012 6193 3040
rect 6052 3000 6058 3012
rect 6181 3009 6193 3012
rect 6227 3009 6239 3043
rect 6181 3003 6239 3009
rect 7006 3000 7012 3052
rect 7064 3040 7070 3052
rect 7469 3043 7527 3049
rect 7469 3040 7481 3043
rect 7064 3012 7481 3040
rect 7064 3000 7070 3012
rect 7469 3009 7481 3012
rect 7515 3009 7527 3043
rect 7469 3003 7527 3009
rect 8110 3000 8116 3052
rect 8168 3040 8174 3052
rect 8297 3043 8355 3049
rect 8297 3040 8309 3043
rect 8168 3012 8309 3040
rect 8168 3000 8174 3012
rect 8297 3009 8309 3012
rect 8343 3009 8355 3043
rect 8846 3040 8852 3052
rect 8297 3003 8355 3009
rect 8404 3012 8852 3040
rect 4890 2972 4896 2984
rect 3896 2944 4896 2972
rect 4890 2932 4896 2944
rect 4948 2932 4954 2984
rect 6270 2932 6276 2984
rect 6328 2972 6334 2984
rect 8404 2972 8432 3012
rect 8846 3000 8852 3012
rect 8904 3000 8910 3052
rect 9646 3012 9680 3052
rect 9674 3000 9680 3012
rect 9732 3000 9738 3052
rect 6328 2944 8432 2972
rect 8864 2944 9168 2972
rect 6328 2932 6334 2944
rect 8481 2907 8539 2913
rect 8481 2873 8493 2907
rect 8527 2904 8539 2907
rect 8864 2904 8892 2944
rect 8527 2876 8892 2904
rect 8527 2873 8539 2876
rect 8481 2867 8539 2873
rect 3878 2836 3884 2848
rect 2915 2808 3884 2836
rect 2915 2805 2927 2808
rect 2869 2799 2927 2805
rect 3878 2796 3884 2808
rect 3936 2796 3942 2848
rect 4062 2796 4068 2848
rect 4120 2836 4126 2848
rect 5258 2836 5264 2848
rect 4120 2808 5264 2836
rect 4120 2796 4126 2808
rect 5258 2796 5264 2808
rect 5316 2796 5322 2848
rect 6641 2839 6699 2845
rect 6641 2805 6653 2839
rect 6687 2836 6699 2839
rect 7650 2836 7656 2848
rect 6687 2808 7656 2836
rect 6687 2805 6699 2808
rect 6641 2799 6699 2805
rect 7650 2796 7656 2808
rect 7708 2796 7714 2848
rect 7929 2839 7987 2845
rect 7929 2805 7941 2839
rect 7975 2836 7987 2839
rect 8202 2836 8208 2848
rect 7975 2808 8208 2836
rect 7975 2805 7987 2808
rect 7929 2799 7987 2805
rect 8202 2796 8208 2808
rect 8260 2796 8266 2848
rect 9140 2836 9168 2944
rect 9214 2932 9220 2984
rect 9272 2972 9278 2984
rect 9272 2944 9317 2972
rect 9272 2932 9278 2944
rect 16574 2836 16580 2848
rect 9140 2808 16580 2836
rect 16574 2796 16580 2808
rect 16632 2796 16638 2848
rect 3036 2746 9844 2768
rect 3036 2694 5666 2746
rect 5718 2694 5730 2746
rect 5782 2694 5794 2746
rect 5846 2694 5858 2746
rect 5910 2694 5922 2746
rect 5974 2694 8766 2746
rect 8818 2694 8830 2746
rect 8882 2694 8894 2746
rect 8946 2694 8958 2746
rect 9010 2694 9022 2746
rect 9074 2694 9844 2746
rect 3036 2672 9844 2694
rect 2682 2592 2688 2644
rect 2740 2632 2746 2644
rect 3418 2632 3424 2644
rect 2740 2604 3424 2632
rect 2740 2592 2746 2604
rect 3418 2592 3424 2604
rect 3476 2592 3482 2644
rect 3513 2635 3571 2641
rect 3513 2601 3525 2635
rect 3559 2632 3571 2635
rect 3694 2632 3700 2644
rect 3559 2604 3700 2632
rect 3559 2601 3571 2604
rect 3513 2595 3571 2601
rect 3694 2592 3700 2604
rect 3752 2592 3758 2644
rect 3970 2592 3976 2644
rect 4028 2632 4034 2644
rect 4157 2635 4215 2641
rect 4157 2632 4169 2635
rect 4028 2604 4169 2632
rect 4028 2592 4034 2604
rect 4157 2601 4169 2604
rect 4203 2601 4215 2635
rect 4157 2595 4215 2601
rect 5445 2635 5503 2641
rect 5445 2601 5457 2635
rect 5491 2632 5503 2635
rect 5534 2632 5540 2644
rect 5491 2604 5540 2632
rect 5491 2601 5503 2604
rect 5445 2595 5503 2601
rect 5534 2592 5540 2604
rect 5592 2592 5598 2644
rect 6086 2632 6092 2644
rect 5644 2604 6092 2632
rect 3234 2524 3240 2576
rect 3292 2564 3298 2576
rect 3605 2567 3663 2573
rect 3605 2564 3617 2567
rect 3292 2536 3617 2564
rect 3292 2524 3298 2536
rect 3605 2533 3617 2536
rect 3651 2533 3663 2567
rect 4062 2564 4068 2576
rect 4023 2536 4068 2564
rect 3605 2527 3663 2533
rect 4062 2524 4068 2536
rect 4120 2524 4126 2576
rect 4522 2524 4528 2576
rect 4580 2524 4586 2576
rect 5077 2567 5135 2573
rect 5077 2533 5089 2567
rect 5123 2564 5135 2567
rect 5644 2564 5672 2604
rect 6086 2592 6092 2604
rect 6144 2592 6150 2644
rect 6457 2635 6515 2641
rect 6457 2601 6469 2635
rect 6503 2632 6515 2635
rect 6546 2632 6552 2644
rect 6503 2604 6552 2632
rect 6503 2601 6515 2604
rect 6457 2595 6515 2601
rect 6546 2592 6552 2604
rect 6604 2592 6610 2644
rect 6914 2632 6920 2644
rect 6875 2604 6920 2632
rect 6914 2592 6920 2604
rect 6972 2592 6978 2644
rect 7098 2632 7104 2644
rect 7059 2604 7104 2632
rect 7098 2592 7104 2604
rect 7156 2592 7162 2644
rect 7926 2592 7932 2644
rect 7984 2632 7990 2644
rect 8113 2635 8171 2641
rect 8113 2632 8125 2635
rect 7984 2604 8125 2632
rect 7984 2592 7990 2604
rect 8113 2601 8125 2604
rect 8159 2601 8171 2635
rect 8113 2595 8171 2601
rect 9033 2635 9091 2641
rect 9033 2601 9045 2635
rect 9079 2632 9091 2635
rect 9079 2604 9260 2632
rect 9079 2601 9091 2604
rect 9033 2595 9091 2601
rect 5123 2536 5672 2564
rect 5721 2567 5779 2573
rect 5123 2533 5135 2536
rect 5077 2527 5135 2533
rect 5721 2533 5733 2567
rect 5767 2533 5779 2567
rect 5721 2527 5779 2533
rect 7469 2567 7527 2573
rect 7469 2533 7481 2567
rect 7515 2564 7527 2567
rect 7742 2564 7748 2576
rect 7515 2536 7748 2564
rect 7515 2533 7527 2536
rect 7469 2527 7527 2533
rect 2682 2456 2688 2508
rect 2740 2496 2746 2508
rect 4540 2496 4568 2524
rect 5537 2499 5595 2505
rect 5537 2496 5549 2499
rect 2740 2468 3924 2496
rect 4540 2468 5549 2496
rect 2740 2456 2746 2468
rect 3326 2428 3332 2440
rect 3287 2400 3332 2428
rect 3326 2388 3332 2400
rect 3384 2388 3390 2440
rect 3418 2388 3424 2440
rect 3476 2428 3482 2440
rect 3786 2428 3792 2440
rect 3476 2400 3792 2428
rect 3476 2388 3482 2400
rect 3786 2388 3792 2400
rect 3844 2388 3850 2440
rect 3896 2437 3924 2468
rect 5537 2465 5549 2468
rect 5583 2465 5595 2499
rect 5537 2459 5595 2465
rect 3881 2431 3939 2437
rect 3881 2397 3893 2431
rect 3927 2428 3939 2431
rect 3970 2428 3976 2440
rect 3927 2400 3976 2428
rect 3927 2397 3939 2400
rect 3881 2391 3939 2397
rect 3970 2388 3976 2400
rect 4028 2388 4034 2440
rect 4341 2431 4399 2437
rect 4341 2397 4353 2431
rect 4387 2428 4399 2431
rect 4522 2428 4528 2440
rect 4387 2400 4528 2428
rect 4387 2397 4399 2400
rect 4341 2391 4399 2397
rect 4522 2388 4528 2400
rect 4580 2388 4586 2440
rect 4706 2388 4712 2440
rect 4764 2428 4770 2440
rect 4801 2431 4859 2437
rect 4801 2428 4813 2431
rect 4764 2400 4813 2428
rect 4764 2388 4770 2400
rect 4801 2397 4813 2400
rect 4847 2397 4859 2431
rect 4801 2391 4859 2397
rect 4893 2431 4951 2437
rect 4893 2397 4905 2431
rect 4939 2428 4951 2431
rect 5166 2428 5172 2440
rect 4939 2400 5172 2428
rect 4939 2397 4951 2400
rect 4893 2391 4951 2397
rect 5166 2388 5172 2400
rect 5224 2388 5230 2440
rect 5261 2431 5319 2437
rect 5261 2397 5273 2431
rect 5307 2428 5319 2431
rect 5736 2428 5764 2527
rect 7742 2524 7748 2536
rect 7800 2524 7806 2576
rect 8573 2567 8631 2573
rect 8573 2533 8585 2567
rect 8619 2564 8631 2567
rect 8846 2564 8852 2576
rect 8619 2536 8852 2564
rect 8619 2533 8631 2536
rect 8573 2527 8631 2533
rect 8846 2524 8852 2536
rect 8904 2524 8910 2576
rect 6822 2456 6828 2508
rect 6880 2496 6886 2508
rect 6880 2468 7328 2496
rect 6880 2456 6886 2468
rect 5307 2400 5764 2428
rect 5905 2431 5963 2437
rect 5307 2397 5319 2400
rect 5261 2391 5319 2397
rect 5905 2397 5917 2431
rect 5951 2428 5963 2431
rect 5997 2431 6055 2437
rect 5997 2428 6009 2431
rect 5951 2400 6009 2428
rect 5951 2397 5963 2400
rect 5905 2391 5963 2397
rect 5997 2397 6009 2400
rect 6043 2397 6055 2431
rect 6273 2431 6331 2437
rect 6273 2428 6285 2431
rect 5997 2391 6055 2397
rect 6196 2400 6285 2428
rect 2777 2363 2835 2369
rect 2777 2329 2789 2363
rect 2823 2360 2835 2363
rect 5537 2363 5595 2369
rect 2823 2332 4660 2360
rect 2823 2329 2835 2332
rect 2777 2323 2835 2329
rect 4632 2301 4660 2332
rect 5537 2329 5549 2363
rect 5583 2360 5595 2363
rect 5920 2360 5948 2391
rect 5583 2332 5948 2360
rect 5583 2329 5595 2332
rect 5537 2323 5595 2329
rect 6196 2301 6224 2400
rect 6273 2397 6285 2400
rect 6319 2397 6331 2431
rect 6730 2428 6736 2440
rect 6691 2400 6736 2428
rect 6273 2391 6331 2397
rect 6730 2388 6736 2400
rect 6788 2388 6794 2440
rect 7190 2428 7196 2440
rect 7151 2400 7196 2428
rect 7190 2388 7196 2400
rect 7248 2388 7254 2440
rect 7300 2437 7328 2468
rect 7374 2456 7380 2508
rect 7432 2496 7438 2508
rect 7561 2499 7619 2505
rect 7561 2496 7573 2499
rect 7432 2468 7573 2496
rect 7432 2456 7438 2468
rect 7561 2465 7573 2468
rect 7607 2465 7619 2499
rect 9030 2496 9036 2508
rect 7561 2459 7619 2465
rect 8312 2468 9036 2496
rect 7285 2431 7343 2437
rect 7285 2397 7297 2431
rect 7331 2397 7343 2431
rect 7285 2391 7343 2397
rect 7745 2431 7803 2437
rect 7745 2397 7757 2431
rect 7791 2428 7803 2431
rect 7834 2428 7840 2440
rect 7791 2400 7840 2428
rect 7791 2397 7803 2400
rect 7745 2391 7803 2397
rect 7834 2388 7840 2400
rect 7892 2388 7898 2440
rect 7926 2388 7932 2440
rect 7984 2428 7990 2440
rect 8312 2437 8340 2468
rect 9030 2456 9036 2468
rect 9088 2496 9094 2508
rect 9232 2496 9260 2604
rect 9088 2468 9260 2496
rect 9953 2499 10011 2505
rect 9088 2456 9094 2468
rect 9953 2465 9965 2499
rect 9999 2496 10011 2499
rect 17770 2496 17776 2508
rect 9999 2468 17776 2496
rect 9999 2465 10011 2468
rect 9953 2459 10011 2465
rect 17770 2456 17776 2468
rect 17828 2456 17834 2508
rect 8297 2431 8355 2437
rect 7984 2400 8029 2428
rect 7984 2388 7990 2400
rect 8297 2397 8309 2431
rect 8343 2397 8355 2431
rect 8297 2391 8355 2397
rect 8389 2431 8447 2437
rect 8389 2397 8401 2431
rect 8435 2397 8447 2431
rect 8389 2391 8447 2397
rect 8757 2431 8815 2437
rect 8757 2397 8769 2431
rect 8803 2428 8815 2431
rect 9398 2428 9404 2440
rect 8803 2400 9404 2428
rect 8803 2397 8815 2400
rect 8757 2391 8815 2397
rect 2685 2295 2743 2301
rect 2685 2261 2697 2295
rect 2731 2292 2743 2295
rect 4525 2295 4583 2301
rect 4525 2292 4537 2295
rect 2731 2264 4537 2292
rect 2731 2261 2743 2264
rect 2685 2255 2743 2261
rect 4525 2261 4537 2264
rect 4571 2261 4583 2295
rect 4525 2255 4583 2261
rect 4617 2295 4675 2301
rect 4617 2261 4629 2295
rect 4663 2261 4675 2295
rect 4617 2255 4675 2261
rect 6181 2295 6239 2301
rect 6181 2261 6193 2295
rect 6227 2261 6239 2295
rect 7208 2292 7236 2388
rect 7650 2320 7656 2372
rect 7708 2360 7714 2372
rect 8404 2360 8432 2391
rect 9398 2388 9404 2400
rect 9456 2388 9462 2440
rect 9493 2431 9551 2437
rect 9493 2397 9505 2431
rect 9539 2428 9551 2431
rect 9858 2428 9864 2440
rect 9539 2400 9864 2428
rect 9539 2397 9551 2400
rect 9493 2391 9551 2397
rect 9858 2388 9864 2400
rect 9916 2388 9922 2440
rect 7708 2332 8432 2360
rect 8680 2332 9352 2360
rect 7708 2320 7714 2332
rect 7834 2292 7840 2304
rect 7208 2264 7840 2292
rect 6181 2255 6239 2261
rect 7834 2252 7840 2264
rect 7892 2252 7898 2304
rect 8018 2252 8024 2304
rect 8076 2292 8082 2304
rect 8680 2292 8708 2332
rect 8076 2264 8708 2292
rect 8076 2252 8082 2264
rect 8938 2252 8944 2304
rect 8996 2292 9002 2304
rect 9324 2301 9352 2332
rect 9217 2295 9275 2301
rect 9217 2292 9229 2295
rect 8996 2264 9229 2292
rect 8996 2252 9002 2264
rect 9217 2261 9229 2264
rect 9263 2261 9275 2295
rect 9217 2255 9275 2261
rect 9309 2295 9367 2301
rect 9309 2261 9321 2295
rect 9355 2261 9367 2295
rect 9309 2255 9367 2261
rect 3036 2202 9844 2224
rect 3036 2150 4116 2202
rect 4168 2150 4180 2202
rect 4232 2150 4244 2202
rect 4296 2150 4308 2202
rect 4360 2150 4372 2202
rect 4424 2150 7216 2202
rect 7268 2150 7280 2202
rect 7332 2150 7344 2202
rect 7396 2150 7408 2202
rect 7460 2150 7472 2202
rect 7524 2150 9844 2202
rect 3036 2128 9844 2150
rect 2958 2048 2964 2100
rect 3016 2088 3022 2100
rect 3605 2091 3663 2097
rect 3605 2088 3617 2091
rect 3016 2060 3617 2088
rect 3016 2048 3022 2060
rect 3605 2057 3617 2060
rect 3651 2057 3663 2091
rect 3605 2051 3663 2057
rect 3878 2048 3884 2100
rect 3936 2088 3942 2100
rect 3936 2060 4200 2088
rect 3936 2048 3942 2060
rect 3050 1980 3056 2032
rect 3108 2020 3114 2032
rect 4172 2020 4200 2060
rect 5166 2048 5172 2100
rect 5224 2088 5230 2100
rect 5261 2091 5319 2097
rect 5261 2088 5273 2091
rect 5224 2060 5273 2088
rect 5224 2048 5230 2060
rect 5261 2057 5273 2060
rect 5307 2088 5319 2091
rect 6454 2088 6460 2100
rect 5307 2060 6460 2088
rect 5307 2057 5319 2060
rect 5261 2051 5319 2057
rect 6454 2048 6460 2060
rect 6512 2048 6518 2100
rect 7561 2091 7619 2097
rect 7561 2057 7573 2091
rect 7607 2088 7619 2091
rect 7742 2088 7748 2100
rect 7607 2060 7748 2088
rect 7607 2057 7619 2060
rect 7561 2051 7619 2057
rect 4617 2023 4675 2029
rect 4617 2020 4629 2023
rect 3108 1992 3924 2020
rect 4172 1992 4629 2020
rect 3108 1980 3114 1992
rect 3896 1964 3924 1992
rect 4617 1989 4629 1992
rect 4663 1989 4675 2023
rect 4890 2020 4896 2032
rect 4803 1992 4896 2020
rect 4617 1983 4675 1989
rect 4890 1980 4896 1992
rect 4948 2020 4954 2032
rect 6270 2020 6276 2032
rect 4948 1992 6276 2020
rect 4948 1980 4954 1992
rect 6270 1980 6276 1992
rect 6328 1980 6334 2032
rect 2682 1912 2688 1964
rect 2740 1952 2746 1964
rect 3329 1955 3387 1961
rect 3329 1952 3341 1955
rect 2740 1924 3341 1952
rect 2740 1912 2746 1924
rect 3329 1921 3341 1924
rect 3375 1952 3387 1955
rect 3418 1952 3424 1964
rect 3375 1924 3424 1952
rect 3375 1921 3387 1924
rect 3329 1915 3387 1921
rect 3418 1912 3424 1924
rect 3476 1912 3482 1964
rect 3510 1912 3516 1964
rect 3568 1952 3574 1964
rect 3789 1955 3847 1961
rect 3789 1952 3801 1955
rect 3568 1924 3801 1952
rect 3568 1912 3574 1924
rect 3789 1921 3801 1924
rect 3835 1921 3847 1955
rect 3789 1915 3847 1921
rect 3878 1912 3884 1964
rect 3936 1952 3942 1964
rect 4157 1955 4215 1961
rect 3936 1924 4029 1952
rect 3936 1912 3942 1924
rect 4157 1921 4169 1955
rect 4203 1952 4215 1955
rect 6178 1952 6184 1964
rect 4203 1924 6184 1952
rect 4203 1921 4215 1924
rect 4157 1915 4215 1921
rect 6178 1912 6184 1924
rect 6236 1912 6242 1964
rect 7668 1961 7696 2060
rect 7742 2048 7748 2060
rect 7800 2048 7806 2100
rect 7834 2048 7840 2100
rect 7892 2088 7898 2100
rect 8110 2088 8116 2100
rect 7892 2060 7937 2088
rect 8071 2060 8116 2088
rect 7892 2048 7898 2060
rect 8110 2048 8116 2060
rect 8168 2048 8174 2100
rect 8478 2048 8484 2100
rect 8536 2088 8542 2100
rect 8573 2091 8631 2097
rect 8573 2088 8585 2091
rect 8536 2060 8585 2088
rect 8536 2048 8542 2060
rect 8573 2057 8585 2060
rect 8619 2057 8631 2091
rect 8573 2051 8631 2057
rect 8849 2091 8907 2097
rect 8849 2057 8861 2091
rect 8895 2088 8907 2091
rect 9214 2088 9220 2100
rect 8895 2060 9220 2088
rect 8895 2057 8907 2060
rect 8849 2051 8907 2057
rect 9214 2048 9220 2060
rect 9272 2048 9278 2100
rect 9401 2091 9459 2097
rect 9401 2057 9413 2091
rect 9447 2088 9459 2091
rect 9447 2060 16574 2088
rect 9447 2057 9459 2060
rect 9401 2051 9459 2057
rect 8202 1980 8208 2032
rect 8260 2020 8266 2032
rect 8260 1992 9168 2020
rect 8260 1980 8266 1992
rect 7653 1955 7711 1961
rect 7653 1921 7665 1955
rect 7699 1921 7711 1955
rect 7653 1915 7711 1921
rect 7929 1955 7987 1961
rect 7929 1921 7941 1955
rect 7975 1921 7987 1955
rect 7929 1915 7987 1921
rect 2869 1887 2927 1893
rect 2869 1853 2881 1887
rect 2915 1884 2927 1887
rect 4433 1887 4491 1893
rect 4433 1884 4445 1887
rect 2915 1856 4445 1884
rect 2915 1853 2927 1856
rect 2869 1847 2927 1853
rect 4433 1853 4445 1856
rect 4479 1853 4491 1887
rect 4433 1847 4491 1853
rect 4522 1844 4528 1896
rect 4580 1884 4586 1896
rect 4982 1884 4988 1896
rect 4580 1856 4988 1884
rect 4580 1844 4586 1856
rect 4982 1844 4988 1856
rect 5040 1884 5046 1896
rect 5353 1887 5411 1893
rect 5353 1884 5365 1887
rect 5040 1856 5365 1884
rect 5040 1844 5046 1856
rect 5353 1853 5365 1856
rect 5399 1853 5411 1887
rect 7944 1884 7972 1915
rect 8294 1912 8300 1964
rect 8352 1952 8358 1964
rect 8389 1955 8447 1961
rect 8389 1952 8401 1955
rect 8352 1924 8401 1952
rect 8352 1912 8358 1924
rect 8389 1921 8401 1924
rect 8435 1921 8447 1955
rect 8389 1915 8447 1921
rect 8665 1955 8723 1961
rect 8665 1921 8677 1955
rect 8711 1952 8723 1955
rect 8938 1952 8944 1964
rect 8711 1924 8944 1952
rect 8711 1921 8723 1924
rect 8665 1915 8723 1921
rect 8938 1912 8944 1924
rect 8996 1912 9002 1964
rect 9140 1961 9168 1992
rect 9125 1955 9183 1961
rect 9125 1921 9137 1955
rect 9171 1921 9183 1955
rect 9125 1915 9183 1921
rect 9217 1955 9275 1961
rect 9217 1921 9229 1955
rect 9263 1921 9275 1955
rect 9217 1915 9275 1921
rect 8478 1884 8484 1896
rect 7944 1856 8484 1884
rect 5353 1847 5411 1853
rect 8478 1844 8484 1856
rect 8536 1844 8542 1896
rect 8570 1844 8576 1896
rect 8628 1884 8634 1896
rect 9232 1884 9260 1915
rect 8628 1856 9260 1884
rect 8628 1844 8634 1856
rect 16546 1828 16574 2060
rect 3142 1776 3148 1828
rect 3200 1816 3206 1828
rect 4065 1819 4123 1825
rect 4065 1816 4077 1819
rect 3200 1788 4077 1816
rect 3200 1776 3206 1788
rect 4065 1785 4077 1788
rect 4111 1785 4123 1819
rect 4065 1779 4123 1785
rect 4341 1819 4399 1825
rect 4341 1785 4353 1819
rect 4387 1816 4399 1819
rect 4387 1788 12434 1816
rect 16546 1788 16580 1828
rect 4387 1785 4399 1788
rect 4341 1779 4399 1785
rect 3513 1751 3571 1757
rect 3513 1717 3525 1751
rect 3559 1748 3571 1751
rect 4246 1748 4252 1760
rect 3559 1720 4252 1748
rect 3559 1717 3571 1720
rect 3513 1711 3571 1717
rect 4246 1708 4252 1720
rect 4304 1708 4310 1760
rect 4706 1708 4712 1760
rect 4764 1748 4770 1760
rect 5077 1751 5135 1757
rect 5077 1748 5089 1751
rect 4764 1720 5089 1748
rect 4764 1708 4770 1720
rect 5077 1717 5089 1720
rect 5123 1748 5135 1751
rect 6362 1748 6368 1760
rect 5123 1720 6368 1748
rect 5123 1717 5135 1720
rect 5077 1711 5135 1717
rect 6362 1708 6368 1720
rect 6420 1708 6426 1760
rect 8386 1708 8392 1760
rect 8444 1748 8450 1760
rect 8941 1751 8999 1757
rect 8941 1748 8953 1751
rect 8444 1720 8953 1748
rect 8444 1708 8450 1720
rect 8941 1717 8953 1720
rect 8987 1717 8999 1751
rect 12406 1748 12434 1788
rect 16574 1776 16580 1788
rect 16632 1776 16638 1828
rect 21358 1748 21364 1760
rect 12406 1720 21364 1748
rect 8941 1711 8999 1717
rect 21358 1708 21364 1720
rect 21416 1708 21422 1760
rect 3036 1658 9844 1680
rect 3036 1606 5666 1658
rect 5718 1606 5730 1658
rect 5782 1606 5794 1658
rect 5846 1606 5858 1658
rect 5910 1606 5922 1658
rect 5974 1606 8766 1658
rect 8818 1606 8830 1658
rect 8882 1606 8894 1658
rect 8946 1606 8958 1658
rect 9010 1606 9022 1658
rect 9074 1606 9844 1658
rect 3036 1584 9844 1606
rect 1026 1504 1032 1556
rect 1084 1544 1090 1556
rect 2869 1547 2927 1553
rect 2869 1544 2881 1547
rect 1084 1516 2881 1544
rect 1084 1504 1090 1516
rect 2869 1513 2881 1516
rect 2915 1513 2927 1547
rect 2869 1507 2927 1513
rect 3418 1504 3424 1556
rect 3476 1544 3482 1556
rect 3973 1547 4031 1553
rect 3973 1544 3985 1547
rect 3476 1516 3985 1544
rect 3476 1504 3482 1516
rect 3973 1513 3985 1516
rect 4019 1513 4031 1547
rect 3973 1507 4031 1513
rect 4062 1504 4068 1556
rect 4120 1544 4126 1556
rect 4157 1547 4215 1553
rect 4157 1544 4169 1547
rect 4120 1516 4169 1544
rect 4120 1504 4126 1516
rect 4157 1513 4169 1516
rect 4203 1513 4215 1547
rect 4157 1507 4215 1513
rect 4246 1504 4252 1556
rect 4304 1544 4310 1556
rect 5074 1544 5080 1556
rect 4304 1516 5080 1544
rect 4304 1504 4310 1516
rect 5074 1504 5080 1516
rect 5132 1504 5138 1556
rect 8389 1547 8447 1553
rect 8389 1513 8401 1547
rect 8435 1544 8447 1547
rect 8478 1544 8484 1556
rect 8435 1516 8484 1544
rect 8435 1513 8447 1516
rect 8389 1507 8447 1513
rect 8478 1504 8484 1516
rect 8536 1544 8542 1556
rect 9122 1544 9128 1556
rect 8536 1516 9128 1544
rect 8536 1504 8542 1516
rect 9122 1504 9128 1516
rect 9180 1504 9186 1556
rect 3326 1436 3332 1488
rect 3384 1476 3390 1488
rect 3605 1479 3663 1485
rect 3605 1476 3617 1479
rect 3384 1448 3617 1476
rect 3384 1436 3390 1448
rect 3605 1445 3617 1448
rect 3651 1476 3663 1479
rect 3651 1448 4476 1476
rect 3651 1445 3663 1448
rect 3605 1439 3663 1445
rect 3510 1368 3516 1420
rect 3568 1408 3574 1420
rect 4341 1411 4399 1417
rect 4341 1408 4353 1411
rect 3568 1380 4353 1408
rect 3568 1368 3574 1380
rect 4341 1377 4353 1380
rect 4387 1377 4399 1411
rect 4448 1408 4476 1448
rect 7926 1436 7932 1488
rect 7984 1476 7990 1488
rect 8938 1476 8944 1488
rect 7984 1448 8944 1476
rect 7984 1436 7990 1448
rect 8938 1436 8944 1448
rect 8996 1436 9002 1488
rect 9953 1479 10011 1485
rect 9953 1476 9965 1479
rect 9048 1448 9965 1476
rect 9048 1408 9076 1448
rect 9953 1445 9965 1448
rect 9999 1445 10011 1479
rect 9953 1439 10011 1445
rect 4448 1380 9076 1408
rect 9125 1411 9183 1417
rect 4341 1371 4399 1377
rect 9125 1377 9137 1411
rect 9171 1408 9183 1411
rect 9214 1408 9220 1420
rect 9171 1380 9220 1408
rect 9171 1377 9183 1380
rect 9125 1371 9183 1377
rect 9214 1368 9220 1380
rect 9272 1368 9278 1420
rect 9324 1380 9628 1408
rect 3329 1343 3387 1349
rect 3329 1309 3341 1343
rect 3375 1340 3387 1343
rect 7558 1340 7564 1352
rect 3375 1312 7564 1340
rect 3375 1309 3387 1312
rect 3329 1303 3387 1309
rect 7558 1300 7564 1312
rect 7616 1300 7622 1352
rect 8573 1343 8631 1349
rect 8573 1309 8585 1343
rect 8619 1340 8631 1343
rect 8665 1343 8723 1349
rect 8665 1340 8677 1343
rect 8619 1312 8677 1340
rect 8619 1309 8631 1312
rect 8573 1303 8631 1309
rect 8665 1309 8677 1312
rect 8711 1340 8723 1343
rect 9324 1340 9352 1380
rect 9490 1340 9496 1352
rect 8711 1312 9352 1340
rect 9451 1312 9496 1340
rect 8711 1309 8723 1312
rect 8665 1303 8723 1309
rect 9490 1300 9496 1312
rect 9548 1300 9554 1352
rect 9600 1340 9628 1380
rect 13814 1340 13820 1352
rect 9600 1312 13820 1340
rect 13814 1300 13820 1312
rect 13872 1300 13878 1352
rect 10870 1272 10876 1284
rect 3528 1244 10876 1272
rect 3528 1213 3556 1244
rect 10870 1232 10876 1244
rect 10928 1232 10934 1284
rect 3513 1207 3571 1213
rect 3513 1173 3525 1207
rect 3559 1173 3571 1207
rect 3786 1204 3792 1216
rect 3747 1176 3792 1204
rect 3513 1167 3571 1173
rect 3786 1164 3792 1176
rect 3844 1164 3850 1216
rect 3878 1164 3884 1216
rect 3936 1204 3942 1216
rect 4525 1207 4583 1213
rect 4525 1204 4537 1207
rect 3936 1176 4537 1204
rect 3936 1164 3942 1176
rect 4525 1173 4537 1176
rect 4571 1173 4583 1207
rect 4525 1167 4583 1173
rect 8662 1164 8668 1216
rect 8720 1204 8726 1216
rect 8849 1207 8907 1213
rect 8849 1204 8861 1207
rect 8720 1176 8861 1204
rect 8720 1164 8726 1176
rect 8849 1173 8861 1176
rect 8895 1173 8907 1207
rect 8849 1167 8907 1173
rect 8938 1164 8944 1216
rect 8996 1204 9002 1216
rect 9309 1207 9367 1213
rect 8996 1176 9041 1204
rect 8996 1164 9002 1176
rect 9309 1173 9321 1207
rect 9355 1204 9367 1207
rect 9582 1204 9588 1216
rect 9355 1176 9588 1204
rect 9355 1173 9367 1176
rect 9309 1167 9367 1173
rect 9582 1164 9588 1176
rect 9640 1164 9646 1216
rect 3036 1114 9844 1136
rect 3036 1062 4116 1114
rect 4168 1062 4180 1114
rect 4232 1062 4244 1114
rect 4296 1062 4308 1114
rect 4360 1062 4372 1114
rect 4424 1062 7216 1114
rect 7268 1062 7280 1114
rect 7332 1062 7344 1114
rect 7396 1062 7408 1114
rect 7460 1062 7472 1114
rect 7524 1062 9844 1114
rect 3036 1040 9844 1062
<< via1 >>
rect 1952 12112 2004 12164
rect 2320 12112 2372 12164
rect 6000 12112 6052 12164
rect 6368 12112 6420 12164
rect 4160 12044 4212 12096
rect 5356 12044 5408 12096
rect 6092 12044 6144 12096
rect 6460 12044 6512 12096
rect 2320 11976 2372 12028
rect 7840 11976 7892 12028
rect 2412 11840 2464 11892
rect 8576 11908 8628 11960
rect 2964 11840 3016 11892
rect 8392 11840 8444 11892
rect 4344 11772 4396 11824
rect 6092 11772 6144 11824
rect 6828 11772 6880 11824
rect 8208 11772 8260 11824
rect 1492 11704 1544 11756
rect 6920 11704 6972 11756
rect 2228 11636 2280 11688
rect 4712 11636 4764 11688
rect 1308 11568 1360 11620
rect 6184 11568 6236 11620
rect 7104 11568 7156 11620
rect 9680 11568 9732 11620
rect 5264 11500 5316 11552
rect 8300 11500 8352 11552
rect 8484 11500 8536 11552
rect 10416 11500 10468 11552
rect 2566 11398 2618 11450
rect 2630 11398 2682 11450
rect 2694 11398 2746 11450
rect 2758 11398 2810 11450
rect 2822 11398 2874 11450
rect 5666 11398 5718 11450
rect 5730 11398 5782 11450
rect 5794 11398 5846 11450
rect 5858 11398 5910 11450
rect 5922 11398 5974 11450
rect 8766 11398 8818 11450
rect 8830 11398 8882 11450
rect 8894 11398 8946 11450
rect 8958 11398 9010 11450
rect 9022 11398 9074 11450
rect 1492 11339 1544 11348
rect 1492 11305 1501 11339
rect 1501 11305 1535 11339
rect 1535 11305 1544 11339
rect 1492 11296 1544 11305
rect 2228 11296 2280 11348
rect 2320 11296 2372 11348
rect 2964 11296 3016 11348
rect 6460 11339 6512 11348
rect 1308 11135 1360 11144
rect 1308 11101 1317 11135
rect 1317 11101 1351 11135
rect 1351 11101 1360 11135
rect 1308 11092 1360 11101
rect 1952 11228 2004 11280
rect 4344 11271 4396 11280
rect 4344 11237 4353 11271
rect 4353 11237 4387 11271
rect 4387 11237 4396 11271
rect 4344 11228 4396 11237
rect 4804 11228 4856 11280
rect 5264 11228 5316 11280
rect 5448 11271 5500 11280
rect 5448 11237 5457 11271
rect 5457 11237 5491 11271
rect 5491 11237 5500 11271
rect 5448 11228 5500 11237
rect 6184 11271 6236 11280
rect 6184 11237 6193 11271
rect 6193 11237 6227 11271
rect 6227 11237 6236 11271
rect 6184 11228 6236 11237
rect 6460 11305 6469 11339
rect 6469 11305 6503 11339
rect 6503 11305 6512 11339
rect 6460 11296 6512 11305
rect 7104 11296 7156 11348
rect 7196 11296 7248 11348
rect 7932 11339 7984 11348
rect 7932 11305 7941 11339
rect 7941 11305 7975 11339
rect 7975 11305 7984 11339
rect 7932 11296 7984 11305
rect 8484 11339 8536 11348
rect 8484 11305 8493 11339
rect 8493 11305 8527 11339
rect 8527 11305 8536 11339
rect 8484 11296 8536 11305
rect 8668 11296 8720 11348
rect 6644 11228 6696 11280
rect 2044 11135 2096 11144
rect 2044 11101 2053 11135
rect 2053 11101 2087 11135
rect 2087 11101 2096 11135
rect 2044 11092 2096 11101
rect 2228 11092 2280 11144
rect 2412 11135 2464 11144
rect 2412 11101 2421 11135
rect 2421 11101 2455 11135
rect 2455 11101 2464 11135
rect 2412 11092 2464 11101
rect 2688 11135 2740 11144
rect 2688 11101 2697 11135
rect 2697 11101 2731 11135
rect 2731 11101 2740 11135
rect 2688 11092 2740 11101
rect 2964 11135 3016 11144
rect 2964 11101 2973 11135
rect 2973 11101 3007 11135
rect 3007 11101 3016 11135
rect 2964 11092 3016 11101
rect 3424 11135 3476 11144
rect 3424 11101 3433 11135
rect 3433 11101 3467 11135
rect 3467 11101 3476 11135
rect 3424 11092 3476 11101
rect 3516 11092 3568 11144
rect 3884 11092 3936 11144
rect 4528 11092 4580 11144
rect 5080 11092 5132 11144
rect 7288 11160 7340 11212
rect 9864 11160 9916 11212
rect 3608 11067 3660 11076
rect 3608 11033 3617 11067
rect 3617 11033 3651 11067
rect 3651 11033 3660 11067
rect 3608 11024 3660 11033
rect 3976 11024 4028 11076
rect 5816 11092 5868 11144
rect 6736 11092 6788 11144
rect 7104 11135 7156 11144
rect 7104 11101 7113 11135
rect 7113 11101 7147 11135
rect 7147 11101 7156 11135
rect 7104 11092 7156 11101
rect 7656 11092 7708 11144
rect 8116 11135 8168 11144
rect 8116 11101 8125 11135
rect 8125 11101 8159 11135
rect 8159 11101 8168 11135
rect 8116 11092 8168 11101
rect 8208 11092 8260 11144
rect 9128 11092 9180 11144
rect 1860 10956 1912 11008
rect 2136 10956 2188 11008
rect 2412 10956 2464 11008
rect 2964 10956 3016 11008
rect 6460 11024 6512 11076
rect 7932 11024 7984 11076
rect 5080 10999 5132 11008
rect 5080 10965 5089 10999
rect 5089 10965 5123 10999
rect 5123 10965 5132 10999
rect 5080 10956 5132 10965
rect 5908 10999 5960 11008
rect 5908 10965 5917 10999
rect 5917 10965 5951 10999
rect 5951 10965 5960 10999
rect 5908 10956 5960 10965
rect 6276 10956 6328 11008
rect 9588 10956 9640 11008
rect 4116 10854 4168 10906
rect 4180 10854 4232 10906
rect 4244 10854 4296 10906
rect 4308 10854 4360 10906
rect 4372 10854 4424 10906
rect 7216 10854 7268 10906
rect 7280 10854 7332 10906
rect 7344 10854 7396 10906
rect 7408 10854 7460 10906
rect 7472 10854 7524 10906
rect 1492 10795 1544 10804
rect 1492 10761 1501 10795
rect 1501 10761 1535 10795
rect 1535 10761 1544 10795
rect 1492 10752 1544 10761
rect 2228 10752 2280 10804
rect 3056 10795 3108 10804
rect 3056 10761 3065 10795
rect 3065 10761 3099 10795
rect 3099 10761 3108 10795
rect 3056 10752 3108 10761
rect 3332 10752 3384 10804
rect 3516 10752 3568 10804
rect 7012 10752 7064 10804
rect 8484 10752 8536 10804
rect 8576 10752 8628 10804
rect 5816 10727 5868 10736
rect 5816 10693 5825 10727
rect 5825 10693 5859 10727
rect 5859 10693 5868 10727
rect 5816 10684 5868 10693
rect 6920 10684 6972 10736
rect 1584 10659 1636 10668
rect 1584 10625 1593 10659
rect 1593 10625 1627 10659
rect 1627 10625 1636 10659
rect 1584 10616 1636 10625
rect 1952 10616 2004 10668
rect 2228 10616 2280 10668
rect 2872 10616 2924 10668
rect 3516 10616 3568 10668
rect 3608 10659 3660 10668
rect 3608 10625 3617 10659
rect 3617 10625 3651 10659
rect 3651 10625 3660 10659
rect 4252 10659 4304 10668
rect 3608 10616 3660 10625
rect 4252 10625 4261 10659
rect 4261 10625 4295 10659
rect 4295 10625 4304 10659
rect 4252 10616 4304 10625
rect 2872 10480 2924 10532
rect 2964 10480 3016 10532
rect 3976 10548 4028 10600
rect 4896 10616 4948 10668
rect 4988 10616 5040 10668
rect 6460 10616 6512 10668
rect 8024 10659 8076 10668
rect 8024 10625 8033 10659
rect 8033 10625 8067 10659
rect 8067 10625 8076 10659
rect 8024 10616 8076 10625
rect 8116 10616 8168 10668
rect 4712 10548 4764 10600
rect 6552 10591 6604 10600
rect 6552 10557 6561 10591
rect 6561 10557 6595 10591
rect 6595 10557 6604 10591
rect 6552 10548 6604 10557
rect 9312 10616 9364 10668
rect 4344 10480 4396 10532
rect 8024 10480 8076 10532
rect 9588 10548 9640 10600
rect 9220 10480 9272 10532
rect 4988 10455 5040 10464
rect 4988 10421 4997 10455
rect 4997 10421 5031 10455
rect 5031 10421 5040 10455
rect 4988 10412 5040 10421
rect 7012 10412 7064 10464
rect 15200 10412 15252 10464
rect 16580 10412 16632 10464
rect 2566 10310 2618 10362
rect 2630 10310 2682 10362
rect 2694 10310 2746 10362
rect 2758 10310 2810 10362
rect 2822 10310 2874 10362
rect 5666 10310 5718 10362
rect 5730 10310 5782 10362
rect 5794 10310 5846 10362
rect 5858 10310 5910 10362
rect 5922 10310 5974 10362
rect 8766 10310 8818 10362
rect 8830 10310 8882 10362
rect 8894 10310 8946 10362
rect 8958 10310 9010 10362
rect 9022 10310 9074 10362
rect 6184 10208 6236 10260
rect 7564 10208 7616 10260
rect 8024 10208 8076 10260
rect 5080 10140 5132 10192
rect 5632 10140 5684 10192
rect 2412 10072 2464 10124
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 2688 9936 2740 9988
rect 3608 10004 3660 10056
rect 3884 10004 3936 10056
rect 3976 10004 4028 10056
rect 4436 9936 4488 9988
rect 1584 9911 1636 9920
rect 1584 9877 1593 9911
rect 1593 9877 1627 9911
rect 1627 9877 1636 9911
rect 1584 9868 1636 9877
rect 1860 9868 1912 9920
rect 3332 9868 3384 9920
rect 3516 9868 3568 9920
rect 5816 9936 5868 9988
rect 6460 10140 6512 10192
rect 8576 10183 8628 10192
rect 8576 10149 8585 10183
rect 8585 10149 8619 10183
rect 8619 10149 8628 10183
rect 8576 10140 8628 10149
rect 8944 10140 8996 10192
rect 9128 10183 9180 10192
rect 9128 10149 9137 10183
rect 9137 10149 9171 10183
rect 9171 10149 9180 10183
rect 9128 10140 9180 10149
rect 7564 10072 7616 10124
rect 8024 10004 8076 10056
rect 8116 10004 8168 10056
rect 8852 10004 8904 10056
rect 7932 9936 7984 9988
rect 8944 9979 8996 9988
rect 6644 9868 6696 9920
rect 8024 9868 8076 9920
rect 8944 9945 8953 9979
rect 8953 9945 8987 9979
rect 8987 9945 8996 9979
rect 8944 9936 8996 9945
rect 4116 9766 4168 9818
rect 4180 9766 4232 9818
rect 4244 9766 4296 9818
rect 4308 9766 4360 9818
rect 4372 9766 4424 9818
rect 7216 9766 7268 9818
rect 7280 9766 7332 9818
rect 7344 9766 7396 9818
rect 7408 9766 7460 9818
rect 7472 9766 7524 9818
rect 1952 9664 2004 9716
rect 2044 9664 2096 9716
rect 2596 9664 2648 9716
rect 3608 9664 3660 9716
rect 3792 9664 3844 9716
rect 1308 9571 1360 9580
rect 1308 9537 1317 9571
rect 1317 9537 1351 9571
rect 1351 9537 1360 9571
rect 1308 9528 1360 9537
rect 1860 9528 1912 9580
rect 3516 9596 3568 9648
rect 2320 9460 2372 9512
rect 3056 9503 3108 9512
rect 3056 9469 3065 9503
rect 3065 9469 3099 9503
rect 3099 9469 3108 9503
rect 3056 9460 3108 9469
rect 4068 9528 4120 9580
rect 3700 9460 3752 9512
rect 4896 9460 4948 9512
rect 5632 9571 5684 9580
rect 5632 9537 5641 9571
rect 5641 9537 5675 9571
rect 5675 9537 5684 9571
rect 5632 9528 5684 9537
rect 5816 9571 5868 9580
rect 5816 9537 5825 9571
rect 5825 9537 5859 9571
rect 5859 9537 5868 9571
rect 6184 9571 6236 9580
rect 5816 9528 5868 9537
rect 6184 9537 6193 9571
rect 6193 9537 6227 9571
rect 6227 9537 6236 9571
rect 6184 9528 6236 9537
rect 5724 9460 5776 9512
rect 2596 9392 2648 9444
rect 5172 9392 5224 9444
rect 6552 9664 6604 9716
rect 8576 9664 8628 9716
rect 8392 9596 8444 9648
rect 7104 9571 7156 9580
rect 7104 9537 7113 9571
rect 7113 9537 7147 9571
rect 7147 9537 7156 9571
rect 7104 9528 7156 9537
rect 7840 9528 7892 9580
rect 9496 9571 9548 9580
rect 9496 9537 9505 9571
rect 9505 9537 9539 9571
rect 9539 9537 9548 9571
rect 9496 9528 9548 9537
rect 2228 9324 2280 9376
rect 3056 9324 3108 9376
rect 4068 9324 4120 9376
rect 4620 9324 4672 9376
rect 5448 9324 5500 9376
rect 5540 9324 5592 9376
rect 6920 9324 6972 9376
rect 7196 9367 7248 9376
rect 7196 9333 7205 9367
rect 7205 9333 7239 9367
rect 7239 9333 7248 9367
rect 7196 9324 7248 9333
rect 9404 9460 9456 9512
rect 9588 9324 9640 9376
rect 2566 9222 2618 9274
rect 2630 9222 2682 9274
rect 2694 9222 2746 9274
rect 2758 9222 2810 9274
rect 2822 9222 2874 9274
rect 5666 9222 5718 9274
rect 5730 9222 5782 9274
rect 5794 9222 5846 9274
rect 5858 9222 5910 9274
rect 5922 9222 5974 9274
rect 8766 9222 8818 9274
rect 8830 9222 8882 9274
rect 8894 9222 8946 9274
rect 8958 9222 9010 9274
rect 9022 9222 9074 9274
rect 1492 9163 1544 9172
rect 1492 9129 1501 9163
rect 1501 9129 1535 9163
rect 1535 9129 1544 9163
rect 1492 9120 1544 9129
rect 2320 9163 2372 9172
rect 2320 9129 2329 9163
rect 2329 9129 2363 9163
rect 2363 9129 2372 9163
rect 2320 9120 2372 9129
rect 3240 9120 3292 9172
rect 3424 9163 3476 9172
rect 3424 9129 3433 9163
rect 3433 9129 3467 9163
rect 3467 9129 3476 9163
rect 3424 9120 3476 9129
rect 3700 9163 3752 9172
rect 3700 9129 3709 9163
rect 3709 9129 3743 9163
rect 3743 9129 3752 9163
rect 3700 9120 3752 9129
rect 7104 9120 7156 9172
rect 9404 9163 9456 9172
rect 9404 9129 9413 9163
rect 9413 9129 9447 9163
rect 9447 9129 9456 9163
rect 9404 9120 9456 9129
rect 3056 9052 3108 9104
rect 3516 9052 3568 9104
rect 3976 9052 4028 9104
rect 1216 8916 1268 8968
rect 5080 8984 5132 9036
rect 5172 8984 5224 9036
rect 2044 8916 2096 8968
rect 1676 8848 1728 8900
rect 2320 8848 2372 8900
rect 1768 8823 1820 8832
rect 1768 8789 1777 8823
rect 1777 8789 1811 8823
rect 1811 8789 1820 8823
rect 1768 8780 1820 8789
rect 2504 8848 2556 8900
rect 2688 8959 2740 8968
rect 2688 8925 2697 8959
rect 2697 8925 2731 8959
rect 2731 8925 2740 8959
rect 2964 8959 3016 8968
rect 2688 8916 2740 8925
rect 2964 8925 2973 8959
rect 2973 8925 3007 8959
rect 3007 8925 3016 8959
rect 2964 8916 3016 8925
rect 3056 8916 3108 8968
rect 3424 8848 3476 8900
rect 3884 8823 3936 8832
rect 3884 8789 3893 8823
rect 3893 8789 3927 8823
rect 3927 8789 3936 8823
rect 3884 8780 3936 8789
rect 4160 8959 4212 8968
rect 4160 8925 4169 8959
rect 4169 8925 4203 8959
rect 4203 8925 4212 8959
rect 4160 8916 4212 8925
rect 4620 8916 4672 8968
rect 8300 8984 8352 9036
rect 8576 8984 8628 9036
rect 5080 8891 5132 8900
rect 4620 8780 4672 8832
rect 5080 8857 5089 8891
rect 5089 8857 5123 8891
rect 5123 8857 5132 8891
rect 5080 8848 5132 8857
rect 5172 8780 5224 8832
rect 7012 8916 7064 8968
rect 5908 8848 5960 8900
rect 8392 8916 8444 8968
rect 9404 8848 9456 8900
rect 7012 8780 7064 8832
rect 8300 8780 8352 8832
rect 9128 8780 9180 8832
rect 4116 8678 4168 8730
rect 4180 8678 4232 8730
rect 4244 8678 4296 8730
rect 4308 8678 4360 8730
rect 4372 8678 4424 8730
rect 7216 8678 7268 8730
rect 7280 8678 7332 8730
rect 7344 8678 7396 8730
rect 7408 8678 7460 8730
rect 7472 8678 7524 8730
rect 1768 8576 1820 8628
rect 1860 8508 1912 8560
rect 4436 8508 4488 8560
rect 5080 8508 5132 8560
rect 6092 8508 6144 8560
rect 1584 8440 1636 8492
rect 2228 8483 2280 8492
rect 2228 8449 2237 8483
rect 2237 8449 2271 8483
rect 2271 8449 2280 8483
rect 2228 8440 2280 8449
rect 6552 8440 6604 8492
rect 6736 8440 6788 8492
rect 6920 8483 6972 8492
rect 6920 8449 6929 8483
rect 6929 8449 6963 8483
rect 6963 8449 6972 8483
rect 6920 8440 6972 8449
rect 8208 8508 8260 8560
rect 1492 8279 1544 8288
rect 1492 8245 1501 8279
rect 1501 8245 1535 8279
rect 1535 8245 1544 8279
rect 1492 8236 1544 8245
rect 1768 8236 1820 8288
rect 3332 8236 3384 8288
rect 5080 8372 5132 8424
rect 5908 8415 5960 8424
rect 5908 8381 5917 8415
rect 5917 8381 5951 8415
rect 5951 8381 5960 8415
rect 5908 8372 5960 8381
rect 9128 8415 9180 8424
rect 9128 8381 9137 8415
rect 9137 8381 9171 8415
rect 9171 8381 9180 8415
rect 9128 8372 9180 8381
rect 7656 8304 7708 8356
rect 3976 8236 4028 8288
rect 4528 8236 4580 8288
rect 5448 8236 5500 8288
rect 6000 8236 6052 8288
rect 7012 8236 7064 8288
rect 2566 8134 2618 8186
rect 2630 8134 2682 8186
rect 2694 8134 2746 8186
rect 2758 8134 2810 8186
rect 2822 8134 2874 8186
rect 5666 8134 5718 8186
rect 5730 8134 5782 8186
rect 5794 8134 5846 8186
rect 5858 8134 5910 8186
rect 5922 8134 5974 8186
rect 8766 8134 8818 8186
rect 8830 8134 8882 8186
rect 8894 8134 8946 8186
rect 8958 8134 9010 8186
rect 9022 8134 9074 8186
rect 1308 8075 1360 8084
rect 1308 8041 1317 8075
rect 1317 8041 1351 8075
rect 1351 8041 1360 8075
rect 1308 8032 1360 8041
rect 3056 8032 3108 8084
rect 3976 8032 4028 8084
rect 4068 8032 4120 8084
rect 4528 8075 4580 8084
rect 4528 8041 4537 8075
rect 4537 8041 4571 8075
rect 4571 8041 4580 8075
rect 4528 8032 4580 8041
rect 8392 8032 8444 8084
rect 8576 8007 8628 8016
rect 8576 7973 8585 8007
rect 8585 7973 8619 8007
rect 8619 7973 8628 8007
rect 8576 7964 8628 7973
rect 1676 7896 1728 7948
rect 6000 7896 6052 7948
rect 1308 7828 1360 7880
rect 3424 7871 3476 7880
rect 3424 7837 3433 7871
rect 3433 7837 3467 7871
rect 3467 7837 3476 7871
rect 3424 7828 3476 7837
rect 2688 7760 2740 7812
rect 3516 7760 3568 7812
rect 2228 7692 2280 7744
rect 3424 7692 3476 7744
rect 4344 7828 4396 7880
rect 4620 7760 4672 7812
rect 4896 7871 4948 7880
rect 4896 7837 4905 7871
rect 4905 7837 4939 7871
rect 4939 7837 4948 7871
rect 7012 7871 7064 7880
rect 4896 7828 4948 7837
rect 7012 7837 7021 7871
rect 7021 7837 7055 7871
rect 7055 7837 7064 7871
rect 7012 7828 7064 7837
rect 4528 7692 4580 7744
rect 5172 7692 5224 7744
rect 6920 7760 6972 7812
rect 8300 7828 8352 7880
rect 8392 7803 8444 7812
rect 8392 7769 8401 7803
rect 8401 7769 8435 7803
rect 8435 7769 8444 7803
rect 8392 7760 8444 7769
rect 7012 7692 7064 7744
rect 8116 7692 8168 7744
rect 9404 7735 9456 7744
rect 9404 7701 9413 7735
rect 9413 7701 9447 7735
rect 9447 7701 9456 7735
rect 9404 7692 9456 7701
rect 4116 7590 4168 7642
rect 4180 7590 4232 7642
rect 4244 7590 4296 7642
rect 4308 7590 4360 7642
rect 4372 7590 4424 7642
rect 7216 7590 7268 7642
rect 7280 7590 7332 7642
rect 7344 7590 7396 7642
rect 7408 7590 7460 7642
rect 7472 7590 7524 7642
rect 3240 7420 3292 7472
rect 4712 7420 4764 7472
rect 5172 7420 5224 7472
rect 8392 7488 8444 7540
rect 7932 7463 7984 7472
rect 7932 7429 7941 7463
rect 7941 7429 7975 7463
rect 7975 7429 7984 7463
rect 7932 7420 7984 7429
rect 1768 7352 1820 7404
rect 4804 7352 4856 7404
rect 1492 7284 1544 7336
rect 4712 7284 4764 7336
rect 6092 7352 6144 7404
rect 6828 7352 6880 7404
rect 7748 7352 7800 7404
rect 9312 7352 9364 7404
rect 1308 7216 1360 7268
rect 2136 7216 2188 7268
rect 8392 7284 8444 7336
rect 9220 7327 9272 7336
rect 9220 7293 9229 7327
rect 9229 7293 9263 7327
rect 9263 7293 9272 7327
rect 9220 7284 9272 7293
rect 9588 7284 9640 7336
rect 1676 7148 1728 7200
rect 4344 7148 4396 7200
rect 5816 7216 5868 7268
rect 6828 7216 6880 7268
rect 7104 7216 7156 7268
rect 7288 7148 7340 7200
rect 9588 7148 9640 7200
rect 2566 7046 2618 7098
rect 2630 7046 2682 7098
rect 2694 7046 2746 7098
rect 2758 7046 2810 7098
rect 2822 7046 2874 7098
rect 5666 7046 5718 7098
rect 5730 7046 5782 7098
rect 5794 7046 5846 7098
rect 5858 7046 5910 7098
rect 5922 7046 5974 7098
rect 8766 7046 8818 7098
rect 8830 7046 8882 7098
rect 8894 7046 8946 7098
rect 8958 7046 9010 7098
rect 9022 7046 9074 7098
rect 940 6944 992 6996
rect 1768 6944 1820 6996
rect 2412 6944 2464 6996
rect 4344 6944 4396 6996
rect 5632 6876 5684 6928
rect 5816 6876 5868 6928
rect 6184 6944 6236 6996
rect 6920 6944 6972 6996
rect 7012 6944 7064 6996
rect 8300 6987 8352 6996
rect 1952 6808 2004 6860
rect 4528 6808 4580 6860
rect 6092 6808 6144 6860
rect 1676 6783 1728 6792
rect 1676 6749 1685 6783
rect 1685 6749 1719 6783
rect 1719 6749 1728 6783
rect 1676 6740 1728 6749
rect 3056 6740 3108 6792
rect 3608 6783 3660 6792
rect 3608 6749 3617 6783
rect 3617 6749 3651 6783
rect 3651 6749 3660 6783
rect 3608 6740 3660 6749
rect 3976 6783 4028 6792
rect 3976 6749 3985 6783
rect 3985 6749 4019 6783
rect 4019 6749 4028 6783
rect 3976 6740 4028 6749
rect 4988 6740 5040 6792
rect 2228 6672 2280 6724
rect 2044 6604 2096 6656
rect 2688 6604 2740 6656
rect 3516 6604 3568 6656
rect 3792 6604 3844 6656
rect 6092 6672 6144 6724
rect 4988 6604 5040 6656
rect 8300 6953 8309 6987
rect 8309 6953 8343 6987
rect 8343 6953 8352 6987
rect 8300 6944 8352 6953
rect 8484 6876 8536 6928
rect 9220 6808 9272 6860
rect 9956 6808 10008 6860
rect 15200 6876 15252 6928
rect 6276 6604 6328 6656
rect 8668 6740 8720 6792
rect 6920 6672 6972 6724
rect 7288 6672 7340 6724
rect 8208 6672 8260 6724
rect 6736 6604 6788 6656
rect 9220 6647 9272 6656
rect 9220 6613 9229 6647
rect 9229 6613 9263 6647
rect 9263 6613 9272 6647
rect 9220 6604 9272 6613
rect 4116 6502 4168 6554
rect 4180 6502 4232 6554
rect 4244 6502 4296 6554
rect 4308 6502 4360 6554
rect 4372 6502 4424 6554
rect 7216 6502 7268 6554
rect 7280 6502 7332 6554
rect 7344 6502 7396 6554
rect 7408 6502 7460 6554
rect 7472 6502 7524 6554
rect 1400 6400 1452 6452
rect 1584 6443 1636 6452
rect 1584 6409 1593 6443
rect 1593 6409 1627 6443
rect 1627 6409 1636 6443
rect 1584 6400 1636 6409
rect 4896 6400 4948 6452
rect 2688 6375 2740 6384
rect 2688 6341 2697 6375
rect 2697 6341 2731 6375
rect 2731 6341 2740 6375
rect 2688 6332 2740 6341
rect 2964 6332 3016 6384
rect 3976 6332 4028 6384
rect 1768 6307 1820 6316
rect 1768 6273 1777 6307
rect 1777 6273 1811 6307
rect 1811 6273 1820 6307
rect 1768 6264 1820 6273
rect 1952 6264 2004 6316
rect 2136 6307 2188 6316
rect 2136 6273 2145 6307
rect 2145 6273 2179 6307
rect 2179 6273 2188 6307
rect 2136 6264 2188 6273
rect 4620 6264 4672 6316
rect 5908 6264 5960 6316
rect 7104 6400 7156 6452
rect 7840 6400 7892 6452
rect 8208 6400 8260 6452
rect 6736 6264 6788 6316
rect 8760 6307 8812 6316
rect 8760 6273 8769 6307
rect 8769 6273 8803 6307
rect 8803 6273 8812 6307
rect 8760 6264 8812 6273
rect 1676 6196 1728 6248
rect 2412 6239 2464 6248
rect 2412 6205 2421 6239
rect 2421 6205 2455 6239
rect 2455 6205 2464 6239
rect 2412 6196 2464 6205
rect 3056 6196 3108 6248
rect 2136 6060 2188 6112
rect 5540 6128 5592 6180
rect 6552 6128 6604 6180
rect 4712 6060 4764 6112
rect 4988 6103 5040 6112
rect 4988 6069 4997 6103
rect 4997 6069 5031 6103
rect 5031 6069 5040 6103
rect 4988 6060 5040 6069
rect 6092 6060 6144 6112
rect 8208 6128 8260 6180
rect 8484 6060 8536 6112
rect 9312 6060 9364 6112
rect 2566 5958 2618 6010
rect 2630 5958 2682 6010
rect 2694 5958 2746 6010
rect 2758 5958 2810 6010
rect 2822 5958 2874 6010
rect 5666 5958 5718 6010
rect 5730 5958 5782 6010
rect 5794 5958 5846 6010
rect 5858 5958 5910 6010
rect 5922 5958 5974 6010
rect 8766 5958 8818 6010
rect 8830 5958 8882 6010
rect 8894 5958 8946 6010
rect 8958 5958 9010 6010
rect 9022 5958 9074 6010
rect 1492 5856 1544 5908
rect 1952 5899 2004 5908
rect 1952 5865 1961 5899
rect 1961 5865 1995 5899
rect 1995 5865 2004 5899
rect 1952 5856 2004 5865
rect 2228 5899 2280 5908
rect 2228 5865 2237 5899
rect 2237 5865 2271 5899
rect 2271 5865 2280 5899
rect 2228 5856 2280 5865
rect 3056 5856 3108 5908
rect 3792 5899 3844 5908
rect 1124 5788 1176 5840
rect 1768 5788 1820 5840
rect 2964 5788 3016 5840
rect 3792 5865 3801 5899
rect 3801 5865 3835 5899
rect 3835 5865 3844 5899
rect 3792 5856 3844 5865
rect 3976 5856 4028 5908
rect 4988 5856 5040 5908
rect 5540 5856 5592 5908
rect 8208 5856 8260 5908
rect 9128 5856 9180 5908
rect 940 5652 992 5704
rect 1676 5652 1728 5704
rect 2044 5695 2096 5704
rect 2044 5661 2053 5695
rect 2053 5661 2087 5695
rect 2087 5661 2096 5695
rect 2044 5652 2096 5661
rect 2136 5652 2188 5704
rect 4160 5788 4212 5840
rect 6828 5831 6880 5840
rect 2872 5648 2924 5700
rect 6828 5797 6837 5831
rect 6837 5797 6871 5831
rect 6871 5797 6880 5831
rect 6828 5788 6880 5797
rect 6276 5720 6328 5772
rect 8576 5763 8628 5772
rect 8576 5729 8585 5763
rect 8585 5729 8619 5763
rect 8619 5729 8628 5763
rect 8576 5720 8628 5729
rect 3608 5652 3660 5704
rect 4252 5695 4304 5704
rect 4252 5661 4261 5695
rect 4261 5661 4295 5695
rect 4295 5661 4304 5695
rect 4252 5652 4304 5661
rect 5908 5652 5960 5704
rect 9404 5695 9456 5704
rect 5540 5584 5592 5636
rect 5816 5584 5868 5636
rect 6092 5584 6144 5636
rect 1768 5516 1820 5568
rect 2872 5516 2924 5568
rect 3148 5516 3200 5568
rect 6552 5516 6604 5568
rect 9404 5661 9413 5695
rect 9413 5661 9447 5695
rect 9447 5661 9456 5695
rect 9404 5652 9456 5661
rect 7012 5584 7064 5636
rect 8300 5627 8352 5636
rect 8300 5593 8309 5627
rect 8309 5593 8343 5627
rect 8343 5593 8352 5627
rect 8300 5584 8352 5593
rect 8024 5516 8076 5568
rect 4116 5414 4168 5466
rect 4180 5414 4232 5466
rect 4244 5414 4296 5466
rect 4308 5414 4360 5466
rect 4372 5414 4424 5466
rect 7216 5414 7268 5466
rect 7280 5414 7332 5466
rect 7344 5414 7396 5466
rect 7408 5414 7460 5466
rect 7472 5414 7524 5466
rect 1860 5312 1912 5364
rect 2596 5312 2648 5364
rect 1216 5244 1268 5296
rect 2412 5244 2464 5296
rect 4620 5312 4672 5364
rect 5080 5355 5132 5364
rect 5080 5321 5089 5355
rect 5089 5321 5123 5355
rect 5123 5321 5132 5355
rect 5080 5312 5132 5321
rect 7748 5312 7800 5364
rect 7932 5312 7984 5364
rect 3332 5219 3384 5228
rect 3332 5185 3341 5219
rect 3341 5185 3375 5219
rect 3375 5185 3384 5219
rect 3332 5176 3384 5185
rect 8024 5244 8076 5296
rect 9128 5244 9180 5296
rect 9312 5244 9364 5296
rect 5540 5219 5592 5228
rect 2964 5108 3016 5160
rect 3608 5108 3660 5160
rect 4068 5108 4120 5160
rect 3332 4972 3384 5024
rect 5540 5185 5549 5219
rect 5549 5185 5583 5219
rect 5583 5185 5592 5219
rect 5540 5176 5592 5185
rect 6000 5176 6052 5228
rect 7748 5176 7800 5228
rect 5908 5108 5960 5160
rect 9404 5176 9456 5228
rect 8668 5151 8720 5160
rect 8668 5117 8677 5151
rect 8677 5117 8711 5151
rect 8711 5117 8720 5151
rect 8668 5108 8720 5117
rect 9588 5108 9640 5160
rect 5540 5040 5592 5092
rect 16580 5040 16632 5092
rect 7104 4972 7156 5024
rect 9312 5015 9364 5024
rect 9312 4981 9321 5015
rect 9321 4981 9355 5015
rect 9355 4981 9364 5015
rect 9312 4972 9364 4981
rect 2780 4947 2832 4956
rect 2780 4913 2789 4947
rect 2789 4913 2823 4947
rect 2823 4913 2832 4947
rect 2780 4904 2832 4913
rect 5666 4870 5718 4922
rect 5730 4870 5782 4922
rect 5794 4870 5846 4922
rect 5858 4870 5910 4922
rect 5922 4870 5974 4922
rect 8766 4870 8818 4922
rect 8830 4870 8882 4922
rect 8894 4870 8946 4922
rect 8958 4870 9010 4922
rect 9022 4870 9074 4922
rect 2780 4768 2832 4820
rect 3424 4768 3476 4820
rect 3792 4811 3844 4820
rect 3792 4777 3801 4811
rect 3801 4777 3835 4811
rect 3835 4777 3844 4811
rect 4436 4811 4488 4820
rect 3792 4768 3844 4777
rect 4436 4777 4445 4811
rect 4445 4777 4479 4811
rect 4479 4777 4488 4811
rect 4436 4768 4488 4777
rect 8484 4768 8536 4820
rect 11060 4700 11112 4752
rect 17776 4700 17828 4752
rect 20628 4700 20680 4752
rect 2688 4675 2740 4684
rect 2688 4641 2697 4675
rect 2697 4641 2731 4675
rect 2731 4641 2740 4675
rect 2688 4632 2740 4641
rect 4436 4632 4488 4684
rect 6276 4675 6328 4684
rect 3424 4607 3476 4616
rect 3424 4573 3433 4607
rect 3433 4573 3467 4607
rect 3467 4573 3476 4607
rect 3424 4564 3476 4573
rect 1032 4496 1084 4548
rect 2688 4496 2740 4548
rect 3148 4496 3200 4548
rect 4068 4564 4120 4616
rect 5080 4564 5132 4616
rect 4712 4496 4764 4548
rect 4988 4496 5040 4548
rect 6276 4641 6285 4675
rect 6285 4641 6319 4675
rect 6319 4641 6328 4675
rect 6276 4632 6328 4641
rect 6552 4675 6604 4684
rect 6552 4641 6561 4675
rect 6561 4641 6595 4675
rect 6595 4641 6604 4675
rect 6552 4632 6604 4641
rect 6276 4496 6328 4548
rect 7104 4496 7156 4548
rect 3608 4471 3660 4480
rect 3608 4437 3617 4471
rect 3617 4437 3651 4471
rect 3651 4437 3660 4471
rect 3608 4428 3660 4437
rect 3792 4428 3844 4480
rect 4804 4471 4856 4480
rect 4804 4437 4813 4471
rect 4813 4437 4847 4471
rect 4847 4437 4856 4471
rect 4804 4428 4856 4437
rect 6092 4471 6144 4480
rect 6092 4437 6101 4471
rect 6101 4437 6135 4471
rect 6135 4437 6144 4471
rect 6092 4428 6144 4437
rect 7840 4428 7892 4480
rect 4116 4326 4168 4378
rect 4180 4326 4232 4378
rect 4244 4326 4296 4378
rect 4308 4326 4360 4378
rect 4372 4326 4424 4378
rect 7216 4326 7268 4378
rect 7280 4326 7332 4378
rect 7344 4326 7396 4378
rect 7408 4326 7460 4378
rect 7472 4326 7524 4378
rect 4988 4224 5040 4276
rect 9496 4224 9548 4276
rect 4344 4156 4396 4208
rect 8208 4156 8260 4208
rect 3608 4131 3660 4140
rect 3608 4097 3617 4131
rect 3617 4097 3651 4131
rect 3651 4097 3660 4131
rect 3608 4088 3660 4097
rect 3976 4131 4028 4140
rect 3976 4097 3985 4131
rect 3985 4097 4019 4131
rect 4019 4097 4028 4131
rect 3976 4088 4028 4097
rect 4988 4088 5040 4140
rect 6552 4088 6604 4140
rect 6828 4131 6880 4140
rect 6828 4097 6837 4131
rect 6837 4097 6871 4131
rect 6871 4097 6880 4131
rect 6828 4088 6880 4097
rect 6920 4088 6972 4140
rect 8576 4131 8628 4140
rect 8576 4097 8585 4131
rect 8585 4097 8619 4131
rect 8619 4097 8628 4131
rect 8576 4088 8628 4097
rect 3700 4020 3752 4072
rect 3608 3884 3660 3936
rect 6000 4020 6052 4072
rect 7104 4020 7156 4072
rect 7656 4063 7708 4072
rect 7656 4029 7665 4063
rect 7665 4029 7699 4063
rect 7699 4029 7708 4063
rect 7656 4020 7708 4029
rect 8300 4020 8352 4072
rect 9404 4020 9456 4072
rect 6276 3952 6328 4004
rect 7196 3952 7248 4004
rect 6552 3884 6604 3936
rect 6736 3927 6788 3936
rect 6736 3893 6745 3927
rect 6745 3893 6779 3927
rect 6779 3893 6788 3927
rect 6736 3884 6788 3893
rect 6920 3884 6972 3936
rect 7656 3884 7708 3936
rect 9220 3884 9272 3936
rect 5666 3782 5718 3834
rect 5730 3782 5782 3834
rect 5794 3782 5846 3834
rect 5858 3782 5910 3834
rect 5922 3782 5974 3834
rect 8766 3782 8818 3834
rect 8830 3782 8882 3834
rect 8894 3782 8946 3834
rect 8958 3782 9010 3834
rect 9022 3782 9074 3834
rect 3424 3680 3476 3732
rect 4344 3680 4396 3732
rect 5172 3723 5224 3732
rect 5172 3689 5181 3723
rect 5181 3689 5215 3723
rect 5215 3689 5224 3723
rect 5172 3680 5224 3689
rect 6276 3723 6328 3732
rect 3608 3612 3660 3664
rect 3700 3612 3752 3664
rect 3792 3544 3844 3596
rect 3424 3476 3476 3528
rect 3976 3476 4028 3528
rect 4528 3544 4580 3596
rect 6000 3612 6052 3664
rect 6276 3689 6285 3723
rect 6285 3689 6319 3723
rect 6319 3689 6328 3723
rect 6276 3680 6328 3689
rect 6552 3680 6604 3732
rect 8300 3680 8352 3732
rect 8576 3680 8628 3732
rect 9220 3723 9272 3732
rect 9220 3689 9229 3723
rect 9229 3689 9263 3723
rect 9263 3689 9272 3723
rect 9220 3680 9272 3689
rect 16580 3680 16632 3732
rect 4804 3476 4856 3528
rect 5632 3476 5684 3528
rect 6092 3544 6144 3596
rect 6276 3476 6328 3528
rect 6552 3519 6604 3528
rect 6552 3485 6561 3519
rect 6561 3485 6595 3519
rect 6595 3485 6604 3519
rect 6552 3476 6604 3485
rect 8392 3612 8444 3664
rect 6920 3587 6972 3596
rect 6920 3553 6929 3587
rect 6929 3553 6963 3587
rect 6963 3553 6972 3587
rect 6920 3544 6972 3553
rect 7380 3544 7432 3596
rect 8392 3519 8444 3528
rect 8392 3485 8401 3519
rect 8401 3485 8435 3519
rect 8435 3485 8444 3519
rect 8392 3476 8444 3485
rect 9404 3612 9456 3664
rect 8576 3544 8628 3596
rect 8852 3544 8904 3596
rect 9956 3544 10008 3596
rect 8760 3476 8812 3528
rect 4620 3408 4672 3460
rect 3516 3340 3568 3392
rect 3700 3340 3752 3392
rect 4988 3340 5040 3392
rect 6000 3340 6052 3392
rect 6736 3340 6788 3392
rect 6920 3340 6972 3392
rect 7932 3340 7984 3392
rect 13820 3408 13872 3460
rect 9036 3340 9088 3392
rect 9496 3340 9548 3392
rect 4116 3238 4168 3290
rect 4180 3238 4232 3290
rect 4244 3238 4296 3290
rect 4308 3238 4360 3290
rect 4372 3238 4424 3290
rect 7216 3238 7268 3290
rect 7280 3238 7332 3290
rect 7344 3238 7396 3290
rect 7408 3238 7460 3290
rect 7472 3238 7524 3290
rect 3332 3136 3384 3188
rect 3884 3136 3936 3188
rect 3424 3068 3476 3120
rect 4620 3136 4672 3188
rect 6828 3179 6880 3188
rect 6828 3145 6837 3179
rect 6837 3145 6871 3179
rect 6871 3145 6880 3179
rect 6828 3136 6880 3145
rect 8208 3136 8260 3188
rect 8576 3136 8628 3188
rect 9036 3179 9088 3188
rect 9036 3145 9045 3179
rect 9045 3145 9079 3179
rect 9079 3145 9088 3179
rect 9036 3136 9088 3145
rect 5172 3068 5224 3120
rect 6092 3068 6144 3120
rect 6276 3068 6328 3120
rect 7656 3068 7708 3120
rect 9220 3068 9272 3120
rect 2780 2864 2832 2916
rect 4528 3000 4580 3052
rect 4712 3043 4764 3052
rect 4712 3009 4721 3043
rect 4721 3009 4755 3043
rect 4755 3009 4764 3043
rect 4712 3000 4764 3009
rect 6000 3000 6052 3052
rect 7012 3000 7064 3052
rect 8116 3000 8168 3052
rect 4896 2932 4948 2984
rect 6276 2932 6328 2984
rect 8852 3000 8904 3052
rect 9680 3000 9732 3052
rect 3884 2796 3936 2848
rect 4068 2796 4120 2848
rect 5264 2796 5316 2848
rect 7656 2796 7708 2848
rect 8208 2796 8260 2848
rect 9220 2975 9272 2984
rect 9220 2941 9229 2975
rect 9229 2941 9263 2975
rect 9263 2941 9272 2975
rect 9220 2932 9272 2941
rect 16580 2796 16632 2848
rect 5666 2694 5718 2746
rect 5730 2694 5782 2746
rect 5794 2694 5846 2746
rect 5858 2694 5910 2746
rect 5922 2694 5974 2746
rect 8766 2694 8818 2746
rect 8830 2694 8882 2746
rect 8894 2694 8946 2746
rect 8958 2694 9010 2746
rect 9022 2694 9074 2746
rect 2688 2592 2740 2644
rect 3424 2592 3476 2644
rect 3700 2592 3752 2644
rect 3976 2592 4028 2644
rect 5540 2592 5592 2644
rect 3240 2524 3292 2576
rect 4068 2567 4120 2576
rect 4068 2533 4077 2567
rect 4077 2533 4111 2567
rect 4111 2533 4120 2567
rect 4068 2524 4120 2533
rect 4528 2524 4580 2576
rect 6092 2592 6144 2644
rect 6552 2592 6604 2644
rect 6920 2635 6972 2644
rect 6920 2601 6929 2635
rect 6929 2601 6963 2635
rect 6963 2601 6972 2635
rect 6920 2592 6972 2601
rect 7104 2635 7156 2644
rect 7104 2601 7113 2635
rect 7113 2601 7147 2635
rect 7147 2601 7156 2635
rect 7104 2592 7156 2601
rect 7932 2592 7984 2644
rect 2688 2456 2740 2508
rect 3332 2431 3384 2440
rect 3332 2397 3341 2431
rect 3341 2397 3375 2431
rect 3375 2397 3384 2431
rect 3332 2388 3384 2397
rect 3424 2388 3476 2440
rect 3792 2431 3844 2440
rect 3792 2397 3801 2431
rect 3801 2397 3835 2431
rect 3835 2397 3844 2431
rect 3792 2388 3844 2397
rect 3976 2388 4028 2440
rect 4528 2388 4580 2440
rect 4712 2388 4764 2440
rect 5172 2388 5224 2440
rect 7748 2524 7800 2576
rect 8852 2524 8904 2576
rect 6828 2456 6880 2508
rect 6736 2431 6788 2440
rect 6736 2397 6745 2431
rect 6745 2397 6779 2431
rect 6779 2397 6788 2431
rect 6736 2388 6788 2397
rect 7196 2431 7248 2440
rect 7196 2397 7205 2431
rect 7205 2397 7239 2431
rect 7239 2397 7248 2431
rect 7196 2388 7248 2397
rect 7380 2456 7432 2508
rect 7840 2388 7892 2440
rect 7932 2431 7984 2440
rect 7932 2397 7941 2431
rect 7941 2397 7975 2431
rect 7975 2397 7984 2431
rect 9036 2456 9088 2508
rect 17776 2456 17828 2508
rect 7932 2388 7984 2397
rect 7656 2320 7708 2372
rect 9404 2388 9456 2440
rect 9864 2388 9916 2440
rect 7840 2252 7892 2304
rect 8024 2252 8076 2304
rect 8944 2252 8996 2304
rect 4116 2150 4168 2202
rect 4180 2150 4232 2202
rect 4244 2150 4296 2202
rect 4308 2150 4360 2202
rect 4372 2150 4424 2202
rect 7216 2150 7268 2202
rect 7280 2150 7332 2202
rect 7344 2150 7396 2202
rect 7408 2150 7460 2202
rect 7472 2150 7524 2202
rect 2964 2048 3016 2100
rect 3884 2048 3936 2100
rect 3056 1980 3108 2032
rect 5172 2048 5224 2100
rect 6460 2048 6512 2100
rect 4896 2023 4948 2032
rect 4896 1989 4905 2023
rect 4905 1989 4939 2023
rect 4939 1989 4948 2023
rect 4896 1980 4948 1989
rect 6276 1980 6328 2032
rect 2688 1912 2740 1964
rect 3424 1912 3476 1964
rect 3516 1912 3568 1964
rect 3884 1955 3936 1964
rect 3884 1921 3893 1955
rect 3893 1921 3927 1955
rect 3927 1921 3936 1955
rect 3884 1912 3936 1921
rect 6184 1912 6236 1964
rect 7748 2048 7800 2100
rect 7840 2091 7892 2100
rect 7840 2057 7849 2091
rect 7849 2057 7883 2091
rect 7883 2057 7892 2091
rect 8116 2091 8168 2100
rect 7840 2048 7892 2057
rect 8116 2057 8125 2091
rect 8125 2057 8159 2091
rect 8159 2057 8168 2091
rect 8116 2048 8168 2057
rect 8484 2048 8536 2100
rect 9220 2048 9272 2100
rect 8208 1980 8260 2032
rect 4528 1844 4580 1896
rect 4988 1844 5040 1896
rect 8300 1912 8352 1964
rect 8944 1912 8996 1964
rect 8484 1844 8536 1896
rect 8576 1844 8628 1896
rect 3148 1776 3200 1828
rect 4252 1708 4304 1760
rect 4712 1708 4764 1760
rect 6368 1708 6420 1760
rect 8392 1708 8444 1760
rect 16580 1776 16632 1828
rect 21364 1708 21416 1760
rect 5666 1606 5718 1658
rect 5730 1606 5782 1658
rect 5794 1606 5846 1658
rect 5858 1606 5910 1658
rect 5922 1606 5974 1658
rect 8766 1606 8818 1658
rect 8830 1606 8882 1658
rect 8894 1606 8946 1658
rect 8958 1606 9010 1658
rect 9022 1606 9074 1658
rect 1032 1504 1084 1556
rect 3424 1504 3476 1556
rect 4068 1504 4120 1556
rect 4252 1504 4304 1556
rect 5080 1504 5132 1556
rect 8484 1504 8536 1556
rect 9128 1504 9180 1556
rect 3332 1436 3384 1488
rect 3516 1368 3568 1420
rect 7932 1436 7984 1488
rect 8944 1436 8996 1488
rect 9220 1368 9272 1420
rect 7564 1300 7616 1352
rect 9496 1343 9548 1352
rect 9496 1309 9505 1343
rect 9505 1309 9539 1343
rect 9539 1309 9548 1343
rect 9496 1300 9548 1309
rect 13820 1300 13872 1352
rect 10876 1232 10928 1284
rect 3792 1207 3844 1216
rect 3792 1173 3801 1207
rect 3801 1173 3835 1207
rect 3835 1173 3844 1207
rect 3792 1164 3844 1173
rect 3884 1164 3936 1216
rect 8668 1164 8720 1216
rect 8944 1207 8996 1216
rect 8944 1173 8953 1207
rect 8953 1173 8987 1207
rect 8987 1173 8996 1207
rect 8944 1164 8996 1173
rect 9588 1164 9640 1216
rect 4116 1062 4168 1114
rect 4180 1062 4232 1114
rect 4244 1062 4296 1114
rect 4308 1062 4360 1114
rect 4372 1062 4424 1114
rect 7216 1062 7268 1114
rect 7280 1062 7332 1114
rect 7344 1062 7396 1114
rect 7408 1062 7460 1114
rect 7472 1062 7524 1114
<< metal2 >>
rect 938 12200 994 13000
rect 1398 12200 1454 13000
rect 1858 12200 1914 13000
rect 2318 12200 2374 13000
rect 2778 12200 2834 13000
rect 3238 12200 3294 13000
rect 3698 12200 3754 13000
rect 4158 12200 4214 13000
rect 4618 12200 4674 13000
rect 5078 12200 5134 13000
rect 5538 12200 5594 13000
rect 5998 12200 6054 13000
rect 6458 12200 6514 13000
rect 16578 12336 16634 12345
rect 16578 12271 16634 12280
rect 846 7848 902 7857
rect 846 7783 902 7792
rect 860 4154 888 7783
rect 952 7002 980 12200
rect 1308 11620 1360 11626
rect 1308 11562 1360 11568
rect 1320 11150 1348 11562
rect 1308 11144 1360 11150
rect 1308 11086 1360 11092
rect 1412 11054 1440 12200
rect 1492 11756 1544 11762
rect 1492 11698 1544 11704
rect 1504 11354 1532 11698
rect 1872 11506 1900 12200
rect 2332 12170 2360 12200
rect 1952 12164 2004 12170
rect 1952 12106 2004 12112
rect 2320 12164 2372 12170
rect 2320 12106 2372 12112
rect 1780 11478 1900 11506
rect 1492 11348 1544 11354
rect 1492 11290 1544 11296
rect 1780 11054 1808 11478
rect 1964 11370 1992 12106
rect 2320 12028 2372 12034
rect 2792 12016 2820 12200
rect 2792 11988 3188 12016
rect 2320 11970 2372 11976
rect 2228 11688 2280 11694
rect 2228 11630 2280 11636
rect 1044 11026 1440 11054
rect 1688 11026 1808 11054
rect 1872 11342 1992 11370
rect 2240 11354 2268 11630
rect 2332 11354 2360 11970
rect 2412 11892 2464 11898
rect 2412 11834 2464 11840
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2228 11348 2280 11354
rect 940 6996 992 7002
rect 940 6938 992 6944
rect 952 5710 980 6938
rect 940 5704 992 5710
rect 940 5646 992 5652
rect 1044 4554 1072 11026
rect 1122 10976 1178 10985
rect 1122 10911 1178 10920
rect 1136 5846 1164 10911
rect 1398 10840 1454 10849
rect 1398 10775 1454 10784
rect 1492 10804 1544 10810
rect 1412 10146 1440 10775
rect 1492 10746 1544 10752
rect 1504 10713 1532 10746
rect 1490 10704 1546 10713
rect 1490 10639 1546 10648
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 1596 10577 1624 10610
rect 1582 10568 1638 10577
rect 1582 10503 1638 10512
rect 1412 10118 1532 10146
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1308 9580 1360 9586
rect 1308 9522 1360 9528
rect 1216 8968 1268 8974
rect 1216 8910 1268 8916
rect 1124 5840 1176 5846
rect 1124 5782 1176 5788
rect 1228 5302 1256 8910
rect 1320 8090 1348 9522
rect 1308 8084 1360 8090
rect 1308 8026 1360 8032
rect 1320 7886 1348 8026
rect 1308 7880 1360 7886
rect 1308 7822 1360 7828
rect 1320 7274 1348 7822
rect 1308 7268 1360 7274
rect 1308 7210 1360 7216
rect 1412 6458 1440 9998
rect 1504 9178 1532 10118
rect 1584 9920 1636 9926
rect 1584 9862 1636 9868
rect 1492 9172 1544 9178
rect 1492 9114 1544 9120
rect 1596 8650 1624 9862
rect 1688 8906 1716 11026
rect 1872 11014 1900 11342
rect 2228 11290 2280 11296
rect 2320 11348 2372 11354
rect 2320 11290 2372 11296
rect 1952 11280 2004 11286
rect 1952 11222 2004 11228
rect 1860 11008 1912 11014
rect 1860 10950 1912 10956
rect 1964 10826 1992 11222
rect 2424 11150 2452 11834
rect 2566 11452 2874 11472
rect 2566 11450 2572 11452
rect 2628 11450 2652 11452
rect 2708 11450 2732 11452
rect 2788 11450 2812 11452
rect 2868 11450 2874 11452
rect 2628 11398 2630 11450
rect 2810 11398 2812 11450
rect 2566 11396 2572 11398
rect 2628 11396 2652 11398
rect 2708 11396 2732 11398
rect 2788 11396 2812 11398
rect 2868 11396 2874 11398
rect 2566 11376 2874 11396
rect 2976 11354 3004 11834
rect 2964 11348 3016 11354
rect 2964 11290 3016 11296
rect 2686 11248 2742 11257
rect 2686 11183 2742 11192
rect 2700 11150 2728 11183
rect 2044 11144 2096 11150
rect 2044 11086 2096 11092
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 2412 11144 2464 11150
rect 2412 11086 2464 11092
rect 2688 11144 2740 11150
rect 2688 11086 2740 11092
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 1780 10798 1992 10826
rect 1780 9081 1808 10798
rect 1952 10668 2004 10674
rect 1952 10610 2004 10616
rect 1860 9920 1912 9926
rect 1860 9862 1912 9868
rect 1872 9586 1900 9862
rect 1964 9722 1992 10610
rect 2056 9722 2084 11086
rect 2136 11008 2188 11014
rect 2136 10950 2188 10956
rect 1952 9716 2004 9722
rect 1952 9658 2004 9664
rect 2044 9716 2096 9722
rect 2044 9658 2096 9664
rect 1860 9580 1912 9586
rect 1860 9522 1912 9528
rect 1766 9072 1822 9081
rect 1766 9007 1822 9016
rect 1676 8900 1728 8906
rect 1676 8842 1728 8848
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 1596 8622 1716 8650
rect 1780 8634 1808 8774
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1492 8288 1544 8294
rect 1492 8230 1544 8236
rect 1504 7342 1532 8230
rect 1492 7336 1544 7342
rect 1492 7278 1544 7284
rect 1490 7168 1546 7177
rect 1490 7103 1546 7112
rect 1400 6452 1452 6458
rect 1400 6394 1452 6400
rect 1504 5914 1532 7103
rect 1596 6458 1624 8434
rect 1688 7954 1716 8622
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 1872 8566 1900 9522
rect 2044 8968 2096 8974
rect 2044 8910 2096 8916
rect 1860 8560 1912 8566
rect 1860 8502 1912 8508
rect 2056 8401 2084 8910
rect 2042 8392 2098 8401
rect 2042 8327 2098 8336
rect 1768 8288 1820 8294
rect 2148 8276 2176 10950
rect 2240 10810 2268 11086
rect 2976 11014 3004 11086
rect 2412 11008 2464 11014
rect 2412 10950 2464 10956
rect 2964 11008 3016 11014
rect 2964 10950 3016 10956
rect 2228 10804 2280 10810
rect 2228 10746 2280 10752
rect 2228 10668 2280 10674
rect 2228 10610 2280 10616
rect 2240 9382 2268 10610
rect 2424 10130 2452 10950
rect 3056 10804 3108 10810
rect 3056 10746 3108 10752
rect 2872 10668 2924 10674
rect 2872 10610 2924 10616
rect 2884 10538 2912 10610
rect 2872 10532 2924 10538
rect 2872 10474 2924 10480
rect 2964 10532 3016 10538
rect 2964 10474 3016 10480
rect 2566 10364 2874 10384
rect 2566 10362 2572 10364
rect 2628 10362 2652 10364
rect 2708 10362 2732 10364
rect 2788 10362 2812 10364
rect 2868 10362 2874 10364
rect 2628 10310 2630 10362
rect 2810 10310 2812 10362
rect 2566 10308 2572 10310
rect 2628 10308 2652 10310
rect 2708 10308 2732 10310
rect 2788 10308 2812 10310
rect 2868 10308 2874 10310
rect 2566 10288 2874 10308
rect 2412 10124 2464 10130
rect 2412 10066 2464 10072
rect 2686 10024 2742 10033
rect 2686 9959 2688 9968
rect 2740 9959 2742 9968
rect 2688 9930 2740 9936
rect 2596 9716 2648 9722
rect 2596 9658 2648 9664
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 2228 9376 2280 9382
rect 2228 9318 2280 9324
rect 2332 9178 2360 9454
rect 2608 9450 2636 9658
rect 2596 9444 2648 9450
rect 2596 9386 2648 9392
rect 2566 9276 2874 9296
rect 2566 9274 2572 9276
rect 2628 9274 2652 9276
rect 2708 9274 2732 9276
rect 2788 9274 2812 9276
rect 2868 9274 2874 9276
rect 2628 9222 2630 9274
rect 2810 9222 2812 9274
rect 2566 9220 2572 9222
rect 2628 9220 2652 9222
rect 2708 9220 2732 9222
rect 2788 9220 2812 9222
rect 2868 9220 2874 9222
rect 2566 9200 2874 9220
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 2686 9072 2742 9081
rect 2686 9007 2742 9016
rect 2870 9072 2926 9081
rect 2870 9007 2926 9016
rect 2700 8974 2728 9007
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2320 8900 2372 8906
rect 2320 8842 2372 8848
rect 2504 8900 2556 8906
rect 2504 8842 2556 8848
rect 2228 8492 2280 8498
rect 2228 8434 2280 8440
rect 1768 8230 1820 8236
rect 1872 8248 2176 8276
rect 1676 7948 1728 7954
rect 1676 7890 1728 7896
rect 1780 7410 1808 8230
rect 1768 7404 1820 7410
rect 1768 7346 1820 7352
rect 1676 7200 1728 7206
rect 1676 7142 1728 7148
rect 1688 6798 1716 7142
rect 1768 6996 1820 7002
rect 1768 6938 1820 6944
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 1584 6452 1636 6458
rect 1584 6394 1636 6400
rect 1688 6254 1716 6734
rect 1780 6322 1808 6938
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 1492 5908 1544 5914
rect 1492 5850 1544 5856
rect 1768 5840 1820 5846
rect 1768 5782 1820 5788
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 1688 5545 1716 5646
rect 1780 5574 1808 5782
rect 1768 5568 1820 5574
rect 1674 5536 1730 5545
rect 1768 5510 1820 5516
rect 1674 5471 1730 5480
rect 1872 5370 1900 8248
rect 2240 7750 2268 8434
rect 2228 7744 2280 7750
rect 2228 7686 2280 7692
rect 2136 7268 2188 7274
rect 2136 7210 2188 7216
rect 1952 6860 2004 6866
rect 1952 6802 2004 6808
rect 1964 6322 1992 6802
rect 2044 6656 2096 6662
rect 2044 6598 2096 6604
rect 1952 6316 2004 6322
rect 1952 6258 2004 6264
rect 1950 6216 2006 6225
rect 1950 6151 2006 6160
rect 1964 5914 1992 6151
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 2056 5710 2084 6598
rect 2148 6322 2176 7210
rect 2240 6730 2268 7686
rect 2228 6724 2280 6730
rect 2228 6666 2280 6672
rect 2226 6352 2282 6361
rect 2136 6316 2188 6322
rect 2226 6287 2282 6296
rect 2136 6258 2188 6264
rect 2136 6112 2188 6118
rect 2136 6054 2188 6060
rect 2148 5710 2176 6054
rect 2240 5914 2268 6287
rect 2228 5908 2280 5914
rect 2228 5850 2280 5856
rect 2044 5704 2096 5710
rect 2044 5646 2096 5652
rect 2136 5704 2188 5710
rect 2136 5646 2188 5652
rect 2332 5522 2360 8842
rect 2516 8276 2544 8842
rect 2884 8786 2912 9007
rect 2976 8974 3004 10474
rect 3068 9518 3096 10746
rect 3056 9512 3108 9518
rect 3160 9489 3188 11988
rect 3056 9454 3108 9460
rect 3146 9480 3202 9489
rect 3146 9415 3202 9424
rect 3056 9376 3108 9382
rect 3252 9330 3280 12200
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 3516 11144 3568 11150
rect 3516 11086 3568 11092
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 3344 10033 3372 10746
rect 3330 10024 3386 10033
rect 3330 9959 3386 9968
rect 3332 9920 3384 9926
rect 3332 9862 3384 9868
rect 3056 9318 3108 9324
rect 3068 9110 3096 9318
rect 3160 9302 3280 9330
rect 3056 9104 3108 9110
rect 3056 9046 3108 9052
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 2884 8758 3004 8786
rect 2424 8248 2544 8276
rect 2424 7002 2452 8248
rect 2566 8188 2874 8208
rect 2566 8186 2572 8188
rect 2628 8186 2652 8188
rect 2708 8186 2732 8188
rect 2788 8186 2812 8188
rect 2868 8186 2874 8188
rect 2628 8134 2630 8186
rect 2810 8134 2812 8186
rect 2566 8132 2572 8134
rect 2628 8132 2652 8134
rect 2708 8132 2732 8134
rect 2788 8132 2812 8134
rect 2868 8132 2874 8134
rect 2566 8112 2874 8132
rect 2686 7984 2742 7993
rect 2686 7919 2742 7928
rect 2700 7818 2728 7919
rect 2688 7812 2740 7818
rect 2688 7754 2740 7760
rect 2566 7100 2874 7120
rect 2566 7098 2572 7100
rect 2628 7098 2652 7100
rect 2708 7098 2732 7100
rect 2788 7098 2812 7100
rect 2868 7098 2874 7100
rect 2628 7046 2630 7098
rect 2810 7046 2812 7098
rect 2566 7044 2572 7046
rect 2628 7044 2652 7046
rect 2708 7044 2732 7046
rect 2788 7044 2812 7046
rect 2868 7044 2874 7046
rect 2566 7024 2874 7044
rect 2412 6996 2464 7002
rect 2412 6938 2464 6944
rect 2976 6769 3004 8758
rect 3068 8090 3096 8910
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 3054 7984 3110 7993
rect 3054 7919 3110 7928
rect 3068 6798 3096 7919
rect 3056 6792 3108 6798
rect 2962 6760 3018 6769
rect 3056 6734 3108 6740
rect 2962 6695 3018 6704
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2700 6390 2728 6598
rect 3068 6474 3096 6734
rect 2976 6446 3096 6474
rect 2976 6390 3004 6446
rect 2688 6384 2740 6390
rect 2688 6326 2740 6332
rect 2964 6384 3016 6390
rect 2964 6326 3016 6332
rect 2412 6248 2464 6254
rect 2412 6190 2464 6196
rect 2424 5681 2452 6190
rect 2566 6012 2874 6032
rect 2566 6010 2572 6012
rect 2628 6010 2652 6012
rect 2708 6010 2732 6012
rect 2788 6010 2812 6012
rect 2868 6010 2874 6012
rect 2628 5958 2630 6010
rect 2810 5958 2812 6010
rect 2566 5956 2572 5958
rect 2628 5956 2652 5958
rect 2708 5956 2732 5958
rect 2788 5956 2812 5958
rect 2868 5956 2874 5958
rect 2566 5936 2874 5956
rect 2976 5846 3004 6326
rect 3056 6248 3108 6254
rect 3056 6190 3108 6196
rect 3068 5914 3096 6190
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 2964 5840 3016 5846
rect 2778 5808 2834 5817
rect 3160 5794 3188 9302
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 3252 7478 3280 9114
rect 3344 8294 3372 9862
rect 3436 9178 3464 11086
rect 3528 10810 3556 11086
rect 3608 11076 3660 11082
rect 3608 11018 3660 11024
rect 3516 10804 3568 10810
rect 3516 10746 3568 10752
rect 3620 10674 3648 11018
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 3608 10668 3660 10674
rect 3608 10610 3660 10616
rect 3528 9926 3556 10610
rect 3620 10062 3648 10610
rect 3608 10056 3660 10062
rect 3608 9998 3660 10004
rect 3516 9920 3568 9926
rect 3516 9862 3568 9868
rect 3606 9888 3662 9897
rect 3606 9823 3662 9832
rect 3620 9722 3648 9823
rect 3608 9716 3660 9722
rect 3608 9658 3660 9664
rect 3516 9648 3568 9654
rect 3712 9602 3740 12200
rect 4172 12102 4200 12200
rect 4160 12096 4212 12102
rect 4160 12038 4212 12044
rect 4344 11824 4396 11830
rect 4344 11766 4396 11772
rect 4356 11286 4384 11766
rect 4344 11280 4396 11286
rect 4344 11222 4396 11228
rect 3884 11144 3936 11150
rect 3804 11104 3884 11132
rect 3804 9722 3832 11104
rect 3884 11086 3936 11092
rect 4528 11144 4580 11150
rect 4528 11086 4580 11092
rect 3976 11076 4028 11082
rect 3976 11018 4028 11024
rect 3882 10976 3938 10985
rect 3882 10911 3938 10920
rect 3896 10305 3924 10911
rect 3988 10849 4016 11018
rect 4116 10908 4424 10928
rect 4116 10906 4122 10908
rect 4178 10906 4202 10908
rect 4258 10906 4282 10908
rect 4338 10906 4362 10908
rect 4418 10906 4424 10908
rect 4178 10854 4180 10906
rect 4360 10854 4362 10906
rect 4116 10852 4122 10854
rect 4178 10852 4202 10854
rect 4258 10852 4282 10854
rect 4338 10852 4362 10854
rect 4418 10852 4424 10854
rect 3974 10840 4030 10849
rect 4116 10832 4424 10852
rect 4540 10849 4568 11086
rect 4526 10840 4582 10849
rect 3974 10775 4030 10784
rect 4526 10775 4582 10784
rect 4252 10668 4304 10674
rect 4252 10610 4304 10616
rect 3976 10600 4028 10606
rect 3976 10542 4028 10548
rect 3882 10296 3938 10305
rect 3882 10231 3938 10240
rect 3988 10169 4016 10542
rect 3974 10160 4030 10169
rect 3974 10095 4030 10104
rect 3884 10056 3936 10062
rect 3884 9998 3936 10004
rect 3976 10056 4028 10062
rect 4264 10033 4292 10610
rect 4342 10568 4398 10577
rect 4342 10503 4344 10512
rect 4396 10503 4398 10512
rect 4344 10474 4396 10480
rect 4632 10169 4660 12200
rect 4712 11688 4764 11694
rect 4712 11630 4764 11636
rect 4724 10606 4752 11630
rect 4804 11280 4856 11286
rect 4804 11222 4856 11228
rect 5092 11234 5120 12200
rect 5356 12096 5408 12102
rect 5356 12038 5408 12044
rect 5264 11552 5316 11558
rect 5264 11494 5316 11500
rect 5276 11286 5304 11494
rect 5264 11280 5316 11286
rect 4712 10600 4764 10606
rect 4712 10542 4764 10548
rect 4816 10418 4844 11222
rect 5092 11206 5212 11234
rect 5264 11222 5316 11228
rect 5080 11144 5132 11150
rect 5078 11112 5080 11121
rect 5132 11112 5134 11121
rect 5078 11047 5134 11056
rect 5080 11008 5132 11014
rect 5080 10950 5132 10956
rect 4896 10668 4948 10674
rect 4896 10610 4948 10616
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 4724 10390 4844 10418
rect 4434 10160 4490 10169
rect 4434 10095 4490 10104
rect 4618 10160 4674 10169
rect 4618 10095 4674 10104
rect 4724 10112 4752 10390
rect 4802 10296 4858 10305
rect 4908 10282 4936 10610
rect 5000 10577 5028 10610
rect 4986 10568 5042 10577
rect 4986 10503 5042 10512
rect 4988 10464 5040 10470
rect 4988 10406 5040 10412
rect 4858 10254 4936 10282
rect 4802 10231 4858 10240
rect 3976 9998 4028 10004
rect 4250 10024 4306 10033
rect 3792 9716 3844 9722
rect 3792 9658 3844 9664
rect 3896 9602 3924 9998
rect 3516 9590 3568 9596
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3436 8906 3464 9114
rect 3528 9110 3556 9590
rect 3620 9574 3740 9602
rect 3804 9574 3924 9602
rect 3516 9104 3568 9110
rect 3516 9046 3568 9052
rect 3424 8900 3476 8906
rect 3424 8842 3476 8848
rect 3332 8288 3384 8294
rect 3332 8230 3384 8236
rect 3344 7868 3372 8230
rect 3424 7880 3476 7886
rect 3344 7840 3424 7868
rect 3240 7472 3292 7478
rect 3240 7414 3292 7420
rect 3238 7304 3294 7313
rect 3238 7239 3294 7248
rect 2964 5782 3016 5788
rect 2778 5743 2834 5752
rect 3068 5766 3188 5794
rect 2410 5672 2466 5681
rect 2410 5607 2466 5616
rect 2332 5494 2544 5522
rect 1860 5364 1912 5370
rect 1860 5306 1912 5312
rect 1216 5296 1268 5302
rect 1216 5238 1268 5244
rect 2412 5296 2464 5302
rect 2412 5238 2464 5244
rect 1032 4548 1084 4554
rect 1032 4490 1084 4496
rect 860 4126 1072 4154
rect 1044 1562 1072 4126
rect 2424 2553 2452 5238
rect 2410 2544 2466 2553
rect 2410 2479 2466 2488
rect 2516 1952 2544 5494
rect 2596 5364 2648 5370
rect 2596 5306 2648 5312
rect 2608 2496 2636 5306
rect 2686 5264 2742 5273
rect 2686 5199 2742 5208
rect 2700 4690 2728 5199
rect 2792 4962 2820 5743
rect 2872 5700 2924 5706
rect 2924 5648 3004 5658
rect 2872 5642 3004 5648
rect 2884 5630 3004 5642
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 2780 4956 2832 4962
rect 2780 4898 2832 4904
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 2688 4684 2740 4690
rect 2688 4626 2740 4632
rect 2688 4548 2740 4554
rect 2688 4490 2740 4496
rect 2700 2650 2728 4490
rect 2792 2922 2820 4762
rect 2884 3097 2912 5510
rect 2976 5166 3004 5630
rect 2964 5160 3016 5166
rect 2964 5102 3016 5108
rect 2870 3088 2926 3097
rect 2870 3023 2926 3032
rect 2780 2916 2832 2922
rect 2780 2858 2832 2864
rect 2688 2644 2740 2650
rect 2688 2586 2740 2592
rect 2688 2508 2740 2514
rect 2608 2468 2688 2496
rect 2688 2450 2740 2456
rect 2976 2106 3004 5102
rect 2964 2100 3016 2106
rect 2964 2042 3016 2048
rect 3068 2038 3096 5766
rect 3148 5568 3200 5574
rect 3146 5536 3148 5545
rect 3200 5536 3202 5545
rect 3146 5471 3202 5480
rect 3148 4548 3200 4554
rect 3148 4490 3200 4496
rect 3056 2032 3108 2038
rect 3056 1974 3108 1980
rect 2688 1964 2740 1970
rect 2516 1924 2688 1952
rect 2688 1906 2740 1912
rect 3160 1834 3188 4490
rect 3252 2582 3280 7239
rect 3344 5681 3372 7840
rect 3424 7822 3476 7828
rect 3516 7812 3568 7818
rect 3516 7754 3568 7760
rect 3424 7744 3476 7750
rect 3424 7686 3476 7692
rect 3330 5672 3386 5681
rect 3330 5607 3386 5616
rect 3344 5234 3372 5607
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 3332 5024 3384 5030
rect 3332 4966 3384 4972
rect 3344 3194 3372 4966
rect 3436 4826 3464 7686
rect 3528 6662 3556 7754
rect 3620 7562 3648 9574
rect 3700 9512 3752 9518
rect 3700 9454 3752 9460
rect 3712 9178 3740 9454
rect 3700 9172 3752 9178
rect 3700 9114 3752 9120
rect 3620 7534 3740 7562
rect 3608 6792 3660 6798
rect 3608 6734 3660 6740
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3620 6361 3648 6734
rect 3606 6352 3662 6361
rect 3606 6287 3662 6296
rect 3608 5704 3660 5710
rect 3608 5646 3660 5652
rect 3620 5166 3648 5646
rect 3608 5160 3660 5166
rect 3608 5102 3660 5108
rect 3424 4820 3476 4826
rect 3424 4762 3476 4768
rect 3514 4720 3570 4729
rect 3514 4655 3570 4664
rect 3424 4616 3476 4622
rect 3424 4558 3476 4564
rect 3436 3738 3464 4558
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3424 3528 3476 3534
rect 3424 3470 3476 3476
rect 3528 3482 3556 4655
rect 3608 4480 3660 4486
rect 3608 4422 3660 4428
rect 3620 4146 3648 4422
rect 3608 4140 3660 4146
rect 3608 4082 3660 4088
rect 3712 4078 3740 7534
rect 3804 7313 3832 9574
rect 3988 9110 4016 9998
rect 4448 9994 4476 10095
rect 4724 10084 4844 10112
rect 4250 9959 4306 9968
rect 4436 9988 4488 9994
rect 4436 9930 4488 9936
rect 4116 9820 4424 9840
rect 4116 9818 4122 9820
rect 4178 9818 4202 9820
rect 4258 9818 4282 9820
rect 4338 9818 4362 9820
rect 4418 9818 4424 9820
rect 4178 9766 4180 9818
rect 4360 9766 4362 9818
rect 4116 9764 4122 9766
rect 4178 9764 4202 9766
rect 4258 9764 4282 9766
rect 4338 9764 4362 9766
rect 4418 9764 4424 9766
rect 4116 9744 4424 9764
rect 4618 9752 4674 9761
rect 4618 9687 4674 9696
rect 4632 9636 4660 9687
rect 4540 9608 4660 9636
rect 4710 9616 4766 9625
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 4080 9382 4108 9522
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 3976 9104 4028 9110
rect 3976 9046 4028 9052
rect 4160 8968 4212 8974
rect 3988 8928 4160 8956
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 3790 7304 3846 7313
rect 3790 7239 3846 7248
rect 3896 6905 3924 8774
rect 3988 8294 4016 8928
rect 4160 8910 4212 8916
rect 4116 8732 4424 8752
rect 4116 8730 4122 8732
rect 4178 8730 4202 8732
rect 4258 8730 4282 8732
rect 4338 8730 4362 8732
rect 4418 8730 4424 8732
rect 4178 8678 4180 8730
rect 4360 8678 4362 8730
rect 4116 8676 4122 8678
rect 4178 8676 4202 8678
rect 4258 8676 4282 8678
rect 4338 8676 4362 8678
rect 4418 8676 4424 8678
rect 4116 8656 4424 8676
rect 4436 8560 4488 8566
rect 4342 8528 4398 8537
rect 4436 8502 4488 8508
rect 4342 8463 4398 8472
rect 4066 8392 4122 8401
rect 4066 8327 4122 8336
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 3988 8090 4016 8230
rect 4080 8090 4108 8327
rect 3976 8084 4028 8090
rect 3976 8026 4028 8032
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 4356 7886 4384 8463
rect 4448 8072 4476 8502
rect 4540 8294 4568 9608
rect 4710 9551 4766 9560
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4632 8974 4660 9318
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 4632 8401 4660 8774
rect 4618 8392 4674 8401
rect 4618 8327 4674 8336
rect 4528 8288 4580 8294
rect 4528 8230 4580 8236
rect 4528 8084 4580 8090
rect 4448 8044 4528 8072
rect 4528 8026 4580 8032
rect 4540 7993 4568 8026
rect 4526 7984 4582 7993
rect 4526 7919 4582 7928
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4620 7812 4672 7818
rect 4620 7754 4672 7760
rect 4528 7744 4580 7750
rect 4528 7686 4580 7692
rect 4116 7644 4424 7664
rect 4116 7642 4122 7644
rect 4178 7642 4202 7644
rect 4258 7642 4282 7644
rect 4338 7642 4362 7644
rect 4418 7642 4424 7644
rect 4178 7590 4180 7642
rect 4360 7590 4362 7642
rect 4116 7588 4122 7590
rect 4178 7588 4202 7590
rect 4258 7588 4282 7590
rect 4338 7588 4362 7590
rect 4418 7588 4424 7590
rect 4116 7568 4424 7588
rect 4344 7200 4396 7206
rect 4344 7142 4396 7148
rect 4356 7002 4384 7142
rect 4344 6996 4396 7002
rect 4344 6938 4396 6944
rect 3882 6896 3938 6905
rect 4540 6866 4568 7686
rect 3882 6831 3938 6840
rect 4528 6860 4580 6866
rect 4528 6802 4580 6808
rect 3976 6792 4028 6798
rect 3882 6760 3938 6769
rect 3976 6734 4028 6740
rect 3882 6695 3938 6704
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3804 6225 3832 6598
rect 3790 6216 3846 6225
rect 3790 6151 3846 6160
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 3804 4826 3832 5850
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 3792 4480 3844 4486
rect 3792 4422 3844 4428
rect 3700 4072 3752 4078
rect 3700 4014 3752 4020
rect 3608 3936 3660 3942
rect 3608 3878 3660 3884
rect 3620 3670 3648 3878
rect 3712 3670 3740 4014
rect 3608 3664 3660 3670
rect 3608 3606 3660 3612
rect 3700 3664 3752 3670
rect 3700 3606 3752 3612
rect 3804 3602 3832 4422
rect 3792 3596 3844 3602
rect 3792 3538 3844 3544
rect 3896 3482 3924 6695
rect 3988 6390 4016 6734
rect 4116 6556 4424 6576
rect 4116 6554 4122 6556
rect 4178 6554 4202 6556
rect 4258 6554 4282 6556
rect 4338 6554 4362 6556
rect 4418 6554 4424 6556
rect 4178 6502 4180 6554
rect 4360 6502 4362 6554
rect 4116 6500 4122 6502
rect 4178 6500 4202 6502
rect 4258 6500 4282 6502
rect 4338 6500 4362 6502
rect 4418 6500 4424 6502
rect 4116 6480 4424 6500
rect 3976 6384 4028 6390
rect 3976 6326 4028 6332
rect 4158 6352 4214 6361
rect 4158 6287 4214 6296
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 3988 4146 4016 5850
rect 4172 5846 4200 6287
rect 4160 5840 4212 5846
rect 4158 5808 4160 5817
rect 4212 5808 4214 5817
rect 4158 5743 4214 5752
rect 4252 5704 4304 5710
rect 4250 5672 4252 5681
rect 4304 5672 4306 5681
rect 4250 5607 4306 5616
rect 4116 5468 4424 5488
rect 4116 5466 4122 5468
rect 4178 5466 4202 5468
rect 4258 5466 4282 5468
rect 4338 5466 4362 5468
rect 4418 5466 4424 5468
rect 4178 5414 4180 5466
rect 4360 5414 4362 5466
rect 4116 5412 4122 5414
rect 4178 5412 4202 5414
rect 4258 5412 4282 5414
rect 4338 5412 4362 5414
rect 4418 5412 4424 5414
rect 4116 5392 4424 5412
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 4080 4622 4108 5102
rect 4436 4820 4488 4826
rect 4436 4762 4488 4768
rect 4448 4690 4476 4762
rect 4436 4684 4488 4690
rect 4436 4626 4488 4632
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 4116 4380 4424 4400
rect 4116 4378 4122 4380
rect 4178 4378 4202 4380
rect 4258 4378 4282 4380
rect 4338 4378 4362 4380
rect 4418 4378 4424 4380
rect 4178 4326 4180 4378
rect 4360 4326 4362 4378
rect 4116 4324 4122 4326
rect 4178 4324 4202 4326
rect 4258 4324 4282 4326
rect 4338 4324 4362 4326
rect 4418 4324 4424 4326
rect 4116 4304 4424 4324
rect 4344 4208 4396 4214
rect 4344 4150 4396 4156
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 4356 3738 4384 4150
rect 4344 3732 4396 3738
rect 4344 3674 4396 3680
rect 3974 3632 4030 3641
rect 4540 3602 4568 6802
rect 4632 6322 4660 7754
rect 4724 7478 4752 9551
rect 4712 7472 4764 7478
rect 4712 7414 4764 7420
rect 4816 7410 4844 10084
rect 5000 9976 5028 10406
rect 5092 10198 5120 10950
rect 5080 10192 5132 10198
rect 5080 10134 5132 10140
rect 4908 9948 5028 9976
rect 4908 9674 4936 9948
rect 5184 9738 5212 11206
rect 5184 9710 5329 9738
rect 5078 9688 5134 9697
rect 4908 9646 5028 9674
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 4908 8537 4936 9454
rect 4894 8528 4950 8537
rect 4894 8463 4950 8472
rect 4896 7880 4948 7886
rect 4896 7822 4948 7828
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 4802 7304 4858 7313
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 4724 6118 4752 7278
rect 4802 7239 4858 7248
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 4620 5364 4672 5370
rect 4724 5352 4752 6054
rect 4672 5324 4752 5352
rect 4620 5306 4672 5312
rect 4816 4672 4844 7239
rect 4908 6458 4936 7822
rect 5000 6798 5028 9646
rect 5301 9636 5329 9710
rect 5078 9623 5134 9632
rect 5092 9042 5120 9623
rect 5276 9608 5329 9636
rect 5170 9480 5226 9489
rect 5170 9415 5172 9424
rect 5224 9415 5226 9424
rect 5172 9386 5224 9392
rect 5184 9042 5212 9386
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 5172 9036 5224 9042
rect 5172 8978 5224 8984
rect 5184 8922 5212 8978
rect 5092 8906 5212 8922
rect 5080 8900 5212 8906
rect 5132 8894 5212 8900
rect 5080 8842 5132 8848
rect 5092 8566 5120 8842
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 5080 8560 5132 8566
rect 5080 8502 5132 8508
rect 5080 8424 5132 8430
rect 5080 8366 5132 8372
rect 4988 6792 5040 6798
rect 4988 6734 5040 6740
rect 4988 6656 5040 6662
rect 4988 6598 5040 6604
rect 4896 6452 4948 6458
rect 4896 6394 4948 6400
rect 5000 6202 5028 6598
rect 4632 4644 4844 4672
rect 4908 6174 5028 6202
rect 3974 3567 4030 3576
rect 4528 3596 4580 3602
rect 3988 3534 4016 3567
rect 4528 3538 4580 3544
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3436 3126 3464 3470
rect 3528 3454 3648 3482
rect 3516 3392 3568 3398
rect 3516 3334 3568 3340
rect 3424 3120 3476 3126
rect 3424 3062 3476 3068
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 3240 2576 3292 2582
rect 3240 2518 3292 2524
rect 3436 2446 3464 2586
rect 3332 2440 3384 2446
rect 3332 2382 3384 2388
rect 3424 2440 3476 2446
rect 3424 2382 3476 2388
rect 3148 1828 3200 1834
rect 3148 1770 3200 1776
rect 1032 1556 1084 1562
rect 1032 1498 1084 1504
rect 3344 1494 3372 2382
rect 3528 1970 3556 3334
rect 3620 2632 3648 3454
rect 3712 3454 3924 3482
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 3712 3398 3740 3454
rect 3700 3392 3752 3398
rect 3700 3334 3752 3340
rect 3882 3224 3938 3233
rect 3882 3159 3884 3168
rect 3936 3159 3938 3168
rect 3884 3130 3936 3136
rect 3884 2848 3936 2854
rect 3884 2790 3936 2796
rect 3700 2644 3752 2650
rect 3620 2604 3700 2632
rect 3700 2586 3752 2592
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 3424 1964 3476 1970
rect 3424 1906 3476 1912
rect 3516 1964 3568 1970
rect 3516 1906 3568 1912
rect 3436 1562 3464 1906
rect 3424 1556 3476 1562
rect 3424 1498 3476 1504
rect 3332 1488 3384 1494
rect 3332 1430 3384 1436
rect 3528 1426 3556 1906
rect 3516 1420 3568 1426
rect 3516 1362 3568 1368
rect 3804 1222 3832 2382
rect 3896 2106 3924 2790
rect 3988 2650 4016 3470
rect 4116 3292 4424 3312
rect 4116 3290 4122 3292
rect 4178 3290 4202 3292
rect 4258 3290 4282 3292
rect 4338 3290 4362 3292
rect 4418 3290 4424 3292
rect 4178 3238 4180 3290
rect 4360 3238 4362 3290
rect 4116 3236 4122 3238
rect 4178 3236 4202 3238
rect 4258 3236 4282 3238
rect 4338 3236 4362 3238
rect 4418 3236 4424 3238
rect 4116 3216 4424 3236
rect 4540 3058 4568 3538
rect 4632 3466 4660 4644
rect 4712 4548 4764 4554
rect 4712 4490 4764 4496
rect 4620 3460 4672 3466
rect 4620 3402 4672 3408
rect 4618 3360 4674 3369
rect 4618 3295 4674 3304
rect 4632 3194 4660 3295
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4724 3058 4752 4490
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 4816 3534 4844 4422
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 4908 3074 4936 6174
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 5000 5914 5028 6054
rect 4988 5908 5040 5914
rect 4988 5850 5040 5856
rect 5092 5370 5120 8366
rect 5184 7750 5212 8774
rect 5276 7857 5304 9608
rect 5262 7848 5318 7857
rect 5262 7783 5318 7792
rect 5172 7744 5224 7750
rect 5224 7704 5304 7732
rect 5172 7686 5224 7692
rect 5172 7472 5224 7478
rect 5172 7414 5224 7420
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 5092 4622 5120 5306
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 4988 4548 5040 4554
rect 4988 4490 5040 4496
rect 5000 4282 5028 4490
rect 5184 4434 5212 7414
rect 5092 4406 5212 4434
rect 4988 4276 5040 4282
rect 4988 4218 5040 4224
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 5000 3398 5028 4082
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 4528 3052 4580 3058
rect 4528 2994 4580 3000
rect 4712 3052 4764 3058
rect 4908 3046 5028 3074
rect 4712 2994 4764 3000
rect 4068 2848 4120 2854
rect 4068 2790 4120 2796
rect 3976 2644 4028 2650
rect 3976 2586 4028 2592
rect 4080 2582 4108 2790
rect 4540 2582 4568 2994
rect 4896 2984 4948 2990
rect 4896 2926 4948 2932
rect 4068 2576 4120 2582
rect 4068 2518 4120 2524
rect 4528 2576 4580 2582
rect 4528 2518 4580 2524
rect 3976 2440 4028 2446
rect 3976 2382 4028 2388
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 3884 2100 3936 2106
rect 3884 2042 3936 2048
rect 3884 1964 3936 1970
rect 3884 1906 3936 1912
rect 3896 1222 3924 1906
rect 3988 1544 4016 2382
rect 4116 2204 4424 2224
rect 4116 2202 4122 2204
rect 4178 2202 4202 2204
rect 4258 2202 4282 2204
rect 4338 2202 4362 2204
rect 4418 2202 4424 2204
rect 4178 2150 4180 2202
rect 4360 2150 4362 2202
rect 4116 2148 4122 2150
rect 4178 2148 4202 2150
rect 4258 2148 4282 2150
rect 4338 2148 4362 2150
rect 4418 2148 4424 2150
rect 4116 2128 4424 2148
rect 4540 1902 4568 2382
rect 4528 1896 4580 1902
rect 4528 1838 4580 1844
rect 4724 1766 4752 2382
rect 4908 2038 4936 2926
rect 4896 2032 4948 2038
rect 4896 1974 4948 1980
rect 5000 1902 5028 3046
rect 4988 1896 5040 1902
rect 4988 1838 5040 1844
rect 4252 1760 4304 1766
rect 4252 1702 4304 1708
rect 4712 1760 4764 1766
rect 4712 1702 4764 1708
rect 4264 1562 4292 1702
rect 5092 1562 5120 4406
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5184 3126 5212 3674
rect 5172 3120 5224 3126
rect 5172 3062 5224 3068
rect 5276 2854 5304 7704
rect 5368 3369 5396 12038
rect 5446 11656 5502 11665
rect 5446 11591 5502 11600
rect 5460 11286 5488 11591
rect 5448 11280 5500 11286
rect 5448 11222 5500 11228
rect 5446 10840 5502 10849
rect 5446 10775 5502 10784
rect 5460 9738 5488 10775
rect 5552 10577 5580 12200
rect 6012 12170 6040 12200
rect 6000 12164 6052 12170
rect 6000 12106 6052 12112
rect 6368 12164 6420 12170
rect 6368 12106 6420 12112
rect 6092 12096 6144 12102
rect 6092 12038 6144 12044
rect 6104 11914 6132 12038
rect 6012 11886 6132 11914
rect 5666 11452 5974 11472
rect 5666 11450 5672 11452
rect 5728 11450 5752 11452
rect 5808 11450 5832 11452
rect 5888 11450 5912 11452
rect 5968 11450 5974 11452
rect 5728 11398 5730 11450
rect 5910 11398 5912 11450
rect 5666 11396 5672 11398
rect 5728 11396 5752 11398
rect 5808 11396 5832 11398
rect 5888 11396 5912 11398
rect 5968 11396 5974 11398
rect 5666 11376 5974 11396
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 5828 10742 5856 11086
rect 5908 11008 5960 11014
rect 5908 10950 5960 10956
rect 5816 10736 5868 10742
rect 5816 10678 5868 10684
rect 5920 10577 5948 10950
rect 5538 10568 5594 10577
rect 5538 10503 5594 10512
rect 5906 10568 5962 10577
rect 5906 10503 5962 10512
rect 5666 10364 5974 10384
rect 5666 10362 5672 10364
rect 5728 10362 5752 10364
rect 5808 10362 5832 10364
rect 5888 10362 5912 10364
rect 5968 10362 5974 10364
rect 5728 10310 5730 10362
rect 5910 10310 5912 10362
rect 5666 10308 5672 10310
rect 5728 10308 5752 10310
rect 5808 10308 5832 10310
rect 5888 10308 5912 10310
rect 5968 10308 5974 10310
rect 5666 10288 5974 10308
rect 5632 10192 5684 10198
rect 5632 10134 5684 10140
rect 5644 9761 5672 10134
rect 5816 9988 5868 9994
rect 5816 9930 5868 9936
rect 5630 9752 5686 9761
rect 5460 9710 5580 9738
rect 5552 9674 5580 9710
rect 5630 9687 5686 9696
rect 5460 9646 5580 9674
rect 5460 9382 5488 9646
rect 5722 9616 5778 9625
rect 5632 9580 5684 9586
rect 5828 9586 5856 9930
rect 5722 9551 5778 9560
rect 5816 9580 5868 9586
rect 5632 9522 5684 9528
rect 5644 9489 5672 9522
rect 5736 9518 5764 9551
rect 5816 9522 5868 9528
rect 5724 9512 5776 9518
rect 5630 9480 5686 9489
rect 5724 9454 5776 9460
rect 5630 9415 5686 9424
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5460 3641 5488 8230
rect 5552 6186 5580 9318
rect 5666 9276 5974 9296
rect 5666 9274 5672 9276
rect 5728 9274 5752 9276
rect 5808 9274 5832 9276
rect 5888 9274 5912 9276
rect 5968 9274 5974 9276
rect 5728 9222 5730 9274
rect 5910 9222 5912 9274
rect 5666 9220 5672 9222
rect 5728 9220 5752 9222
rect 5808 9220 5832 9222
rect 5888 9220 5912 9222
rect 5968 9220 5974 9222
rect 5666 9200 5974 9220
rect 5908 8900 5960 8906
rect 5908 8842 5960 8848
rect 5920 8430 5948 8842
rect 5908 8424 5960 8430
rect 5908 8366 5960 8372
rect 6012 8378 6040 11886
rect 6092 11824 6144 11830
rect 6092 11766 6144 11772
rect 6104 8566 6132 11766
rect 6184 11620 6236 11626
rect 6184 11562 6236 11568
rect 6196 11286 6224 11562
rect 6184 11280 6236 11286
rect 6184 11222 6236 11228
rect 6276 11008 6328 11014
rect 6276 10950 6328 10956
rect 6184 10260 6236 10266
rect 6184 10202 6236 10208
rect 6196 9586 6224 10202
rect 6184 9580 6236 9586
rect 6184 9522 6236 9528
rect 6182 9480 6238 9489
rect 6182 9415 6238 9424
rect 6092 8560 6144 8566
rect 6196 8537 6224 9415
rect 6092 8502 6144 8508
rect 6182 8528 6238 8537
rect 6182 8463 6238 8472
rect 6012 8350 6132 8378
rect 6000 8288 6052 8294
rect 6000 8230 6052 8236
rect 5666 8188 5974 8208
rect 5666 8186 5672 8188
rect 5728 8186 5752 8188
rect 5808 8186 5832 8188
rect 5888 8186 5912 8188
rect 5968 8186 5974 8188
rect 5728 8134 5730 8186
rect 5910 8134 5912 8186
rect 5666 8132 5672 8134
rect 5728 8132 5752 8134
rect 5808 8132 5832 8134
rect 5888 8132 5912 8134
rect 5968 8132 5974 8134
rect 5666 8112 5974 8132
rect 6012 7954 6040 8230
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 6104 7528 6132 8350
rect 6104 7500 6224 7528
rect 6092 7404 6144 7410
rect 6092 7346 6144 7352
rect 5828 7274 6040 7290
rect 5816 7268 6040 7274
rect 5868 7262 6040 7268
rect 5816 7210 5868 7216
rect 5666 7100 5974 7120
rect 5666 7098 5672 7100
rect 5728 7098 5752 7100
rect 5808 7098 5832 7100
rect 5888 7098 5912 7100
rect 5968 7098 5974 7100
rect 5728 7046 5730 7098
rect 5910 7046 5912 7098
rect 5666 7044 5672 7046
rect 5728 7044 5752 7046
rect 5808 7044 5832 7046
rect 5888 7044 5912 7046
rect 5968 7044 5974 7046
rect 5666 7024 5974 7044
rect 5632 6928 5684 6934
rect 5632 6870 5684 6876
rect 5816 6928 5868 6934
rect 5816 6870 5868 6876
rect 5644 6225 5672 6870
rect 5828 6633 5856 6870
rect 5814 6624 5870 6633
rect 5814 6559 5870 6568
rect 6012 6338 6040 7262
rect 6104 6866 6132 7346
rect 6196 7002 6224 7500
rect 6184 6996 6236 7002
rect 6184 6938 6236 6944
rect 6288 6882 6316 10950
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 6196 6854 6316 6882
rect 6090 6760 6146 6769
rect 6090 6695 6092 6704
rect 6144 6695 6146 6704
rect 6092 6666 6144 6672
rect 5920 6322 6040 6338
rect 5908 6316 6040 6322
rect 5960 6310 6040 6316
rect 5908 6258 5960 6264
rect 6104 6236 6132 6666
rect 5630 6216 5686 6225
rect 5540 6180 5592 6186
rect 5630 6151 5686 6160
rect 6012 6208 6132 6236
rect 5540 6122 5592 6128
rect 5666 6012 5974 6032
rect 5666 6010 5672 6012
rect 5728 6010 5752 6012
rect 5808 6010 5832 6012
rect 5888 6010 5912 6012
rect 5968 6010 5974 6012
rect 5728 5958 5730 6010
rect 5910 5958 5912 6010
rect 5666 5956 5672 5958
rect 5728 5956 5752 5958
rect 5808 5956 5832 5958
rect 5888 5956 5912 5958
rect 5968 5956 5974 5958
rect 5666 5936 5974 5956
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5552 5642 5580 5850
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 5540 5636 5592 5642
rect 5540 5578 5592 5584
rect 5816 5636 5868 5642
rect 5816 5578 5868 5584
rect 5552 5234 5580 5578
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 5828 5148 5856 5578
rect 5920 5273 5948 5646
rect 6012 5522 6040 6208
rect 6092 6112 6144 6118
rect 6092 6054 6144 6060
rect 6104 5642 6132 6054
rect 6092 5636 6144 5642
rect 6092 5578 6144 5584
rect 6012 5494 6132 5522
rect 5906 5264 5962 5273
rect 5906 5199 5962 5208
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 5908 5160 5960 5166
rect 5828 5120 5908 5148
rect 5908 5102 5960 5108
rect 5540 5092 5592 5098
rect 5540 5034 5592 5040
rect 5446 3632 5502 3641
rect 5446 3567 5502 3576
rect 5354 3360 5410 3369
rect 5354 3295 5410 3304
rect 5264 2848 5316 2854
rect 5264 2790 5316 2796
rect 5552 2650 5580 5034
rect 5666 4924 5974 4944
rect 5666 4922 5672 4924
rect 5728 4922 5752 4924
rect 5808 4922 5832 4924
rect 5888 4922 5912 4924
rect 5968 4922 5974 4924
rect 5728 4870 5730 4922
rect 5910 4870 5912 4922
rect 5666 4868 5672 4870
rect 5728 4868 5752 4870
rect 5808 4868 5832 4870
rect 5888 4868 5912 4870
rect 5968 4868 5974 4870
rect 5666 4848 5974 4868
rect 6012 4808 6040 5170
rect 5828 4780 6040 4808
rect 5828 3924 5856 4780
rect 6104 4706 6132 5494
rect 6012 4678 6132 4706
rect 6012 4078 6040 4678
rect 6092 4480 6144 4486
rect 6092 4422 6144 4428
rect 6000 4072 6052 4078
rect 6000 4014 6052 4020
rect 5828 3896 6040 3924
rect 5666 3836 5974 3856
rect 5666 3834 5672 3836
rect 5728 3834 5752 3836
rect 5808 3834 5832 3836
rect 5888 3834 5912 3836
rect 5968 3834 5974 3836
rect 5728 3782 5730 3834
rect 5910 3782 5912 3834
rect 5666 3780 5672 3782
rect 5728 3780 5752 3782
rect 5808 3780 5832 3782
rect 5888 3780 5912 3782
rect 5968 3780 5974 3782
rect 5666 3760 5974 3780
rect 6012 3670 6040 3896
rect 6000 3664 6052 3670
rect 5630 3632 5686 3641
rect 6000 3606 6052 3612
rect 6104 3602 6132 4422
rect 5630 3567 5686 3576
rect 6092 3596 6144 3602
rect 5644 3534 5672 3567
rect 6092 3538 6144 3544
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 6000 3392 6052 3398
rect 6000 3334 6052 3340
rect 6012 3058 6040 3334
rect 6092 3120 6144 3126
rect 6092 3062 6144 3068
rect 6000 3052 6052 3058
rect 6000 2994 6052 3000
rect 5666 2748 5974 2768
rect 5666 2746 5672 2748
rect 5728 2746 5752 2748
rect 5808 2746 5832 2748
rect 5888 2746 5912 2748
rect 5968 2746 5974 2748
rect 5728 2694 5730 2746
rect 5910 2694 5912 2746
rect 5666 2692 5672 2694
rect 5728 2692 5752 2694
rect 5808 2692 5832 2694
rect 5888 2692 5912 2694
rect 5968 2692 5974 2694
rect 5666 2672 5974 2692
rect 6104 2650 6132 3062
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 6092 2644 6144 2650
rect 6092 2586 6144 2592
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 5184 2106 5212 2382
rect 5172 2100 5224 2106
rect 5172 2042 5224 2048
rect 6196 1970 6224 6854
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6288 5778 6316 6598
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 6288 4690 6316 5714
rect 6276 4684 6328 4690
rect 6276 4626 6328 4632
rect 6276 4548 6328 4554
rect 6276 4490 6328 4496
rect 6288 4010 6316 4490
rect 6276 4004 6328 4010
rect 6276 3946 6328 3952
rect 6288 3738 6316 3946
rect 6276 3732 6328 3738
rect 6276 3674 6328 3680
rect 6276 3528 6328 3534
rect 6276 3470 6328 3476
rect 6288 3126 6316 3470
rect 6276 3120 6328 3126
rect 6276 3062 6328 3068
rect 6276 2984 6328 2990
rect 6276 2926 6328 2932
rect 6288 2038 6316 2926
rect 6276 2032 6328 2038
rect 6276 1974 6328 1980
rect 6184 1964 6236 1970
rect 6184 1906 6236 1912
rect 6380 1766 6408 12106
rect 6472 12102 6500 12200
rect 6460 12096 6512 12102
rect 6460 12038 6512 12044
rect 7840 12028 7892 12034
rect 7840 11970 7892 11976
rect 6828 11824 6880 11830
rect 6828 11766 6880 11772
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 6472 11082 6500 11290
rect 6644 11280 6696 11286
rect 6644 11222 6696 11228
rect 6460 11076 6512 11082
rect 6460 11018 6512 11024
rect 6472 10674 6500 11018
rect 6460 10668 6512 10674
rect 6460 10610 6512 10616
rect 6472 10198 6500 10610
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 6460 10192 6512 10198
rect 6460 10134 6512 10140
rect 6458 10024 6514 10033
rect 6458 9959 6514 9968
rect 6472 2106 6500 9959
rect 6564 9722 6592 10542
rect 6656 10033 6684 11222
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6642 10024 6698 10033
rect 6642 9959 6698 9968
rect 6644 9920 6696 9926
rect 6644 9862 6696 9868
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6552 8492 6604 8498
rect 6552 8434 6604 8440
rect 6564 7449 6592 8434
rect 6550 7440 6606 7449
rect 6550 7375 6606 7384
rect 6550 7304 6606 7313
rect 6550 7239 6606 7248
rect 6564 6186 6592 7239
rect 6552 6180 6604 6186
rect 6552 6122 6604 6128
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6564 4690 6592 5510
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6564 4146 6592 4626
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 6564 3738 6592 3878
rect 6552 3732 6604 3738
rect 6552 3674 6604 3680
rect 6656 3641 6684 9862
rect 6748 8498 6776 11086
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6734 8392 6790 8401
rect 6734 8327 6790 8336
rect 6748 6662 6776 8327
rect 6840 7410 6868 11766
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6932 10742 6960 11698
rect 7104 11620 7156 11626
rect 7104 11562 7156 11568
rect 7116 11354 7144 11562
rect 7104 11348 7156 11354
rect 7104 11290 7156 11296
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7208 11257 7236 11290
rect 7194 11248 7250 11257
rect 7300 11218 7788 11234
rect 7194 11183 7250 11192
rect 7288 11212 7788 11218
rect 7340 11206 7788 11212
rect 7288 11154 7340 11160
rect 7104 11144 7156 11150
rect 7656 11144 7708 11150
rect 7104 11086 7156 11092
rect 7562 11112 7618 11121
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 6920 10736 6972 10742
rect 6920 10678 6972 10684
rect 7024 10554 7052 10746
rect 6932 10526 7052 10554
rect 6932 9489 6960 10526
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 6918 9480 6974 9489
rect 6918 9415 6974 9424
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6932 8498 6960 9318
rect 7024 8974 7052 10406
rect 7116 9704 7144 11086
rect 7656 11086 7708 11092
rect 7562 11047 7618 11056
rect 7216 10908 7524 10928
rect 7216 10906 7222 10908
rect 7278 10906 7302 10908
rect 7358 10906 7382 10908
rect 7438 10906 7462 10908
rect 7518 10906 7524 10908
rect 7278 10854 7280 10906
rect 7460 10854 7462 10906
rect 7216 10852 7222 10854
rect 7278 10852 7302 10854
rect 7358 10852 7382 10854
rect 7438 10852 7462 10854
rect 7518 10852 7524 10854
rect 7216 10832 7524 10852
rect 7576 10266 7604 11047
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7216 9820 7524 9840
rect 7216 9818 7222 9820
rect 7278 9818 7302 9820
rect 7358 9818 7382 9820
rect 7438 9818 7462 9820
rect 7518 9818 7524 9820
rect 7278 9766 7280 9818
rect 7460 9766 7462 9818
rect 7216 9764 7222 9766
rect 7278 9764 7302 9766
rect 7358 9764 7382 9766
rect 7438 9764 7462 9766
rect 7518 9764 7524 9766
rect 7216 9744 7524 9764
rect 7116 9676 7236 9704
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 7116 9178 7144 9522
rect 7208 9382 7236 9676
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 7012 8832 7064 8838
rect 7012 8774 7064 8780
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 7024 8378 7052 8774
rect 7216 8732 7524 8752
rect 7216 8730 7222 8732
rect 7278 8730 7302 8732
rect 7358 8730 7382 8732
rect 7438 8730 7462 8732
rect 7518 8730 7524 8732
rect 7278 8678 7280 8730
rect 7460 8678 7462 8730
rect 7216 8676 7222 8678
rect 7278 8676 7302 8678
rect 7358 8676 7382 8678
rect 7438 8676 7462 8678
rect 7518 8676 7524 8678
rect 7216 8656 7524 8676
rect 7194 8528 7250 8537
rect 7194 8463 7250 8472
rect 6932 8350 7052 8378
rect 6932 7818 6960 8350
rect 7012 8288 7064 8294
rect 7012 8230 7064 8236
rect 7024 7886 7052 8230
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 6828 7268 6880 7274
rect 6828 7210 6880 7216
rect 6736 6656 6788 6662
rect 6736 6598 6788 6604
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6748 3942 6776 6258
rect 6840 5930 6868 7210
rect 6932 7002 6960 7754
rect 7012 7744 7064 7750
rect 7208 7732 7236 8463
rect 7012 7686 7064 7692
rect 7116 7704 7236 7732
rect 7024 7002 7052 7686
rect 7116 7528 7144 7704
rect 7216 7644 7524 7664
rect 7216 7642 7222 7644
rect 7278 7642 7302 7644
rect 7358 7642 7382 7644
rect 7438 7642 7462 7644
rect 7518 7642 7524 7644
rect 7278 7590 7280 7642
rect 7460 7590 7462 7642
rect 7216 7588 7222 7590
rect 7278 7588 7302 7590
rect 7358 7588 7382 7590
rect 7438 7588 7462 7590
rect 7518 7588 7524 7590
rect 7216 7568 7524 7588
rect 7116 7500 7236 7528
rect 7104 7268 7156 7274
rect 7104 7210 7156 7216
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 7012 6996 7064 7002
rect 7012 6938 7064 6944
rect 6920 6724 6972 6730
rect 6972 6684 7052 6712
rect 6920 6666 6972 6672
rect 7024 6633 7052 6684
rect 7010 6624 7066 6633
rect 7010 6559 7066 6568
rect 6840 5902 6960 5930
rect 6828 5840 6880 5846
rect 6828 5782 6880 5788
rect 6840 4298 6868 5782
rect 6932 5273 6960 5902
rect 7024 5642 7052 6559
rect 7116 6458 7144 7210
rect 7208 6769 7236 7500
rect 7288 7200 7340 7206
rect 7288 7142 7340 7148
rect 7194 6760 7250 6769
rect 7300 6730 7328 7142
rect 7194 6695 7250 6704
rect 7288 6724 7340 6730
rect 7288 6666 7340 6672
rect 7216 6556 7524 6576
rect 7216 6554 7222 6556
rect 7278 6554 7302 6556
rect 7358 6554 7382 6556
rect 7438 6554 7462 6556
rect 7518 6554 7524 6556
rect 7278 6502 7280 6554
rect 7460 6502 7462 6554
rect 7216 6500 7222 6502
rect 7278 6500 7302 6502
rect 7358 6500 7382 6502
rect 7438 6500 7462 6502
rect 7518 6500 7524 6502
rect 7216 6480 7524 6500
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 7102 6216 7158 6225
rect 7102 6151 7158 6160
rect 7012 5636 7064 5642
rect 7012 5578 7064 5584
rect 6918 5264 6974 5273
rect 6918 5199 6974 5208
rect 7024 5012 7052 5578
rect 7116 5216 7144 6151
rect 7216 5468 7524 5488
rect 7216 5466 7222 5468
rect 7278 5466 7302 5468
rect 7358 5466 7382 5468
rect 7438 5466 7462 5468
rect 7518 5466 7524 5468
rect 7278 5414 7280 5466
rect 7460 5414 7462 5466
rect 7216 5412 7222 5414
rect 7278 5412 7302 5414
rect 7358 5412 7382 5414
rect 7438 5412 7462 5414
rect 7518 5412 7524 5414
rect 7216 5392 7524 5412
rect 7116 5188 7236 5216
rect 7104 5024 7156 5030
rect 7024 4984 7104 5012
rect 7104 4966 7156 4972
rect 7116 4554 7144 4966
rect 7208 4729 7236 5188
rect 7194 4720 7250 4729
rect 7194 4655 7250 4664
rect 7104 4548 7156 4554
rect 7104 4490 7156 4496
rect 6840 4270 7052 4298
rect 6918 4176 6974 4185
rect 6828 4140 6880 4146
rect 6918 4111 6920 4120
rect 6828 4082 6880 4088
rect 6972 4111 6974 4120
rect 6920 4082 6972 4088
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6642 3632 6698 3641
rect 6642 3567 6698 3576
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6564 2650 6592 3470
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 6748 2446 6776 3334
rect 6840 3194 6868 4082
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 6932 3602 6960 3878
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 6826 3088 6882 3097
rect 6826 3023 6882 3032
rect 6840 2514 6868 3023
rect 6932 2650 6960 3334
rect 7024 3058 7052 4270
rect 7116 4264 7144 4490
rect 7216 4380 7524 4400
rect 7216 4378 7222 4380
rect 7278 4378 7302 4380
rect 7358 4378 7382 4380
rect 7438 4378 7462 4380
rect 7518 4378 7524 4380
rect 7278 4326 7280 4378
rect 7460 4326 7462 4378
rect 7216 4324 7222 4326
rect 7278 4324 7302 4326
rect 7358 4324 7382 4326
rect 7438 4324 7462 4326
rect 7518 4324 7524 4326
rect 7216 4304 7524 4324
rect 7116 4236 7236 4264
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 7012 3052 7064 3058
rect 7012 2994 7064 3000
rect 7116 2650 7144 4014
rect 7208 4010 7236 4236
rect 7196 4004 7248 4010
rect 7196 3946 7248 3952
rect 7378 3632 7434 3641
rect 7378 3567 7380 3576
rect 7432 3567 7434 3576
rect 7380 3538 7432 3544
rect 7216 3292 7524 3312
rect 7216 3290 7222 3292
rect 7278 3290 7302 3292
rect 7358 3290 7382 3292
rect 7438 3290 7462 3292
rect 7518 3290 7524 3292
rect 7278 3238 7280 3290
rect 7460 3238 7462 3290
rect 7216 3236 7222 3238
rect 7278 3236 7302 3238
rect 7358 3236 7382 3238
rect 7438 3236 7462 3238
rect 7518 3236 7524 3238
rect 7216 3216 7524 3236
rect 7194 3088 7250 3097
rect 7194 3023 7250 3032
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 6828 2508 6880 2514
rect 6828 2450 6880 2456
rect 7208 2446 7236 3023
rect 7378 2544 7434 2553
rect 7378 2479 7380 2488
rect 7432 2479 7434 2488
rect 7380 2450 7432 2456
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7216 2204 7524 2224
rect 7216 2202 7222 2204
rect 7278 2202 7302 2204
rect 7358 2202 7382 2204
rect 7438 2202 7462 2204
rect 7518 2202 7524 2204
rect 7278 2150 7280 2202
rect 7460 2150 7462 2202
rect 7216 2148 7222 2150
rect 7278 2148 7302 2150
rect 7358 2148 7382 2150
rect 7438 2148 7462 2150
rect 7518 2148 7524 2150
rect 7216 2128 7524 2148
rect 6460 2100 6512 2106
rect 6460 2042 6512 2048
rect 6368 1760 6420 1766
rect 6368 1702 6420 1708
rect 5666 1660 5974 1680
rect 5666 1658 5672 1660
rect 5728 1658 5752 1660
rect 5808 1658 5832 1660
rect 5888 1658 5912 1660
rect 5968 1658 5974 1660
rect 5728 1606 5730 1658
rect 5910 1606 5912 1658
rect 5666 1604 5672 1606
rect 5728 1604 5752 1606
rect 5808 1604 5832 1606
rect 5888 1604 5912 1606
rect 5968 1604 5974 1606
rect 5666 1584 5974 1604
rect 4068 1556 4120 1562
rect 3988 1516 4068 1544
rect 4068 1498 4120 1504
rect 4252 1556 4304 1562
rect 4252 1498 4304 1504
rect 5080 1556 5132 1562
rect 5080 1498 5132 1504
rect 7576 1358 7604 10066
rect 7668 8362 7696 11086
rect 7656 8356 7708 8362
rect 7656 8298 7708 8304
rect 7760 7562 7788 11206
rect 7852 9586 7880 11970
rect 8576 11960 8628 11966
rect 8576 11902 8628 11908
rect 8392 11892 8444 11898
rect 8392 11834 8444 11840
rect 8208 11824 8260 11830
rect 8208 11766 8260 11772
rect 7932 11348 7984 11354
rect 7932 11290 7984 11296
rect 7944 11082 7972 11290
rect 8220 11150 8248 11766
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 7932 11076 7984 11082
rect 7932 11018 7984 11024
rect 7944 10248 7972 11018
rect 8022 10704 8078 10713
rect 8128 10674 8156 11086
rect 8022 10639 8024 10648
rect 8076 10639 8078 10648
rect 8116 10668 8168 10674
rect 8024 10610 8076 10616
rect 8116 10610 8168 10616
rect 8024 10532 8076 10538
rect 8024 10474 8076 10480
rect 8036 10266 8064 10474
rect 8024 10260 8076 10266
rect 7944 10220 8024 10248
rect 8024 10202 8076 10208
rect 8128 10169 8156 10610
rect 8114 10160 8170 10169
rect 8312 10146 8340 11494
rect 8114 10095 8170 10104
rect 8220 10118 8340 10146
rect 8024 10056 8076 10062
rect 8022 10024 8024 10033
rect 8116 10056 8168 10062
rect 8076 10024 8078 10033
rect 7932 9988 7984 9994
rect 8116 9998 8168 10004
rect 8022 9959 8078 9968
rect 7932 9930 7984 9936
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 7944 9160 7972 9930
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 7668 7534 7788 7562
rect 7852 9132 7972 9160
rect 7668 4078 7696 7534
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 7760 6769 7788 7346
rect 7746 6760 7802 6769
rect 7746 6695 7802 6704
rect 7852 6610 7880 9132
rect 7930 9072 7986 9081
rect 7930 9007 7986 9016
rect 7944 7478 7972 9007
rect 7932 7472 7984 7478
rect 7932 7414 7984 7420
rect 7760 6582 7880 6610
rect 7760 5370 7788 6582
rect 7840 6452 7892 6458
rect 7840 6394 7892 6400
rect 7748 5364 7800 5370
rect 7748 5306 7800 5312
rect 7748 5228 7800 5234
rect 7748 5170 7800 5176
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 7668 3126 7696 3878
rect 7656 3120 7708 3126
rect 7656 3062 7708 3068
rect 7656 2848 7708 2854
rect 7656 2790 7708 2796
rect 7668 2378 7696 2790
rect 7760 2582 7788 5170
rect 7852 4570 7880 6394
rect 7944 5370 7972 7414
rect 8036 5574 8064 9862
rect 8128 9625 8156 9998
rect 8114 9616 8170 9625
rect 8114 9551 8170 9560
rect 8220 8566 8248 10118
rect 8298 10024 8354 10033
rect 8298 9959 8354 9968
rect 8312 9042 8340 9959
rect 8404 9654 8432 11834
rect 8484 11552 8536 11558
rect 8484 11494 8536 11500
rect 8496 11354 8524 11494
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8588 10810 8616 11902
rect 9680 11620 9732 11626
rect 9680 11562 9732 11568
rect 8766 11452 9074 11472
rect 8766 11450 8772 11452
rect 8828 11450 8852 11452
rect 8908 11450 8932 11452
rect 8988 11450 9012 11452
rect 9068 11450 9074 11452
rect 8828 11398 8830 11450
rect 9010 11398 9012 11450
rect 8766 11396 8772 11398
rect 8828 11396 8852 11398
rect 8908 11396 8932 11398
rect 8988 11396 9012 11398
rect 9068 11396 9074 11398
rect 8766 11376 9074 11396
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 8576 10804 8628 10810
rect 8576 10746 8628 10752
rect 8392 9648 8444 9654
rect 8392 9590 8444 9596
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 8208 8560 8260 8566
rect 8208 8502 8260 8508
rect 8312 7970 8340 8774
rect 8404 8090 8432 8910
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8220 7942 8340 7970
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 8024 5568 8076 5574
rect 8024 5510 8076 5516
rect 7932 5364 7984 5370
rect 7932 5306 7984 5312
rect 8024 5296 8076 5302
rect 8024 5238 8076 5244
rect 7852 4542 7972 4570
rect 7840 4480 7892 4486
rect 7840 4422 7892 4428
rect 7748 2576 7800 2582
rect 7748 2518 7800 2524
rect 7852 2446 7880 4422
rect 7944 3505 7972 4542
rect 7930 3496 7986 3505
rect 7930 3431 7986 3440
rect 7932 3392 7984 3398
rect 7932 3334 7984 3340
rect 7944 2650 7972 3334
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 7840 2440 7892 2446
rect 7746 2408 7802 2417
rect 7656 2372 7708 2378
rect 7840 2382 7892 2388
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 7746 2343 7802 2352
rect 7656 2314 7708 2320
rect 7760 2106 7788 2343
rect 7840 2304 7892 2310
rect 7840 2246 7892 2252
rect 7852 2106 7880 2246
rect 7748 2100 7800 2106
rect 7748 2042 7800 2048
rect 7840 2100 7892 2106
rect 7840 2042 7892 2048
rect 7944 1494 7972 2382
rect 8036 2310 8064 5238
rect 8128 3058 8156 7686
rect 8220 7177 8248 7942
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 8206 7168 8262 7177
rect 8206 7103 8262 7112
rect 8312 7002 8340 7822
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 8404 7546 8432 7754
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8392 7336 8444 7342
rect 8392 7278 8444 7284
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 8208 6724 8260 6730
rect 8208 6666 8260 6672
rect 8220 6458 8248 6666
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8208 6180 8260 6186
rect 8208 6122 8260 6128
rect 8220 5914 8248 6122
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 8206 5808 8262 5817
rect 8206 5743 8262 5752
rect 8220 4321 8248 5743
rect 8312 5642 8340 6938
rect 8300 5636 8352 5642
rect 8300 5578 8352 5584
rect 8404 4434 8432 7278
rect 8496 6934 8524 10746
rect 8574 10704 8630 10713
rect 8574 10639 8630 10648
rect 8588 10198 8616 10639
rect 8576 10192 8628 10198
rect 8576 10134 8628 10140
rect 8588 9722 8616 10134
rect 8576 9716 8628 9722
rect 8576 9658 8628 9664
rect 8576 9036 8628 9042
rect 8576 8978 8628 8984
rect 8588 8022 8616 8978
rect 8576 8016 8628 8022
rect 8576 7958 8628 7964
rect 8484 6928 8536 6934
rect 8484 6870 8536 6876
rect 8484 6112 8536 6118
rect 8484 6054 8536 6060
rect 8496 4826 8524 6054
rect 8588 5778 8616 7958
rect 8680 6882 8708 11290
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 8766 10364 9074 10384
rect 8766 10362 8772 10364
rect 8828 10362 8852 10364
rect 8908 10362 8932 10364
rect 8988 10362 9012 10364
rect 9068 10362 9074 10364
rect 8828 10310 8830 10362
rect 9010 10310 9012 10362
rect 8766 10308 8772 10310
rect 8828 10308 8852 10310
rect 8908 10308 8932 10310
rect 8988 10308 9012 10310
rect 9068 10308 9074 10310
rect 8766 10288 9074 10308
rect 9140 10198 9168 11086
rect 9588 11008 9640 11014
rect 9588 10950 9640 10956
rect 9600 10713 9628 10950
rect 9586 10704 9642 10713
rect 9312 10668 9364 10674
rect 9586 10639 9642 10648
rect 9312 10610 9364 10616
rect 9220 10532 9272 10538
rect 9220 10474 9272 10480
rect 8944 10192 8996 10198
rect 9128 10192 9180 10198
rect 8944 10134 8996 10140
rect 9034 10160 9090 10169
rect 8852 10056 8904 10062
rect 8850 10024 8852 10033
rect 8904 10024 8906 10033
rect 8956 9994 8984 10134
rect 9128 10134 9180 10140
rect 9034 10095 9090 10104
rect 8850 9959 8906 9968
rect 8944 9988 8996 9994
rect 8944 9930 8996 9936
rect 9048 9674 9076 10095
rect 9048 9646 9168 9674
rect 8766 9276 9074 9296
rect 8766 9274 8772 9276
rect 8828 9274 8852 9276
rect 8908 9274 8932 9276
rect 8988 9274 9012 9276
rect 9068 9274 9074 9276
rect 8828 9222 8830 9274
rect 9010 9222 9012 9274
rect 8766 9220 8772 9222
rect 8828 9220 8852 9222
rect 8908 9220 8932 9222
rect 8988 9220 9012 9222
rect 9068 9220 9074 9222
rect 8766 9200 9074 9220
rect 9140 8838 9168 9646
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 8766 8188 9074 8208
rect 8766 8186 8772 8188
rect 8828 8186 8852 8188
rect 8908 8186 8932 8188
rect 8988 8186 9012 8188
rect 9068 8186 9074 8188
rect 8828 8134 8830 8186
rect 9010 8134 9012 8186
rect 8766 8132 8772 8134
rect 8828 8132 8852 8134
rect 8908 8132 8932 8134
rect 8988 8132 9012 8134
rect 9068 8132 9074 8134
rect 8766 8112 9074 8132
rect 8766 7100 9074 7120
rect 8766 7098 8772 7100
rect 8828 7098 8852 7100
rect 8908 7098 8932 7100
rect 8988 7098 9012 7100
rect 9068 7098 9074 7100
rect 8828 7046 8830 7098
rect 9010 7046 9012 7098
rect 8766 7044 8772 7046
rect 8828 7044 8852 7046
rect 8908 7044 8932 7046
rect 8988 7044 9012 7046
rect 9068 7044 9074 7046
rect 8766 7024 9074 7044
rect 8680 6854 8800 6882
rect 8668 6792 8720 6798
rect 8668 6734 8720 6740
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8680 5658 8708 6734
rect 8772 6322 8800 6854
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 8766 6012 9074 6032
rect 8766 6010 8772 6012
rect 8828 6010 8852 6012
rect 8908 6010 8932 6012
rect 8988 6010 9012 6012
rect 9068 6010 9074 6012
rect 8828 5958 8830 6010
rect 9010 5958 9012 6010
rect 8766 5956 8772 5958
rect 8828 5956 8852 5958
rect 8908 5956 8932 5958
rect 8988 5956 9012 5958
rect 9068 5956 9074 5958
rect 8766 5936 9074 5956
rect 9140 5914 9168 8366
rect 9232 7342 9260 10474
rect 9324 7834 9352 10610
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 9494 9888 9550 9897
rect 9494 9823 9550 9832
rect 9508 9586 9536 9823
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 9416 9178 9444 9454
rect 9600 9382 9628 10542
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 9404 8900 9456 8906
rect 9404 8842 9456 8848
rect 9416 8265 9444 8842
rect 9402 8256 9458 8265
rect 9402 8191 9458 8200
rect 9324 7806 9536 7834
rect 9404 7744 9456 7750
rect 9404 7686 9456 7692
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9220 7336 9272 7342
rect 9220 7278 9272 7284
rect 9232 6866 9260 7278
rect 9220 6860 9272 6866
rect 9220 6802 9272 6808
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 8588 5630 8708 5658
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8588 4457 8616 5630
rect 9128 5296 9180 5302
rect 9128 5238 9180 5244
rect 8668 5160 8720 5166
rect 8668 5102 8720 5108
rect 8312 4406 8432 4434
rect 8574 4448 8630 4457
rect 8206 4312 8262 4321
rect 8206 4247 8262 4256
rect 8208 4208 8260 4214
rect 8208 4150 8260 4156
rect 8312 4162 8340 4406
rect 8574 4383 8630 4392
rect 8220 3194 8248 4150
rect 8312 4134 8524 4162
rect 8300 4072 8352 4078
rect 8352 4032 8432 4060
rect 8300 4014 8352 4020
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8116 3052 8168 3058
rect 8116 2994 8168 3000
rect 8220 2938 8248 3130
rect 8312 3097 8340 3674
rect 8404 3670 8432 4032
rect 8392 3664 8444 3670
rect 8392 3606 8444 3612
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 8298 3088 8354 3097
rect 8298 3023 8354 3032
rect 8128 2910 8248 2938
rect 8298 2952 8354 2961
rect 8024 2304 8076 2310
rect 8024 2246 8076 2252
rect 8128 2106 8156 2910
rect 8298 2887 8354 2896
rect 8208 2848 8260 2854
rect 8208 2790 8260 2796
rect 8116 2100 8168 2106
rect 8116 2042 8168 2048
rect 8220 2038 8248 2790
rect 8208 2032 8260 2038
rect 8208 1974 8260 1980
rect 8312 1970 8340 2887
rect 8300 1964 8352 1970
rect 8300 1906 8352 1912
rect 8404 1766 8432 3470
rect 8496 2106 8524 4134
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 8588 3738 8616 4082
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 8588 3194 8616 3538
rect 8680 3233 8708 5102
rect 8766 4924 9074 4944
rect 8766 4922 8772 4924
rect 8828 4922 8852 4924
rect 8908 4922 8932 4924
rect 8988 4922 9012 4924
rect 9068 4922 9074 4924
rect 8828 4870 8830 4922
rect 9010 4870 9012 4922
rect 8766 4868 8772 4870
rect 8828 4868 8852 4870
rect 8908 4868 8932 4870
rect 8988 4868 9012 4870
rect 9068 4868 9074 4870
rect 8766 4848 9074 4868
rect 8766 3836 9074 3856
rect 8766 3834 8772 3836
rect 8828 3834 8852 3836
rect 8908 3834 8932 3836
rect 8988 3834 9012 3836
rect 9068 3834 9074 3836
rect 8828 3782 8830 3834
rect 9010 3782 9012 3834
rect 8766 3780 8772 3782
rect 8828 3780 8852 3782
rect 8908 3780 8932 3782
rect 8988 3780 9012 3782
rect 9068 3780 9074 3782
rect 8766 3760 9074 3780
rect 8852 3596 8904 3602
rect 8852 3538 8904 3544
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 8666 3224 8722 3233
rect 8576 3188 8628 3194
rect 8666 3159 8722 3168
rect 8576 3130 8628 3136
rect 8574 3088 8630 3097
rect 8574 3023 8630 3032
rect 8484 2100 8536 2106
rect 8484 2042 8536 2048
rect 8588 1902 8616 3023
rect 8772 2836 8800 3470
rect 8864 3058 8892 3538
rect 9036 3392 9088 3398
rect 9036 3334 9088 3340
rect 9048 3194 9076 3334
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 8852 3052 8904 3058
rect 9140 3040 9168 5238
rect 9232 3942 9260 6598
rect 9324 6225 9352 7346
rect 9310 6216 9366 6225
rect 9310 6151 9366 6160
rect 9312 6112 9364 6118
rect 9312 6054 9364 6060
rect 9324 5302 9352 6054
rect 9416 5710 9444 7686
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 9312 5296 9364 5302
rect 9312 5238 9364 5244
rect 9404 5228 9456 5234
rect 9404 5170 9456 5176
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9218 3768 9274 3777
rect 9218 3703 9220 3712
rect 9272 3703 9274 3712
rect 9220 3674 9272 3680
rect 9218 3632 9274 3641
rect 9218 3567 9274 3576
rect 9232 3126 9260 3567
rect 9220 3120 9272 3126
rect 9220 3062 9272 3068
rect 8852 2994 8904 3000
rect 9048 3012 9168 3040
rect 8680 2808 8800 2836
rect 9048 2836 9076 3012
rect 9220 2984 9272 2990
rect 9220 2926 9272 2932
rect 9048 2808 9168 2836
rect 8680 2632 8708 2808
rect 8766 2748 9074 2768
rect 8766 2746 8772 2748
rect 8828 2746 8852 2748
rect 8908 2746 8932 2748
rect 8988 2746 9012 2748
rect 9068 2746 9074 2748
rect 8828 2694 8830 2746
rect 9010 2694 9012 2746
rect 8766 2692 8772 2694
rect 8828 2692 8852 2694
rect 8908 2692 8932 2694
rect 8988 2692 9012 2694
rect 9068 2692 9074 2694
rect 8766 2672 9074 2692
rect 9140 2632 9168 2808
rect 8680 2604 8800 2632
rect 8484 1896 8536 1902
rect 8484 1838 8536 1844
rect 8576 1896 8628 1902
rect 8576 1838 8628 1844
rect 8392 1760 8444 1766
rect 8392 1702 8444 1708
rect 8496 1562 8524 1838
rect 8772 1748 8800 2604
rect 9048 2604 9168 2632
rect 8852 2576 8904 2582
rect 8850 2544 8852 2553
rect 8904 2544 8906 2553
rect 9048 2514 9076 2604
rect 8850 2479 8906 2488
rect 9036 2508 9088 2514
rect 9036 2450 9088 2456
rect 8944 2304 8996 2310
rect 8944 2246 8996 2252
rect 8956 1970 8984 2246
rect 9126 2136 9182 2145
rect 9232 2106 9260 2926
rect 9126 2071 9182 2080
rect 9220 2100 9272 2106
rect 8944 1964 8996 1970
rect 8944 1906 8996 1912
rect 8680 1720 8800 1748
rect 8484 1556 8536 1562
rect 8484 1498 8536 1504
rect 7932 1488 7984 1494
rect 7932 1430 7984 1436
rect 7564 1352 7616 1358
rect 7564 1294 7616 1300
rect 8680 1222 8708 1720
rect 8766 1660 9074 1680
rect 8766 1658 8772 1660
rect 8828 1658 8852 1660
rect 8908 1658 8932 1660
rect 8988 1658 9012 1660
rect 9068 1658 9074 1660
rect 8828 1606 8830 1658
rect 9010 1606 9012 1658
rect 8766 1604 8772 1606
rect 8828 1604 8852 1606
rect 8908 1604 8932 1606
rect 8988 1604 9012 1606
rect 9068 1604 9074 1606
rect 8766 1584 9074 1604
rect 9140 1562 9168 2071
rect 9220 2042 9272 2048
rect 9128 1556 9180 1562
rect 9128 1498 9180 1504
rect 8944 1488 8996 1494
rect 8944 1430 8996 1436
rect 8956 1329 8984 1430
rect 9220 1420 9272 1426
rect 9220 1362 9272 1368
rect 8942 1320 8998 1329
rect 8942 1255 8998 1264
rect 8956 1222 8984 1255
rect 3792 1216 3844 1222
rect 3792 1158 3844 1164
rect 3884 1216 3936 1222
rect 3884 1158 3936 1164
rect 8668 1216 8720 1222
rect 8668 1158 8720 1164
rect 8944 1216 8996 1222
rect 8944 1158 8996 1164
rect 4116 1116 4424 1136
rect 4116 1114 4122 1116
rect 4178 1114 4202 1116
rect 4258 1114 4282 1116
rect 4338 1114 4362 1116
rect 4418 1114 4424 1116
rect 4178 1062 4180 1114
rect 4360 1062 4362 1114
rect 4116 1060 4122 1062
rect 4178 1060 4202 1062
rect 4258 1060 4282 1062
rect 4338 1060 4362 1062
rect 4418 1060 4424 1062
rect 4116 1040 4424 1060
rect 7216 1116 7524 1136
rect 7216 1114 7222 1116
rect 7278 1114 7302 1116
rect 7358 1114 7382 1116
rect 7438 1114 7462 1116
rect 7518 1114 7524 1116
rect 7278 1062 7280 1114
rect 7460 1062 7462 1114
rect 7216 1060 7222 1062
rect 7278 1060 7302 1062
rect 7358 1060 7382 1062
rect 7438 1060 7462 1062
rect 7518 1060 7524 1062
rect 7216 1040 7524 1060
rect 9232 513 9260 1362
rect 9324 921 9352 4966
rect 9416 4162 9444 5170
rect 9508 4282 9536 7806
rect 9600 7342 9628 9318
rect 9692 7449 9720 11562
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 9864 11212 9916 11218
rect 9864 11154 9916 11160
rect 9876 7857 9904 11154
rect 9862 7848 9918 7857
rect 9862 7783 9918 7792
rect 9678 7440 9734 7449
rect 9678 7375 9734 7384
rect 9588 7336 9640 7342
rect 9588 7278 9640 7284
rect 9588 7200 9640 7206
rect 9588 7142 9640 7148
rect 9600 5930 9628 7142
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 9600 5902 9904 5930
rect 9770 5808 9826 5817
rect 9770 5743 9826 5752
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9496 4276 9548 4282
rect 9496 4218 9548 4224
rect 9416 4134 9536 4162
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 9416 3670 9444 4014
rect 9404 3664 9456 3670
rect 9404 3606 9456 3612
rect 9508 3482 9536 4134
rect 9416 3454 9536 3482
rect 9416 2446 9444 3454
rect 9496 3392 9548 3398
rect 9496 3334 9548 3340
rect 9404 2440 9456 2446
rect 9404 2382 9456 2388
rect 9508 1358 9536 3334
rect 9600 2666 9628 5102
rect 9678 4992 9734 5001
rect 9678 4927 9734 4936
rect 9692 3058 9720 4927
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9600 2638 9720 2666
rect 9692 2258 9720 2638
rect 9784 2417 9812 5743
rect 9876 2446 9904 5902
rect 9968 3602 9996 6802
rect 10428 6225 10456 11494
rect 16592 10470 16620 12271
rect 20718 11928 20774 11937
rect 20718 11863 20774 11872
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 11058 9888 11114 9897
rect 11058 9823 11114 9832
rect 10874 9480 10930 9489
rect 10874 9415 10930 9424
rect 10414 6216 10470 6225
rect 10414 6151 10470 6160
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 9864 2440 9916 2446
rect 9770 2408 9826 2417
rect 9864 2382 9916 2388
rect 9770 2343 9826 2352
rect 9600 2230 9720 2258
rect 9496 1352 9548 1358
rect 9496 1294 9548 1300
rect 9600 1222 9628 2230
rect 10888 1290 10916 9415
rect 11072 4758 11100 9823
rect 15212 6934 15240 10406
rect 15200 6928 15252 6934
rect 20732 6914 20760 11863
rect 21362 11112 21418 11121
rect 21362 11047 21418 11056
rect 15200 6870 15252 6876
rect 20640 6886 20760 6914
rect 16580 5092 16632 5098
rect 16580 5034 16632 5040
rect 11060 4752 11112 4758
rect 11060 4694 11112 4700
rect 13818 4584 13874 4593
rect 13818 4519 13874 4528
rect 13832 3466 13860 4519
rect 16592 4185 16620 5034
rect 20640 4758 20668 6886
rect 17776 4752 17828 4758
rect 17776 4694 17828 4700
rect 20628 4752 20680 4758
rect 20628 4694 20680 4700
rect 16578 4176 16634 4185
rect 16578 4111 16634 4120
rect 16578 3768 16634 3777
rect 16578 3703 16580 3712
rect 16632 3703 16634 3712
rect 16580 3674 16632 3680
rect 13820 3460 13872 3466
rect 13820 3402 13872 3408
rect 16578 2952 16634 2961
rect 16578 2887 16634 2896
rect 16592 2854 16620 2887
rect 16580 2848 16632 2854
rect 16580 2790 16632 2796
rect 16578 2544 16634 2553
rect 17788 2514 17816 4694
rect 16578 2479 16634 2488
rect 17776 2508 17828 2514
rect 16592 1834 16620 2479
rect 17776 2450 17828 2456
rect 16580 1828 16632 1834
rect 16580 1770 16632 1776
rect 21376 1766 21404 11047
rect 21364 1760 21416 1766
rect 13818 1728 13874 1737
rect 21364 1702 21416 1708
rect 13818 1663 13874 1672
rect 13832 1358 13860 1663
rect 13820 1352 13872 1358
rect 13820 1294 13872 1300
rect 10876 1284 10928 1290
rect 10876 1226 10928 1232
rect 9588 1216 9640 1222
rect 9588 1158 9640 1164
rect 9310 912 9366 921
rect 9310 847 9366 856
rect 9218 504 9274 513
rect 9218 439 9274 448
<< via2 >>
rect 16578 12280 16634 12336
rect 846 7792 902 7848
rect 1122 10920 1178 10976
rect 1398 10784 1454 10840
rect 1490 10648 1546 10704
rect 1582 10512 1638 10568
rect 2572 11450 2628 11452
rect 2652 11450 2708 11452
rect 2732 11450 2788 11452
rect 2812 11450 2868 11452
rect 2572 11398 2618 11450
rect 2618 11398 2628 11450
rect 2652 11398 2682 11450
rect 2682 11398 2694 11450
rect 2694 11398 2708 11450
rect 2732 11398 2746 11450
rect 2746 11398 2758 11450
rect 2758 11398 2788 11450
rect 2812 11398 2822 11450
rect 2822 11398 2868 11450
rect 2572 11396 2628 11398
rect 2652 11396 2708 11398
rect 2732 11396 2788 11398
rect 2812 11396 2868 11398
rect 2686 11192 2742 11248
rect 1766 9016 1822 9072
rect 1490 7112 1546 7168
rect 2042 8336 2098 8392
rect 2572 10362 2628 10364
rect 2652 10362 2708 10364
rect 2732 10362 2788 10364
rect 2812 10362 2868 10364
rect 2572 10310 2618 10362
rect 2618 10310 2628 10362
rect 2652 10310 2682 10362
rect 2682 10310 2694 10362
rect 2694 10310 2708 10362
rect 2732 10310 2746 10362
rect 2746 10310 2758 10362
rect 2758 10310 2788 10362
rect 2812 10310 2822 10362
rect 2822 10310 2868 10362
rect 2572 10308 2628 10310
rect 2652 10308 2708 10310
rect 2732 10308 2788 10310
rect 2812 10308 2868 10310
rect 2686 9988 2742 10024
rect 2686 9968 2688 9988
rect 2688 9968 2740 9988
rect 2740 9968 2742 9988
rect 2572 9274 2628 9276
rect 2652 9274 2708 9276
rect 2732 9274 2788 9276
rect 2812 9274 2868 9276
rect 2572 9222 2618 9274
rect 2618 9222 2628 9274
rect 2652 9222 2682 9274
rect 2682 9222 2694 9274
rect 2694 9222 2708 9274
rect 2732 9222 2746 9274
rect 2746 9222 2758 9274
rect 2758 9222 2788 9274
rect 2812 9222 2822 9274
rect 2822 9222 2868 9274
rect 2572 9220 2628 9222
rect 2652 9220 2708 9222
rect 2732 9220 2788 9222
rect 2812 9220 2868 9222
rect 2686 9016 2742 9072
rect 2870 9016 2926 9072
rect 1674 5480 1730 5536
rect 1950 6160 2006 6216
rect 2226 6296 2282 6352
rect 3146 9424 3202 9480
rect 3330 9968 3386 10024
rect 2572 8186 2628 8188
rect 2652 8186 2708 8188
rect 2732 8186 2788 8188
rect 2812 8186 2868 8188
rect 2572 8134 2618 8186
rect 2618 8134 2628 8186
rect 2652 8134 2682 8186
rect 2682 8134 2694 8186
rect 2694 8134 2708 8186
rect 2732 8134 2746 8186
rect 2746 8134 2758 8186
rect 2758 8134 2788 8186
rect 2812 8134 2822 8186
rect 2822 8134 2868 8186
rect 2572 8132 2628 8134
rect 2652 8132 2708 8134
rect 2732 8132 2788 8134
rect 2812 8132 2868 8134
rect 2686 7928 2742 7984
rect 2572 7098 2628 7100
rect 2652 7098 2708 7100
rect 2732 7098 2788 7100
rect 2812 7098 2868 7100
rect 2572 7046 2618 7098
rect 2618 7046 2628 7098
rect 2652 7046 2682 7098
rect 2682 7046 2694 7098
rect 2694 7046 2708 7098
rect 2732 7046 2746 7098
rect 2746 7046 2758 7098
rect 2758 7046 2788 7098
rect 2812 7046 2822 7098
rect 2822 7046 2868 7098
rect 2572 7044 2628 7046
rect 2652 7044 2708 7046
rect 2732 7044 2788 7046
rect 2812 7044 2868 7046
rect 3054 7928 3110 7984
rect 2962 6704 3018 6760
rect 2572 6010 2628 6012
rect 2652 6010 2708 6012
rect 2732 6010 2788 6012
rect 2812 6010 2868 6012
rect 2572 5958 2618 6010
rect 2618 5958 2628 6010
rect 2652 5958 2682 6010
rect 2682 5958 2694 6010
rect 2694 5958 2708 6010
rect 2732 5958 2746 6010
rect 2746 5958 2758 6010
rect 2758 5958 2788 6010
rect 2812 5958 2822 6010
rect 2822 5958 2868 6010
rect 2572 5956 2628 5958
rect 2652 5956 2708 5958
rect 2732 5956 2788 5958
rect 2812 5956 2868 5958
rect 2778 5752 2834 5808
rect 3606 9832 3662 9888
rect 3882 10920 3938 10976
rect 4122 10906 4178 10908
rect 4202 10906 4258 10908
rect 4282 10906 4338 10908
rect 4362 10906 4418 10908
rect 4122 10854 4168 10906
rect 4168 10854 4178 10906
rect 4202 10854 4232 10906
rect 4232 10854 4244 10906
rect 4244 10854 4258 10906
rect 4282 10854 4296 10906
rect 4296 10854 4308 10906
rect 4308 10854 4338 10906
rect 4362 10854 4372 10906
rect 4372 10854 4418 10906
rect 4122 10852 4178 10854
rect 4202 10852 4258 10854
rect 4282 10852 4338 10854
rect 4362 10852 4418 10854
rect 3974 10784 4030 10840
rect 4526 10784 4582 10840
rect 3882 10240 3938 10296
rect 3974 10104 4030 10160
rect 4342 10532 4398 10568
rect 4342 10512 4344 10532
rect 4344 10512 4396 10532
rect 4396 10512 4398 10532
rect 5078 11092 5080 11112
rect 5080 11092 5132 11112
rect 5132 11092 5134 11112
rect 5078 11056 5134 11092
rect 4434 10104 4490 10160
rect 4618 10104 4674 10160
rect 4802 10240 4858 10296
rect 4986 10512 5042 10568
rect 3238 7248 3294 7304
rect 2410 5616 2466 5672
rect 2410 2488 2466 2544
rect 2686 5208 2742 5264
rect 2870 3032 2926 3088
rect 3146 5516 3148 5536
rect 3148 5516 3200 5536
rect 3200 5516 3202 5536
rect 3146 5480 3202 5516
rect 3330 5616 3386 5672
rect 3606 6296 3662 6352
rect 3514 4664 3570 4720
rect 4250 9968 4306 10024
rect 4122 9818 4178 9820
rect 4202 9818 4258 9820
rect 4282 9818 4338 9820
rect 4362 9818 4418 9820
rect 4122 9766 4168 9818
rect 4168 9766 4178 9818
rect 4202 9766 4232 9818
rect 4232 9766 4244 9818
rect 4244 9766 4258 9818
rect 4282 9766 4296 9818
rect 4296 9766 4308 9818
rect 4308 9766 4338 9818
rect 4362 9766 4372 9818
rect 4372 9766 4418 9818
rect 4122 9764 4178 9766
rect 4202 9764 4258 9766
rect 4282 9764 4338 9766
rect 4362 9764 4418 9766
rect 4618 9696 4674 9752
rect 3790 7248 3846 7304
rect 4122 8730 4178 8732
rect 4202 8730 4258 8732
rect 4282 8730 4338 8732
rect 4362 8730 4418 8732
rect 4122 8678 4168 8730
rect 4168 8678 4178 8730
rect 4202 8678 4232 8730
rect 4232 8678 4244 8730
rect 4244 8678 4258 8730
rect 4282 8678 4296 8730
rect 4296 8678 4308 8730
rect 4308 8678 4338 8730
rect 4362 8678 4372 8730
rect 4372 8678 4418 8730
rect 4122 8676 4178 8678
rect 4202 8676 4258 8678
rect 4282 8676 4338 8678
rect 4362 8676 4418 8678
rect 4342 8472 4398 8528
rect 4066 8336 4122 8392
rect 4710 9560 4766 9616
rect 4618 8336 4674 8392
rect 4526 7928 4582 7984
rect 4122 7642 4178 7644
rect 4202 7642 4258 7644
rect 4282 7642 4338 7644
rect 4362 7642 4418 7644
rect 4122 7590 4168 7642
rect 4168 7590 4178 7642
rect 4202 7590 4232 7642
rect 4232 7590 4244 7642
rect 4244 7590 4258 7642
rect 4282 7590 4296 7642
rect 4296 7590 4308 7642
rect 4308 7590 4338 7642
rect 4362 7590 4372 7642
rect 4372 7590 4418 7642
rect 4122 7588 4178 7590
rect 4202 7588 4258 7590
rect 4282 7588 4338 7590
rect 4362 7588 4418 7590
rect 3882 6840 3938 6896
rect 3882 6704 3938 6760
rect 3790 6160 3846 6216
rect 4122 6554 4178 6556
rect 4202 6554 4258 6556
rect 4282 6554 4338 6556
rect 4362 6554 4418 6556
rect 4122 6502 4168 6554
rect 4168 6502 4178 6554
rect 4202 6502 4232 6554
rect 4232 6502 4244 6554
rect 4244 6502 4258 6554
rect 4282 6502 4296 6554
rect 4296 6502 4308 6554
rect 4308 6502 4338 6554
rect 4362 6502 4372 6554
rect 4372 6502 4418 6554
rect 4122 6500 4178 6502
rect 4202 6500 4258 6502
rect 4282 6500 4338 6502
rect 4362 6500 4418 6502
rect 4158 6296 4214 6352
rect 4158 5788 4160 5808
rect 4160 5788 4212 5808
rect 4212 5788 4214 5808
rect 4158 5752 4214 5788
rect 4250 5652 4252 5672
rect 4252 5652 4304 5672
rect 4304 5652 4306 5672
rect 4250 5616 4306 5652
rect 4122 5466 4178 5468
rect 4202 5466 4258 5468
rect 4282 5466 4338 5468
rect 4362 5466 4418 5468
rect 4122 5414 4168 5466
rect 4168 5414 4178 5466
rect 4202 5414 4232 5466
rect 4232 5414 4244 5466
rect 4244 5414 4258 5466
rect 4282 5414 4296 5466
rect 4296 5414 4308 5466
rect 4308 5414 4338 5466
rect 4362 5414 4372 5466
rect 4372 5414 4418 5466
rect 4122 5412 4178 5414
rect 4202 5412 4258 5414
rect 4282 5412 4338 5414
rect 4362 5412 4418 5414
rect 4122 4378 4178 4380
rect 4202 4378 4258 4380
rect 4282 4378 4338 4380
rect 4362 4378 4418 4380
rect 4122 4326 4168 4378
rect 4168 4326 4178 4378
rect 4202 4326 4232 4378
rect 4232 4326 4244 4378
rect 4244 4326 4258 4378
rect 4282 4326 4296 4378
rect 4296 4326 4308 4378
rect 4308 4326 4338 4378
rect 4362 4326 4372 4378
rect 4372 4326 4418 4378
rect 4122 4324 4178 4326
rect 4202 4324 4258 4326
rect 4282 4324 4338 4326
rect 4362 4324 4418 4326
rect 3974 3576 4030 3632
rect 4894 8472 4950 8528
rect 4802 7248 4858 7304
rect 5078 9632 5134 9688
rect 5170 9444 5226 9480
rect 5170 9424 5172 9444
rect 5172 9424 5224 9444
rect 5224 9424 5226 9444
rect 3882 3188 3938 3224
rect 3882 3168 3884 3188
rect 3884 3168 3936 3188
rect 3936 3168 3938 3188
rect 4122 3290 4178 3292
rect 4202 3290 4258 3292
rect 4282 3290 4338 3292
rect 4362 3290 4418 3292
rect 4122 3238 4168 3290
rect 4168 3238 4178 3290
rect 4202 3238 4232 3290
rect 4232 3238 4244 3290
rect 4244 3238 4258 3290
rect 4282 3238 4296 3290
rect 4296 3238 4308 3290
rect 4308 3238 4338 3290
rect 4362 3238 4372 3290
rect 4372 3238 4418 3290
rect 4122 3236 4178 3238
rect 4202 3236 4258 3238
rect 4282 3236 4338 3238
rect 4362 3236 4418 3238
rect 4618 3304 4674 3360
rect 5262 7792 5318 7848
rect 4122 2202 4178 2204
rect 4202 2202 4258 2204
rect 4282 2202 4338 2204
rect 4362 2202 4418 2204
rect 4122 2150 4168 2202
rect 4168 2150 4178 2202
rect 4202 2150 4232 2202
rect 4232 2150 4244 2202
rect 4244 2150 4258 2202
rect 4282 2150 4296 2202
rect 4296 2150 4308 2202
rect 4308 2150 4338 2202
rect 4362 2150 4372 2202
rect 4372 2150 4418 2202
rect 4122 2148 4178 2150
rect 4202 2148 4258 2150
rect 4282 2148 4338 2150
rect 4362 2148 4418 2150
rect 5446 11600 5502 11656
rect 5446 10784 5502 10840
rect 5672 11450 5728 11452
rect 5752 11450 5808 11452
rect 5832 11450 5888 11452
rect 5912 11450 5968 11452
rect 5672 11398 5718 11450
rect 5718 11398 5728 11450
rect 5752 11398 5782 11450
rect 5782 11398 5794 11450
rect 5794 11398 5808 11450
rect 5832 11398 5846 11450
rect 5846 11398 5858 11450
rect 5858 11398 5888 11450
rect 5912 11398 5922 11450
rect 5922 11398 5968 11450
rect 5672 11396 5728 11398
rect 5752 11396 5808 11398
rect 5832 11396 5888 11398
rect 5912 11396 5968 11398
rect 5538 10512 5594 10568
rect 5906 10512 5962 10568
rect 5672 10362 5728 10364
rect 5752 10362 5808 10364
rect 5832 10362 5888 10364
rect 5912 10362 5968 10364
rect 5672 10310 5718 10362
rect 5718 10310 5728 10362
rect 5752 10310 5782 10362
rect 5782 10310 5794 10362
rect 5794 10310 5808 10362
rect 5832 10310 5846 10362
rect 5846 10310 5858 10362
rect 5858 10310 5888 10362
rect 5912 10310 5922 10362
rect 5922 10310 5968 10362
rect 5672 10308 5728 10310
rect 5752 10308 5808 10310
rect 5832 10308 5888 10310
rect 5912 10308 5968 10310
rect 5630 9696 5686 9752
rect 5722 9560 5778 9616
rect 5630 9424 5686 9480
rect 5672 9274 5728 9276
rect 5752 9274 5808 9276
rect 5832 9274 5888 9276
rect 5912 9274 5968 9276
rect 5672 9222 5718 9274
rect 5718 9222 5728 9274
rect 5752 9222 5782 9274
rect 5782 9222 5794 9274
rect 5794 9222 5808 9274
rect 5832 9222 5846 9274
rect 5846 9222 5858 9274
rect 5858 9222 5888 9274
rect 5912 9222 5922 9274
rect 5922 9222 5968 9274
rect 5672 9220 5728 9222
rect 5752 9220 5808 9222
rect 5832 9220 5888 9222
rect 5912 9220 5968 9222
rect 6182 9424 6238 9480
rect 6182 8472 6238 8528
rect 5672 8186 5728 8188
rect 5752 8186 5808 8188
rect 5832 8186 5888 8188
rect 5912 8186 5968 8188
rect 5672 8134 5718 8186
rect 5718 8134 5728 8186
rect 5752 8134 5782 8186
rect 5782 8134 5794 8186
rect 5794 8134 5808 8186
rect 5832 8134 5846 8186
rect 5846 8134 5858 8186
rect 5858 8134 5888 8186
rect 5912 8134 5922 8186
rect 5922 8134 5968 8186
rect 5672 8132 5728 8134
rect 5752 8132 5808 8134
rect 5832 8132 5888 8134
rect 5912 8132 5968 8134
rect 5672 7098 5728 7100
rect 5752 7098 5808 7100
rect 5832 7098 5888 7100
rect 5912 7098 5968 7100
rect 5672 7046 5718 7098
rect 5718 7046 5728 7098
rect 5752 7046 5782 7098
rect 5782 7046 5794 7098
rect 5794 7046 5808 7098
rect 5832 7046 5846 7098
rect 5846 7046 5858 7098
rect 5858 7046 5888 7098
rect 5912 7046 5922 7098
rect 5922 7046 5968 7098
rect 5672 7044 5728 7046
rect 5752 7044 5808 7046
rect 5832 7044 5888 7046
rect 5912 7044 5968 7046
rect 5814 6568 5870 6624
rect 6090 6724 6146 6760
rect 6090 6704 6092 6724
rect 6092 6704 6144 6724
rect 6144 6704 6146 6724
rect 5630 6160 5686 6216
rect 5672 6010 5728 6012
rect 5752 6010 5808 6012
rect 5832 6010 5888 6012
rect 5912 6010 5968 6012
rect 5672 5958 5718 6010
rect 5718 5958 5728 6010
rect 5752 5958 5782 6010
rect 5782 5958 5794 6010
rect 5794 5958 5808 6010
rect 5832 5958 5846 6010
rect 5846 5958 5858 6010
rect 5858 5958 5888 6010
rect 5912 5958 5922 6010
rect 5922 5958 5968 6010
rect 5672 5956 5728 5958
rect 5752 5956 5808 5958
rect 5832 5956 5888 5958
rect 5912 5956 5968 5958
rect 5906 5208 5962 5264
rect 5446 3576 5502 3632
rect 5354 3304 5410 3360
rect 5672 4922 5728 4924
rect 5752 4922 5808 4924
rect 5832 4922 5888 4924
rect 5912 4922 5968 4924
rect 5672 4870 5718 4922
rect 5718 4870 5728 4922
rect 5752 4870 5782 4922
rect 5782 4870 5794 4922
rect 5794 4870 5808 4922
rect 5832 4870 5846 4922
rect 5846 4870 5858 4922
rect 5858 4870 5888 4922
rect 5912 4870 5922 4922
rect 5922 4870 5968 4922
rect 5672 4868 5728 4870
rect 5752 4868 5808 4870
rect 5832 4868 5888 4870
rect 5912 4868 5968 4870
rect 5672 3834 5728 3836
rect 5752 3834 5808 3836
rect 5832 3834 5888 3836
rect 5912 3834 5968 3836
rect 5672 3782 5718 3834
rect 5718 3782 5728 3834
rect 5752 3782 5782 3834
rect 5782 3782 5794 3834
rect 5794 3782 5808 3834
rect 5832 3782 5846 3834
rect 5846 3782 5858 3834
rect 5858 3782 5888 3834
rect 5912 3782 5922 3834
rect 5922 3782 5968 3834
rect 5672 3780 5728 3782
rect 5752 3780 5808 3782
rect 5832 3780 5888 3782
rect 5912 3780 5968 3782
rect 5630 3576 5686 3632
rect 5672 2746 5728 2748
rect 5752 2746 5808 2748
rect 5832 2746 5888 2748
rect 5912 2746 5968 2748
rect 5672 2694 5718 2746
rect 5718 2694 5728 2746
rect 5752 2694 5782 2746
rect 5782 2694 5794 2746
rect 5794 2694 5808 2746
rect 5832 2694 5846 2746
rect 5846 2694 5858 2746
rect 5858 2694 5888 2746
rect 5912 2694 5922 2746
rect 5922 2694 5968 2746
rect 5672 2692 5728 2694
rect 5752 2692 5808 2694
rect 5832 2692 5888 2694
rect 5912 2692 5968 2694
rect 6458 9968 6514 10024
rect 6642 9968 6698 10024
rect 6550 7384 6606 7440
rect 6550 7248 6606 7304
rect 6734 8336 6790 8392
rect 7194 11192 7250 11248
rect 6918 9424 6974 9480
rect 7562 11056 7618 11112
rect 7222 10906 7278 10908
rect 7302 10906 7358 10908
rect 7382 10906 7438 10908
rect 7462 10906 7518 10908
rect 7222 10854 7268 10906
rect 7268 10854 7278 10906
rect 7302 10854 7332 10906
rect 7332 10854 7344 10906
rect 7344 10854 7358 10906
rect 7382 10854 7396 10906
rect 7396 10854 7408 10906
rect 7408 10854 7438 10906
rect 7462 10854 7472 10906
rect 7472 10854 7518 10906
rect 7222 10852 7278 10854
rect 7302 10852 7358 10854
rect 7382 10852 7438 10854
rect 7462 10852 7518 10854
rect 7222 9818 7278 9820
rect 7302 9818 7358 9820
rect 7382 9818 7438 9820
rect 7462 9818 7518 9820
rect 7222 9766 7268 9818
rect 7268 9766 7278 9818
rect 7302 9766 7332 9818
rect 7332 9766 7344 9818
rect 7344 9766 7358 9818
rect 7382 9766 7396 9818
rect 7396 9766 7408 9818
rect 7408 9766 7438 9818
rect 7462 9766 7472 9818
rect 7472 9766 7518 9818
rect 7222 9764 7278 9766
rect 7302 9764 7358 9766
rect 7382 9764 7438 9766
rect 7462 9764 7518 9766
rect 7222 8730 7278 8732
rect 7302 8730 7358 8732
rect 7382 8730 7438 8732
rect 7462 8730 7518 8732
rect 7222 8678 7268 8730
rect 7268 8678 7278 8730
rect 7302 8678 7332 8730
rect 7332 8678 7344 8730
rect 7344 8678 7358 8730
rect 7382 8678 7396 8730
rect 7396 8678 7408 8730
rect 7408 8678 7438 8730
rect 7462 8678 7472 8730
rect 7472 8678 7518 8730
rect 7222 8676 7278 8678
rect 7302 8676 7358 8678
rect 7382 8676 7438 8678
rect 7462 8676 7518 8678
rect 7194 8472 7250 8528
rect 7222 7642 7278 7644
rect 7302 7642 7358 7644
rect 7382 7642 7438 7644
rect 7462 7642 7518 7644
rect 7222 7590 7268 7642
rect 7268 7590 7278 7642
rect 7302 7590 7332 7642
rect 7332 7590 7344 7642
rect 7344 7590 7358 7642
rect 7382 7590 7396 7642
rect 7396 7590 7408 7642
rect 7408 7590 7438 7642
rect 7462 7590 7472 7642
rect 7472 7590 7518 7642
rect 7222 7588 7278 7590
rect 7302 7588 7358 7590
rect 7382 7588 7438 7590
rect 7462 7588 7518 7590
rect 7010 6568 7066 6624
rect 7194 6704 7250 6760
rect 7222 6554 7278 6556
rect 7302 6554 7358 6556
rect 7382 6554 7438 6556
rect 7462 6554 7518 6556
rect 7222 6502 7268 6554
rect 7268 6502 7278 6554
rect 7302 6502 7332 6554
rect 7332 6502 7344 6554
rect 7344 6502 7358 6554
rect 7382 6502 7396 6554
rect 7396 6502 7408 6554
rect 7408 6502 7438 6554
rect 7462 6502 7472 6554
rect 7472 6502 7518 6554
rect 7222 6500 7278 6502
rect 7302 6500 7358 6502
rect 7382 6500 7438 6502
rect 7462 6500 7518 6502
rect 7102 6160 7158 6216
rect 6918 5208 6974 5264
rect 7222 5466 7278 5468
rect 7302 5466 7358 5468
rect 7382 5466 7438 5468
rect 7462 5466 7518 5468
rect 7222 5414 7268 5466
rect 7268 5414 7278 5466
rect 7302 5414 7332 5466
rect 7332 5414 7344 5466
rect 7344 5414 7358 5466
rect 7382 5414 7396 5466
rect 7396 5414 7408 5466
rect 7408 5414 7438 5466
rect 7462 5414 7472 5466
rect 7472 5414 7518 5466
rect 7222 5412 7278 5414
rect 7302 5412 7358 5414
rect 7382 5412 7438 5414
rect 7462 5412 7518 5414
rect 7194 4664 7250 4720
rect 6918 4140 6974 4176
rect 6918 4120 6920 4140
rect 6920 4120 6972 4140
rect 6972 4120 6974 4140
rect 6642 3576 6698 3632
rect 6826 3032 6882 3088
rect 7222 4378 7278 4380
rect 7302 4378 7358 4380
rect 7382 4378 7438 4380
rect 7462 4378 7518 4380
rect 7222 4326 7268 4378
rect 7268 4326 7278 4378
rect 7302 4326 7332 4378
rect 7332 4326 7344 4378
rect 7344 4326 7358 4378
rect 7382 4326 7396 4378
rect 7396 4326 7408 4378
rect 7408 4326 7438 4378
rect 7462 4326 7472 4378
rect 7472 4326 7518 4378
rect 7222 4324 7278 4326
rect 7302 4324 7358 4326
rect 7382 4324 7438 4326
rect 7462 4324 7518 4326
rect 7378 3596 7434 3632
rect 7378 3576 7380 3596
rect 7380 3576 7432 3596
rect 7432 3576 7434 3596
rect 7222 3290 7278 3292
rect 7302 3290 7358 3292
rect 7382 3290 7438 3292
rect 7462 3290 7518 3292
rect 7222 3238 7268 3290
rect 7268 3238 7278 3290
rect 7302 3238 7332 3290
rect 7332 3238 7344 3290
rect 7344 3238 7358 3290
rect 7382 3238 7396 3290
rect 7396 3238 7408 3290
rect 7408 3238 7438 3290
rect 7462 3238 7472 3290
rect 7472 3238 7518 3290
rect 7222 3236 7278 3238
rect 7302 3236 7358 3238
rect 7382 3236 7438 3238
rect 7462 3236 7518 3238
rect 7194 3032 7250 3088
rect 7378 2508 7434 2544
rect 7378 2488 7380 2508
rect 7380 2488 7432 2508
rect 7432 2488 7434 2508
rect 7222 2202 7278 2204
rect 7302 2202 7358 2204
rect 7382 2202 7438 2204
rect 7462 2202 7518 2204
rect 7222 2150 7268 2202
rect 7268 2150 7278 2202
rect 7302 2150 7332 2202
rect 7332 2150 7344 2202
rect 7344 2150 7358 2202
rect 7382 2150 7396 2202
rect 7396 2150 7408 2202
rect 7408 2150 7438 2202
rect 7462 2150 7472 2202
rect 7472 2150 7518 2202
rect 7222 2148 7278 2150
rect 7302 2148 7358 2150
rect 7382 2148 7438 2150
rect 7462 2148 7518 2150
rect 5672 1658 5728 1660
rect 5752 1658 5808 1660
rect 5832 1658 5888 1660
rect 5912 1658 5968 1660
rect 5672 1606 5718 1658
rect 5718 1606 5728 1658
rect 5752 1606 5782 1658
rect 5782 1606 5794 1658
rect 5794 1606 5808 1658
rect 5832 1606 5846 1658
rect 5846 1606 5858 1658
rect 5858 1606 5888 1658
rect 5912 1606 5922 1658
rect 5922 1606 5968 1658
rect 5672 1604 5728 1606
rect 5752 1604 5808 1606
rect 5832 1604 5888 1606
rect 5912 1604 5968 1606
rect 8022 10668 8078 10704
rect 8022 10648 8024 10668
rect 8024 10648 8076 10668
rect 8076 10648 8078 10668
rect 8114 10104 8170 10160
rect 8022 10004 8024 10024
rect 8024 10004 8076 10024
rect 8076 10004 8078 10024
rect 8022 9968 8078 10004
rect 7746 6704 7802 6760
rect 7930 9016 7986 9072
rect 8114 9560 8170 9616
rect 8298 9968 8354 10024
rect 8772 11450 8828 11452
rect 8852 11450 8908 11452
rect 8932 11450 8988 11452
rect 9012 11450 9068 11452
rect 8772 11398 8818 11450
rect 8818 11398 8828 11450
rect 8852 11398 8882 11450
rect 8882 11398 8894 11450
rect 8894 11398 8908 11450
rect 8932 11398 8946 11450
rect 8946 11398 8958 11450
rect 8958 11398 8988 11450
rect 9012 11398 9022 11450
rect 9022 11398 9068 11450
rect 8772 11396 8828 11398
rect 8852 11396 8908 11398
rect 8932 11396 8988 11398
rect 9012 11396 9068 11398
rect 7930 3440 7986 3496
rect 7746 2352 7802 2408
rect 8206 7112 8262 7168
rect 8206 5752 8262 5808
rect 8574 10648 8630 10704
rect 8772 10362 8828 10364
rect 8852 10362 8908 10364
rect 8932 10362 8988 10364
rect 9012 10362 9068 10364
rect 8772 10310 8818 10362
rect 8818 10310 8828 10362
rect 8852 10310 8882 10362
rect 8882 10310 8894 10362
rect 8894 10310 8908 10362
rect 8932 10310 8946 10362
rect 8946 10310 8958 10362
rect 8958 10310 8988 10362
rect 9012 10310 9022 10362
rect 9022 10310 9068 10362
rect 8772 10308 8828 10310
rect 8852 10308 8908 10310
rect 8932 10308 8988 10310
rect 9012 10308 9068 10310
rect 9586 10648 9642 10704
rect 8850 10004 8852 10024
rect 8852 10004 8904 10024
rect 8904 10004 8906 10024
rect 8850 9968 8906 10004
rect 9034 10104 9090 10160
rect 8772 9274 8828 9276
rect 8852 9274 8908 9276
rect 8932 9274 8988 9276
rect 9012 9274 9068 9276
rect 8772 9222 8818 9274
rect 8818 9222 8828 9274
rect 8852 9222 8882 9274
rect 8882 9222 8894 9274
rect 8894 9222 8908 9274
rect 8932 9222 8946 9274
rect 8946 9222 8958 9274
rect 8958 9222 8988 9274
rect 9012 9222 9022 9274
rect 9022 9222 9068 9274
rect 8772 9220 8828 9222
rect 8852 9220 8908 9222
rect 8932 9220 8988 9222
rect 9012 9220 9068 9222
rect 8772 8186 8828 8188
rect 8852 8186 8908 8188
rect 8932 8186 8988 8188
rect 9012 8186 9068 8188
rect 8772 8134 8818 8186
rect 8818 8134 8828 8186
rect 8852 8134 8882 8186
rect 8882 8134 8894 8186
rect 8894 8134 8908 8186
rect 8932 8134 8946 8186
rect 8946 8134 8958 8186
rect 8958 8134 8988 8186
rect 9012 8134 9022 8186
rect 9022 8134 9068 8186
rect 8772 8132 8828 8134
rect 8852 8132 8908 8134
rect 8932 8132 8988 8134
rect 9012 8132 9068 8134
rect 8772 7098 8828 7100
rect 8852 7098 8908 7100
rect 8932 7098 8988 7100
rect 9012 7098 9068 7100
rect 8772 7046 8818 7098
rect 8818 7046 8828 7098
rect 8852 7046 8882 7098
rect 8882 7046 8894 7098
rect 8894 7046 8908 7098
rect 8932 7046 8946 7098
rect 8946 7046 8958 7098
rect 8958 7046 8988 7098
rect 9012 7046 9022 7098
rect 9022 7046 9068 7098
rect 8772 7044 8828 7046
rect 8852 7044 8908 7046
rect 8932 7044 8988 7046
rect 9012 7044 9068 7046
rect 8772 6010 8828 6012
rect 8852 6010 8908 6012
rect 8932 6010 8988 6012
rect 9012 6010 9068 6012
rect 8772 5958 8818 6010
rect 8818 5958 8828 6010
rect 8852 5958 8882 6010
rect 8882 5958 8894 6010
rect 8894 5958 8908 6010
rect 8932 5958 8946 6010
rect 8946 5958 8958 6010
rect 8958 5958 8988 6010
rect 9012 5958 9022 6010
rect 9022 5958 9068 6010
rect 8772 5956 8828 5958
rect 8852 5956 8908 5958
rect 8932 5956 8988 5958
rect 9012 5956 9068 5958
rect 9494 9832 9550 9888
rect 9402 8200 9458 8256
rect 8206 4256 8262 4312
rect 8574 4392 8630 4448
rect 8298 3032 8354 3088
rect 8298 2896 8354 2952
rect 8772 4922 8828 4924
rect 8852 4922 8908 4924
rect 8932 4922 8988 4924
rect 9012 4922 9068 4924
rect 8772 4870 8818 4922
rect 8818 4870 8828 4922
rect 8852 4870 8882 4922
rect 8882 4870 8894 4922
rect 8894 4870 8908 4922
rect 8932 4870 8946 4922
rect 8946 4870 8958 4922
rect 8958 4870 8988 4922
rect 9012 4870 9022 4922
rect 9022 4870 9068 4922
rect 8772 4868 8828 4870
rect 8852 4868 8908 4870
rect 8932 4868 8988 4870
rect 9012 4868 9068 4870
rect 8772 3834 8828 3836
rect 8852 3834 8908 3836
rect 8932 3834 8988 3836
rect 9012 3834 9068 3836
rect 8772 3782 8818 3834
rect 8818 3782 8828 3834
rect 8852 3782 8882 3834
rect 8882 3782 8894 3834
rect 8894 3782 8908 3834
rect 8932 3782 8946 3834
rect 8946 3782 8958 3834
rect 8958 3782 8988 3834
rect 9012 3782 9022 3834
rect 9022 3782 9068 3834
rect 8772 3780 8828 3782
rect 8852 3780 8908 3782
rect 8932 3780 8988 3782
rect 9012 3780 9068 3782
rect 8666 3168 8722 3224
rect 8574 3032 8630 3088
rect 9310 6160 9366 6216
rect 9218 3732 9274 3768
rect 9218 3712 9220 3732
rect 9220 3712 9272 3732
rect 9272 3712 9274 3732
rect 9218 3576 9274 3632
rect 8772 2746 8828 2748
rect 8852 2746 8908 2748
rect 8932 2746 8988 2748
rect 9012 2746 9068 2748
rect 8772 2694 8818 2746
rect 8818 2694 8828 2746
rect 8852 2694 8882 2746
rect 8882 2694 8894 2746
rect 8894 2694 8908 2746
rect 8932 2694 8946 2746
rect 8946 2694 8958 2746
rect 8958 2694 8988 2746
rect 9012 2694 9022 2746
rect 9022 2694 9068 2746
rect 8772 2692 8828 2694
rect 8852 2692 8908 2694
rect 8932 2692 8988 2694
rect 9012 2692 9068 2694
rect 8850 2524 8852 2544
rect 8852 2524 8904 2544
rect 8904 2524 8906 2544
rect 8850 2488 8906 2524
rect 9126 2080 9182 2136
rect 8772 1658 8828 1660
rect 8852 1658 8908 1660
rect 8932 1658 8988 1660
rect 9012 1658 9068 1660
rect 8772 1606 8818 1658
rect 8818 1606 8828 1658
rect 8852 1606 8882 1658
rect 8882 1606 8894 1658
rect 8894 1606 8908 1658
rect 8932 1606 8946 1658
rect 8946 1606 8958 1658
rect 8958 1606 8988 1658
rect 9012 1606 9022 1658
rect 9022 1606 9068 1658
rect 8772 1604 8828 1606
rect 8852 1604 8908 1606
rect 8932 1604 8988 1606
rect 9012 1604 9068 1606
rect 8942 1264 8998 1320
rect 4122 1114 4178 1116
rect 4202 1114 4258 1116
rect 4282 1114 4338 1116
rect 4362 1114 4418 1116
rect 4122 1062 4168 1114
rect 4168 1062 4178 1114
rect 4202 1062 4232 1114
rect 4232 1062 4244 1114
rect 4244 1062 4258 1114
rect 4282 1062 4296 1114
rect 4296 1062 4308 1114
rect 4308 1062 4338 1114
rect 4362 1062 4372 1114
rect 4372 1062 4418 1114
rect 4122 1060 4178 1062
rect 4202 1060 4258 1062
rect 4282 1060 4338 1062
rect 4362 1060 4418 1062
rect 7222 1114 7278 1116
rect 7302 1114 7358 1116
rect 7382 1114 7438 1116
rect 7462 1114 7518 1116
rect 7222 1062 7268 1114
rect 7268 1062 7278 1114
rect 7302 1062 7332 1114
rect 7332 1062 7344 1114
rect 7344 1062 7358 1114
rect 7382 1062 7396 1114
rect 7396 1062 7408 1114
rect 7408 1062 7438 1114
rect 7462 1062 7472 1114
rect 7472 1062 7518 1114
rect 7222 1060 7278 1062
rect 7302 1060 7358 1062
rect 7382 1060 7438 1062
rect 7462 1060 7518 1062
rect 9862 7792 9918 7848
rect 9678 7384 9734 7440
rect 9770 5752 9826 5808
rect 9678 4936 9734 4992
rect 20718 11872 20774 11928
rect 11058 9832 11114 9888
rect 10874 9424 10930 9480
rect 10414 6160 10470 6216
rect 9770 2352 9826 2408
rect 21362 11056 21418 11112
rect 13818 4528 13874 4584
rect 16578 4120 16634 4176
rect 16578 3732 16634 3768
rect 16578 3712 16580 3732
rect 16580 3712 16632 3732
rect 16632 3712 16634 3732
rect 16578 2896 16634 2952
rect 16578 2488 16634 2544
rect 13818 1672 13874 1728
rect 9310 856 9366 912
rect 9218 448 9274 504
<< metal3 >>
rect 14000 12336 34000 12368
rect 14000 12280 16578 12336
rect 16634 12280 34000 12336
rect 14000 12248 34000 12280
rect 14000 11928 34000 11960
rect 14000 11872 20718 11928
rect 20774 11872 34000 11928
rect 14000 11840 34000 11872
rect 5441 11658 5507 11661
rect 5441 11656 12450 11658
rect 5441 11600 5446 11656
rect 5502 11600 12450 11656
rect 5441 11598 12450 11600
rect 5441 11595 5507 11598
rect 12390 11522 12450 11598
rect 14000 11522 34000 11552
rect 12390 11462 34000 11522
rect 2560 11456 2880 11457
rect 2560 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2880 11456
rect 2560 11391 2880 11392
rect 5660 11456 5980 11457
rect 5660 11392 5668 11456
rect 5732 11392 5748 11456
rect 5812 11392 5828 11456
rect 5892 11392 5908 11456
rect 5972 11392 5980 11456
rect 5660 11391 5980 11392
rect 8760 11456 9080 11457
rect 8760 11392 8768 11456
rect 8832 11392 8848 11456
rect 8912 11392 8928 11456
rect 8992 11392 9008 11456
rect 9072 11392 9080 11456
rect 14000 11432 34000 11462
rect 8760 11391 9080 11392
rect 2681 11250 2747 11253
rect 7189 11250 7255 11253
rect 2681 11248 7255 11250
rect 2681 11192 2686 11248
rect 2742 11192 7194 11248
rect 7250 11192 7255 11248
rect 2681 11190 7255 11192
rect 2681 11187 2747 11190
rect 7189 11187 7255 11190
rect 5073 11114 5139 11117
rect 7557 11114 7623 11117
rect 5073 11112 7623 11114
rect 5073 11056 5078 11112
rect 5134 11056 7562 11112
rect 7618 11056 7623 11112
rect 5073 11054 7623 11056
rect 5073 11051 5139 11054
rect 7557 11051 7623 11054
rect 14000 11112 34000 11144
rect 14000 11056 21362 11112
rect 21418 11056 34000 11112
rect 14000 11024 34000 11056
rect 1117 10978 1183 10981
rect 3877 10978 3943 10981
rect 1117 10976 3943 10978
rect 1117 10920 1122 10976
rect 1178 10920 3882 10976
rect 3938 10920 3943 10976
rect 1117 10918 3943 10920
rect 1117 10915 1183 10918
rect 3877 10915 3943 10918
rect 4110 10912 4430 10913
rect 4110 10848 4118 10912
rect 4182 10848 4198 10912
rect 4262 10848 4278 10912
rect 4342 10848 4358 10912
rect 4422 10848 4430 10912
rect 4110 10847 4430 10848
rect 7210 10912 7530 10913
rect 7210 10848 7218 10912
rect 7282 10848 7298 10912
rect 7362 10848 7378 10912
rect 7442 10848 7458 10912
rect 7522 10848 7530 10912
rect 7210 10847 7530 10848
rect 1393 10842 1459 10845
rect 3969 10842 4035 10845
rect 1393 10840 4035 10842
rect 1393 10784 1398 10840
rect 1454 10784 3974 10840
rect 4030 10784 4035 10840
rect 1393 10782 4035 10784
rect 1393 10779 1459 10782
rect 3969 10779 4035 10782
rect 4521 10842 4587 10845
rect 5441 10842 5507 10845
rect 4521 10840 5507 10842
rect 4521 10784 4526 10840
rect 4582 10784 5446 10840
rect 5502 10784 5507 10840
rect 4521 10782 5507 10784
rect 4521 10779 4587 10782
rect 5441 10779 5507 10782
rect 1485 10706 1551 10709
rect 8017 10706 8083 10709
rect 1485 10704 8083 10706
rect 1485 10648 1490 10704
rect 1546 10648 8022 10704
rect 8078 10648 8083 10704
rect 1485 10646 8083 10648
rect 1485 10643 1551 10646
rect 8017 10643 8083 10646
rect 8569 10706 8635 10709
rect 9581 10706 9647 10709
rect 14000 10706 34000 10736
rect 8569 10704 34000 10706
rect 8569 10648 8574 10704
rect 8630 10648 9586 10704
rect 9642 10648 34000 10704
rect 8569 10646 34000 10648
rect 8569 10643 8635 10646
rect 9581 10643 9647 10646
rect 14000 10616 34000 10646
rect 1577 10570 1643 10573
rect 4337 10570 4403 10573
rect 1577 10568 4403 10570
rect 1577 10512 1582 10568
rect 1638 10512 4342 10568
rect 4398 10512 4403 10568
rect 1577 10510 4403 10512
rect 1577 10507 1643 10510
rect 4337 10507 4403 10510
rect 4981 10568 5047 10573
rect 4981 10512 4986 10568
rect 5042 10512 5047 10568
rect 4981 10507 5047 10512
rect 5533 10568 5599 10573
rect 5533 10512 5538 10568
rect 5594 10512 5599 10568
rect 5533 10507 5599 10512
rect 5901 10570 5967 10573
rect 5901 10568 12450 10570
rect 5901 10512 5906 10568
rect 5962 10512 12450 10568
rect 5901 10510 12450 10512
rect 5901 10507 5967 10510
rect 4984 10434 5044 10507
rect 3558 10374 5044 10434
rect 2560 10368 2880 10369
rect 2560 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2880 10368
rect 2560 10303 2880 10304
rect 2681 10026 2747 10029
rect 3325 10026 3391 10029
rect 2681 10024 3434 10026
rect 2681 9968 2686 10024
rect 2742 9968 3330 10024
rect 3386 9968 3434 10024
rect 2681 9966 3434 9968
rect 2681 9963 2747 9966
rect 3325 9963 3434 9966
rect 3141 9482 3207 9485
rect 3006 9480 3207 9482
rect 3006 9424 3146 9480
rect 3202 9424 3207 9480
rect 3006 9422 3207 9424
rect 3374 9482 3434 9963
rect 3558 9893 3618 10374
rect 3877 10298 3943 10301
rect 4797 10298 4863 10301
rect 3877 10296 4863 10298
rect 3877 10240 3882 10296
rect 3938 10240 4802 10296
rect 4858 10240 4863 10296
rect 3877 10238 4863 10240
rect 3877 10235 3943 10238
rect 4797 10235 4863 10238
rect 3969 10162 4035 10165
rect 4429 10162 4495 10165
rect 3969 10160 4495 10162
rect 3969 10104 3974 10160
rect 4030 10104 4434 10160
rect 4490 10104 4495 10160
rect 3969 10102 4495 10104
rect 3969 10099 4035 10102
rect 4429 10099 4495 10102
rect 4613 10160 4679 10165
rect 4613 10104 4618 10160
rect 4674 10104 4679 10160
rect 4613 10099 4679 10104
rect 4245 10026 4311 10029
rect 3926 10024 4311 10026
rect 3926 9968 4250 10024
rect 4306 9968 4311 10024
rect 3926 9966 4311 9968
rect 3558 9888 3667 9893
rect 3558 9832 3606 9888
rect 3662 9832 3667 9888
rect 3558 9830 3667 9832
rect 3601 9827 3667 9830
rect 3926 9618 3986 9966
rect 4245 9963 4311 9966
rect 4110 9824 4430 9825
rect 4110 9760 4118 9824
rect 4182 9760 4198 9824
rect 4262 9760 4278 9824
rect 4342 9760 4358 9824
rect 4422 9760 4430 9824
rect 4110 9759 4430 9760
rect 4616 9757 4676 10099
rect 5536 10026 5596 10507
rect 5660 10368 5980 10369
rect 5660 10304 5668 10368
rect 5732 10304 5748 10368
rect 5812 10304 5828 10368
rect 5892 10304 5908 10368
rect 5972 10304 5980 10368
rect 5660 10303 5980 10304
rect 8760 10368 9080 10369
rect 8760 10304 8768 10368
rect 8832 10304 8848 10368
rect 8912 10304 8928 10368
rect 8992 10304 9008 10368
rect 9072 10304 9080 10368
rect 8760 10303 9080 10304
rect 12390 10298 12450 10510
rect 14000 10298 34000 10328
rect 12390 10238 34000 10298
rect 14000 10208 34000 10238
rect 8109 10162 8175 10165
rect 9029 10162 9095 10165
rect 8109 10160 9095 10162
rect 8109 10104 8114 10160
rect 8170 10104 9034 10160
rect 9090 10104 9095 10160
rect 8109 10102 9095 10104
rect 8109 10099 8175 10102
rect 9029 10099 9095 10102
rect 6453 10026 6519 10029
rect 5536 10024 6519 10026
rect 5536 9968 6458 10024
rect 6514 9968 6519 10024
rect 5536 9966 6519 9968
rect 6453 9963 6519 9966
rect 6637 10026 6703 10029
rect 8017 10026 8083 10029
rect 8293 10026 8359 10029
rect 8845 10026 8911 10029
rect 6637 10024 7850 10026
rect 6637 9968 6642 10024
rect 6698 9968 7850 10024
rect 6637 9966 7850 9968
rect 6637 9963 6703 9966
rect 7790 9890 7850 9966
rect 8017 10024 8911 10026
rect 8017 9968 8022 10024
rect 8078 9968 8298 10024
rect 8354 9968 8850 10024
rect 8906 9968 8911 10024
rect 8017 9966 8911 9968
rect 8017 9963 8083 9966
rect 8293 9963 8359 9966
rect 8845 9963 8911 9966
rect 9489 9890 9555 9893
rect 7790 9888 9555 9890
rect 7790 9832 9494 9888
rect 9550 9832 9555 9888
rect 7790 9830 9555 9832
rect 9489 9827 9555 9830
rect 11053 9890 11119 9893
rect 14000 9890 34000 9920
rect 11053 9888 34000 9890
rect 11053 9832 11058 9888
rect 11114 9832 34000 9888
rect 11053 9830 34000 9832
rect 11053 9827 11119 9830
rect 7210 9824 7530 9825
rect 7210 9760 7218 9824
rect 7282 9760 7298 9824
rect 7362 9760 7378 9824
rect 7442 9760 7458 9824
rect 7522 9760 7530 9824
rect 14000 9800 34000 9830
rect 7210 9759 7530 9760
rect 4613 9752 4679 9757
rect 5625 9754 5691 9757
rect 4613 9696 4618 9752
rect 4674 9696 4679 9752
rect 4613 9691 4679 9696
rect 5398 9752 5691 9754
rect 5398 9696 5630 9752
rect 5686 9696 5691 9752
rect 5398 9694 5691 9696
rect 5073 9690 5139 9693
rect 5398 9690 5458 9694
rect 5625 9691 5691 9694
rect 5073 9688 5458 9690
rect 5073 9632 5078 9688
rect 5134 9632 5458 9688
rect 5073 9630 5458 9632
rect 5073 9627 5139 9630
rect 4705 9618 4771 9621
rect 3926 9616 4771 9618
rect 3926 9560 4710 9616
rect 4766 9560 4771 9616
rect 3926 9558 4771 9560
rect 4705 9555 4771 9558
rect 5717 9618 5783 9621
rect 8109 9618 8175 9621
rect 5717 9616 8175 9618
rect 5717 9560 5722 9616
rect 5778 9560 8114 9616
rect 8170 9560 8175 9616
rect 5717 9558 8175 9560
rect 5717 9555 5783 9558
rect 8109 9555 8175 9558
rect 5165 9482 5231 9485
rect 3374 9480 5231 9482
rect 3374 9424 5170 9480
rect 5226 9424 5231 9480
rect 3374 9422 5231 9424
rect 2560 9280 2880 9281
rect 2560 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2880 9280
rect 2560 9215 2880 9216
rect 1761 9074 1827 9077
rect 2681 9074 2747 9077
rect 1761 9072 2747 9074
rect 1761 9016 1766 9072
rect 1822 9016 2686 9072
rect 2742 9016 2747 9072
rect 1761 9014 2747 9016
rect 1761 9011 1827 9014
rect 2681 9011 2747 9014
rect 2865 9074 2931 9077
rect 3006 9074 3066 9422
rect 3141 9419 3207 9422
rect 5165 9419 5231 9422
rect 5625 9482 5691 9485
rect 6177 9482 6243 9485
rect 5625 9480 6243 9482
rect 5625 9424 5630 9480
rect 5686 9424 6182 9480
rect 6238 9424 6243 9480
rect 5625 9422 6243 9424
rect 5625 9419 5691 9422
rect 6177 9419 6243 9422
rect 6913 9482 6979 9485
rect 10869 9482 10935 9485
rect 14000 9482 34000 9512
rect 6913 9480 7114 9482
rect 6913 9424 6918 9480
rect 6974 9424 7114 9480
rect 6913 9422 7114 9424
rect 6913 9419 6979 9422
rect 5660 9280 5980 9281
rect 5660 9216 5668 9280
rect 5732 9216 5748 9280
rect 5812 9216 5828 9280
rect 5892 9216 5908 9280
rect 5972 9216 5980 9280
rect 5660 9215 5980 9216
rect 2865 9072 3066 9074
rect 2865 9016 2870 9072
rect 2926 9016 3066 9072
rect 2865 9014 3066 9016
rect 2865 9011 2931 9014
rect 7054 8938 7114 9422
rect 10869 9480 34000 9482
rect 10869 9424 10874 9480
rect 10930 9424 34000 9480
rect 10869 9422 34000 9424
rect 10869 9419 10935 9422
rect 14000 9392 34000 9422
rect 8760 9280 9080 9281
rect 8760 9216 8768 9280
rect 8832 9216 8848 9280
rect 8912 9216 8928 9280
rect 8992 9216 9008 9280
rect 9072 9216 9080 9280
rect 8760 9215 9080 9216
rect 7925 9074 7991 9077
rect 14000 9074 34000 9104
rect 7925 9072 34000 9074
rect 7925 9016 7930 9072
rect 7986 9016 34000 9072
rect 7925 9014 34000 9016
rect 7925 9011 7991 9014
rect 14000 8984 34000 9014
rect 7054 8878 12450 8938
rect 4110 8736 4430 8737
rect 4110 8672 4118 8736
rect 4182 8672 4198 8736
rect 4262 8672 4278 8736
rect 4342 8672 4358 8736
rect 4422 8672 4430 8736
rect 4110 8671 4430 8672
rect 7210 8736 7530 8737
rect 7210 8672 7218 8736
rect 7282 8672 7298 8736
rect 7362 8672 7378 8736
rect 7442 8672 7458 8736
rect 7522 8672 7530 8736
rect 7210 8671 7530 8672
rect 12390 8666 12450 8878
rect 14000 8666 34000 8696
rect 12390 8606 34000 8666
rect 14000 8576 34000 8606
rect 4337 8530 4403 8533
rect 4889 8530 4955 8533
rect 4337 8528 4955 8530
rect 4337 8472 4342 8528
rect 4398 8472 4894 8528
rect 4950 8472 4955 8528
rect 4337 8470 4955 8472
rect 4337 8467 4403 8470
rect 4889 8467 4955 8470
rect 6177 8530 6243 8533
rect 7189 8530 7255 8533
rect 6177 8528 7255 8530
rect 6177 8472 6182 8528
rect 6238 8472 7194 8528
rect 7250 8472 7255 8528
rect 6177 8470 7255 8472
rect 6177 8467 6243 8470
rect 7189 8467 7255 8470
rect 2037 8394 2103 8397
rect 4061 8394 4127 8397
rect 2037 8392 4127 8394
rect 2037 8336 2042 8392
rect 2098 8336 4066 8392
rect 4122 8336 4127 8392
rect 2037 8334 4127 8336
rect 2037 8331 2103 8334
rect 4061 8331 4127 8334
rect 4613 8394 4679 8397
rect 6729 8394 6795 8397
rect 4613 8392 6795 8394
rect 4613 8336 4618 8392
rect 4674 8336 6734 8392
rect 6790 8336 6795 8392
rect 4613 8334 6795 8336
rect 4613 8331 4679 8334
rect 6729 8331 6795 8334
rect 9397 8258 9463 8261
rect 14000 8258 34000 8288
rect 9397 8256 34000 8258
rect 9397 8200 9402 8256
rect 9458 8200 34000 8256
rect 9397 8198 34000 8200
rect 9397 8195 9463 8198
rect 2560 8192 2880 8193
rect 2560 8128 2568 8192
rect 2632 8128 2648 8192
rect 2712 8128 2728 8192
rect 2792 8128 2808 8192
rect 2872 8128 2880 8192
rect 2560 8127 2880 8128
rect 5660 8192 5980 8193
rect 5660 8128 5668 8192
rect 5732 8128 5748 8192
rect 5812 8128 5828 8192
rect 5892 8128 5908 8192
rect 5972 8128 5980 8192
rect 5660 8127 5980 8128
rect 8760 8192 9080 8193
rect 8760 8128 8768 8192
rect 8832 8128 8848 8192
rect 8912 8128 8928 8192
rect 8992 8128 9008 8192
rect 9072 8128 9080 8192
rect 14000 8168 34000 8198
rect 8760 8127 9080 8128
rect 2681 7986 2747 7989
rect 3049 7986 3115 7989
rect 4521 7986 4587 7989
rect 2681 7984 4587 7986
rect 2681 7928 2686 7984
rect 2742 7928 3054 7984
rect 3110 7928 4526 7984
rect 4582 7928 4587 7984
rect 2681 7926 4587 7928
rect 2681 7923 2747 7926
rect 3049 7923 3115 7926
rect 4521 7923 4587 7926
rect 841 7850 907 7853
rect 5257 7850 5323 7853
rect 841 7848 5323 7850
rect 841 7792 846 7848
rect 902 7792 5262 7848
rect 5318 7792 5323 7848
rect 841 7790 5323 7792
rect 841 7787 907 7790
rect 5257 7787 5323 7790
rect 9857 7850 9923 7853
rect 14000 7850 34000 7880
rect 9857 7848 34000 7850
rect 9857 7792 9862 7848
rect 9918 7792 34000 7848
rect 9857 7790 34000 7792
rect 9857 7787 9923 7790
rect 14000 7760 34000 7790
rect 4110 7648 4430 7649
rect 4110 7584 4118 7648
rect 4182 7584 4198 7648
rect 4262 7584 4278 7648
rect 4342 7584 4358 7648
rect 4422 7584 4430 7648
rect 4110 7583 4430 7584
rect 7210 7648 7530 7649
rect 7210 7584 7218 7648
rect 7282 7584 7298 7648
rect 7362 7584 7378 7648
rect 7442 7584 7458 7648
rect 7522 7584 7530 7648
rect 7210 7583 7530 7584
rect 6545 7442 6611 7445
rect 1534 7440 6611 7442
rect 1534 7384 6550 7440
rect 6606 7384 6611 7440
rect 1534 7382 6611 7384
rect 1534 7173 1594 7382
rect 6545 7379 6611 7382
rect 9673 7442 9739 7445
rect 14000 7442 34000 7472
rect 9673 7440 34000 7442
rect 9673 7384 9678 7440
rect 9734 7384 34000 7440
rect 9673 7382 34000 7384
rect 9673 7379 9739 7382
rect 14000 7352 34000 7382
rect 3233 7306 3299 7309
rect 3785 7306 3851 7309
rect 3233 7304 3851 7306
rect 3233 7248 3238 7304
rect 3294 7248 3790 7304
rect 3846 7248 3851 7304
rect 3233 7246 3851 7248
rect 3233 7243 3299 7246
rect 3785 7243 3851 7246
rect 4797 7306 4863 7309
rect 6545 7306 6611 7309
rect 4797 7304 6194 7306
rect 4797 7248 4802 7304
rect 4858 7248 6194 7304
rect 4797 7246 6194 7248
rect 4797 7243 4863 7246
rect 1485 7168 1594 7173
rect 1485 7112 1490 7168
rect 1546 7112 1594 7168
rect 1485 7110 1594 7112
rect 6134 7170 6194 7246
rect 6545 7304 12450 7306
rect 6545 7248 6550 7304
rect 6606 7248 12450 7304
rect 6545 7246 12450 7248
rect 6545 7243 6611 7246
rect 8201 7170 8267 7173
rect 6134 7168 8267 7170
rect 6134 7112 8206 7168
rect 8262 7112 8267 7168
rect 6134 7110 8267 7112
rect 1485 7107 1551 7110
rect 8201 7107 8267 7110
rect 2560 7104 2880 7105
rect 2560 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2880 7104
rect 2560 7039 2880 7040
rect 5660 7104 5980 7105
rect 5660 7040 5668 7104
rect 5732 7040 5748 7104
rect 5812 7040 5828 7104
rect 5892 7040 5908 7104
rect 5972 7040 5980 7104
rect 5660 7039 5980 7040
rect 8760 7104 9080 7105
rect 8760 7040 8768 7104
rect 8832 7040 8848 7104
rect 8912 7040 8928 7104
rect 8992 7040 9008 7104
rect 9072 7040 9080 7104
rect 8760 7039 9080 7040
rect 12390 7034 12450 7246
rect 14000 7034 34000 7064
rect 12390 6974 34000 7034
rect 14000 6944 34000 6974
rect 3877 6898 3943 6901
rect 3877 6896 12450 6898
rect 3877 6840 3882 6896
rect 3938 6840 12450 6896
rect 3877 6838 12450 6840
rect 3877 6835 3943 6838
rect 2957 6762 3023 6765
rect 3877 6762 3943 6765
rect 2957 6760 3943 6762
rect 2957 6704 2962 6760
rect 3018 6704 3882 6760
rect 3938 6704 3943 6760
rect 2957 6702 3943 6704
rect 2957 6699 3023 6702
rect 3877 6699 3943 6702
rect 6085 6762 6151 6765
rect 7189 6762 7255 6765
rect 6085 6760 7255 6762
rect 6085 6704 6090 6760
rect 6146 6704 7194 6760
rect 7250 6704 7255 6760
rect 6085 6702 7255 6704
rect 6085 6699 6151 6702
rect 7189 6699 7255 6702
rect 7741 6760 7807 6765
rect 7741 6704 7746 6760
rect 7802 6704 7807 6760
rect 7741 6699 7807 6704
rect 5809 6626 5875 6629
rect 7005 6626 7071 6629
rect 5809 6624 7071 6626
rect 5809 6568 5814 6624
rect 5870 6568 7010 6624
rect 7066 6568 7071 6624
rect 5809 6566 7071 6568
rect 5809 6563 5875 6566
rect 7005 6563 7071 6566
rect 4110 6560 4430 6561
rect 4110 6496 4118 6560
rect 4182 6496 4198 6560
rect 4262 6496 4278 6560
rect 4342 6496 4358 6560
rect 4422 6496 4430 6560
rect 4110 6495 4430 6496
rect 7210 6560 7530 6561
rect 7210 6496 7218 6560
rect 7282 6496 7298 6560
rect 7362 6496 7378 6560
rect 7442 6496 7458 6560
rect 7522 6496 7530 6560
rect 7210 6495 7530 6496
rect 2221 6354 2287 6357
rect 3601 6354 3667 6357
rect 2221 6352 3667 6354
rect 2221 6296 2226 6352
rect 2282 6296 3606 6352
rect 3662 6296 3667 6352
rect 2221 6294 3667 6296
rect 2221 6291 2287 6294
rect 3601 6291 3667 6294
rect 4153 6354 4219 6357
rect 7744 6354 7804 6699
rect 12390 6626 12450 6838
rect 14000 6626 34000 6656
rect 12390 6566 34000 6626
rect 14000 6536 34000 6566
rect 4153 6352 7804 6354
rect 4153 6296 4158 6352
rect 4214 6296 7804 6352
rect 4153 6294 7804 6296
rect 4153 6291 4219 6294
rect 1945 6218 2011 6221
rect 3785 6218 3851 6221
rect 1945 6216 3851 6218
rect 1945 6160 1950 6216
rect 2006 6160 3790 6216
rect 3846 6160 3851 6216
rect 1945 6158 3851 6160
rect 1945 6155 2011 6158
rect 3785 6155 3851 6158
rect 5625 6218 5691 6221
rect 7097 6218 7163 6221
rect 9305 6218 9371 6221
rect 5625 6216 6194 6218
rect 5625 6160 5630 6216
rect 5686 6160 6194 6216
rect 5625 6158 6194 6160
rect 5625 6155 5691 6158
rect 6134 6082 6194 6158
rect 7097 6216 9371 6218
rect 7097 6160 7102 6216
rect 7158 6160 9310 6216
rect 9366 6160 9371 6216
rect 7097 6158 9371 6160
rect 7097 6155 7163 6158
rect 9305 6155 9371 6158
rect 10409 6218 10475 6221
rect 14000 6218 34000 6248
rect 10409 6216 34000 6218
rect 10409 6160 10414 6216
rect 10470 6160 34000 6216
rect 10409 6158 34000 6160
rect 10409 6155 10475 6158
rect 14000 6128 34000 6158
rect 6134 6022 7298 6082
rect 2560 6016 2880 6017
rect 2560 5952 2568 6016
rect 2632 5952 2648 6016
rect 2712 5952 2728 6016
rect 2792 5952 2808 6016
rect 2872 5952 2880 6016
rect 2560 5951 2880 5952
rect 5660 6016 5980 6017
rect 5660 5952 5668 6016
rect 5732 5952 5748 6016
rect 5812 5952 5828 6016
rect 5892 5952 5908 6016
rect 5972 5952 5980 6016
rect 5660 5951 5980 5952
rect 2773 5810 2839 5813
rect 4153 5810 4219 5813
rect 2773 5808 4219 5810
rect 2773 5752 2778 5808
rect 2834 5752 4158 5808
rect 4214 5752 4219 5808
rect 2773 5750 4219 5752
rect 7238 5810 7298 6022
rect 8760 6016 9080 6017
rect 8760 5952 8768 6016
rect 8832 5952 8848 6016
rect 8912 5952 8928 6016
rect 8992 5952 9008 6016
rect 9072 5952 9080 6016
rect 8760 5951 9080 5952
rect 8201 5810 8267 5813
rect 7238 5808 8267 5810
rect 7238 5752 8206 5808
rect 8262 5752 8267 5808
rect 7238 5750 8267 5752
rect 2773 5747 2839 5750
rect 4153 5747 4219 5750
rect 8201 5747 8267 5750
rect 9765 5810 9831 5813
rect 14000 5810 34000 5840
rect 9765 5808 34000 5810
rect 9765 5752 9770 5808
rect 9826 5752 34000 5808
rect 9765 5750 34000 5752
rect 9765 5747 9831 5750
rect 14000 5720 34000 5750
rect 2405 5674 2471 5677
rect 3325 5674 3391 5677
rect 4245 5674 4311 5677
rect 2405 5672 4311 5674
rect 2405 5616 2410 5672
rect 2466 5616 3330 5672
rect 3386 5616 4250 5672
rect 4306 5616 4311 5672
rect 2405 5614 4311 5616
rect 2405 5611 2471 5614
rect 3325 5611 3391 5614
rect 4245 5611 4311 5614
rect 1669 5538 1735 5541
rect 3141 5538 3207 5541
rect 1669 5536 3207 5538
rect 1669 5480 1674 5536
rect 1730 5480 3146 5536
rect 3202 5480 3207 5536
rect 1669 5478 3207 5480
rect 1669 5475 1735 5478
rect 3141 5475 3207 5478
rect 4110 5472 4430 5473
rect 4110 5408 4118 5472
rect 4182 5408 4198 5472
rect 4262 5408 4278 5472
rect 4342 5408 4358 5472
rect 4422 5408 4430 5472
rect 4110 5407 4430 5408
rect 7210 5472 7530 5473
rect 7210 5408 7218 5472
rect 7282 5408 7298 5472
rect 7362 5408 7378 5472
rect 7442 5408 7458 5472
rect 7522 5408 7530 5472
rect 7210 5407 7530 5408
rect 14000 5402 34000 5432
rect 12390 5342 34000 5402
rect 2681 5266 2747 5269
rect 5901 5266 5967 5269
rect 2681 5264 5967 5266
rect 2681 5208 2686 5264
rect 2742 5208 5906 5264
rect 5962 5208 5967 5264
rect 2681 5206 5967 5208
rect 2681 5203 2747 5206
rect 5901 5203 5967 5206
rect 6913 5266 6979 5269
rect 12390 5266 12450 5342
rect 14000 5312 34000 5342
rect 6913 5264 12450 5266
rect 6913 5208 6918 5264
rect 6974 5208 12450 5264
rect 6913 5206 12450 5208
rect 6913 5203 6979 5206
rect 9673 4994 9739 4997
rect 14000 4994 34000 5024
rect 9673 4992 34000 4994
rect 9673 4936 9678 4992
rect 9734 4936 34000 4992
rect 9673 4934 34000 4936
rect 9673 4931 9739 4934
rect 5660 4928 5980 4929
rect 5660 4864 5668 4928
rect 5732 4864 5748 4928
rect 5812 4864 5828 4928
rect 5892 4864 5908 4928
rect 5972 4864 5980 4928
rect 5660 4863 5980 4864
rect 8760 4928 9080 4929
rect 8760 4864 8768 4928
rect 8832 4864 8848 4928
rect 8912 4864 8928 4928
rect 8992 4864 9008 4928
rect 9072 4864 9080 4928
rect 14000 4904 34000 4934
rect 8760 4863 9080 4864
rect 3509 4722 3575 4725
rect 7189 4722 7255 4725
rect 3509 4720 7255 4722
rect 3509 4664 3514 4720
rect 3570 4664 7194 4720
rect 7250 4664 7255 4720
rect 3509 4662 7255 4664
rect 3509 4659 3575 4662
rect 7189 4659 7255 4662
rect 13813 4586 13879 4589
rect 14000 4586 34000 4616
rect 13813 4584 34000 4586
rect 13813 4528 13818 4584
rect 13874 4528 34000 4584
rect 13813 4526 34000 4528
rect 13813 4523 13879 4526
rect 14000 4496 34000 4526
rect 8569 4450 8635 4453
rect 8569 4448 9460 4450
rect 8569 4392 8574 4448
rect 8630 4392 9460 4448
rect 8569 4390 9460 4392
rect 8569 4387 8635 4390
rect 4110 4384 4430 4385
rect 4110 4320 4118 4384
rect 4182 4320 4198 4384
rect 4262 4320 4278 4384
rect 4342 4320 4358 4384
rect 4422 4320 4430 4384
rect 4110 4319 4430 4320
rect 7210 4384 7530 4385
rect 7210 4320 7218 4384
rect 7282 4320 7298 4384
rect 7362 4320 7378 4384
rect 7442 4320 7458 4384
rect 7522 4320 7530 4384
rect 7210 4319 7530 4320
rect 8201 4314 8267 4317
rect 8201 4312 9276 4314
rect 8201 4256 8206 4312
rect 8262 4256 9276 4312
rect 8201 4254 9276 4256
rect 8201 4251 8267 4254
rect 6913 4178 6979 4181
rect 2454 4176 6979 4178
rect 2454 4120 6918 4176
rect 6974 4120 6979 4176
rect 2454 4118 6979 4120
rect 2454 3332 2514 4118
rect 6913 4115 6979 4118
rect 5660 3840 5980 3841
rect 5660 3776 5668 3840
rect 5732 3776 5748 3840
rect 5812 3776 5828 3840
rect 5892 3776 5908 3840
rect 5972 3776 5980 3840
rect 5660 3775 5980 3776
rect 8760 3840 9080 3841
rect 8760 3776 8768 3840
rect 8832 3776 8848 3840
rect 8912 3776 8928 3840
rect 8992 3776 9008 3840
rect 9072 3776 9080 3840
rect 8760 3775 9080 3776
rect 9216 3773 9276 4254
rect 9213 3768 9279 3773
rect 9213 3712 9218 3768
rect 9274 3712 9279 3768
rect 9213 3707 9279 3712
rect 3969 3634 4035 3637
rect 5441 3634 5507 3637
rect 3969 3632 5507 3634
rect 3969 3576 3974 3632
rect 4030 3576 5446 3632
rect 5502 3576 5507 3632
rect 3969 3574 5507 3576
rect 3969 3571 4035 3574
rect 5441 3571 5507 3574
rect 5625 3634 5691 3637
rect 6637 3634 6703 3637
rect 5625 3632 6703 3634
rect 5625 3576 5630 3632
rect 5686 3576 6642 3632
rect 6698 3576 6703 3632
rect 5625 3574 6703 3576
rect 5625 3571 5691 3574
rect 6637 3571 6703 3574
rect 7373 3634 7439 3637
rect 9213 3634 9279 3637
rect 7373 3632 9279 3634
rect 7373 3576 7378 3632
rect 7434 3576 9218 3632
rect 9274 3576 9279 3632
rect 7373 3574 9279 3576
rect 7373 3571 7439 3574
rect 9213 3571 9279 3574
rect 7925 3498 7991 3501
rect 3926 3496 7991 3498
rect 3926 3440 7930 3496
rect 7986 3440 7991 3496
rect 3926 3438 7991 3440
rect 3926 3229 3986 3438
rect 7925 3435 7991 3438
rect 4613 3362 4679 3365
rect 5349 3362 5415 3365
rect 9400 3362 9460 4390
rect 14000 4176 34000 4208
rect 14000 4120 16578 4176
rect 16634 4120 34000 4176
rect 14000 4088 34000 4120
rect 14000 3768 34000 3800
rect 14000 3712 16578 3768
rect 16634 3712 34000 3768
rect 14000 3680 34000 3712
rect 14000 3362 34000 3392
rect 4613 3360 5415 3362
rect 4613 3304 4618 3360
rect 4674 3304 5354 3360
rect 5410 3304 5415 3360
rect 4613 3302 5415 3304
rect 4613 3299 4679 3302
rect 5349 3299 5415 3302
rect 9308 3302 9460 3362
rect 12390 3302 34000 3362
rect 4110 3296 4430 3297
rect 4110 3232 4118 3296
rect 4182 3232 4198 3296
rect 4262 3232 4278 3296
rect 4342 3232 4358 3296
rect 4422 3232 4430 3296
rect 4110 3231 4430 3232
rect 7210 3296 7530 3297
rect 7210 3232 7218 3296
rect 7282 3232 7298 3296
rect 7362 3232 7378 3296
rect 7442 3232 7458 3296
rect 7522 3232 7530 3296
rect 7210 3231 7530 3232
rect 3877 3224 3986 3229
rect 8661 3226 8727 3229
rect 3877 3168 3882 3224
rect 3938 3168 3986 3224
rect 3877 3166 3986 3168
rect 7790 3224 8727 3226
rect 7790 3168 8666 3224
rect 8722 3168 8727 3224
rect 7790 3166 8727 3168
rect 3877 3163 3943 3166
rect 2865 3090 2931 3093
rect 6821 3090 6887 3093
rect 2865 3088 6887 3090
rect 2865 3032 2870 3088
rect 2926 3032 6826 3088
rect 6882 3032 6887 3088
rect 2865 3030 6887 3032
rect 2865 3027 2931 3030
rect 6821 3027 6887 3030
rect 7189 3090 7255 3093
rect 7790 3090 7850 3166
rect 8661 3163 8727 3166
rect 7189 3088 7850 3090
rect 7189 3032 7194 3088
rect 7250 3032 7850 3088
rect 7189 3030 7850 3032
rect 8293 3090 8359 3093
rect 8569 3090 8635 3093
rect 9308 3090 9368 3302
rect 8293 3088 8635 3090
rect 8293 3032 8298 3088
rect 8354 3032 8574 3088
rect 8630 3032 8635 3088
rect 8293 3030 8635 3032
rect 7189 3027 7255 3030
rect 8293 3027 8359 3030
rect 8569 3027 8635 3030
rect 8894 3030 9368 3090
rect 8293 2954 8359 2957
rect 8894 2954 8954 3030
rect 12390 2954 12450 3302
rect 14000 3272 34000 3302
rect 8293 2952 8954 2954
rect 8293 2896 8298 2952
rect 8354 2896 8954 2952
rect 8293 2894 8954 2896
rect 9630 2894 12450 2954
rect 14000 2952 34000 2984
rect 14000 2896 16578 2952
rect 16634 2896 34000 2952
rect 8293 2891 8359 2894
rect 5660 2752 5980 2753
rect 5660 2688 5668 2752
rect 5732 2688 5748 2752
rect 5812 2688 5828 2752
rect 5892 2688 5908 2752
rect 5972 2688 5980 2752
rect 5660 2687 5980 2688
rect 8760 2752 9080 2753
rect 8760 2688 8768 2752
rect 8832 2688 8848 2752
rect 8912 2688 8928 2752
rect 8992 2688 9008 2752
rect 9072 2688 9080 2752
rect 8760 2687 9080 2688
rect 2405 2546 2471 2549
rect 7373 2546 7439 2549
rect 2405 2544 7439 2546
rect 2405 2488 2410 2544
rect 2466 2488 7378 2544
rect 7434 2488 7439 2544
rect 2405 2486 7439 2488
rect 2405 2483 2471 2486
rect 7373 2483 7439 2486
rect 8845 2546 8911 2549
rect 9630 2546 9690 2894
rect 14000 2864 34000 2896
rect 8845 2544 9690 2546
rect 8845 2488 8850 2544
rect 8906 2488 9690 2544
rect 8845 2486 9690 2488
rect 14000 2544 34000 2576
rect 14000 2488 16578 2544
rect 16634 2488 34000 2544
rect 8845 2483 8911 2486
rect 14000 2456 34000 2488
rect 7741 2410 7807 2413
rect 9765 2410 9831 2413
rect 7741 2408 9831 2410
rect 7741 2352 7746 2408
rect 7802 2352 9770 2408
rect 9826 2352 9831 2408
rect 7741 2350 9831 2352
rect 7741 2347 7807 2350
rect 9765 2347 9831 2350
rect 4110 2208 4430 2209
rect 4110 2144 4118 2208
rect 4182 2144 4198 2208
rect 4262 2144 4278 2208
rect 4342 2144 4358 2208
rect 4422 2144 4430 2208
rect 4110 2143 4430 2144
rect 7210 2208 7530 2209
rect 7210 2144 7218 2208
rect 7282 2144 7298 2208
rect 7362 2144 7378 2208
rect 7442 2144 7458 2208
rect 7522 2144 7530 2208
rect 7210 2143 7530 2144
rect 9121 2138 9187 2141
rect 14000 2138 34000 2168
rect 9121 2136 34000 2138
rect 9121 2080 9126 2136
rect 9182 2080 34000 2136
rect 9121 2078 34000 2080
rect 9121 2075 9187 2078
rect 14000 2048 34000 2078
rect 13813 1730 13879 1733
rect 14000 1730 34000 1760
rect 13813 1728 34000 1730
rect 13813 1672 13818 1728
rect 13874 1672 34000 1728
rect 13813 1670 34000 1672
rect 13813 1667 13879 1670
rect 5660 1664 5980 1665
rect 5660 1600 5668 1664
rect 5732 1600 5748 1664
rect 5812 1600 5828 1664
rect 5892 1600 5908 1664
rect 5972 1600 5980 1664
rect 5660 1599 5980 1600
rect 8760 1664 9080 1665
rect 8760 1600 8768 1664
rect 8832 1600 8848 1664
rect 8912 1600 8928 1664
rect 8992 1600 9008 1664
rect 9072 1600 9080 1664
rect 14000 1640 34000 1670
rect 8760 1599 9080 1600
rect 8937 1322 9003 1325
rect 14000 1322 34000 1352
rect 8937 1320 34000 1322
rect 8937 1264 8942 1320
rect 8998 1264 34000 1320
rect 8937 1262 34000 1264
rect 8937 1259 9003 1262
rect 14000 1232 34000 1262
rect 4110 1120 4430 1121
rect 4110 1056 4118 1120
rect 4182 1056 4198 1120
rect 4262 1056 4278 1120
rect 4342 1056 4358 1120
rect 4422 1056 4430 1120
rect 4110 1055 4430 1056
rect 7210 1120 7530 1121
rect 7210 1056 7218 1120
rect 7282 1056 7298 1120
rect 7362 1056 7378 1120
rect 7442 1056 7458 1120
rect 7522 1056 7530 1120
rect 7210 1055 7530 1056
rect 9305 914 9371 917
rect 14000 914 34000 944
rect 9305 912 34000 914
rect 9305 856 9310 912
rect 9366 856 34000 912
rect 9305 854 34000 856
rect 9305 851 9371 854
rect 14000 824 34000 854
rect 9213 506 9279 509
rect 14000 506 34000 536
rect 9213 504 34000 506
rect 9213 448 9218 504
rect 9274 448 34000 504
rect 9213 446 34000 448
rect 9213 443 9279 446
rect 14000 416 34000 446
<< via3 >>
rect 2568 11452 2632 11456
rect 2568 11396 2572 11452
rect 2572 11396 2628 11452
rect 2628 11396 2632 11452
rect 2568 11392 2632 11396
rect 2648 11452 2712 11456
rect 2648 11396 2652 11452
rect 2652 11396 2708 11452
rect 2708 11396 2712 11452
rect 2648 11392 2712 11396
rect 2728 11452 2792 11456
rect 2728 11396 2732 11452
rect 2732 11396 2788 11452
rect 2788 11396 2792 11452
rect 2728 11392 2792 11396
rect 2808 11452 2872 11456
rect 2808 11396 2812 11452
rect 2812 11396 2868 11452
rect 2868 11396 2872 11452
rect 2808 11392 2872 11396
rect 5668 11452 5732 11456
rect 5668 11396 5672 11452
rect 5672 11396 5728 11452
rect 5728 11396 5732 11452
rect 5668 11392 5732 11396
rect 5748 11452 5812 11456
rect 5748 11396 5752 11452
rect 5752 11396 5808 11452
rect 5808 11396 5812 11452
rect 5748 11392 5812 11396
rect 5828 11452 5892 11456
rect 5828 11396 5832 11452
rect 5832 11396 5888 11452
rect 5888 11396 5892 11452
rect 5828 11392 5892 11396
rect 5908 11452 5972 11456
rect 5908 11396 5912 11452
rect 5912 11396 5968 11452
rect 5968 11396 5972 11452
rect 5908 11392 5972 11396
rect 8768 11452 8832 11456
rect 8768 11396 8772 11452
rect 8772 11396 8828 11452
rect 8828 11396 8832 11452
rect 8768 11392 8832 11396
rect 8848 11452 8912 11456
rect 8848 11396 8852 11452
rect 8852 11396 8908 11452
rect 8908 11396 8912 11452
rect 8848 11392 8912 11396
rect 8928 11452 8992 11456
rect 8928 11396 8932 11452
rect 8932 11396 8988 11452
rect 8988 11396 8992 11452
rect 8928 11392 8992 11396
rect 9008 11452 9072 11456
rect 9008 11396 9012 11452
rect 9012 11396 9068 11452
rect 9068 11396 9072 11452
rect 9008 11392 9072 11396
rect 4118 10908 4182 10912
rect 4118 10852 4122 10908
rect 4122 10852 4178 10908
rect 4178 10852 4182 10908
rect 4118 10848 4182 10852
rect 4198 10908 4262 10912
rect 4198 10852 4202 10908
rect 4202 10852 4258 10908
rect 4258 10852 4262 10908
rect 4198 10848 4262 10852
rect 4278 10908 4342 10912
rect 4278 10852 4282 10908
rect 4282 10852 4338 10908
rect 4338 10852 4342 10908
rect 4278 10848 4342 10852
rect 4358 10908 4422 10912
rect 4358 10852 4362 10908
rect 4362 10852 4418 10908
rect 4418 10852 4422 10908
rect 4358 10848 4422 10852
rect 7218 10908 7282 10912
rect 7218 10852 7222 10908
rect 7222 10852 7278 10908
rect 7278 10852 7282 10908
rect 7218 10848 7282 10852
rect 7298 10908 7362 10912
rect 7298 10852 7302 10908
rect 7302 10852 7358 10908
rect 7358 10852 7362 10908
rect 7298 10848 7362 10852
rect 7378 10908 7442 10912
rect 7378 10852 7382 10908
rect 7382 10852 7438 10908
rect 7438 10852 7442 10908
rect 7378 10848 7442 10852
rect 7458 10908 7522 10912
rect 7458 10852 7462 10908
rect 7462 10852 7518 10908
rect 7518 10852 7522 10908
rect 7458 10848 7522 10852
rect 2568 10364 2632 10368
rect 2568 10308 2572 10364
rect 2572 10308 2628 10364
rect 2628 10308 2632 10364
rect 2568 10304 2632 10308
rect 2648 10364 2712 10368
rect 2648 10308 2652 10364
rect 2652 10308 2708 10364
rect 2708 10308 2712 10364
rect 2648 10304 2712 10308
rect 2728 10364 2792 10368
rect 2728 10308 2732 10364
rect 2732 10308 2788 10364
rect 2788 10308 2792 10364
rect 2728 10304 2792 10308
rect 2808 10364 2872 10368
rect 2808 10308 2812 10364
rect 2812 10308 2868 10364
rect 2868 10308 2872 10364
rect 2808 10304 2872 10308
rect 4118 9820 4182 9824
rect 4118 9764 4122 9820
rect 4122 9764 4178 9820
rect 4178 9764 4182 9820
rect 4118 9760 4182 9764
rect 4198 9820 4262 9824
rect 4198 9764 4202 9820
rect 4202 9764 4258 9820
rect 4258 9764 4262 9820
rect 4198 9760 4262 9764
rect 4278 9820 4342 9824
rect 4278 9764 4282 9820
rect 4282 9764 4338 9820
rect 4338 9764 4342 9820
rect 4278 9760 4342 9764
rect 4358 9820 4422 9824
rect 4358 9764 4362 9820
rect 4362 9764 4418 9820
rect 4418 9764 4422 9820
rect 4358 9760 4422 9764
rect 5668 10364 5732 10368
rect 5668 10308 5672 10364
rect 5672 10308 5728 10364
rect 5728 10308 5732 10364
rect 5668 10304 5732 10308
rect 5748 10364 5812 10368
rect 5748 10308 5752 10364
rect 5752 10308 5808 10364
rect 5808 10308 5812 10364
rect 5748 10304 5812 10308
rect 5828 10364 5892 10368
rect 5828 10308 5832 10364
rect 5832 10308 5888 10364
rect 5888 10308 5892 10364
rect 5828 10304 5892 10308
rect 5908 10364 5972 10368
rect 5908 10308 5912 10364
rect 5912 10308 5968 10364
rect 5968 10308 5972 10364
rect 5908 10304 5972 10308
rect 8768 10364 8832 10368
rect 8768 10308 8772 10364
rect 8772 10308 8828 10364
rect 8828 10308 8832 10364
rect 8768 10304 8832 10308
rect 8848 10364 8912 10368
rect 8848 10308 8852 10364
rect 8852 10308 8908 10364
rect 8908 10308 8912 10364
rect 8848 10304 8912 10308
rect 8928 10364 8992 10368
rect 8928 10308 8932 10364
rect 8932 10308 8988 10364
rect 8988 10308 8992 10364
rect 8928 10304 8992 10308
rect 9008 10364 9072 10368
rect 9008 10308 9012 10364
rect 9012 10308 9068 10364
rect 9068 10308 9072 10364
rect 9008 10304 9072 10308
rect 7218 9820 7282 9824
rect 7218 9764 7222 9820
rect 7222 9764 7278 9820
rect 7278 9764 7282 9820
rect 7218 9760 7282 9764
rect 7298 9820 7362 9824
rect 7298 9764 7302 9820
rect 7302 9764 7358 9820
rect 7358 9764 7362 9820
rect 7298 9760 7362 9764
rect 7378 9820 7442 9824
rect 7378 9764 7382 9820
rect 7382 9764 7438 9820
rect 7438 9764 7442 9820
rect 7378 9760 7442 9764
rect 7458 9820 7522 9824
rect 7458 9764 7462 9820
rect 7462 9764 7518 9820
rect 7518 9764 7522 9820
rect 7458 9760 7522 9764
rect 2568 9276 2632 9280
rect 2568 9220 2572 9276
rect 2572 9220 2628 9276
rect 2628 9220 2632 9276
rect 2568 9216 2632 9220
rect 2648 9276 2712 9280
rect 2648 9220 2652 9276
rect 2652 9220 2708 9276
rect 2708 9220 2712 9276
rect 2648 9216 2712 9220
rect 2728 9276 2792 9280
rect 2728 9220 2732 9276
rect 2732 9220 2788 9276
rect 2788 9220 2792 9276
rect 2728 9216 2792 9220
rect 2808 9276 2872 9280
rect 2808 9220 2812 9276
rect 2812 9220 2868 9276
rect 2868 9220 2872 9276
rect 2808 9216 2872 9220
rect 5668 9276 5732 9280
rect 5668 9220 5672 9276
rect 5672 9220 5728 9276
rect 5728 9220 5732 9276
rect 5668 9216 5732 9220
rect 5748 9276 5812 9280
rect 5748 9220 5752 9276
rect 5752 9220 5808 9276
rect 5808 9220 5812 9276
rect 5748 9216 5812 9220
rect 5828 9276 5892 9280
rect 5828 9220 5832 9276
rect 5832 9220 5888 9276
rect 5888 9220 5892 9276
rect 5828 9216 5892 9220
rect 5908 9276 5972 9280
rect 5908 9220 5912 9276
rect 5912 9220 5968 9276
rect 5968 9220 5972 9276
rect 5908 9216 5972 9220
rect 8768 9276 8832 9280
rect 8768 9220 8772 9276
rect 8772 9220 8828 9276
rect 8828 9220 8832 9276
rect 8768 9216 8832 9220
rect 8848 9276 8912 9280
rect 8848 9220 8852 9276
rect 8852 9220 8908 9276
rect 8908 9220 8912 9276
rect 8848 9216 8912 9220
rect 8928 9276 8992 9280
rect 8928 9220 8932 9276
rect 8932 9220 8988 9276
rect 8988 9220 8992 9276
rect 8928 9216 8992 9220
rect 9008 9276 9072 9280
rect 9008 9220 9012 9276
rect 9012 9220 9068 9276
rect 9068 9220 9072 9276
rect 9008 9216 9072 9220
rect 4118 8732 4182 8736
rect 4118 8676 4122 8732
rect 4122 8676 4178 8732
rect 4178 8676 4182 8732
rect 4118 8672 4182 8676
rect 4198 8732 4262 8736
rect 4198 8676 4202 8732
rect 4202 8676 4258 8732
rect 4258 8676 4262 8732
rect 4198 8672 4262 8676
rect 4278 8732 4342 8736
rect 4278 8676 4282 8732
rect 4282 8676 4338 8732
rect 4338 8676 4342 8732
rect 4278 8672 4342 8676
rect 4358 8732 4422 8736
rect 4358 8676 4362 8732
rect 4362 8676 4418 8732
rect 4418 8676 4422 8732
rect 4358 8672 4422 8676
rect 7218 8732 7282 8736
rect 7218 8676 7222 8732
rect 7222 8676 7278 8732
rect 7278 8676 7282 8732
rect 7218 8672 7282 8676
rect 7298 8732 7362 8736
rect 7298 8676 7302 8732
rect 7302 8676 7358 8732
rect 7358 8676 7362 8732
rect 7298 8672 7362 8676
rect 7378 8732 7442 8736
rect 7378 8676 7382 8732
rect 7382 8676 7438 8732
rect 7438 8676 7442 8732
rect 7378 8672 7442 8676
rect 7458 8732 7522 8736
rect 7458 8676 7462 8732
rect 7462 8676 7518 8732
rect 7518 8676 7522 8732
rect 7458 8672 7522 8676
rect 2568 8188 2632 8192
rect 2568 8132 2572 8188
rect 2572 8132 2628 8188
rect 2628 8132 2632 8188
rect 2568 8128 2632 8132
rect 2648 8188 2712 8192
rect 2648 8132 2652 8188
rect 2652 8132 2708 8188
rect 2708 8132 2712 8188
rect 2648 8128 2712 8132
rect 2728 8188 2792 8192
rect 2728 8132 2732 8188
rect 2732 8132 2788 8188
rect 2788 8132 2792 8188
rect 2728 8128 2792 8132
rect 2808 8188 2872 8192
rect 2808 8132 2812 8188
rect 2812 8132 2868 8188
rect 2868 8132 2872 8188
rect 2808 8128 2872 8132
rect 5668 8188 5732 8192
rect 5668 8132 5672 8188
rect 5672 8132 5728 8188
rect 5728 8132 5732 8188
rect 5668 8128 5732 8132
rect 5748 8188 5812 8192
rect 5748 8132 5752 8188
rect 5752 8132 5808 8188
rect 5808 8132 5812 8188
rect 5748 8128 5812 8132
rect 5828 8188 5892 8192
rect 5828 8132 5832 8188
rect 5832 8132 5888 8188
rect 5888 8132 5892 8188
rect 5828 8128 5892 8132
rect 5908 8188 5972 8192
rect 5908 8132 5912 8188
rect 5912 8132 5968 8188
rect 5968 8132 5972 8188
rect 5908 8128 5972 8132
rect 8768 8188 8832 8192
rect 8768 8132 8772 8188
rect 8772 8132 8828 8188
rect 8828 8132 8832 8188
rect 8768 8128 8832 8132
rect 8848 8188 8912 8192
rect 8848 8132 8852 8188
rect 8852 8132 8908 8188
rect 8908 8132 8912 8188
rect 8848 8128 8912 8132
rect 8928 8188 8992 8192
rect 8928 8132 8932 8188
rect 8932 8132 8988 8188
rect 8988 8132 8992 8188
rect 8928 8128 8992 8132
rect 9008 8188 9072 8192
rect 9008 8132 9012 8188
rect 9012 8132 9068 8188
rect 9068 8132 9072 8188
rect 9008 8128 9072 8132
rect 4118 7644 4182 7648
rect 4118 7588 4122 7644
rect 4122 7588 4178 7644
rect 4178 7588 4182 7644
rect 4118 7584 4182 7588
rect 4198 7644 4262 7648
rect 4198 7588 4202 7644
rect 4202 7588 4258 7644
rect 4258 7588 4262 7644
rect 4198 7584 4262 7588
rect 4278 7644 4342 7648
rect 4278 7588 4282 7644
rect 4282 7588 4338 7644
rect 4338 7588 4342 7644
rect 4278 7584 4342 7588
rect 4358 7644 4422 7648
rect 4358 7588 4362 7644
rect 4362 7588 4418 7644
rect 4418 7588 4422 7644
rect 4358 7584 4422 7588
rect 7218 7644 7282 7648
rect 7218 7588 7222 7644
rect 7222 7588 7278 7644
rect 7278 7588 7282 7644
rect 7218 7584 7282 7588
rect 7298 7644 7362 7648
rect 7298 7588 7302 7644
rect 7302 7588 7358 7644
rect 7358 7588 7362 7644
rect 7298 7584 7362 7588
rect 7378 7644 7442 7648
rect 7378 7588 7382 7644
rect 7382 7588 7438 7644
rect 7438 7588 7442 7644
rect 7378 7584 7442 7588
rect 7458 7644 7522 7648
rect 7458 7588 7462 7644
rect 7462 7588 7518 7644
rect 7518 7588 7522 7644
rect 7458 7584 7522 7588
rect 2568 7100 2632 7104
rect 2568 7044 2572 7100
rect 2572 7044 2628 7100
rect 2628 7044 2632 7100
rect 2568 7040 2632 7044
rect 2648 7100 2712 7104
rect 2648 7044 2652 7100
rect 2652 7044 2708 7100
rect 2708 7044 2712 7100
rect 2648 7040 2712 7044
rect 2728 7100 2792 7104
rect 2728 7044 2732 7100
rect 2732 7044 2788 7100
rect 2788 7044 2792 7100
rect 2728 7040 2792 7044
rect 2808 7100 2872 7104
rect 2808 7044 2812 7100
rect 2812 7044 2868 7100
rect 2868 7044 2872 7100
rect 2808 7040 2872 7044
rect 5668 7100 5732 7104
rect 5668 7044 5672 7100
rect 5672 7044 5728 7100
rect 5728 7044 5732 7100
rect 5668 7040 5732 7044
rect 5748 7100 5812 7104
rect 5748 7044 5752 7100
rect 5752 7044 5808 7100
rect 5808 7044 5812 7100
rect 5748 7040 5812 7044
rect 5828 7100 5892 7104
rect 5828 7044 5832 7100
rect 5832 7044 5888 7100
rect 5888 7044 5892 7100
rect 5828 7040 5892 7044
rect 5908 7100 5972 7104
rect 5908 7044 5912 7100
rect 5912 7044 5968 7100
rect 5968 7044 5972 7100
rect 5908 7040 5972 7044
rect 8768 7100 8832 7104
rect 8768 7044 8772 7100
rect 8772 7044 8828 7100
rect 8828 7044 8832 7100
rect 8768 7040 8832 7044
rect 8848 7100 8912 7104
rect 8848 7044 8852 7100
rect 8852 7044 8908 7100
rect 8908 7044 8912 7100
rect 8848 7040 8912 7044
rect 8928 7100 8992 7104
rect 8928 7044 8932 7100
rect 8932 7044 8988 7100
rect 8988 7044 8992 7100
rect 8928 7040 8992 7044
rect 9008 7100 9072 7104
rect 9008 7044 9012 7100
rect 9012 7044 9068 7100
rect 9068 7044 9072 7100
rect 9008 7040 9072 7044
rect 4118 6556 4182 6560
rect 4118 6500 4122 6556
rect 4122 6500 4178 6556
rect 4178 6500 4182 6556
rect 4118 6496 4182 6500
rect 4198 6556 4262 6560
rect 4198 6500 4202 6556
rect 4202 6500 4258 6556
rect 4258 6500 4262 6556
rect 4198 6496 4262 6500
rect 4278 6556 4342 6560
rect 4278 6500 4282 6556
rect 4282 6500 4338 6556
rect 4338 6500 4342 6556
rect 4278 6496 4342 6500
rect 4358 6556 4422 6560
rect 4358 6500 4362 6556
rect 4362 6500 4418 6556
rect 4418 6500 4422 6556
rect 4358 6496 4422 6500
rect 7218 6556 7282 6560
rect 7218 6500 7222 6556
rect 7222 6500 7278 6556
rect 7278 6500 7282 6556
rect 7218 6496 7282 6500
rect 7298 6556 7362 6560
rect 7298 6500 7302 6556
rect 7302 6500 7358 6556
rect 7358 6500 7362 6556
rect 7298 6496 7362 6500
rect 7378 6556 7442 6560
rect 7378 6500 7382 6556
rect 7382 6500 7438 6556
rect 7438 6500 7442 6556
rect 7378 6496 7442 6500
rect 7458 6556 7522 6560
rect 7458 6500 7462 6556
rect 7462 6500 7518 6556
rect 7518 6500 7522 6556
rect 7458 6496 7522 6500
rect 2568 6012 2632 6016
rect 2568 5956 2572 6012
rect 2572 5956 2628 6012
rect 2628 5956 2632 6012
rect 2568 5952 2632 5956
rect 2648 6012 2712 6016
rect 2648 5956 2652 6012
rect 2652 5956 2708 6012
rect 2708 5956 2712 6012
rect 2648 5952 2712 5956
rect 2728 6012 2792 6016
rect 2728 5956 2732 6012
rect 2732 5956 2788 6012
rect 2788 5956 2792 6012
rect 2728 5952 2792 5956
rect 2808 6012 2872 6016
rect 2808 5956 2812 6012
rect 2812 5956 2868 6012
rect 2868 5956 2872 6012
rect 2808 5952 2872 5956
rect 5668 6012 5732 6016
rect 5668 5956 5672 6012
rect 5672 5956 5728 6012
rect 5728 5956 5732 6012
rect 5668 5952 5732 5956
rect 5748 6012 5812 6016
rect 5748 5956 5752 6012
rect 5752 5956 5808 6012
rect 5808 5956 5812 6012
rect 5748 5952 5812 5956
rect 5828 6012 5892 6016
rect 5828 5956 5832 6012
rect 5832 5956 5888 6012
rect 5888 5956 5892 6012
rect 5828 5952 5892 5956
rect 5908 6012 5972 6016
rect 5908 5956 5912 6012
rect 5912 5956 5968 6012
rect 5968 5956 5972 6012
rect 5908 5952 5972 5956
rect 8768 6012 8832 6016
rect 8768 5956 8772 6012
rect 8772 5956 8828 6012
rect 8828 5956 8832 6012
rect 8768 5952 8832 5956
rect 8848 6012 8912 6016
rect 8848 5956 8852 6012
rect 8852 5956 8908 6012
rect 8908 5956 8912 6012
rect 8848 5952 8912 5956
rect 8928 6012 8992 6016
rect 8928 5956 8932 6012
rect 8932 5956 8988 6012
rect 8988 5956 8992 6012
rect 8928 5952 8992 5956
rect 9008 6012 9072 6016
rect 9008 5956 9012 6012
rect 9012 5956 9068 6012
rect 9068 5956 9072 6012
rect 9008 5952 9072 5956
rect 4118 5468 4182 5472
rect 4118 5412 4122 5468
rect 4122 5412 4178 5468
rect 4178 5412 4182 5468
rect 4118 5408 4182 5412
rect 4198 5468 4262 5472
rect 4198 5412 4202 5468
rect 4202 5412 4258 5468
rect 4258 5412 4262 5468
rect 4198 5408 4262 5412
rect 4278 5468 4342 5472
rect 4278 5412 4282 5468
rect 4282 5412 4338 5468
rect 4338 5412 4342 5468
rect 4278 5408 4342 5412
rect 4358 5468 4422 5472
rect 4358 5412 4362 5468
rect 4362 5412 4418 5468
rect 4418 5412 4422 5468
rect 4358 5408 4422 5412
rect 7218 5468 7282 5472
rect 7218 5412 7222 5468
rect 7222 5412 7278 5468
rect 7278 5412 7282 5468
rect 7218 5408 7282 5412
rect 7298 5468 7362 5472
rect 7298 5412 7302 5468
rect 7302 5412 7358 5468
rect 7358 5412 7362 5468
rect 7298 5408 7362 5412
rect 7378 5468 7442 5472
rect 7378 5412 7382 5468
rect 7382 5412 7438 5468
rect 7438 5412 7442 5468
rect 7378 5408 7442 5412
rect 7458 5468 7522 5472
rect 7458 5412 7462 5468
rect 7462 5412 7518 5468
rect 7518 5412 7522 5468
rect 7458 5408 7522 5412
rect 5668 4924 5732 4928
rect 5668 4868 5672 4924
rect 5672 4868 5728 4924
rect 5728 4868 5732 4924
rect 5668 4864 5732 4868
rect 5748 4924 5812 4928
rect 5748 4868 5752 4924
rect 5752 4868 5808 4924
rect 5808 4868 5812 4924
rect 5748 4864 5812 4868
rect 5828 4924 5892 4928
rect 5828 4868 5832 4924
rect 5832 4868 5888 4924
rect 5888 4868 5892 4924
rect 5828 4864 5892 4868
rect 5908 4924 5972 4928
rect 5908 4868 5912 4924
rect 5912 4868 5968 4924
rect 5968 4868 5972 4924
rect 5908 4864 5972 4868
rect 8768 4924 8832 4928
rect 8768 4868 8772 4924
rect 8772 4868 8828 4924
rect 8828 4868 8832 4924
rect 8768 4864 8832 4868
rect 8848 4924 8912 4928
rect 8848 4868 8852 4924
rect 8852 4868 8908 4924
rect 8908 4868 8912 4924
rect 8848 4864 8912 4868
rect 8928 4924 8992 4928
rect 8928 4868 8932 4924
rect 8932 4868 8988 4924
rect 8988 4868 8992 4924
rect 8928 4864 8992 4868
rect 9008 4924 9072 4928
rect 9008 4868 9012 4924
rect 9012 4868 9068 4924
rect 9068 4868 9072 4924
rect 9008 4864 9072 4868
rect 4118 4380 4182 4384
rect 4118 4324 4122 4380
rect 4122 4324 4178 4380
rect 4178 4324 4182 4380
rect 4118 4320 4182 4324
rect 4198 4380 4262 4384
rect 4198 4324 4202 4380
rect 4202 4324 4258 4380
rect 4258 4324 4262 4380
rect 4198 4320 4262 4324
rect 4278 4380 4342 4384
rect 4278 4324 4282 4380
rect 4282 4324 4338 4380
rect 4338 4324 4342 4380
rect 4278 4320 4342 4324
rect 4358 4380 4422 4384
rect 4358 4324 4362 4380
rect 4362 4324 4418 4380
rect 4418 4324 4422 4380
rect 4358 4320 4422 4324
rect 7218 4380 7282 4384
rect 7218 4324 7222 4380
rect 7222 4324 7278 4380
rect 7278 4324 7282 4380
rect 7218 4320 7282 4324
rect 7298 4380 7362 4384
rect 7298 4324 7302 4380
rect 7302 4324 7358 4380
rect 7358 4324 7362 4380
rect 7298 4320 7362 4324
rect 7378 4380 7442 4384
rect 7378 4324 7382 4380
rect 7382 4324 7438 4380
rect 7438 4324 7442 4380
rect 7378 4320 7442 4324
rect 7458 4380 7522 4384
rect 7458 4324 7462 4380
rect 7462 4324 7518 4380
rect 7518 4324 7522 4380
rect 7458 4320 7522 4324
rect 5668 3836 5732 3840
rect 5668 3780 5672 3836
rect 5672 3780 5728 3836
rect 5728 3780 5732 3836
rect 5668 3776 5732 3780
rect 5748 3836 5812 3840
rect 5748 3780 5752 3836
rect 5752 3780 5808 3836
rect 5808 3780 5812 3836
rect 5748 3776 5812 3780
rect 5828 3836 5892 3840
rect 5828 3780 5832 3836
rect 5832 3780 5888 3836
rect 5888 3780 5892 3836
rect 5828 3776 5892 3780
rect 5908 3836 5972 3840
rect 5908 3780 5912 3836
rect 5912 3780 5968 3836
rect 5968 3780 5972 3836
rect 5908 3776 5972 3780
rect 8768 3836 8832 3840
rect 8768 3780 8772 3836
rect 8772 3780 8828 3836
rect 8828 3780 8832 3836
rect 8768 3776 8832 3780
rect 8848 3836 8912 3840
rect 8848 3780 8852 3836
rect 8852 3780 8908 3836
rect 8908 3780 8912 3836
rect 8848 3776 8912 3780
rect 8928 3836 8992 3840
rect 8928 3780 8932 3836
rect 8932 3780 8988 3836
rect 8988 3780 8992 3836
rect 8928 3776 8992 3780
rect 9008 3836 9072 3840
rect 9008 3780 9012 3836
rect 9012 3780 9068 3836
rect 9068 3780 9072 3836
rect 9008 3776 9072 3780
rect 4118 3292 4182 3296
rect 4118 3236 4122 3292
rect 4122 3236 4178 3292
rect 4178 3236 4182 3292
rect 4118 3232 4182 3236
rect 4198 3292 4262 3296
rect 4198 3236 4202 3292
rect 4202 3236 4258 3292
rect 4258 3236 4262 3292
rect 4198 3232 4262 3236
rect 4278 3292 4342 3296
rect 4278 3236 4282 3292
rect 4282 3236 4338 3292
rect 4338 3236 4342 3292
rect 4278 3232 4342 3236
rect 4358 3292 4422 3296
rect 4358 3236 4362 3292
rect 4362 3236 4418 3292
rect 4418 3236 4422 3292
rect 4358 3232 4422 3236
rect 7218 3292 7282 3296
rect 7218 3236 7222 3292
rect 7222 3236 7278 3292
rect 7278 3236 7282 3292
rect 7218 3232 7282 3236
rect 7298 3292 7362 3296
rect 7298 3236 7302 3292
rect 7302 3236 7358 3292
rect 7358 3236 7362 3292
rect 7298 3232 7362 3236
rect 7378 3292 7442 3296
rect 7378 3236 7382 3292
rect 7382 3236 7438 3292
rect 7438 3236 7442 3292
rect 7378 3232 7442 3236
rect 7458 3292 7522 3296
rect 7458 3236 7462 3292
rect 7462 3236 7518 3292
rect 7518 3236 7522 3292
rect 7458 3232 7522 3236
rect 5668 2748 5732 2752
rect 5668 2692 5672 2748
rect 5672 2692 5728 2748
rect 5728 2692 5732 2748
rect 5668 2688 5732 2692
rect 5748 2748 5812 2752
rect 5748 2692 5752 2748
rect 5752 2692 5808 2748
rect 5808 2692 5812 2748
rect 5748 2688 5812 2692
rect 5828 2748 5892 2752
rect 5828 2692 5832 2748
rect 5832 2692 5888 2748
rect 5888 2692 5892 2748
rect 5828 2688 5892 2692
rect 5908 2748 5972 2752
rect 5908 2692 5912 2748
rect 5912 2692 5968 2748
rect 5968 2692 5972 2748
rect 5908 2688 5972 2692
rect 8768 2748 8832 2752
rect 8768 2692 8772 2748
rect 8772 2692 8828 2748
rect 8828 2692 8832 2748
rect 8768 2688 8832 2692
rect 8848 2748 8912 2752
rect 8848 2692 8852 2748
rect 8852 2692 8908 2748
rect 8908 2692 8912 2748
rect 8848 2688 8912 2692
rect 8928 2748 8992 2752
rect 8928 2692 8932 2748
rect 8932 2692 8988 2748
rect 8988 2692 8992 2748
rect 8928 2688 8992 2692
rect 9008 2748 9072 2752
rect 9008 2692 9012 2748
rect 9012 2692 9068 2748
rect 9068 2692 9072 2748
rect 9008 2688 9072 2692
rect 4118 2204 4182 2208
rect 4118 2148 4122 2204
rect 4122 2148 4178 2204
rect 4178 2148 4182 2204
rect 4118 2144 4182 2148
rect 4198 2204 4262 2208
rect 4198 2148 4202 2204
rect 4202 2148 4258 2204
rect 4258 2148 4262 2204
rect 4198 2144 4262 2148
rect 4278 2204 4342 2208
rect 4278 2148 4282 2204
rect 4282 2148 4338 2204
rect 4338 2148 4342 2204
rect 4278 2144 4342 2148
rect 4358 2204 4422 2208
rect 4358 2148 4362 2204
rect 4362 2148 4418 2204
rect 4418 2148 4422 2204
rect 4358 2144 4422 2148
rect 7218 2204 7282 2208
rect 7218 2148 7222 2204
rect 7222 2148 7278 2204
rect 7278 2148 7282 2204
rect 7218 2144 7282 2148
rect 7298 2204 7362 2208
rect 7298 2148 7302 2204
rect 7302 2148 7358 2204
rect 7358 2148 7362 2204
rect 7298 2144 7362 2148
rect 7378 2204 7442 2208
rect 7378 2148 7382 2204
rect 7382 2148 7438 2204
rect 7438 2148 7442 2204
rect 7378 2144 7442 2148
rect 7458 2204 7522 2208
rect 7458 2148 7462 2204
rect 7462 2148 7518 2204
rect 7518 2148 7522 2204
rect 7458 2144 7522 2148
rect 5668 1660 5732 1664
rect 5668 1604 5672 1660
rect 5672 1604 5728 1660
rect 5728 1604 5732 1660
rect 5668 1600 5732 1604
rect 5748 1660 5812 1664
rect 5748 1604 5752 1660
rect 5752 1604 5808 1660
rect 5808 1604 5812 1660
rect 5748 1600 5812 1604
rect 5828 1660 5892 1664
rect 5828 1604 5832 1660
rect 5832 1604 5888 1660
rect 5888 1604 5892 1660
rect 5828 1600 5892 1604
rect 5908 1660 5972 1664
rect 5908 1604 5912 1660
rect 5912 1604 5968 1660
rect 5968 1604 5972 1660
rect 5908 1600 5972 1604
rect 8768 1660 8832 1664
rect 8768 1604 8772 1660
rect 8772 1604 8828 1660
rect 8828 1604 8832 1660
rect 8768 1600 8832 1604
rect 8848 1660 8912 1664
rect 8848 1604 8852 1660
rect 8852 1604 8908 1660
rect 8908 1604 8912 1660
rect 8848 1600 8912 1604
rect 8928 1660 8992 1664
rect 8928 1604 8932 1660
rect 8932 1604 8988 1660
rect 8988 1604 8992 1660
rect 8928 1600 8992 1604
rect 9008 1660 9072 1664
rect 9008 1604 9012 1660
rect 9012 1604 9068 1660
rect 9068 1604 9072 1660
rect 9008 1600 9072 1604
rect 4118 1116 4182 1120
rect 4118 1060 4122 1116
rect 4122 1060 4178 1116
rect 4178 1060 4182 1116
rect 4118 1056 4182 1060
rect 4198 1116 4262 1120
rect 4198 1060 4202 1116
rect 4202 1060 4258 1116
rect 4258 1060 4262 1116
rect 4198 1056 4262 1060
rect 4278 1116 4342 1120
rect 4278 1060 4282 1116
rect 4282 1060 4338 1116
rect 4338 1060 4342 1116
rect 4278 1056 4342 1060
rect 4358 1116 4422 1120
rect 4358 1060 4362 1116
rect 4362 1060 4418 1116
rect 4418 1060 4422 1116
rect 4358 1056 4422 1060
rect 7218 1116 7282 1120
rect 7218 1060 7222 1116
rect 7222 1060 7278 1116
rect 7278 1060 7282 1116
rect 7218 1056 7282 1060
rect 7298 1116 7362 1120
rect 7298 1060 7302 1116
rect 7302 1060 7358 1116
rect 7358 1060 7362 1116
rect 7298 1056 7362 1060
rect 7378 1116 7442 1120
rect 7378 1060 7382 1116
rect 7382 1060 7438 1116
rect 7438 1060 7442 1116
rect 7378 1056 7442 1060
rect 7458 1116 7522 1120
rect 7458 1060 7462 1116
rect 7462 1060 7518 1116
rect 7518 1060 7522 1116
rect 7458 1056 7522 1060
<< metal4 >>
rect 2560 11456 2880 11472
rect 2560 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2880 11456
rect 2560 10368 2880 11392
rect 2560 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2880 10368
rect 2560 9280 2880 10304
rect 2560 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2880 9280
rect 2560 8218 2880 9216
rect 2560 8192 2602 8218
rect 2838 8192 2880 8218
rect 2560 8128 2568 8192
rect 2872 8128 2880 8192
rect 2560 7982 2602 8128
rect 2838 7982 2880 8128
rect 2560 7104 2880 7982
rect 2560 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2880 7104
rect 2560 6016 2880 7040
rect 2560 5952 2568 6016
rect 2632 5952 2648 6016
rect 2712 5952 2728 6016
rect 2792 5952 2808 6016
rect 2872 5952 2880 6016
rect 2560 4838 2880 5952
rect 2560 4602 2602 4838
rect 2838 4602 2880 4838
rect 1996 4196 2276 4238
rect 1996 3960 2018 4196
rect 2254 3960 2276 4196
rect 1996 3918 2276 3960
rect 1256 2506 1536 2548
rect 1256 2270 1278 2506
rect 1514 2270 1536 2506
rect 1256 2228 1536 2270
rect 2560 1458 2880 4602
rect 2560 1222 2602 1458
rect 2838 1222 2880 1458
rect 2560 1088 2880 1222
rect 3560 9266 3880 11424
rect 3560 9030 3602 9266
rect 3838 9030 3880 9266
rect 3560 5886 3880 9030
rect 3560 5650 3602 5886
rect 3838 5650 3880 5886
rect 3560 2506 3880 5650
rect 3560 2270 3602 2506
rect 3838 2270 3880 2506
rect 3560 1088 3880 2270
rect 4110 10912 4430 11472
rect 5660 11456 5980 11472
rect 4110 10848 4118 10912
rect 4182 10848 4198 10912
rect 4262 10848 4278 10912
rect 4342 10848 4358 10912
rect 4422 10848 4430 10912
rect 4110 9908 4430 10848
rect 4110 9824 4152 9908
rect 4388 9824 4430 9908
rect 4110 9760 4118 9824
rect 4422 9760 4430 9824
rect 4110 9672 4152 9760
rect 4388 9672 4430 9760
rect 4110 8736 4430 9672
rect 4110 8672 4118 8736
rect 4182 8672 4198 8736
rect 4262 8672 4278 8736
rect 4342 8672 4358 8736
rect 4422 8672 4430 8736
rect 4110 7648 4430 8672
rect 4110 7584 4118 7648
rect 4182 7584 4198 7648
rect 4262 7584 4278 7648
rect 4342 7584 4358 7648
rect 4422 7584 4430 7648
rect 4110 6560 4430 7584
rect 4110 6496 4118 6560
rect 4182 6528 4198 6560
rect 4262 6528 4278 6560
rect 4342 6528 4358 6560
rect 4422 6496 4430 6560
rect 4110 6292 4152 6496
rect 4388 6292 4430 6496
rect 4110 5472 4430 6292
rect 4110 5408 4118 5472
rect 4182 5408 4198 5472
rect 4262 5408 4278 5472
rect 4342 5408 4358 5472
rect 4422 5408 4430 5472
rect 4110 4384 4430 5408
rect 4110 4320 4118 4384
rect 4182 4320 4198 4384
rect 4262 4320 4278 4384
rect 4342 4320 4358 4384
rect 4422 4320 4430 4384
rect 4110 3296 4430 4320
rect 4110 3232 4118 3296
rect 4182 3232 4198 3296
rect 4262 3232 4278 3296
rect 4342 3232 4358 3296
rect 4422 3232 4430 3296
rect 4110 3148 4430 3232
rect 4110 2912 4152 3148
rect 4388 2912 4430 3148
rect 4110 2208 4430 2912
rect 4110 2144 4118 2208
rect 4182 2144 4198 2208
rect 4262 2144 4278 2208
rect 4342 2144 4358 2208
rect 4422 2144 4430 2208
rect 4110 1120 4430 2144
rect 4110 1056 4118 1120
rect 4182 1056 4198 1120
rect 4262 1056 4278 1120
rect 4342 1056 4358 1120
rect 4422 1056 4430 1120
rect 5110 10956 5430 11424
rect 5110 10720 5152 10956
rect 5388 10720 5430 10956
rect 5110 7576 5430 10720
rect 5110 7340 5152 7576
rect 5388 7340 5430 7576
rect 5110 4196 5430 7340
rect 5110 3960 5152 4196
rect 5388 3960 5430 4196
rect 5110 1088 5430 3960
rect 5660 11392 5668 11456
rect 5732 11392 5748 11456
rect 5812 11392 5828 11456
rect 5892 11392 5908 11456
rect 5972 11392 5980 11456
rect 5660 10368 5980 11392
rect 5660 10304 5668 10368
rect 5732 10304 5748 10368
rect 5812 10304 5828 10368
rect 5892 10304 5908 10368
rect 5972 10304 5980 10368
rect 5660 9280 5980 10304
rect 5660 9216 5668 9280
rect 5732 9216 5748 9280
rect 5812 9216 5828 9280
rect 5892 9216 5908 9280
rect 5972 9216 5980 9280
rect 5660 8218 5980 9216
rect 5660 8192 5702 8218
rect 5938 8192 5980 8218
rect 5660 8128 5668 8192
rect 5972 8128 5980 8192
rect 5660 7982 5702 8128
rect 5938 7982 5980 8128
rect 5660 7104 5980 7982
rect 5660 7040 5668 7104
rect 5732 7040 5748 7104
rect 5812 7040 5828 7104
rect 5892 7040 5908 7104
rect 5972 7040 5980 7104
rect 5660 6016 5980 7040
rect 5660 5952 5668 6016
rect 5732 5952 5748 6016
rect 5812 5952 5828 6016
rect 5892 5952 5908 6016
rect 5972 5952 5980 6016
rect 5660 4928 5980 5952
rect 5660 4864 5668 4928
rect 5732 4864 5748 4928
rect 5812 4864 5828 4928
rect 5892 4864 5908 4928
rect 5972 4864 5980 4928
rect 5660 4838 5980 4864
rect 5660 4602 5702 4838
rect 5938 4602 5980 4838
rect 5660 3840 5980 4602
rect 5660 3776 5668 3840
rect 5732 3776 5748 3840
rect 5812 3776 5828 3840
rect 5892 3776 5908 3840
rect 5972 3776 5980 3840
rect 5660 2752 5980 3776
rect 5660 2688 5668 2752
rect 5732 2688 5748 2752
rect 5812 2688 5828 2752
rect 5892 2688 5908 2752
rect 5972 2688 5980 2752
rect 5660 1664 5980 2688
rect 5660 1600 5668 1664
rect 5732 1600 5748 1664
rect 5812 1600 5828 1664
rect 5892 1600 5908 1664
rect 5972 1600 5980 1664
rect 5660 1458 5980 1600
rect 5660 1222 5702 1458
rect 5938 1222 5980 1458
rect 4110 1040 4430 1056
rect 5660 1040 5980 1222
rect 6660 9266 6980 11424
rect 6660 9030 6702 9266
rect 6938 9030 6980 9266
rect 6660 5886 6980 9030
rect 6660 5650 6702 5886
rect 6938 5650 6980 5886
rect 6660 2506 6980 5650
rect 6660 2270 6702 2506
rect 6938 2270 6980 2506
rect 6660 1088 6980 2270
rect 7210 10912 7530 11472
rect 8760 11456 9080 11472
rect 7210 10848 7218 10912
rect 7282 10848 7298 10912
rect 7362 10848 7378 10912
rect 7442 10848 7458 10912
rect 7522 10848 7530 10912
rect 7210 9908 7530 10848
rect 7210 9824 7252 9908
rect 7488 9824 7530 9908
rect 7210 9760 7218 9824
rect 7522 9760 7530 9824
rect 7210 9672 7252 9760
rect 7488 9672 7530 9760
rect 7210 8736 7530 9672
rect 7210 8672 7218 8736
rect 7282 8672 7298 8736
rect 7362 8672 7378 8736
rect 7442 8672 7458 8736
rect 7522 8672 7530 8736
rect 7210 7648 7530 8672
rect 7210 7584 7218 7648
rect 7282 7584 7298 7648
rect 7362 7584 7378 7648
rect 7442 7584 7458 7648
rect 7522 7584 7530 7648
rect 7210 6560 7530 7584
rect 7210 6496 7218 6560
rect 7282 6528 7298 6560
rect 7362 6528 7378 6560
rect 7442 6528 7458 6560
rect 7522 6496 7530 6560
rect 7210 6292 7252 6496
rect 7488 6292 7530 6496
rect 7210 5472 7530 6292
rect 7210 5408 7218 5472
rect 7282 5408 7298 5472
rect 7362 5408 7378 5472
rect 7442 5408 7458 5472
rect 7522 5408 7530 5472
rect 7210 4384 7530 5408
rect 7210 4320 7218 4384
rect 7282 4320 7298 4384
rect 7362 4320 7378 4384
rect 7442 4320 7458 4384
rect 7522 4320 7530 4384
rect 7210 3296 7530 4320
rect 7210 3232 7218 3296
rect 7282 3232 7298 3296
rect 7362 3232 7378 3296
rect 7442 3232 7458 3296
rect 7522 3232 7530 3296
rect 7210 3148 7530 3232
rect 7210 2912 7252 3148
rect 7488 2912 7530 3148
rect 7210 2208 7530 2912
rect 7210 2144 7218 2208
rect 7282 2144 7298 2208
rect 7362 2144 7378 2208
rect 7442 2144 7458 2208
rect 7522 2144 7530 2208
rect 7210 1120 7530 2144
rect 7210 1056 7218 1120
rect 7282 1056 7298 1120
rect 7362 1056 7378 1120
rect 7442 1056 7458 1120
rect 7522 1056 7530 1120
rect 8210 10956 8530 11424
rect 8210 10720 8252 10956
rect 8488 10720 8530 10956
rect 8210 7576 8530 10720
rect 8210 7340 8252 7576
rect 8488 7340 8530 7576
rect 8210 4196 8530 7340
rect 8210 3960 8252 4196
rect 8488 3960 8530 4196
rect 8210 1088 8530 3960
rect 8760 11392 8768 11456
rect 8832 11392 8848 11456
rect 8912 11392 8928 11456
rect 8992 11392 9008 11456
rect 9072 11392 9080 11456
rect 8760 10368 9080 11392
rect 8760 10304 8768 10368
rect 8832 10304 8848 10368
rect 8912 10304 8928 10368
rect 8992 10304 9008 10368
rect 9072 10304 9080 10368
rect 8760 9280 9080 10304
rect 8760 9216 8768 9280
rect 8832 9216 8848 9280
rect 8912 9216 8928 9280
rect 8992 9216 9008 9280
rect 9072 9216 9080 9280
rect 8760 8218 9080 9216
rect 8760 8192 8802 8218
rect 9038 8192 9080 8218
rect 8760 8128 8768 8192
rect 9072 8128 9080 8192
rect 8760 7982 8802 8128
rect 9038 7982 9080 8128
rect 8760 7104 9080 7982
rect 8760 7040 8768 7104
rect 8832 7040 8848 7104
rect 8912 7040 8928 7104
rect 8992 7040 9008 7104
rect 9072 7040 9080 7104
rect 8760 6016 9080 7040
rect 8760 5952 8768 6016
rect 8832 5952 8848 6016
rect 8912 5952 8928 6016
rect 8992 5952 9008 6016
rect 9072 5952 9080 6016
rect 8760 4928 9080 5952
rect 8760 4864 8768 4928
rect 8832 4864 8848 4928
rect 8912 4864 8928 4928
rect 8992 4864 9008 4928
rect 9072 4864 9080 4928
rect 8760 4838 9080 4864
rect 8760 4602 8802 4838
rect 9038 4602 9080 4838
rect 8760 3840 9080 4602
rect 8760 3776 8768 3840
rect 8832 3776 8848 3840
rect 8912 3776 8928 3840
rect 8992 3776 9008 3840
rect 9072 3776 9080 3840
rect 8760 2752 9080 3776
rect 8760 2688 8768 2752
rect 8832 2688 8848 2752
rect 8912 2688 8928 2752
rect 8992 2688 9008 2752
rect 9072 2688 9080 2752
rect 8760 1664 9080 2688
rect 8760 1600 8768 1664
rect 8832 1600 8848 1664
rect 8912 1600 8928 1664
rect 8992 1600 9008 1664
rect 9072 1600 9080 1664
rect 8760 1458 9080 1600
rect 8760 1222 8802 1458
rect 9038 1222 9080 1458
rect 7210 1040 7530 1056
rect 8760 1040 9080 1222
<< via4 >>
rect 2602 8192 2838 8218
rect 2602 8128 2632 8192
rect 2632 8128 2648 8192
rect 2648 8128 2712 8192
rect 2712 8128 2728 8192
rect 2728 8128 2792 8192
rect 2792 8128 2808 8192
rect 2808 8128 2838 8192
rect 2602 7982 2838 8128
rect 2602 4602 2838 4838
rect 2018 3960 2254 4196
rect 1278 2270 1514 2506
rect 2602 1222 2838 1458
rect 3602 9030 3838 9266
rect 3602 5650 3838 5886
rect 3602 2270 3838 2506
rect 4152 9824 4388 9908
rect 4152 9760 4182 9824
rect 4182 9760 4198 9824
rect 4198 9760 4262 9824
rect 4262 9760 4278 9824
rect 4278 9760 4342 9824
rect 4342 9760 4358 9824
rect 4358 9760 4388 9824
rect 4152 9672 4388 9760
rect 4152 6496 4182 6528
rect 4182 6496 4198 6528
rect 4198 6496 4262 6528
rect 4262 6496 4278 6528
rect 4278 6496 4342 6528
rect 4342 6496 4358 6528
rect 4358 6496 4388 6528
rect 4152 6292 4388 6496
rect 4152 2912 4388 3148
rect 5152 10720 5388 10956
rect 5152 7340 5388 7576
rect 5152 3960 5388 4196
rect 5702 8192 5938 8218
rect 5702 8128 5732 8192
rect 5732 8128 5748 8192
rect 5748 8128 5812 8192
rect 5812 8128 5828 8192
rect 5828 8128 5892 8192
rect 5892 8128 5908 8192
rect 5908 8128 5938 8192
rect 5702 7982 5938 8128
rect 5702 4602 5938 4838
rect 5702 1222 5938 1458
rect 6702 9030 6938 9266
rect 6702 5650 6938 5886
rect 6702 2270 6938 2506
rect 7252 9824 7488 9908
rect 7252 9760 7282 9824
rect 7282 9760 7298 9824
rect 7298 9760 7362 9824
rect 7362 9760 7378 9824
rect 7378 9760 7442 9824
rect 7442 9760 7458 9824
rect 7458 9760 7488 9824
rect 7252 9672 7488 9760
rect 7252 6496 7282 6528
rect 7282 6496 7298 6528
rect 7298 6496 7362 6528
rect 7362 6496 7378 6528
rect 7378 6496 7442 6528
rect 7442 6496 7458 6528
rect 7458 6496 7488 6528
rect 7252 6292 7488 6496
rect 7252 2912 7488 3148
rect 8252 10720 8488 10956
rect 8252 7340 8488 7576
rect 8252 3960 8488 4196
rect 8802 8192 9038 8218
rect 8802 8128 8832 8192
rect 8832 8128 8848 8192
rect 8848 8128 8912 8192
rect 8912 8128 8928 8192
rect 8928 8128 8992 8192
rect 8992 8128 9008 8192
rect 9008 8128 9038 8192
rect 8802 7982 9038 8128
rect 8802 4602 9038 4838
rect 8802 1222 9038 1458
<< metal5 >>
rect 920 10956 9844 10998
rect 920 10720 5152 10956
rect 5388 10720 8252 10956
rect 8488 10720 9844 10956
rect 920 10678 9844 10720
rect 920 9908 9844 9950
rect 920 9672 4152 9908
rect 4388 9672 7252 9908
rect 7488 9672 9844 9908
rect 920 9630 9844 9672
rect 920 9266 9844 9308
rect 920 9030 3602 9266
rect 3838 9030 6702 9266
rect 6938 9030 9844 9266
rect 920 8988 9844 9030
rect 920 8218 9844 8260
rect 920 7982 2602 8218
rect 2838 7982 5702 8218
rect 5938 7982 8802 8218
rect 9038 7982 9844 8218
rect 920 7940 9844 7982
rect 920 7576 9844 7618
rect 920 7340 5152 7576
rect 5388 7340 8252 7576
rect 8488 7340 9844 7576
rect 920 7298 9844 7340
rect 920 6528 9844 6570
rect 920 6292 4152 6528
rect 4388 6292 7252 6528
rect 7488 6292 9844 6528
rect 920 6250 9844 6292
rect 920 5886 9844 5928
rect 920 5650 3602 5886
rect 3838 5650 6702 5886
rect 6938 5650 9844 5886
rect 920 5608 9844 5650
rect 920 4838 9844 4880
rect 920 4602 2602 4838
rect 2838 4602 5702 4838
rect 5938 4602 8802 4838
rect 9038 4602 9844 4838
rect 920 4560 9844 4602
rect 920 4196 9844 4238
rect 920 3960 2018 4196
rect 2254 3960 5152 4196
rect 5388 3960 8252 4196
rect 8488 3960 9844 4196
rect 920 3918 9844 3960
rect 920 3148 9844 3190
rect 920 2912 4152 3148
rect 4388 2912 7252 3148
rect 7488 2912 9844 3148
rect 920 2870 9844 2912
rect 920 2506 9844 2548
rect 920 2270 1278 2506
rect 1514 2270 3602 2506
rect 3838 2270 6702 2506
rect 6938 2270 9844 2506
rect 920 2228 9844 2270
rect 920 1458 9844 1500
rect 920 1222 2602 1458
rect 2838 1222 5702 1458
rect 5938 1222 8802 1458
rect 9038 1222 9844 1458
rect 920 1180 9844 1222
use sky130_fd_sc_hd__clkbuf_1  output36 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 3588 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1636915332
transform -1 0 3588 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1636915332
transform -1 0 3588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1636915332
transform 1 0 3036 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1636915332
transform 1 0 3036 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1636915332
transform -1 0 3588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1636915332
transform -1 0 3588 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1636915332
transform -1 0 3588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1636915332
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1636915332
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1636915332
transform 1 0 3036 0 -1 4352
box -38 -48 314 592
use gpio_logic_high  gpio_logic_high
timestamp 1637281321
transform 1 0 1196 0 1 1680
box -38 -48 1418 2768
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1636915332
transform 1 0 3588 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 3772 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1636915332
transform -1 0 4140 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1636915332
transform -1 0 4140 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1636915332
transform -1 0 3956 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  output38
timestamp 1636915332
transform -1 0 4416 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1636915332
transform -1 0 4508 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1636915332
transform -1 0 4324 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1636915332
transform -1 0 4600 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1636915332
transform -1 0 4692 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1636915332
transform -1 0 5152 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1636915332
transform -1 0 5336 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1636915332
transform -1 0 4968 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1636915332
transform -1 0 4784 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 5612 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 5428 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1636915332
transform -1 0 5520 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_50 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 5520 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_52
timestamp 1636915332
transform 1 0 5704 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 4692 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1636915332
transform 1 0 3588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1636915332
transform -1 0 4140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1636915332
transform -1 0 4324 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1636915332
transform -1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1636915332
transform 1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_46 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 5152 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1636915332
transform -1 0 5152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _125_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_50
timestamp 1636915332
transform 1 0 5520 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1636915332
transform 1 0 5612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _124_
timestamp 1636915332
transform -1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1636915332
transform -1 0 4140 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1636915332
transform -1 0 3864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbn_1  _209_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 4324 0 -1 3264
box -38 -48 2430 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1636915332
transform -1 0 4324 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1636915332
transform -1 0 3864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1636915332
transform -1 0 4048 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _112_
timestamp 1636915332
transform -1 0 4324 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_40
timestamp 1636915332
transform 1 0 4600 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1636915332
transform -1 0 4600 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1636915332
transform -1 0 4968 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1636915332
transform -1 0 5244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1636915332
transform 1 0 5612 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output28 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 5612 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1636915332
transform -1 0 5980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbn_1  _208_
timestamp 1636915332
transform 1 0 3588 0 -1 4352
box -38 -48 2430 592
use sky130_fd_sc_hd__decap_12  FILLER_0_64
timestamp 1636915332
transform 1 0 6808 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_62
timestamp 1636915332
transform 1 0 6624 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1636915332
transform -1 0 7636 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_76
timestamp 1636915332
transform 1 0 7912 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_70
timestamp 1636915332
transform 1 0 7360 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1636915332
transform 1 0 8188 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1636915332
transform 1 0 8188 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1636915332
transform -1 0 8188 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1636915332
transform -1 0 7912 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1636915332
transform -1 0 8464 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_80
timestamp 1636915332
transform 1 0 8280 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1636915332
transform -1 0 8372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _186_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 8004 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _185_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 7268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1636915332
transform -1 0 6992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _131_
timestamp 1636915332
transform 1 0 6256 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _130_
timestamp 1636915332
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1636915332
transform -1 0 7544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_61
timestamp 1636915332
transform 1 0 6532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1636915332
transform 1 0 8280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold22 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 7544 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _134_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 7544 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1636915332
transform 1 0 8188 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_77
timestamp 1636915332
transform 1 0 8004 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_63
timestamp 1636915332
transform 1 0 6716 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__dfbbn_1  _205_
timestamp 1636915332
transform 1 0 6532 0 1 3264
box -38 -48 2430 592
use sky130_fd_sc_hd__or2b_1  _132_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 5980 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1636915332
transform -1 0 8648 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1636915332
transform 1 0 6808 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold20
timestamp 1636915332
transform 1 0 6072 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_2  gpio_in_buf OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 8188 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1636915332
transform 1 0 8188 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1636915332
transform 1 0 5980 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1636915332
transform 1 0 9200 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1636915332
transform -1 0 8924 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  const_source OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 8924 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _184_
timestamp 1636915332
transform -1 0 8924 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _182_
timestamp 1636915332
transform -1 0 8648 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 1636915332
transform 1 0 8924 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90
timestamp 1636915332
transform 1 0 9200 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1636915332
transform -1 0 8648 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _180_
timestamp 1636915332
transform 1 0 9292 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1636915332
transform -1 0 9844 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1636915332
transform -1 0 9844 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1636915332
transform 1 0 8372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _183_
timestamp 1636915332
transform 1 0 8740 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1636915332
transform 1 0 9292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1636915332
transform -1 0 9844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _194_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 8648 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1636915332
transform -1 0 9844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_93
timestamp 1636915332
transform 1 0 9476 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _179_
timestamp 1636915332
transform 1 0 8924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1636915332
transform -1 0 9844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_93
timestamp 1636915332
transform 1 0 9476 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _195_
timestamp 1636915332
transform -1 0 9476 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1636915332
transform -1 0 9844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_93
timestamp 1636915332
transform 1 0 9476 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1636915332
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_26
timestamp 1636915332
transform 1 0 3312 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _217_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 3312 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1636915332
transform 1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1636915332
transform -1 0 1472 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _190_
timestamp 1636915332
transform -1 0 1748 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _147_
timestamp 1636915332
transform -1 0 3036 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _146_
timestamp 1636915332
transform -1 0 2024 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _144_
timestamp 1636915332
transform 1 0 2024 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _128_
timestamp 1636915332
transform -1 0 3496 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _119_
timestamp 1636915332
transform 1 0 2300 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1636915332
transform 1 0 920 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _216_
timestamp 1636915332
transform 1 0 2392 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_1  _188_
timestamp 1636915332
transform -1 0 1564 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _149_
timestamp 1636915332
transform -1 0 1840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _118_
timestamp 1636915332
transform 1 0 1840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _106__5
timestamp 1636915332
transform 1 0 2116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1636915332
transform 1 0 920 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1636915332
transform 1 0 1196 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _215_
timestamp 1636915332
transform 1 0 1656 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_1  _143_
timestamp 1636915332
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1636915332
transform 1 0 920 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1636915332
transform 1 0 1196 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold15
timestamp 1636915332
transform -1 0 5612 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _114_
timestamp 1636915332
transform 1 0 3680 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _113_
timestamp 1636915332
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _110_
timestamp 1636915332
transform 1 0 5704 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _108_
timestamp 1636915332
transform 1 0 4324 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1636915332
transform 1 0 5612 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_36
timestamp 1636915332
transform 1 0 4232 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfbbn_1  _206_
timestamp 1636915332
transform 1 0 5796 0 -1 5440
box -38 -48 2430 592
use sky130_fd_sc_hd__or2_1  _116_
timestamp 1636915332
transform 1 0 5336 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_7_46
timestamp 1636915332
transform 1 0 5152 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_1  _222_
timestamp 1636915332
transform 1 0 4232 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__or2b_1  _145_
timestamp 1636915332
transform -1 0 4140 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1636915332
transform 1 0 3496 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_35
timestamp 1636915332
transform 1 0 4140 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1636915332
transform -1 0 6072 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1636915332
transform -1 0 5704 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2
timestamp 1636915332
transform 1 0 4232 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dfbbn_1  _203_
timestamp 1636915332
transform 1 0 3588 0 1 6528
box -38 -48 2430 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1636915332
transform 1 0 3496 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1636915332
transform 1 0 8096 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _223_
timestamp 1636915332
transform 1 0 6256 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_6_57
timestamp 1636915332
transform 1 0 6164 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1636915332
transform 1 0 8280 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1636915332
transform 1 0 8188 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _221_
timestamp 1636915332
transform -1 0 8648 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__or2b_1  _120_
timestamp 1636915332
transform 1 0 6164 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1636915332
transform 1 0 6072 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_63
timestamp 1636915332
transform 1 0 6716 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1636915332
transform -1 0 6900 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dfbbn_1  _207_
timestamp 1636915332
transform 1 0 6900 0 -1 6528
box -38 -48 2430 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1636915332
transform 1 0 6072 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _220_
timestamp 1636915332
transform 1 0 6532 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__or2b_1  _102_
timestamp 1636915332
transform 1 0 5980 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold19
timestamp 1636915332
transform 1 0 8832 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1636915332
transform -1 0 9844 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _197_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 8648 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1636915332
transform -1 0 9844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_serial_clock_A
timestamp 1636915332
transform -1 0 9568 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1
timestamp 1636915332
transform -1 0 9476 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1636915332
transform 1 0 8648 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1636915332
transform -1 0 9844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_93
timestamp 1636915332
transform 1 0 9476 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1636915332
transform 1 0 9292 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1636915332
transform -1 0 9844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _196_
timestamp 1636915332
transform 1 0 8740 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1636915332
transform 1 0 8372 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1636915332
transform 1 0 8648 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1636915332
transform -1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1636915332
transform 1 0 1656 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_serial_clock OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 1288 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dfbbn_1  _202_
timestamp 1636915332
transform 1 0 2576 0 -1 7616
box -38 -48 2430 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1636915332
transform 1 0 920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1636915332
transform 1 0 1196 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__5_A
timestamp 1636915332
transform 1 0 2392 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_1  _214_
timestamp 1636915332
transform -1 0 3496 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _106__4
timestamp 1636915332
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1636915332
transform 1 0 920 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__4_A
timestamp 1636915332
transform -1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold17
timestamp 1636915332
transform -1 0 2300 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _213_
timestamp 1636915332
transform 1 0 2300 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_1  _150_
timestamp 1636915332
transform 1 0 1288 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1636915332
transform 1 0 920 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1636915332
transform 1 0 1196 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _187_
timestamp 1636915332
transform -1 0 1564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _106__3
timestamp 1636915332
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1636915332
transform 1 0 920 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1636915332
transform 1 0 920 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 1636915332
transform 1 0 1196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__3_A
timestamp 1636915332
transform -1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _156_
timestamp 1636915332
transform 1 0 1564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _152_
timestamp 1636915332
transform -1 0 2116 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _138_
timestamp 1636915332
transform 1 0 2116 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1636915332
transform 1 0 1656 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _106__2
timestamp 1636915332
transform -1 0 2668 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _136_
timestamp 1636915332
transform 1 0 3220 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _137_
timestamp 1636915332
transform -1 0 2668 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _140_
timestamp 1636915332
transform -1 0 3220 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _142_
timestamp 1636915332
transform -1 0 2944 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbn_1  _204_
timestamp 1636915332
transform 1 0 2668 0 -1 9792
box -38 -48 2430 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1636915332
transform 1 0 5704 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold21
timestamp 1636915332
transform 1 0 4968 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1636915332
transform 1 0 3588 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dfbbn_1  _210_
timestamp 1636915332
transform 1 0 5152 0 1 7616
box -38 -48 2430 592
use sky130_fd_sc_hd__or2b_1  _151_
timestamp 1636915332
transform -1 0 4876 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _107_
timestamp 1636915332
transform 1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1636915332
transform 1 0 3496 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _218_
timestamp 1636915332
transform 1 0 4140 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1636915332
transform -1 0 4140 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1636915332
transform 1 0 4140 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _219_
timestamp 1636915332
transform 1 0 5336 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__or2_1  _159_
timestamp 1636915332
transform -1 0 5612 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _153_
timestamp 1636915332
transform 1 0 4876 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _104_
timestamp 1636915332
transform 1 0 5612 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1636915332
transform 1 0 3496 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_45
timestamp 1636915332
transform 1 0 5060 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__2_A
timestamp 1636915332
transform 1 0 3588 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_clock OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 8004 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__or2b_1  _126_
timestamp 1636915332
transform 1 0 8004 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1636915332
transform 1 0 6072 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold16
timestamp 1636915332
transform 1 0 7544 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_serial_clock
timestamp 1636915332
transform 1 0 8280 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1636915332
transform 1 0 6164 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dfbbn_1  _201_
timestamp 1636915332
transform -1 0 9568 0 -1 8704
box -38 -48 2430 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1636915332
transform -1 0 7176 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1636915332
transform 1 0 6072 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1636915332
transform 1 0 5980 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_12  input17 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 7176 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1636915332
transform 1 0 6164 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dfbbn_1  _200_
timestamp 1636915332
transform -1 0 9568 0 -1 9792
box -38 -48 2430 592
use sky130_fd_sc_hd__inv_2  _106__1
timestamp 1636915332
transform -1 0 7176 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1636915332
transform 1 0 6072 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _193_
timestamp 1636915332
transform 1 0 8648 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_83
timestamp 1636915332
transform 1 0 8556 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1636915332
transform -1 0 9844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_93
timestamp 1636915332
transform 1 0 9476 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold14
timestamp 1636915332
transform 1 0 8740 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1636915332
transform 1 0 8648 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1636915332
transform -1 0 9844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_93
timestamp 1636915332
transform 1 0 9476 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1636915332
transform 1 0 8740 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1636915332
transform 1 0 8648 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1636915332
transform -1 0 9844 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1636915332
transform -1 0 9844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_93
timestamp 1636915332
transform 1 0 9476 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1636915332
transform -1 0 9844 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _212_
timestamp 1636915332
transform -1 0 3496 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_1  _189_
timestamp 1636915332
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1636915332
transform 1 0 920 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1636915332
transform 1 0 1196 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold18
timestamp 1636915332
transform 1 0 2392 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _178_
timestamp 1636915332
transform -1 0 1564 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _172_
timestamp 1636915332
transform -1 0 1840 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _170_
timestamp 1636915332
transform -1 0 2116 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _167_
timestamp 1636915332
transform 1 0 2116 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _139_
timestamp 1636915332
transform -1 0 3680 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1636915332
transform 1 0 920 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1636915332
transform 1 0 1196 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1636915332
transform 1 0 1196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1636915332
transform 1 0 920 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _174_
timestamp 1636915332
transform 1 0 1564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _176_
timestamp 1636915332
transform -1 0 1564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _173_
timestamp 1636915332
transform -1 0 2116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _168_
timestamp 1636915332
transform 1 0 2116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1636915332
transform -1 0 2944 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp 1636915332
transform -1 0 2668 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _162_
timestamp 1636915332
transform 1 0 2944 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _161_
timestamp 1636915332
transform -1 0 3496 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbn_1  _199_
timestamp 1636915332
transform 1 0 3680 0 1 9792
box -38 -48 2430 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1636915332
transform 1 0 3496 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_29
timestamp 1636915332
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1636915332
transform 1 0 5244 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _177_
timestamp 1636915332
transform -1 0 6072 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _171_
timestamp 1636915332
transform 1 0 4324 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _169_
timestamp 1636915332
transform -1 0 4324 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _148_
timestamp 1636915332
transform -1 0 5060 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_30
timestamp 1636915332
transform 1 0 3680 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1636915332
transform -1 0 5244 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1636915332
transform 1 0 3496 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _141_
timestamp 1636915332
transform 1 0 3588 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_18_34
timestamp 1636915332
transform 1 0 4048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _154_
timestamp 1636915332
transform 1 0 4416 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1636915332
transform -1 0 4416 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_41
timestamp 1636915332
transform 1 0 4692 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _158_
timestamp 1636915332
transform -1 0 5060 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _155_
timestamp 1636915332
transform -1 0 5336 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1636915332
transform -1 0 5704 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1636915332
transform 1 0 5704 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _211_
timestamp 1636915332
transform -1 0 7912 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__or2b_1  _157_
timestamp 1636915332
transform -1 0 8464 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__dfbbn_1  _198_
timestamp 1636915332
transform 1 0 6164 0 -1 10880
box -38 -48 2430 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1636915332
transform 1 0 6072 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1636915332
transform -1 0 7636 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1636915332
transform -1 0 7176 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1636915332
transform 1 0 8280 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _175_
timestamp 1636915332
transform -1 0 6716 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _163_
timestamp 1636915332
transform -1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1636915332
transform 1 0 6072 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_79
timestamp 1636915332
transform 1 0 8188 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_68
timestamp 1636915332
transform 1 0 7176 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_63
timestamp 1636915332
transform 1 0 6716 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _122_
timestamp 1636915332
transform 1 0 8740 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1636915332
transform 1 0 8648 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__1_A
timestamp 1636915332
transform 1 0 8464 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _191_
timestamp 1636915332
transform 1 0 9200 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1636915332
transform -1 0 9844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _192_
timestamp 1636915332
transform -1 0 9384 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _181_
timestamp 1636915332
transform -1 0 9476 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _165_
timestamp 1636915332
transform 1 0 8556 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1636915332
transform 1 0 8740 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1636915332
transform 1 0 8648 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1636915332
transform -1 0 9844 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1636915332
transform -1 0 9844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_93
timestamp 1636915332
transform 1 0 9476 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__A
timestamp 1636915332
transform -1 0 9568 0 1 10880
box -38 -48 222 592
<< labels >>
rlabel metal2 s 938 12200 994 13000 6 gpio_defaults[0]
port 0 nsew signal input
rlabel metal2 s 5538 12200 5594 13000 6 gpio_defaults[10]
port 1 nsew signal input
rlabel metal2 s 5998 12200 6054 13000 6 gpio_defaults[11]
port 2 nsew signal input
rlabel metal2 s 6458 12200 6514 13000 6 gpio_defaults[12]
port 3 nsew signal input
rlabel metal2 s 1398 12200 1454 13000 6 gpio_defaults[1]
port 4 nsew signal input
rlabel metal2 s 1858 12200 1914 13000 6 gpio_defaults[2]
port 5 nsew signal input
rlabel metal2 s 2318 12200 2374 13000 6 gpio_defaults[3]
port 6 nsew signal input
rlabel metal2 s 2778 12200 2834 13000 6 gpio_defaults[4]
port 7 nsew signal input
rlabel metal2 s 3238 12200 3294 13000 6 gpio_defaults[5]
port 8 nsew signal input
rlabel metal2 s 3698 12200 3754 13000 6 gpio_defaults[6]
port 9 nsew signal input
rlabel metal2 s 4158 12200 4214 13000 6 gpio_defaults[7]
port 10 nsew signal input
rlabel metal2 s 4618 12200 4674 13000 6 gpio_defaults[8]
port 11 nsew signal input
rlabel metal2 s 5078 12200 5134 13000 6 gpio_defaults[9]
port 12 nsew signal input
rlabel metal3 s 14000 824 34000 944 6 mgmt_gpio_in
port 13 nsew signal tristate
rlabel metal3 s 14000 1640 34000 1760 6 mgmt_gpio_oeb
port 14 nsew signal input
rlabel metal3 s 14000 2048 34000 2168 6 mgmt_gpio_out
port 15 nsew signal input
rlabel metal3 s 14000 1232 34000 1352 6 one
port 16 nsew signal tristate
rlabel metal3 s 14000 2456 34000 2576 6 pad_gpio_ana_en
port 17 nsew signal tristate
rlabel metal3 s 14000 2864 34000 2984 6 pad_gpio_ana_pol
port 18 nsew signal tristate
rlabel metal3 s 14000 3272 34000 3392 6 pad_gpio_ana_sel
port 19 nsew signal tristate
rlabel metal3 s 14000 3680 34000 3800 6 pad_gpio_dm[0]
port 20 nsew signal tristate
rlabel metal3 s 14000 4088 34000 4208 6 pad_gpio_dm[1]
port 21 nsew signal tristate
rlabel metal3 s 14000 4496 34000 4616 6 pad_gpio_dm[2]
port 22 nsew signal tristate
rlabel metal3 s 14000 4904 34000 5024 6 pad_gpio_holdover
port 23 nsew signal tristate
rlabel metal3 s 14000 5312 34000 5432 6 pad_gpio_ib_mode_sel
port 24 nsew signal tristate
rlabel metal3 s 14000 5720 34000 5840 6 pad_gpio_in
port 25 nsew signal input
rlabel metal3 s 14000 6128 34000 6248 6 pad_gpio_inenb
port 26 nsew signal tristate
rlabel metal3 s 14000 6536 34000 6656 6 pad_gpio_out
port 27 nsew signal tristate
rlabel metal3 s 14000 6944 34000 7064 6 pad_gpio_outenb
port 28 nsew signal tristate
rlabel metal3 s 14000 7352 34000 7472 6 pad_gpio_slow_sel
port 29 nsew signal tristate
rlabel metal3 s 14000 7760 34000 7880 6 pad_gpio_vtrip_sel
port 30 nsew signal tristate
rlabel metal3 s 14000 8168 34000 8288 6 resetn
port 31 nsew signal input
rlabel metal3 s 14000 8576 34000 8696 6 resetn_out
port 32 nsew signal tristate
rlabel metal3 s 14000 8984 34000 9104 6 serial_clock
port 33 nsew signal input
rlabel metal3 s 14000 9392 34000 9512 6 serial_clock_out
port 34 nsew signal tristate
rlabel metal3 s 14000 9800 34000 9920 6 serial_data_in
port 35 nsew signal input
rlabel metal3 s 14000 10208 34000 10328 6 serial_data_out
port 36 nsew signal tristate
rlabel metal3 s 14000 10616 34000 10736 6 serial_load
port 37 nsew signal input
rlabel metal3 s 14000 11024 34000 11144 6 serial_load_out
port 38 nsew signal tristate
rlabel metal3 s 14000 11432 34000 11552 6 user_gpio_in
port 39 nsew signal tristate
rlabel metal3 s 14000 11840 34000 11960 6 user_gpio_oeb
port 40 nsew signal input
rlabel metal3 s 14000 12248 34000 12368 6 user_gpio_out
port 41 nsew signal input
rlabel metal5 s 920 1180 9844 1500 6 vccd
port 42 nsew power input
rlabel metal5 s 920 4560 9844 4880 6 vccd
port 42 nsew power input
rlabel metal5 s 920 7940 9844 8260 6 vccd
port 42 nsew power input
rlabel metal4 s 2560 1088 2880 11472 6 vccd
port 42 nsew power input
rlabel metal4 s 5660 1040 5980 11472 6 vccd
port 42 nsew power input
rlabel metal4 s 8760 1040 9080 11472 6 vccd
port 42 nsew power input
rlabel metal5 s 920 2228 9844 2548 6 vccd1
port 43 nsew power input
rlabel metal5 s 920 5608 9844 5928 6 vccd1
port 43 nsew power input
rlabel metal5 s 920 8988 9844 9308 6 vccd1
port 43 nsew power input
rlabel metal4 s 3560 1088 3880 11424 6 vccd1
port 43 nsew power input
rlabel metal4 s 6660 1088 6980 11424 6 vccd1
port 43 nsew power input
rlabel metal5 s 920 2870 9844 3190 6 vssd
port 44 nsew ground input
rlabel metal5 s 920 6250 9844 6570 6 vssd
port 44 nsew ground input
rlabel metal5 s 920 9630 9844 9950 6 vssd
port 44 nsew ground input
rlabel metal4 s 4110 1040 4430 11472 6 vssd
port 44 nsew ground input
rlabel metal4 s 7210 1040 7530 11472 6 vssd
port 44 nsew ground input
rlabel metal5 s 920 3918 9844 4238 6 vssd1
port 45 nsew ground input
rlabel metal5 s 920 7298 9844 7618 6 vssd1
port 45 nsew ground input
rlabel metal5 s 920 10678 9844 10998 6 vssd1
port 45 nsew ground input
rlabel metal4 s 5110 1088 5430 11424 6 vssd1
port 45 nsew ground input
rlabel metal4 s 8210 1088 8530 11424 6 vssd1
port 45 nsew ground input
rlabel metal3 s 14000 416 34000 536 6 zero
port 46 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 34000 13000
<< end >>
