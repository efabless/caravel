magic
tech sky130A
magscale 1 2
timestamp 1665478365
<< metal1 >>
rect 366174 1027828 366180 1027880
rect 366232 1027868 366238 1027880
rect 366542 1027868 366548 1027880
rect 366232 1027840 366548 1027868
rect 366232 1027828 366238 1027840
rect 366542 1027828 366548 1027840
rect 366600 1027828 366606 1027880
rect 366174 1024360 366180 1024412
rect 366232 1024400 366238 1024412
rect 366542 1024400 366548 1024412
rect 366232 1024372 366548 1024400
rect 366232 1024360 366238 1024372
rect 366542 1024360 366548 1024372
rect 366600 1024360 366606 1024412
rect 504542 1007020 504548 1007072
rect 504600 1007060 504606 1007072
rect 514202 1007060 514208 1007072
rect 504600 1007032 514208 1007060
rect 504600 1007020 504606 1007032
rect 514202 1007020 514208 1007032
rect 514260 1007020 514266 1007072
rect 554130 1006952 554136 1007004
rect 554188 1006992 554194 1007004
rect 559650 1006992 559656 1007004
rect 554188 1006964 559656 1006992
rect 554188 1006952 554194 1006964
rect 559650 1006952 559656 1006964
rect 559708 1006952 559714 1007004
rect 506198 1006884 506204 1006936
rect 506256 1006924 506262 1006936
rect 514018 1006924 514024 1006936
rect 506256 1006896 514024 1006924
rect 506256 1006884 506262 1006896
rect 514018 1006884 514024 1006896
rect 514076 1006884 514082 1006936
rect 145742 1006816 145748 1006868
rect 145800 1006856 145806 1006868
rect 151722 1006856 151728 1006868
rect 145800 1006828 151728 1006856
rect 145800 1006816 145806 1006828
rect 151722 1006816 151728 1006828
rect 151780 1006816 151786 1006868
rect 427998 1006816 428004 1006868
rect 428056 1006856 428062 1006868
rect 439498 1006856 439504 1006868
rect 428056 1006828 439504 1006856
rect 428056 1006816 428062 1006828
rect 439498 1006816 439504 1006828
rect 439556 1006816 439562 1006868
rect 555142 1006816 555148 1006868
rect 555200 1006856 555206 1006868
rect 562318 1006856 562324 1006868
rect 555200 1006828 562324 1006856
rect 555200 1006816 555206 1006828
rect 562318 1006816 562324 1006828
rect 562376 1006816 562382 1006868
rect 300118 1006680 300124 1006732
rect 300176 1006720 300182 1006732
rect 307754 1006720 307760 1006732
rect 300176 1006692 307760 1006720
rect 300176 1006680 300182 1006692
rect 307754 1006680 307760 1006692
rect 307812 1006680 307818 1006732
rect 357710 1006680 357716 1006732
rect 357768 1006720 357774 1006732
rect 373994 1006720 374000 1006732
rect 357768 1006692 374000 1006720
rect 357768 1006680 357774 1006692
rect 373994 1006680 374000 1006692
rect 374052 1006680 374058 1006732
rect 400858 1006680 400864 1006732
rect 400916 1006720 400922 1006732
rect 430850 1006720 430856 1006732
rect 400916 1006692 430856 1006720
rect 400916 1006680 400922 1006692
rect 430850 1006680 430856 1006692
rect 430908 1006680 430914 1006732
rect 557166 1006680 557172 1006732
rect 557224 1006720 557230 1006732
rect 566642 1006720 566648 1006732
rect 557224 1006692 566648 1006720
rect 557224 1006680 557230 1006692
rect 566642 1006680 566648 1006692
rect 566700 1006680 566706 1006732
rect 144546 1006544 144552 1006596
rect 144604 1006584 144610 1006596
rect 151446 1006584 151452 1006596
rect 144604 1006556 151452 1006584
rect 144604 1006544 144610 1006556
rect 151446 1006544 151452 1006556
rect 151504 1006544 151510 1006596
rect 298738 1006544 298744 1006596
rect 298796 1006584 298802 1006596
rect 306098 1006584 306104 1006596
rect 298796 1006556 306104 1006584
rect 298796 1006544 298802 1006556
rect 306098 1006544 306104 1006556
rect 306156 1006544 306162 1006596
rect 427170 1006544 427176 1006596
rect 427228 1006584 427234 1006596
rect 445018 1006584 445024 1006596
rect 427228 1006556 445024 1006584
rect 427228 1006544 427234 1006556
rect 445018 1006544 445024 1006556
rect 445076 1006544 445082 1006596
rect 94682 1006408 94688 1006460
rect 94740 1006448 94746 1006460
rect 101122 1006448 101128 1006460
rect 94740 1006420 101128 1006448
rect 94740 1006408 94746 1006420
rect 101122 1006408 101128 1006420
rect 101180 1006408 101186 1006460
rect 148318 1006408 148324 1006460
rect 148376 1006448 148382 1006460
rect 148376 1006420 151814 1006448
rect 148376 1006408 148382 1006420
rect 151786 1006380 151814 1006420
rect 249058 1006408 249064 1006460
rect 249116 1006448 249122 1006460
rect 255314 1006448 255320 1006460
rect 249116 1006420 255320 1006448
rect 249116 1006408 249122 1006420
rect 255314 1006408 255320 1006420
rect 255372 1006408 255378 1006460
rect 304074 1006408 304080 1006460
rect 304132 1006448 304138 1006460
rect 304132 1006420 311204 1006448
rect 304132 1006408 304138 1006420
rect 152090 1006380 152096 1006392
rect 151786 1006352 152096 1006380
rect 152090 1006340 152096 1006352
rect 152148 1006340 152154 1006392
rect 210418 1006340 210424 1006392
rect 210476 1006380 210482 1006392
rect 228358 1006380 228364 1006392
rect 210476 1006352 228364 1006380
rect 210476 1006340 210482 1006352
rect 228358 1006340 228364 1006352
rect 228416 1006340 228422 1006392
rect 94498 1006272 94504 1006324
rect 94556 1006312 94562 1006324
rect 100294 1006312 100300 1006324
rect 94556 1006284 100300 1006312
rect 94556 1006272 94562 1006284
rect 100294 1006272 100300 1006284
rect 100352 1006272 100358 1006324
rect 144178 1006272 144184 1006324
rect 144236 1006312 144242 1006324
rect 150894 1006312 150900 1006324
rect 144236 1006284 150900 1006312
rect 144236 1006272 144242 1006284
rect 150894 1006272 150900 1006284
rect 150952 1006272 150958 1006324
rect 158254 1006272 158260 1006324
rect 158312 1006312 158318 1006324
rect 158312 1006284 171134 1006312
rect 158312 1006272 158318 1006284
rect 93118 1006136 93124 1006188
rect 93176 1006176 93182 1006188
rect 99466 1006176 99472 1006188
rect 93176 1006148 99472 1006176
rect 93176 1006136 93182 1006148
rect 99466 1006136 99472 1006148
rect 99524 1006136 99530 1006188
rect 102778 1006136 102784 1006188
rect 102836 1006176 102842 1006188
rect 103974 1006176 103980 1006188
rect 102836 1006148 103980 1006176
rect 102836 1006136 102842 1006148
rect 103974 1006136 103980 1006148
rect 104032 1006136 104038 1006188
rect 106826 1006136 106832 1006188
rect 106884 1006176 106890 1006188
rect 124858 1006176 124864 1006188
rect 106884 1006148 124864 1006176
rect 106884 1006136 106890 1006148
rect 124858 1006136 124864 1006148
rect 124916 1006136 124922 1006188
rect 145558 1006136 145564 1006188
rect 145616 1006176 145622 1006188
rect 151262 1006176 151268 1006188
rect 145616 1006148 151268 1006176
rect 145616 1006136 145622 1006148
rect 151262 1006136 151268 1006148
rect 151320 1006136 151326 1006188
rect 151446 1006136 151452 1006188
rect 151504 1006176 151510 1006188
rect 159450 1006176 159456 1006188
rect 151504 1006148 159456 1006176
rect 151504 1006136 151510 1006148
rect 159450 1006136 159456 1006148
rect 159508 1006136 159514 1006188
rect 160278 1006136 160284 1006188
rect 160336 1006176 160342 1006188
rect 164878 1006176 164884 1006188
rect 160336 1006148 164884 1006176
rect 160336 1006136 160342 1006148
rect 164878 1006136 164884 1006148
rect 164936 1006136 164942 1006188
rect 171106 1006176 171134 1006284
rect 250254 1006272 250260 1006324
rect 250312 1006312 250318 1006324
rect 254118 1006312 254124 1006324
rect 250312 1006284 254124 1006312
rect 250312 1006272 250318 1006284
rect 254118 1006272 254124 1006284
rect 254176 1006272 254182 1006324
rect 298922 1006272 298928 1006324
rect 298980 1006312 298986 1006324
rect 305270 1006312 305276 1006324
rect 298980 1006284 305276 1006312
rect 298980 1006272 298986 1006284
rect 305270 1006272 305276 1006284
rect 305328 1006272 305334 1006324
rect 306926 1006312 306932 1006324
rect 305932 1006284 306932 1006312
rect 208394 1006204 208400 1006256
rect 208452 1006244 208458 1006256
rect 208452 1006216 214604 1006244
rect 208452 1006204 208458 1006216
rect 175918 1006176 175924 1006188
rect 171106 1006148 175924 1006176
rect 175918 1006136 175924 1006148
rect 175976 1006136 175982 1006188
rect 214576 1006108 214604 1006216
rect 247862 1006136 247868 1006188
rect 247920 1006176 247926 1006188
rect 253658 1006176 253664 1006188
rect 247920 1006148 253664 1006176
rect 247920 1006136 247926 1006148
rect 253658 1006136 253664 1006148
rect 253716 1006136 253722 1006188
rect 262674 1006136 262680 1006188
rect 262732 1006176 262738 1006188
rect 278038 1006176 278044 1006188
rect 262732 1006148 278044 1006176
rect 262732 1006136 262738 1006148
rect 278038 1006136 278044 1006148
rect 278096 1006136 278102 1006188
rect 300302 1006136 300308 1006188
rect 300360 1006176 300366 1006188
rect 305932 1006176 305960 1006284
rect 306926 1006272 306932 1006284
rect 306984 1006272 306990 1006324
rect 311176 1006312 311204 1006420
rect 314654 1006408 314660 1006460
rect 314712 1006448 314718 1006460
rect 319438 1006448 319444 1006460
rect 314712 1006420 319444 1006448
rect 314712 1006408 314718 1006420
rect 319438 1006408 319444 1006420
rect 319496 1006408 319502 1006460
rect 361390 1006408 361396 1006460
rect 361448 1006448 361454 1006460
rect 371878 1006448 371884 1006460
rect 361448 1006420 371884 1006448
rect 361448 1006408 361454 1006420
rect 371878 1006408 371884 1006420
rect 371936 1006408 371942 1006460
rect 423490 1006408 423496 1006460
rect 423548 1006448 423554 1006460
rect 447134 1006448 447140 1006460
rect 423548 1006420 447140 1006448
rect 423548 1006408 423554 1006420
rect 447134 1006408 447140 1006420
rect 447192 1006408 447198 1006460
rect 501690 1006408 501696 1006460
rect 501748 1006448 501754 1006460
rect 518158 1006448 518164 1006460
rect 501748 1006420 518164 1006448
rect 501748 1006408 501754 1006420
rect 518158 1006408 518164 1006420
rect 518216 1006408 518222 1006460
rect 520918 1006448 520924 1006460
rect 518866 1006420 520924 1006448
rect 331858 1006312 331864 1006324
rect 311176 1006284 331864 1006312
rect 331858 1006272 331864 1006284
rect 331916 1006272 331922 1006324
rect 424318 1006272 424324 1006324
rect 424376 1006312 424382 1006324
rect 438854 1006312 438860 1006324
rect 424376 1006284 438860 1006312
rect 424376 1006272 424382 1006284
rect 438854 1006272 438860 1006284
rect 438912 1006272 438918 1006324
rect 502150 1006272 502156 1006324
rect 502208 1006312 502214 1006324
rect 518866 1006312 518894 1006420
rect 520918 1006408 520924 1006420
rect 520976 1006408 520982 1006460
rect 552290 1006408 552296 1006460
rect 552348 1006448 552354 1006460
rect 554774 1006448 554780 1006460
rect 552348 1006420 554780 1006448
rect 552348 1006408 552354 1006420
rect 554774 1006408 554780 1006420
rect 554832 1006408 554838 1006460
rect 556798 1006408 556804 1006460
rect 556856 1006448 556862 1006460
rect 569218 1006448 569224 1006460
rect 556856 1006420 569224 1006448
rect 556856 1006408 556862 1006420
rect 569218 1006408 569224 1006420
rect 569276 1006408 569282 1006460
rect 502208 1006284 518894 1006312
rect 502208 1006272 502214 1006284
rect 554314 1006272 554320 1006324
rect 554372 1006312 554378 1006324
rect 554372 1006284 557534 1006312
rect 554372 1006272 554378 1006284
rect 300360 1006148 305960 1006176
rect 300360 1006136 300366 1006148
rect 306098 1006136 306104 1006188
rect 306156 1006176 306162 1006188
rect 311802 1006176 311808 1006188
rect 306156 1006148 311808 1006176
rect 306156 1006136 306162 1006148
rect 311802 1006136 311808 1006148
rect 311860 1006136 311866 1006188
rect 314654 1006136 314660 1006188
rect 314712 1006176 314718 1006188
rect 324958 1006176 324964 1006188
rect 314712 1006148 324964 1006176
rect 314712 1006136 314718 1006148
rect 324958 1006136 324964 1006148
rect 325016 1006136 325022 1006188
rect 365070 1006136 365076 1006188
rect 365128 1006176 365134 1006188
rect 367738 1006176 367744 1006188
rect 365128 1006148 367744 1006176
rect 365128 1006136 365134 1006148
rect 367738 1006136 367744 1006148
rect 367796 1006136 367802 1006188
rect 500494 1006136 500500 1006188
rect 500552 1006176 500558 1006188
rect 505738 1006176 505744 1006188
rect 500552 1006148 505744 1006176
rect 500552 1006136 500558 1006148
rect 505738 1006136 505744 1006148
rect 505796 1006136 505802 1006188
rect 516778 1006176 516784 1006188
rect 509206 1006148 516784 1006176
rect 214576 1006080 219434 1006108
rect 93302 1006000 93308 1006052
rect 93360 1006040 93366 1006052
rect 98270 1006040 98276 1006052
rect 93360 1006012 98276 1006040
rect 93360 1006000 93366 1006012
rect 98270 1006000 98276 1006012
rect 98328 1006000 98334 1006052
rect 101398 1006000 101404 1006052
rect 101456 1006040 101462 1006052
rect 104802 1006040 104808 1006052
rect 101456 1006012 104808 1006040
rect 101456 1006000 101462 1006012
rect 104802 1006000 104808 1006012
rect 104860 1006000 104866 1006052
rect 107654 1006000 107660 1006052
rect 107712 1006040 107718 1006052
rect 126238 1006040 126244 1006052
rect 107712 1006012 126244 1006040
rect 107712 1006000 107718 1006012
rect 126238 1006000 126244 1006012
rect 126296 1006000 126302 1006052
rect 148870 1006000 148876 1006052
rect 148928 1006040 148934 1006052
rect 150066 1006040 150072 1006052
rect 148928 1006012 150072 1006040
rect 148928 1006000 148934 1006012
rect 150066 1006000 150072 1006012
rect 150124 1006000 150130 1006052
rect 158622 1006000 158628 1006052
rect 158680 1006040 158686 1006052
rect 177298 1006040 177304 1006052
rect 158680 1006012 177304 1006040
rect 158680 1006000 158686 1006012
rect 177298 1006000 177304 1006012
rect 177356 1006000 177362 1006052
rect 197998 1006000 198004 1006052
rect 198056 1006040 198062 1006052
rect 201034 1006040 201040 1006052
rect 198056 1006012 201040 1006040
rect 198056 1006000 198062 1006012
rect 201034 1006000 201040 1006012
rect 201092 1006000 201098 1006052
rect 219406 1006040 219434 1006080
rect 229738 1006040 229744 1006052
rect 219406 1006012 229744 1006040
rect 229738 1006000 229744 1006012
rect 229796 1006000 229802 1006052
rect 247678 1006000 247684 1006052
rect 247736 1006040 247742 1006052
rect 250254 1006040 250260 1006052
rect 247736 1006012 250260 1006040
rect 247736 1006000 247742 1006012
rect 250254 1006000 250260 1006012
rect 250312 1006000 250318 1006052
rect 250438 1006000 250444 1006052
rect 250496 1006040 250502 1006052
rect 252462 1006040 252468 1006052
rect 250496 1006012 252468 1006040
rect 250496 1006000 250502 1006012
rect 252462 1006000 252468 1006012
rect 252520 1006000 252526 1006052
rect 261846 1006000 261852 1006052
rect 261904 1006040 261910 1006052
rect 280798 1006040 280804 1006052
rect 261904 1006012 280804 1006040
rect 261904 1006000 261910 1006012
rect 280798 1006000 280804 1006012
rect 280856 1006000 280862 1006052
rect 303246 1006000 303252 1006052
rect 303304 1006040 303310 1006052
rect 304074 1006040 304080 1006052
rect 303304 1006012 304080 1006040
rect 303304 1006000 303310 1006012
rect 304074 1006000 304080 1006012
rect 304132 1006000 304138 1006052
rect 305270 1006000 305276 1006052
rect 305328 1006040 305334 1006052
rect 332042 1006040 332048 1006052
rect 305328 1006012 332048 1006040
rect 305328 1006000 305334 1006012
rect 332042 1006000 332048 1006012
rect 332100 1006000 332106 1006052
rect 354858 1006000 354864 1006052
rect 354916 1006040 354922 1006052
rect 356698 1006040 356704 1006052
rect 354916 1006012 356704 1006040
rect 354916 1006000 354922 1006012
rect 356698 1006000 356704 1006012
rect 356756 1006000 356762 1006052
rect 357342 1006000 357348 1006052
rect 357400 1006040 357406 1006052
rect 376018 1006040 376024 1006052
rect 357400 1006012 376024 1006040
rect 357400 1006000 357406 1006012
rect 376018 1006000 376024 1006012
rect 376076 1006000 376082 1006052
rect 423490 1006000 423496 1006052
rect 423548 1006040 423554 1006052
rect 427814 1006040 427820 1006052
rect 423548 1006012 427820 1006040
rect 423548 1006000 423554 1006012
rect 427814 1006000 427820 1006012
rect 427872 1006000 427878 1006052
rect 429194 1006000 429200 1006052
rect 429252 1006040 429258 1006052
rect 471238 1006040 471244 1006052
rect 429252 1006012 471244 1006040
rect 429252 1006000 429258 1006012
rect 471238 1006000 471244 1006012
rect 471296 1006000 471302 1006052
rect 499666 1006000 499672 1006052
rect 499724 1006040 499730 1006052
rect 502978 1006040 502984 1006052
rect 499724 1006012 502984 1006040
rect 499724 1006000 499730 1006012
rect 502978 1006000 502984 1006012
rect 503036 1006000 503042 1006052
rect 505370 1006000 505376 1006052
rect 505428 1006040 505434 1006052
rect 509206 1006040 509234 1006148
rect 516778 1006136 516784 1006148
rect 516836 1006136 516842 1006188
rect 551462 1006136 551468 1006188
rect 551520 1006176 551526 1006188
rect 555418 1006176 555424 1006188
rect 551520 1006148 555424 1006176
rect 551520 1006136 551526 1006148
rect 555418 1006136 555424 1006148
rect 555476 1006136 555482 1006188
rect 505428 1006012 509234 1006040
rect 505428 1006000 505434 1006012
rect 514018 1006000 514024 1006052
rect 514076 1006040 514082 1006052
rect 522298 1006040 522304 1006052
rect 514076 1006012 522304 1006040
rect 514076 1006000 514082 1006012
rect 522298 1006000 522304 1006012
rect 522356 1006000 522362 1006052
rect 553118 1006000 553124 1006052
rect 553176 1006040 553182 1006052
rect 556798 1006040 556804 1006052
rect 553176 1006012 556804 1006040
rect 553176 1006000 553182 1006012
rect 556798 1006000 556804 1006012
rect 556856 1006000 556862 1006052
rect 557506 1006040 557534 1006284
rect 562318 1006272 562324 1006324
rect 562376 1006312 562382 1006324
rect 571978 1006312 571984 1006324
rect 562376 1006284 571984 1006312
rect 562376 1006272 562382 1006284
rect 571978 1006272 571984 1006284
rect 572036 1006272 572042 1006324
rect 560846 1006136 560852 1006188
rect 560904 1006176 560910 1006188
rect 563974 1006176 563980 1006188
rect 560904 1006148 563980 1006176
rect 560904 1006136 560910 1006148
rect 563974 1006136 563980 1006148
rect 564032 1006136 564038 1006188
rect 574738 1006040 574744 1006052
rect 557506 1006012 574744 1006040
rect 574738 1006000 574744 1006012
rect 574796 1006000 574802 1006052
rect 428366 1005796 428372 1005848
rect 428424 1005836 428430 1005848
rect 440878 1005836 440884 1005848
rect 428424 1005808 440884 1005836
rect 428424 1005796 428430 1005808
rect 440878 1005796 440884 1005808
rect 440936 1005796 440942 1005848
rect 509050 1005796 509056 1005848
rect 509108 1005836 509114 1005848
rect 514018 1005836 514024 1005848
rect 509108 1005808 514024 1005836
rect 509108 1005796 509114 1005808
rect 514018 1005796 514024 1005808
rect 514076 1005796 514082 1005848
rect 567838 1005836 567844 1005848
rect 563256 1005808 567844 1005836
rect 360562 1005660 360568 1005712
rect 360620 1005700 360626 1005712
rect 377398 1005700 377404 1005712
rect 360620 1005672 377404 1005700
rect 360620 1005660 360626 1005672
rect 377398 1005660 377404 1005672
rect 377456 1005660 377462 1005712
rect 427538 1005660 427544 1005712
rect 427596 1005700 427602 1005712
rect 427596 1005672 436784 1005700
rect 427596 1005660 427602 1005672
rect 359734 1005524 359740 1005576
rect 359792 1005564 359798 1005576
rect 373258 1005564 373264 1005576
rect 359792 1005536 373264 1005564
rect 359792 1005524 359798 1005536
rect 373258 1005524 373264 1005536
rect 373316 1005524 373322 1005576
rect 430850 1005524 430856 1005576
rect 430908 1005564 430914 1005576
rect 433978 1005564 433984 1005576
rect 430908 1005536 433984 1005564
rect 430908 1005524 430914 1005536
rect 433978 1005524 433984 1005536
rect 434036 1005524 434042 1005576
rect 436756 1005564 436784 1005672
rect 438854 1005660 438860 1005712
rect 438912 1005700 438918 1005712
rect 451918 1005700 451924 1005712
rect 438912 1005672 451924 1005700
rect 438912 1005660 438918 1005672
rect 451918 1005660 451924 1005672
rect 451976 1005660 451982 1005712
rect 555970 1005660 555976 1005712
rect 556028 1005700 556034 1005712
rect 563054 1005700 563060 1005712
rect 556028 1005672 563060 1005700
rect 556028 1005660 556034 1005672
rect 563054 1005660 563060 1005672
rect 563112 1005660 563118 1005712
rect 449158 1005564 449164 1005576
rect 436756 1005536 449164 1005564
rect 449158 1005524 449164 1005536
rect 449216 1005524 449222 1005576
rect 505002 1005524 505008 1005576
rect 505060 1005564 505066 1005576
rect 505060 1005536 518894 1005564
rect 505060 1005524 505066 1005536
rect 356514 1005388 356520 1005440
rect 356572 1005428 356578 1005440
rect 378778 1005428 378784 1005440
rect 356572 1005400 378784 1005428
rect 356572 1005388 356578 1005400
rect 378778 1005388 378784 1005400
rect 378836 1005388 378842 1005440
rect 431954 1005388 431960 1005440
rect 432012 1005428 432018 1005440
rect 443638 1005428 443644 1005440
rect 432012 1005400 443644 1005428
rect 432012 1005388 432018 1005400
rect 443638 1005388 443644 1005400
rect 443696 1005388 443702 1005440
rect 447134 1005388 447140 1005440
rect 447192 1005428 447198 1005440
rect 457438 1005428 457444 1005440
rect 447192 1005400 457444 1005428
rect 447192 1005388 447198 1005400
rect 457438 1005388 457444 1005400
rect 457496 1005388 457502 1005440
rect 508222 1005388 508228 1005440
rect 508280 1005428 508286 1005440
rect 510982 1005428 510988 1005440
rect 508280 1005400 510988 1005428
rect 508280 1005388 508286 1005400
rect 510982 1005388 510988 1005400
rect 511040 1005388 511046 1005440
rect 518866 1005428 518894 1005536
rect 554774 1005524 554780 1005576
rect 554832 1005564 554838 1005576
rect 563256 1005564 563284 1005808
rect 567838 1005796 567844 1005808
rect 567896 1005796 567902 1005848
rect 563974 1005660 563980 1005712
rect 564032 1005700 564038 1005712
rect 570598 1005700 570604 1005712
rect 564032 1005672 570604 1005700
rect 564032 1005660 564038 1005672
rect 570598 1005660 570604 1005672
rect 570656 1005660 570662 1005712
rect 554832 1005536 563284 1005564
rect 554832 1005524 554838 1005536
rect 522482 1005428 522488 1005440
rect 518866 1005400 522488 1005428
rect 522482 1005388 522488 1005400
rect 522540 1005388 522546 1005440
rect 555142 1005388 555148 1005440
rect 555200 1005428 555206 1005440
rect 573542 1005428 573548 1005440
rect 555200 1005400 573548 1005428
rect 555200 1005388 555206 1005400
rect 573542 1005388 573548 1005400
rect 573600 1005388 573606 1005440
rect 425514 1005320 425520 1005372
rect 425572 1005360 425578 1005372
rect 431770 1005360 431776 1005372
rect 425572 1005332 431776 1005360
rect 425572 1005320 425578 1005332
rect 431770 1005320 431776 1005332
rect 431828 1005320 431834 1005372
rect 263042 1005252 263048 1005304
rect 263100 1005292 263106 1005304
rect 279418 1005292 279424 1005304
rect 263100 1005264 279424 1005292
rect 263100 1005252 263106 1005264
rect 279418 1005252 279424 1005264
rect 279476 1005252 279482 1005304
rect 356882 1005252 356888 1005304
rect 356940 1005292 356946 1005304
rect 381538 1005292 381544 1005304
rect 356940 1005264 381544 1005292
rect 356940 1005252 356946 1005264
rect 381538 1005252 381544 1005264
rect 381596 1005252 381602 1005304
rect 431926 1005264 432276 1005292
rect 149698 1005184 149704 1005236
rect 149756 1005224 149762 1005236
rect 152918 1005224 152924 1005236
rect 149756 1005196 152924 1005224
rect 149756 1005184 149762 1005196
rect 152918 1005184 152924 1005196
rect 152976 1005184 152982 1005236
rect 304258 1005184 304264 1005236
rect 304316 1005224 304322 1005236
rect 307294 1005224 307300 1005236
rect 304316 1005196 307300 1005224
rect 304316 1005184 304322 1005196
rect 307294 1005184 307300 1005196
rect 307352 1005184 307358 1005236
rect 430022 1005184 430028 1005236
rect 430080 1005224 430086 1005236
rect 431926 1005224 431954 1005264
rect 430080 1005196 431954 1005224
rect 430080 1005184 430086 1005196
rect 432248 1005156 432276 1005264
rect 432414 1005252 432420 1005304
rect 432472 1005292 432478 1005304
rect 465718 1005292 465724 1005304
rect 432472 1005264 465724 1005292
rect 432472 1005252 432478 1005264
rect 465718 1005252 465724 1005264
rect 465776 1005252 465782 1005304
rect 500494 1005252 500500 1005304
rect 500552 1005292 500558 1005304
rect 519538 1005292 519544 1005304
rect 500552 1005264 519544 1005292
rect 500552 1005252 500558 1005264
rect 519538 1005252 519544 1005264
rect 519596 1005252 519602 1005304
rect 551094 1005252 551100 1005304
rect 551152 1005292 551158 1005304
rect 573358 1005292 573364 1005304
rect 551152 1005264 573364 1005292
rect 551152 1005252 551158 1005264
rect 573358 1005252 573364 1005264
rect 573416 1005252 573422 1005304
rect 432598 1005156 432604 1005168
rect 432248 1005128 432604 1005156
rect 432598 1005116 432604 1005128
rect 432656 1005116 432662 1005168
rect 507026 1005116 507032 1005168
rect 507084 1005156 507090 1005168
rect 509694 1005156 509700 1005168
rect 507084 1005128 509700 1005156
rect 507084 1005116 507090 1005128
rect 509694 1005116 509700 1005128
rect 509752 1005116 509758 1005168
rect 151078 1005048 151084 1005100
rect 151136 1005088 151142 1005100
rect 153746 1005088 153752 1005100
rect 151136 1005060 153752 1005088
rect 151136 1005048 151142 1005060
rect 153746 1005048 153752 1005060
rect 153804 1005048 153810 1005100
rect 363414 1005048 363420 1005100
rect 363472 1005088 363478 1005100
rect 364518 1005088 364524 1005100
rect 363472 1005060 364524 1005088
rect 363472 1005048 363478 1005060
rect 364518 1005048 364524 1005060
rect 364576 1005048 364582 1005100
rect 365070 1005048 365076 1005100
rect 365128 1005088 365134 1005100
rect 370498 1005088 370504 1005100
rect 365128 1005060 370504 1005088
rect 365128 1005048 365134 1005060
rect 370498 1005048 370504 1005060
rect 370556 1005048 370562 1005100
rect 424686 1005048 424692 1005100
rect 424744 1005088 424750 1005100
rect 431494 1005088 431500 1005100
rect 424744 1005060 431500 1005088
rect 424744 1005048 424750 1005060
rect 431494 1005048 431500 1005060
rect 431552 1005048 431558 1005100
rect 431678 1005048 431684 1005100
rect 431736 1005088 431742 1005100
rect 431736 1005060 432092 1005088
rect 431736 1005048 431742 1005060
rect 432064 1005020 432092 1005060
rect 434162 1005020 434168 1005032
rect 432064 1004992 434168 1005020
rect 434162 1004980 434168 1004992
rect 434220 1004980 434226 1005032
rect 508222 1004980 508228 1005032
rect 508280 1005020 508286 1005032
rect 511258 1005020 511264 1005032
rect 508280 1004992 511264 1005020
rect 508280 1004980 508286 1004992
rect 511258 1004980 511264 1004992
rect 511316 1004980 511322 1005032
rect 149882 1004912 149888 1004964
rect 149940 1004952 149946 1004964
rect 152918 1004952 152924 1004964
rect 149940 1004924 152924 1004952
rect 149940 1004912 149946 1004924
rect 152918 1004912 152924 1004924
rect 152976 1004912 152982 1004964
rect 154390 1004912 154396 1004964
rect 154448 1004952 154454 1004964
rect 160646 1004952 160652 1004964
rect 154448 1004924 160652 1004952
rect 154448 1004912 154454 1004924
rect 160646 1004912 160652 1004924
rect 160704 1004912 160710 1004964
rect 209222 1004912 209228 1004964
rect 209280 1004952 209286 1004964
rect 211798 1004952 211804 1004964
rect 209280 1004924 211804 1004952
rect 209280 1004912 209286 1004924
rect 211798 1004912 211804 1004924
rect 211856 1004912 211862 1004964
rect 305822 1004912 305828 1004964
rect 305880 1004952 305886 1004964
rect 308950 1004952 308956 1004964
rect 305880 1004924 308956 1004952
rect 305880 1004912 305886 1004924
rect 308950 1004912 308956 1004924
rect 309008 1004912 309014 1004964
rect 353202 1004912 353208 1004964
rect 353260 1004952 353266 1004964
rect 355686 1004952 355692 1004964
rect 353260 1004924 355692 1004952
rect 353260 1004912 353266 1004924
rect 355686 1004912 355692 1004924
rect 355744 1004912 355750 1004964
rect 361390 1004912 361396 1004964
rect 361448 1004952 361454 1004964
rect 365162 1004952 365168 1004964
rect 361448 1004924 365168 1004952
rect 361448 1004912 361454 1004924
rect 365162 1004912 365168 1004924
rect 365220 1004912 365226 1004964
rect 429194 1004912 429200 1004964
rect 429252 1004952 429258 1004964
rect 431908 1004952 431914 1004964
rect 429252 1004924 431914 1004952
rect 429252 1004912 429258 1004924
rect 431908 1004912 431914 1004924
rect 431966 1004912 431972 1004964
rect 432414 1004844 432420 1004896
rect 432472 1004884 432478 1004896
rect 438118 1004884 438124 1004896
rect 432472 1004856 438124 1004884
rect 432472 1004844 432478 1004856
rect 438118 1004844 438124 1004856
rect 438176 1004844 438182 1004896
rect 507854 1004844 507860 1004896
rect 507912 1004884 507918 1004896
rect 510062 1004884 510068 1004896
rect 507912 1004856 510068 1004884
rect 507912 1004844 507918 1004856
rect 510062 1004844 510068 1004856
rect 510120 1004844 510126 1004896
rect 151262 1004776 151268 1004828
rect 151320 1004816 151326 1004828
rect 154114 1004816 154120 1004828
rect 151320 1004788 154120 1004816
rect 151320 1004776 151326 1004788
rect 154114 1004776 154120 1004788
rect 154172 1004776 154178 1004828
rect 159450 1004776 159456 1004828
rect 159508 1004816 159514 1004828
rect 162118 1004816 162124 1004828
rect 159508 1004788 162124 1004816
rect 159508 1004776 159514 1004788
rect 162118 1004776 162124 1004788
rect 162176 1004776 162182 1004828
rect 207198 1004776 207204 1004828
rect 207256 1004816 207262 1004828
rect 209866 1004816 209872 1004828
rect 207256 1004788 209872 1004816
rect 207256 1004776 207262 1004788
rect 209866 1004776 209872 1004788
rect 209924 1004776 209930 1004828
rect 304442 1004776 304448 1004828
rect 304500 1004816 304506 1004828
rect 306926 1004816 306932 1004828
rect 304500 1004788 306932 1004816
rect 304500 1004776 304506 1004788
rect 306926 1004776 306932 1004788
rect 306984 1004776 306990 1004828
rect 313826 1004776 313832 1004828
rect 313884 1004816 313890 1004828
rect 316034 1004816 316040 1004828
rect 313884 1004788 316040 1004816
rect 313884 1004776 313890 1004788
rect 316034 1004776 316040 1004788
rect 316092 1004776 316098 1004828
rect 364242 1004776 364248 1004828
rect 364300 1004816 364306 1004828
rect 366358 1004816 366364 1004828
rect 364300 1004788 366364 1004816
rect 364300 1004776 364306 1004788
rect 366358 1004776 366364 1004788
rect 366416 1004776 366422 1004828
rect 430022 1004776 430028 1004828
rect 430080 1004816 430086 1004828
rect 432230 1004816 432236 1004828
rect 430080 1004788 432236 1004816
rect 430080 1004776 430086 1004788
rect 432230 1004776 432236 1004788
rect 432288 1004776 432294 1004828
rect 498102 1004776 498108 1004828
rect 498160 1004816 498166 1004828
rect 499666 1004816 499672 1004828
rect 498160 1004788 499672 1004816
rect 498160 1004776 498166 1004788
rect 499666 1004776 499672 1004788
rect 499724 1004776 499730 1004828
rect 555970 1004776 555976 1004828
rect 556028 1004816 556034 1004828
rect 558178 1004816 558184 1004828
rect 556028 1004788 558184 1004816
rect 556028 1004776 556034 1004788
rect 558178 1004776 558184 1004788
rect 558236 1004776 558242 1004828
rect 94866 1004640 94872 1004692
rect 94924 1004680 94930 1004692
rect 103146 1004680 103152 1004692
rect 94924 1004652 103152 1004680
rect 94924 1004640 94930 1004652
rect 103146 1004640 103152 1004652
rect 103204 1004640 103210 1004692
rect 106182 1004640 106188 1004692
rect 106240 1004680 106246 1004692
rect 108482 1004680 108488 1004692
rect 106240 1004652 108488 1004680
rect 106240 1004640 106246 1004652
rect 108482 1004640 108488 1004652
rect 108540 1004640 108546 1004692
rect 160646 1004640 160652 1004692
rect 160704 1004680 160710 1004692
rect 162854 1004680 162860 1004692
rect 160704 1004652 162860 1004680
rect 160704 1004640 160710 1004652
rect 162854 1004640 162860 1004652
rect 162912 1004640 162918 1004692
rect 209222 1004640 209228 1004692
rect 209280 1004680 209286 1004692
rect 211154 1004680 211160 1004692
rect 209280 1004652 211160 1004680
rect 209280 1004640 209286 1004652
rect 211154 1004640 211160 1004652
rect 211212 1004640 211218 1004692
rect 212534 1004640 212540 1004692
rect 212592 1004680 212598 1004692
rect 217318 1004680 217324 1004692
rect 212592 1004652 217324 1004680
rect 212592 1004640 212598 1004652
rect 217318 1004640 217324 1004652
rect 217376 1004640 217382 1004692
rect 305638 1004640 305644 1004692
rect 305696 1004680 305702 1004692
rect 308122 1004680 308128 1004692
rect 305696 1004652 308128 1004680
rect 305696 1004640 305702 1004652
rect 308122 1004640 308128 1004652
rect 308180 1004640 308186 1004692
rect 315482 1004640 315488 1004692
rect 315540 1004680 315546 1004692
rect 318058 1004680 318064 1004692
rect 315540 1004652 318064 1004680
rect 315540 1004640 315546 1004652
rect 318058 1004640 318064 1004652
rect 318116 1004640 318122 1004692
rect 354582 1004640 354588 1004692
rect 354640 1004680 354646 1004692
rect 355686 1004680 355692 1004692
rect 354640 1004652 355692 1004680
rect 354640 1004640 354646 1004652
rect 355686 1004640 355692 1004652
rect 355744 1004640 355750 1004692
rect 362586 1004640 362592 1004692
rect 362644 1004680 362650 1004692
rect 364978 1004680 364984 1004692
rect 362644 1004652 364984 1004680
rect 362644 1004640 362650 1004652
rect 364978 1004640 364984 1004652
rect 365036 1004640 365042 1004692
rect 431678 1004640 431684 1004692
rect 431736 1004680 431742 1004692
rect 433518 1004680 433524 1004692
rect 431736 1004652 433524 1004680
rect 431736 1004640 431742 1004652
rect 433518 1004640 433524 1004652
rect 433576 1004640 433582 1004692
rect 499482 1004640 499488 1004692
rect 499540 1004680 499546 1004692
rect 501322 1004680 501328 1004692
rect 499540 1004652 501328 1004680
rect 499540 1004640 499546 1004652
rect 501322 1004640 501328 1004652
rect 501380 1004640 501386 1004692
rect 509050 1004640 509056 1004692
rect 509108 1004680 509114 1004692
rect 509108 1004652 509234 1004680
rect 509108 1004640 509114 1004652
rect 364518 1004504 364524 1004556
rect 364576 1004544 364582 1004556
rect 366542 1004544 366548 1004556
rect 364576 1004516 366548 1004544
rect 364576 1004504 364582 1004516
rect 366542 1004504 366548 1004516
rect 366600 1004504 366606 1004556
rect 509206 1004544 509234 1004652
rect 510338 1004640 510344 1004692
rect 510396 1004680 510402 1004692
rect 515398 1004680 515404 1004692
rect 510396 1004652 515404 1004680
rect 510396 1004640 510402 1004652
rect 515398 1004640 515404 1004652
rect 515456 1004640 515462 1004692
rect 557626 1004640 557632 1004692
rect 557684 1004680 557690 1004692
rect 559558 1004680 559564 1004692
rect 557684 1004652 559564 1004680
rect 557684 1004640 557690 1004652
rect 559558 1004640 559564 1004652
rect 559616 1004640 559622 1004692
rect 561674 1004640 561680 1004692
rect 561732 1004680 561738 1004692
rect 566458 1004680 566464 1004692
rect 561732 1004652 566464 1004680
rect 561732 1004640 561738 1004652
rect 566458 1004640 566464 1004652
rect 566516 1004640 566522 1004692
rect 510798 1004544 510804 1004556
rect 509206 1004516 510804 1004544
rect 510798 1004504 510804 1004516
rect 510856 1004504 510862 1004556
rect 432874 1004028 432880 1004080
rect 432932 1004068 432938 1004080
rect 462314 1004068 462320 1004080
rect 432932 1004040 462320 1004068
rect 432932 1004028 432938 1004040
rect 462314 1004028 462320 1004040
rect 462372 1004028 462378 1004080
rect 425514 1003892 425520 1003944
rect 425572 1003932 425578 1003944
rect 467834 1003932 467840 1003944
rect 425572 1003904 467840 1003932
rect 425572 1003892 425578 1003904
rect 467834 1003892 467840 1003904
rect 467892 1003892 467898 1003944
rect 505370 1003892 505376 1003944
rect 505428 1003932 505434 1003944
rect 516594 1003932 516600 1003944
rect 505428 1003904 516600 1003932
rect 505428 1003892 505434 1003904
rect 516594 1003892 516600 1003904
rect 516652 1003892 516658 1003944
rect 445018 1002804 445024 1002856
rect 445076 1002844 445082 1002856
rect 454678 1002844 454684 1002856
rect 445076 1002816 454684 1002844
rect 445076 1002804 445082 1002816
rect 454678 1002804 454684 1002816
rect 454736 1002804 454742 1002856
rect 558822 1002736 558828 1002788
rect 558880 1002776 558886 1002788
rect 562318 1002776 562324 1002788
rect 558880 1002748 562324 1002776
rect 558880 1002736 558886 1002748
rect 562318 1002736 562324 1002748
rect 562376 1002736 562382 1002788
rect 424686 1002668 424692 1002720
rect 424744 1002708 424750 1002720
rect 446214 1002708 446220 1002720
rect 424744 1002680 446220 1002708
rect 424744 1002668 424750 1002680
rect 446214 1002668 446220 1002680
rect 446272 1002668 446278 1002720
rect 97258 1002600 97264 1002652
rect 97316 1002640 97322 1002652
rect 102318 1002640 102324 1002652
rect 97316 1002612 102324 1002640
rect 97316 1002600 97322 1002612
rect 102318 1002600 102324 1002612
rect 102376 1002600 102382 1002652
rect 557994 1002600 558000 1002652
rect 558052 1002640 558058 1002652
rect 560294 1002640 560300 1002652
rect 558052 1002612 560300 1002640
rect 558052 1002600 558058 1002612
rect 560294 1002600 560300 1002612
rect 560352 1002600 560358 1002652
rect 105998 1002532 106004 1002584
rect 106056 1002572 106062 1002584
rect 109494 1002572 109500 1002584
rect 106056 1002544 109500 1002572
rect 106056 1002532 106062 1002544
rect 109494 1002532 109500 1002544
rect 109552 1002532 109558 1002584
rect 427814 1002532 427820 1002584
rect 427872 1002572 427878 1002584
rect 468754 1002572 468760 1002584
rect 427872 1002544 468760 1002572
rect 427872 1002532 427878 1002544
rect 468754 1002532 468760 1002544
rect 468812 1002532 468818 1002584
rect 502518 1002532 502524 1002584
rect 502576 1002572 502582 1002584
rect 516042 1002572 516048 1002584
rect 502576 1002544 516048 1002572
rect 502576 1002532 502582 1002544
rect 516042 1002532 516048 1002544
rect 516100 1002532 516106 1002584
rect 563054 1002532 563060 1002584
rect 563112 1002572 563118 1002584
rect 571242 1002572 571248 1002584
rect 563112 1002544 571248 1002572
rect 563112 1002532 563118 1002544
rect 571242 1002532 571248 1002544
rect 571300 1002532 571306 1002584
rect 98638 1002464 98644 1002516
rect 98696 1002504 98702 1002516
rect 101950 1002504 101956 1002516
rect 98696 1002476 101956 1002504
rect 98696 1002464 98702 1002476
rect 101950 1002464 101956 1002476
rect 102008 1002464 102014 1002516
rect 157426 1002464 157432 1002516
rect 157484 1002504 157490 1002516
rect 159358 1002504 159364 1002516
rect 157484 1002476 159364 1002504
rect 157484 1002464 157490 1002476
rect 159358 1002464 159364 1002476
rect 159416 1002464 159422 1002516
rect 203334 1002464 203340 1002516
rect 203392 1002504 203398 1002516
rect 206370 1002504 206376 1002516
rect 203392 1002476 206376 1002504
rect 203392 1002464 203398 1002476
rect 206370 1002464 206376 1002476
rect 206428 1002464 206434 1002516
rect 251818 1002464 251824 1002516
rect 251876 1002504 251882 1002516
rect 255314 1002504 255320 1002516
rect 251876 1002476 255320 1002504
rect 251876 1002464 251882 1002476
rect 255314 1002464 255320 1002476
rect 255372 1002464 255378 1002516
rect 261018 1002464 261024 1002516
rect 261076 1002504 261082 1002516
rect 264238 1002504 264244 1002516
rect 261076 1002476 264244 1002504
rect 261076 1002464 261082 1002476
rect 264238 1002464 264244 1002476
rect 264296 1002464 264302 1002516
rect 108022 1002396 108028 1002448
rect 108080 1002436 108086 1002448
rect 110414 1002436 110420 1002448
rect 108080 1002408 110420 1002436
rect 108080 1002396 108086 1002408
rect 110414 1002396 110420 1002408
rect 110472 1002396 110478 1002448
rect 557994 1002396 558000 1002448
rect 558052 1002436 558058 1002448
rect 561030 1002436 561036 1002448
rect 558052 1002408 561036 1002436
rect 558052 1002396 558058 1002408
rect 561030 1002396 561036 1002408
rect 561088 1002396 561094 1002448
rect 97442 1002328 97448 1002380
rect 97500 1002368 97506 1002380
rect 100294 1002368 100300 1002380
rect 97500 1002340 100300 1002368
rect 97500 1002328 97506 1002340
rect 100294 1002328 100300 1002340
rect 100352 1002328 100358 1002380
rect 158622 1002328 158628 1002380
rect 158680 1002368 158686 1002380
rect 160370 1002368 160376 1002380
rect 158680 1002340 160376 1002368
rect 158680 1002328 158686 1002340
rect 160370 1002328 160376 1002340
rect 160428 1002328 160434 1002380
rect 211246 1002328 211252 1002380
rect 211304 1002368 211310 1002380
rect 215938 1002368 215944 1002380
rect 211304 1002340 215944 1002368
rect 211304 1002328 211310 1002340
rect 215938 1002328 215944 1002340
rect 215996 1002328 216002 1002380
rect 253106 1002328 253112 1002380
rect 253164 1002368 253170 1002380
rect 256142 1002368 256148 1002380
rect 253164 1002340 256148 1002368
rect 253164 1002328 253170 1002340
rect 256142 1002328 256148 1002340
rect 256200 1002328 256206 1002380
rect 310146 1002328 310152 1002380
rect 310204 1002368 310210 1002380
rect 311894 1002368 311900 1002380
rect 310204 1002340 311900 1002368
rect 310204 1002328 310210 1002340
rect 311894 1002328 311900 1002340
rect 311952 1002328 311958 1002380
rect 358538 1002328 358544 1002380
rect 358596 1002368 358602 1002380
rect 360838 1002368 360844 1002380
rect 358596 1002340 360844 1002368
rect 358596 1002328 358602 1002340
rect 360838 1002328 360844 1002340
rect 360896 1002328 360902 1002380
rect 105630 1002260 105636 1002312
rect 105688 1002300 105694 1002312
rect 107838 1002300 107844 1002312
rect 105688 1002272 107844 1002300
rect 105688 1002260 105694 1002272
rect 107838 1002260 107844 1002272
rect 107896 1002260 107902 1002312
rect 108482 1002260 108488 1002312
rect 108540 1002300 108546 1002312
rect 111058 1002300 111064 1002312
rect 108540 1002272 111064 1002300
rect 108540 1002260 108546 1002272
rect 111058 1002260 111064 1002272
rect 111116 1002260 111122 1002312
rect 153930 1002260 153936 1002312
rect 153988 1002300 153994 1002312
rect 155770 1002300 155776 1002312
rect 153988 1002272 155776 1002300
rect 153988 1002260 153994 1002272
rect 155770 1002260 155776 1002272
rect 155828 1002260 155834 1002312
rect 551922 1002260 551928 1002312
rect 551980 1002300 551986 1002312
rect 554314 1002300 554320 1002312
rect 551980 1002272 554320 1002300
rect 551980 1002260 551986 1002272
rect 554314 1002260 554320 1002272
rect 554372 1002260 554378 1002312
rect 560478 1002260 560484 1002312
rect 560536 1002300 560542 1002312
rect 563054 1002300 563060 1002312
rect 560536 1002272 563060 1002300
rect 560536 1002260 560542 1002272
rect 563054 1002260 563060 1002272
rect 563112 1002260 563118 1002312
rect 98822 1002192 98828 1002244
rect 98880 1002232 98886 1002244
rect 101122 1002232 101128 1002244
rect 98880 1002204 101128 1002232
rect 98880 1002192 98886 1002204
rect 101122 1002192 101128 1002204
rect 101180 1002192 101186 1002244
rect 156598 1002192 156604 1002244
rect 156656 1002232 156662 1002244
rect 158714 1002232 158720 1002244
rect 156656 1002204 158720 1002232
rect 156656 1002192 156662 1002204
rect 158714 1002192 158720 1002204
rect 158772 1002192 158778 1002244
rect 204898 1002192 204904 1002244
rect 204956 1002232 204962 1002244
rect 206370 1002232 206376 1002244
rect 204956 1002204 206376 1002232
rect 204956 1002192 204962 1002204
rect 206370 1002192 206376 1002204
rect 206428 1002192 206434 1002244
rect 252002 1002192 252008 1002244
rect 252060 1002232 252066 1002244
rect 254486 1002232 254492 1002244
rect 252060 1002204 254492 1002232
rect 252060 1002192 252066 1002204
rect 254486 1002192 254492 1002204
rect 254544 1002192 254550 1002244
rect 303062 1002192 303068 1002244
rect 303120 1002232 303126 1002244
rect 306098 1002232 306104 1002244
rect 303120 1002204 306104 1002232
rect 303120 1002192 303126 1002204
rect 306098 1002192 306104 1002204
rect 306156 1002192 306162 1002244
rect 359366 1002192 359372 1002244
rect 359424 1002192 359430 1002244
rect 500678 1002192 500684 1002244
rect 500736 1002232 500742 1002244
rect 503346 1002232 503352 1002244
rect 500736 1002204 503352 1002232
rect 500736 1002192 500742 1002204
rect 503346 1002192 503352 1002204
rect 503404 1002192 503410 1002244
rect 104802 1002124 104808 1002176
rect 104860 1002164 104866 1002176
rect 106366 1002164 106372 1002176
rect 104860 1002136 106372 1002164
rect 104860 1002124 104866 1002136
rect 106366 1002124 106372 1002136
rect 106424 1002124 106430 1002176
rect 106826 1002124 106832 1002176
rect 106884 1002164 106890 1002176
rect 109034 1002164 109040 1002176
rect 106884 1002136 109040 1002164
rect 106884 1002124 106890 1002136
rect 109034 1002124 109040 1002136
rect 109092 1002124 109098 1002176
rect 152642 1002124 152648 1002176
rect 152700 1002164 152706 1002176
rect 154574 1002164 154580 1002176
rect 152700 1002136 154580 1002164
rect 152700 1002124 152706 1002136
rect 154574 1002124 154580 1002136
rect 154632 1002124 154638 1002176
rect 96522 1002056 96528 1002108
rect 96580 1002096 96586 1002108
rect 99098 1002096 99104 1002108
rect 96580 1002068 99104 1002096
rect 96580 1002056 96586 1002068
rect 99098 1002056 99104 1002068
rect 99156 1002056 99162 1002108
rect 100202 1002056 100208 1002108
rect 100260 1002096 100266 1002108
rect 103146 1002096 103152 1002108
rect 100260 1002068 103152 1002096
rect 100260 1002056 100266 1002068
rect 103146 1002056 103152 1002068
rect 103204 1002056 103210 1002108
rect 109678 1002056 109684 1002108
rect 109736 1002096 109742 1002108
rect 111886 1002096 111892 1002108
rect 109736 1002068 111892 1002096
rect 109736 1002056 109742 1002068
rect 111886 1002056 111892 1002068
rect 111944 1002056 111950 1002108
rect 148962 1002056 148968 1002108
rect 149020 1002096 149026 1002108
rect 150894 1002096 150900 1002108
rect 149020 1002068 150900 1002096
rect 149020 1002056 149026 1002068
rect 150894 1002056 150900 1002068
rect 150952 1002056 150958 1002108
rect 154942 1002056 154948 1002108
rect 155000 1002096 155006 1002108
rect 157334 1002096 157340 1002108
rect 155000 1002068 157340 1002096
rect 155000 1002056 155006 1002068
rect 157334 1002056 157340 1002068
rect 157392 1002056 157398 1002108
rect 211246 1002056 211252 1002108
rect 211304 1002096 211310 1002108
rect 213178 1002096 213184 1002108
rect 211304 1002068 213184 1002096
rect 211304 1002056 211310 1002068
rect 213178 1002056 213184 1002068
rect 213236 1002056 213242 1002108
rect 250990 1002056 250996 1002108
rect 251048 1002096 251054 1002108
rect 253290 1002096 253296 1002108
rect 251048 1002068 253296 1002096
rect 251048 1002056 251054 1002068
rect 253290 1002056 253296 1002068
rect 253348 1002056 253354 1002108
rect 253474 1002056 253480 1002108
rect 253532 1002096 253538 1002108
rect 256142 1002096 256148 1002108
rect 253532 1002068 256148 1002096
rect 253532 1002056 253538 1002068
rect 256142 1002056 256148 1002068
rect 256200 1002056 256206 1002108
rect 263502 1002056 263508 1002108
rect 263560 1002096 263566 1002108
rect 265618 1002096 265624 1002108
rect 263560 1002068 265624 1002096
rect 263560 1002056 263566 1002068
rect 265618 1002056 265624 1002068
rect 265676 1002056 265682 1002108
rect 307018 1002056 307024 1002108
rect 307076 1002096 307082 1002108
rect 308950 1002096 308956 1002108
rect 307076 1002068 308956 1002096
rect 307076 1002056 307082 1002068
rect 308950 1002056 308956 1002068
rect 309008 1002056 309014 1002108
rect 310974 1002056 310980 1002108
rect 311032 1002096 311038 1002108
rect 313274 1002096 313280 1002108
rect 311032 1002068 313280 1002096
rect 311032 1002056 311038 1002068
rect 313274 1002056 313280 1002068
rect 313332 1002056 313338 1002108
rect 105998 1001988 106004 1002040
rect 106056 1002028 106062 1002040
rect 107746 1002028 107752 1002040
rect 106056 1002000 107752 1002028
rect 106056 1001988 106062 1002000
rect 107746 1001988 107752 1002000
rect 107804 1001988 107810 1002040
rect 152458 1001988 152464 1002040
rect 152516 1002028 152522 1002040
rect 153746 1002028 153752 1002040
rect 152516 1002000 153752 1002028
rect 152516 1001988 152522 1002000
rect 153746 1001988 153752 1002000
rect 153804 1001988 153810 1002040
rect 358722 1001988 358728 1002040
rect 358780 1002028 358786 1002040
rect 359384 1002028 359412 1002192
rect 560018 1002124 560024 1002176
rect 560076 1002164 560082 1002176
rect 562502 1002164 562508 1002176
rect 560076 1002136 562508 1002164
rect 560076 1002124 560082 1002136
rect 562502 1002124 562508 1002136
rect 562560 1002124 562566 1002176
rect 360562 1002056 360568 1002108
rect 360620 1002096 360626 1002108
rect 363598 1002096 363604 1002108
rect 360620 1002068 363604 1002096
rect 360620 1002056 360626 1002068
rect 363598 1002056 363604 1002068
rect 363656 1002056 363662 1002108
rect 433334 1002056 433340 1002108
rect 433392 1002096 433398 1002108
rect 436738 1002096 436744 1002108
rect 433392 1002068 436744 1002096
rect 433392 1002056 433398 1002068
rect 436738 1002056 436744 1002068
rect 436796 1002056 436802 1002108
rect 502242 1002056 502248 1002108
rect 502300 1002096 502306 1002108
rect 504174 1002096 504180 1002108
rect 502300 1002068 504180 1002096
rect 502300 1002056 502306 1002068
rect 504174 1002056 504180 1002068
rect 504232 1002056 504238 1002108
rect 509878 1002056 509884 1002108
rect 509936 1002096 509942 1002108
rect 512638 1002096 512644 1002108
rect 509936 1002068 512644 1002096
rect 509936 1002056 509942 1002068
rect 512638 1002056 512644 1002068
rect 512696 1002056 512702 1002108
rect 358780 1002000 359412 1002028
rect 358780 1001988 358786 1002000
rect 553302 1001988 553308 1002040
rect 553360 1002028 553366 1002040
rect 553946 1002028 553952 1002040
rect 553360 1002000 553952 1002028
rect 553360 1001988 553366 1002000
rect 553946 1001988 553952 1002000
rect 554004 1001988 554010 1002040
rect 560846 1001988 560852 1002040
rect 560904 1002028 560910 1002040
rect 565078 1002028 565084 1002040
rect 560904 1002000 565084 1002028
rect 560904 1001988 560910 1002000
rect 565078 1001988 565084 1002000
rect 565136 1001988 565142 1002040
rect 96338 1001920 96344 1001972
rect 96396 1001960 96402 1001972
rect 98270 1001960 98276 1001972
rect 96396 1001932 98276 1001960
rect 96396 1001920 96402 1001932
rect 98270 1001920 98276 1001932
rect 98328 1001920 98334 1001972
rect 100018 1001920 100024 1001972
rect 100076 1001960 100082 1001972
rect 101950 1001960 101956 1001972
rect 100076 1001932 101956 1001960
rect 100076 1001920 100082 1001932
rect 101950 1001920 101956 1001932
rect 102008 1001920 102014 1001972
rect 108850 1001920 108856 1001972
rect 108908 1001960 108914 1001972
rect 112070 1001960 112076 1001972
rect 108908 1001932 112076 1001960
rect 108908 1001920 108914 1001932
rect 112070 1001920 112076 1001932
rect 112128 1001920 112134 1001972
rect 147582 1001920 147588 1001972
rect 147640 1001960 147646 1001972
rect 149238 1001960 149244 1001972
rect 147640 1001932 149244 1001960
rect 147640 1001920 147646 1001932
rect 149238 1001920 149244 1001932
rect 149296 1001920 149302 1001972
rect 154574 1001920 154580 1001972
rect 154632 1001960 154638 1001972
rect 155770 1001960 155776 1001972
rect 154632 1001932 155776 1001960
rect 154632 1001920 154638 1001932
rect 155770 1001920 155776 1001932
rect 155828 1001920 155834 1001972
rect 157794 1001920 157800 1001972
rect 157852 1001960 157858 1001972
rect 160186 1001960 160192 1001972
rect 157852 1001932 160192 1001960
rect 157852 1001920 157858 1001932
rect 160186 1001920 160192 1001932
rect 160244 1001920 160250 1001972
rect 195330 1001920 195336 1001972
rect 195388 1001960 195394 1001972
rect 203886 1001960 203892 1001972
rect 195388 1001932 203892 1001960
rect 195388 1001920 195394 1001932
rect 203886 1001920 203892 1001932
rect 203944 1001920 203950 1001972
rect 204162 1001920 204168 1001972
rect 204220 1001960 204226 1001972
rect 205542 1001960 205548 1001972
rect 204220 1001932 205548 1001960
rect 204220 1001920 204226 1001932
rect 205542 1001920 205548 1001932
rect 205600 1001920 205606 1001972
rect 212074 1001920 212080 1001972
rect 212132 1001960 212138 1001972
rect 213914 1001960 213920 1001972
rect 212132 1001932 213920 1001960
rect 212132 1001920 212138 1001932
rect 213914 1001920 213920 1001932
rect 213972 1001920 213978 1001972
rect 249702 1001920 249708 1001972
rect 249760 1001960 249766 1001972
rect 252462 1001960 252468 1001972
rect 249760 1001932 252468 1001960
rect 249760 1001920 249766 1001932
rect 252462 1001920 252468 1001932
rect 252520 1001920 252526 1001972
rect 261018 1001920 261024 1001972
rect 261076 1001960 261082 1001972
rect 263594 1001960 263600 1001972
rect 261076 1001932 263600 1001960
rect 261076 1001920 261082 1001932
rect 263594 1001920 263600 1001932
rect 263652 1001920 263658 1001972
rect 263870 1001920 263876 1001972
rect 263928 1001960 263934 1001972
rect 266998 1001960 267004 1001972
rect 263928 1001932 267004 1001960
rect 263928 1001920 263934 1001932
rect 266998 1001920 267004 1001932
rect 267056 1001920 267062 1001972
rect 302878 1001920 302884 1001972
rect 302936 1001960 302942 1001972
rect 306098 1001960 306104 1001972
rect 302936 1001932 306104 1001960
rect 302936 1001920 302942 1001932
rect 306098 1001920 306104 1001932
rect 306156 1001920 306162 1001972
rect 308398 1001920 308404 1001972
rect 308456 1001960 308462 1001972
rect 309778 1001960 309784 1001972
rect 308456 1001932 309784 1001960
rect 308456 1001920 308462 1001932
rect 309778 1001920 309784 1001932
rect 309836 1001920 309842 1001972
rect 312630 1001920 312636 1001972
rect 312688 1001960 312694 1001972
rect 314654 1001960 314660 1001972
rect 312688 1001932 314660 1001960
rect 312688 1001920 312694 1001932
rect 314654 1001920 314660 1001932
rect 314712 1001920 314718 1001972
rect 351822 1001920 351828 1001972
rect 351880 1001960 351886 1001972
rect 354030 1001960 354036 1001972
rect 351880 1001932 354036 1001960
rect 351880 1001920 351886 1001932
rect 354030 1001920 354036 1001932
rect 354088 1001920 354094 1001972
rect 355962 1001920 355968 1001972
rect 356020 1001960 356026 1001972
rect 357342 1001960 357348 1001972
rect 356020 1001932 357348 1001960
rect 356020 1001920 356026 1001932
rect 357342 1001920 357348 1001932
rect 357400 1001920 357406 1001972
rect 360194 1001920 360200 1001972
rect 360252 1001960 360258 1001972
rect 362218 1001960 362224 1001972
rect 360252 1001932 362224 1001960
rect 360252 1001920 360258 1001932
rect 362218 1001920 362224 1001932
rect 362276 1001920 362282 1001972
rect 365898 1001920 365904 1001972
rect 365956 1001960 365962 1001972
rect 369118 1001960 369124 1001972
rect 365956 1001932 369124 1001960
rect 365956 1001920 365962 1001932
rect 369118 1001920 369124 1001932
rect 369176 1001920 369182 1001972
rect 419442 1001920 419448 1001972
rect 419500 1001960 419506 1001972
rect 421466 1001960 421472 1001972
rect 419500 1001932 421472 1001960
rect 419500 1001920 419506 1001932
rect 421466 1001920 421472 1001932
rect 421524 1001920 421530 1001972
rect 425054 1001920 425060 1001972
rect 425112 1001960 425118 1001972
rect 426342 1001960 426348 1001972
rect 425112 1001932 426348 1001960
rect 425112 1001920 425118 1001932
rect 426342 1001920 426348 1001932
rect 426400 1001920 426406 1001972
rect 426526 1001920 426532 1001972
rect 426584 1001960 426590 1001972
rect 427814 1001960 427820 1001972
rect 426584 1001932 427820 1001960
rect 426584 1001920 426590 1001932
rect 427814 1001920 427820 1001932
rect 427872 1001920 427878 1001972
rect 428366 1001920 428372 1001972
rect 428424 1001960 428430 1001972
rect 431218 1001960 431224 1001972
rect 428424 1001932 431224 1001960
rect 428424 1001920 428430 1001932
rect 431218 1001920 431224 1001932
rect 431276 1001920 431282 1001972
rect 467834 1001920 467840 1001972
rect 467892 1001960 467898 1001972
rect 472618 1001960 472624 1001972
rect 467892 1001932 472624 1001960
rect 467892 1001920 467898 1001932
rect 472618 1001920 472624 1001932
rect 472676 1001920 472682 1001972
rect 496722 1001920 496728 1001972
rect 496780 1001960 496786 1001972
rect 498470 1001960 498476 1001972
rect 496780 1001932 498476 1001960
rect 496780 1001920 496786 1001932
rect 498470 1001920 498476 1001932
rect 498528 1001920 498534 1001972
rect 500862 1001920 500868 1001972
rect 500920 1001960 500926 1001972
rect 502518 1001960 502524 1001972
rect 500920 1001932 502524 1001960
rect 500920 1001920 500926 1001932
rect 502518 1001920 502524 1001932
rect 502576 1001920 502582 1001972
rect 503346 1001920 503352 1001972
rect 503404 1001960 503410 1001972
rect 504358 1001960 504364 1001972
rect 503404 1001932 504364 1001960
rect 503404 1001920 503410 1001932
rect 504358 1001920 504364 1001932
rect 504416 1001920 504422 1001972
rect 506198 1001920 506204 1001972
rect 506256 1001960 506262 1001972
rect 507854 1001960 507860 1001972
rect 506256 1001932 507860 1001960
rect 506256 1001920 506262 1001932
rect 507854 1001920 507860 1001932
rect 507912 1001920 507918 1001972
rect 558822 1001920 558828 1001972
rect 558880 1001960 558886 1001972
rect 560386 1001960 560392 1001972
rect 558880 1001932 560392 1001960
rect 558880 1001920 558886 1001932
rect 560386 1001920 560392 1001932
rect 560444 1001920 560450 1001972
rect 439498 1001172 439504 1001224
rect 439556 1001212 439562 1001224
rect 446398 1001212 446404 1001224
rect 439556 1001184 446404 1001212
rect 439556 1001172 439562 1001184
rect 446398 1001172 446404 1001184
rect 446456 1001172 446462 1001224
rect 500678 1001172 500684 1001224
rect 500736 1001212 500742 1001224
rect 519998 1001212 520004 1001224
rect 500736 1001184 520004 1001212
rect 500736 1001172 500742 1001184
rect 519998 1001172 520004 1001184
rect 520056 1001172 520062 1001224
rect 298462 1000424 298468 1000476
rect 298520 1000464 298526 1000476
rect 309134 1000464 309140 1000476
rect 298520 1000436 309140 1000464
rect 298520 1000424 298526 1000436
rect 309134 1000424 309140 1000436
rect 309192 1000424 309198 1000476
rect 92658 999744 92664 999796
rect 92716 999784 92722 999796
rect 98822 999784 98828 999796
rect 92716 999756 98828 999784
rect 92716 999744 92722 999756
rect 98822 999744 98828 999756
rect 98880 999744 98886 999796
rect 427814 999744 427820 999796
rect 427872 999784 427878 999796
rect 437474 999784 437480 999796
rect 427872 999756 437480 999784
rect 427872 999744 427878 999756
rect 437474 999744 437480 999756
rect 437532 999744 437538 999796
rect 446214 999744 446220 999796
rect 446272 999784 446278 999796
rect 459554 999784 459560 999796
rect 446272 999756 459560 999784
rect 446272 999744 446278 999756
rect 459554 999744 459560 999756
rect 459612 999744 459618 999796
rect 195974 999132 195980 999184
rect 196032 999172 196038 999184
rect 203518 999172 203524 999184
rect 196032 999144 203524 999172
rect 196032 999132 196038 999144
rect 203518 999132 203524 999144
rect 203576 999132 203582 999184
rect 249334 999132 249340 999184
rect 249392 999172 249398 999184
rect 250438 999172 250444 999184
rect 249392 999144 250444 999172
rect 249392 999132 249398 999144
rect 250438 999132 250444 999144
rect 250496 999132 250502 999184
rect 301038 999132 301044 999184
rect 301096 999172 301102 999184
rect 303062 999172 303068 999184
rect 301096 999144 303068 999172
rect 301096 999132 301102 999144
rect 303062 999132 303068 999144
rect 303120 999132 303126 999184
rect 373994 999132 374000 999184
rect 374052 999172 374058 999184
rect 381722 999172 381728 999184
rect 374052 999144 381728 999172
rect 374052 999132 374058 999144
rect 381722 999132 381728 999144
rect 381780 999132 381786 999184
rect 438118 999064 438124 999116
rect 438176 999104 438182 999116
rect 443454 999104 443460 999116
rect 438176 999076 443460 999104
rect 438176 999064 438182 999076
rect 443454 999064 443460 999076
rect 443512 999064 443518 999116
rect 449158 999064 449164 999116
rect 449216 999104 449222 999116
rect 451734 999104 451740 999116
rect 449216 999076 451740 999104
rect 449216 999064 449222 999076
rect 451734 999064 451740 999076
rect 451792 999064 451798 999116
rect 516594 999064 516600 999116
rect 516652 999104 516658 999116
rect 520182 999104 520188 999116
rect 516652 999076 520188 999104
rect 516652 999064 516658 999076
rect 520182 999064 520188 999076
rect 520240 999064 520246 999116
rect 300854 998996 300860 999048
rect 300912 999036 300918 999048
rect 304442 999036 304448 999048
rect 300912 999008 304448 999036
rect 300912 998996 300918 999008
rect 304442 998996 304448 999008
rect 304500 998996 304506 999048
rect 451918 998996 451924 999048
rect 451976 999036 451982 999048
rect 456794 999036 456800 999048
rect 451976 999008 456800 999036
rect 451976 998996 451982 999008
rect 456794 998996 456800 999008
rect 456852 998996 456858 999048
rect 199838 998792 199844 998844
rect 199896 998832 199902 998844
rect 199896 998804 205634 998832
rect 199896 998792 199902 998804
rect 199378 998656 199384 998708
rect 199436 998696 199442 998708
rect 204346 998696 204352 998708
rect 199436 998668 204352 998696
rect 199436 998656 199442 998668
rect 204346 998656 204352 998668
rect 204404 998656 204410 998708
rect 196618 998520 196624 998572
rect 196676 998560 196682 998572
rect 202690 998560 202696 998572
rect 196676 998532 202696 998560
rect 196676 998520 196682 998532
rect 202690 998520 202696 998532
rect 202748 998520 202754 998572
rect 205606 998560 205634 998804
rect 371878 998792 371884 998844
rect 371936 998832 371942 998844
rect 383102 998832 383108 998844
rect 371936 998804 383108 998832
rect 371936 998792 371942 998804
rect 383102 998792 383108 998804
rect 383160 998792 383166 998844
rect 443638 998724 443644 998776
rect 443696 998764 443702 998776
rect 445754 998764 445760 998776
rect 443696 998736 445760 998764
rect 443696 998724 443702 998736
rect 445754 998724 445760 998736
rect 445812 998724 445818 998776
rect 353202 998656 353208 998708
rect 353260 998696 353266 998708
rect 372890 998696 372896 998708
rect 353260 998668 372896 998696
rect 353260 998656 353266 998668
rect 372890 998656 372896 998668
rect 372948 998656 372954 998708
rect 553302 998588 553308 998640
rect 553360 998628 553366 998640
rect 555142 998628 555148 998640
rect 553360 998600 555148 998628
rect 553360 998588 553366 998600
rect 555142 998588 555148 998600
rect 555200 998588 555206 998640
rect 206278 998560 206284 998572
rect 205606 998532 206284 998560
rect 206278 998520 206284 998532
rect 206336 998520 206342 998572
rect 355962 998520 355968 998572
rect 356020 998560 356026 998572
rect 376294 998560 376300 998572
rect 356020 998532 376300 998560
rect 356020 998520 356026 998532
rect 376294 998520 376300 998532
rect 376352 998520 376358 998572
rect 516778 998520 516784 998572
rect 516836 998560 516842 998572
rect 522942 998560 522948 998572
rect 516836 998532 522948 998560
rect 516836 998520 516842 998532
rect 522942 998520 522948 998532
rect 523000 998520 523006 998572
rect 555418 998520 555424 998572
rect 555476 998560 555482 998572
rect 568482 998560 568488 998572
rect 555476 998532 568488 998560
rect 555476 998520 555482 998532
rect 568482 998520 568488 998532
rect 568540 998520 568546 998572
rect 195514 998384 195520 998436
rect 195572 998424 195578 998436
rect 204162 998424 204168 998436
rect 195572 998396 204168 998424
rect 195572 998384 195578 998396
rect 204162 998384 204168 998396
rect 204220 998384 204226 998436
rect 360838 998384 360844 998436
rect 360896 998424 360902 998436
rect 383286 998424 383292 998436
rect 360896 998396 383292 998424
rect 360896 998384 360902 998396
rect 383286 998384 383292 998396
rect 383344 998384 383350 998436
rect 446398 998384 446404 998436
rect 446456 998424 446462 998436
rect 472434 998424 472440 998436
rect 446456 998396 472440 998424
rect 446456 998384 446462 998396
rect 472434 998384 472440 998396
rect 472492 998384 472498 998436
rect 502242 998384 502248 998436
rect 502300 998424 502306 998436
rect 517054 998424 517060 998436
rect 502300 998396 517060 998424
rect 502300 998384 502306 998396
rect 517054 998384 517060 998396
rect 517112 998384 517118 998436
rect 553118 998384 553124 998436
rect 553176 998424 553182 998436
rect 569862 998424 569868 998436
rect 553176 998396 569868 998424
rect 553176 998384 553182 998396
rect 569862 998384 569868 998396
rect 569920 998384 569926 998436
rect 92290 998248 92296 998300
rect 92348 998288 92354 998300
rect 94866 998288 94872 998300
rect 92348 998260 94872 998288
rect 92348 998248 92354 998260
rect 94866 998248 94872 998260
rect 94924 998248 94930 998300
rect 202138 998180 202144 998232
rect 202196 998220 202202 998232
rect 205542 998220 205548 998232
rect 202196 998192 205548 998220
rect 202196 998180 202202 998192
rect 205542 998180 205548 998192
rect 205600 998180 205606 998232
rect 258166 998112 258172 998164
rect 258224 998152 258230 998164
rect 259454 998152 259460 998164
rect 258224 998124 259460 998152
rect 258224 998112 258230 998124
rect 259454 998112 259460 998124
rect 259512 998112 259518 998164
rect 378778 998112 378784 998164
rect 378836 998152 378842 998164
rect 381262 998152 381268 998164
rect 378836 998124 381268 998152
rect 378836 998112 378842 998124
rect 381262 998112 381268 998124
rect 381320 998112 381326 998164
rect 202690 998084 202696 998096
rect 195946 998056 202696 998084
rect 195146 997772 195152 997824
rect 195204 997812 195210 997824
rect 195946 997812 195974 998056
rect 202690 998044 202696 998056
rect 202748 998044 202754 998096
rect 260190 998044 260196 998096
rect 260248 998084 260254 998096
rect 262858 998084 262864 998096
rect 260248 998056 262864 998084
rect 260248 998044 260254 998056
rect 262858 998044 262864 998056
rect 262916 998044 262922 998096
rect 376018 998044 376024 998096
rect 376076 998084 376082 998096
rect 378410 998084 378416 998096
rect 376076 998056 378416 998084
rect 376076 998044 376082 998056
rect 378410 998044 378416 998056
rect 378468 998044 378474 998096
rect 591114 998044 591120 998096
rect 591172 998084 591178 998096
rect 625798 998084 625804 998096
rect 591172 998056 625804 998084
rect 591172 998044 591178 998056
rect 625798 998044 625804 998056
rect 625856 998044 625862 998096
rect 254578 997976 254584 998028
rect 254636 998016 254642 998028
rect 257338 998016 257344 998028
rect 254636 997988 257344 998016
rect 254636 997976 254642 997988
rect 257338 997976 257344 997988
rect 257396 997976 257402 998028
rect 198642 997908 198648 997960
rect 198700 997948 198706 997960
rect 200666 997948 200672 997960
rect 198700 997920 200672 997948
rect 198700 997908 198706 997920
rect 200666 997908 200672 997920
rect 200724 997908 200730 997960
rect 200850 997908 200856 997960
rect 200908 997948 200914 997960
rect 203518 997948 203524 997960
rect 200908 997920 203524 997948
rect 200908 997908 200914 997920
rect 203518 997908 203524 997920
rect 203576 997908 203582 997960
rect 259822 997908 259828 997960
rect 259880 997948 259886 997960
rect 262214 997948 262220 997960
rect 259880 997920 262220 997948
rect 259880 997908 259886 997920
rect 262214 997908 262220 997920
rect 262272 997908 262278 997960
rect 519998 997908 520004 997960
rect 520056 997948 520062 997960
rect 523862 997948 523868 997960
rect 520056 997920 523868 997948
rect 520056 997908 520062 997920
rect 523862 997908 523868 997920
rect 523920 997908 523926 997960
rect 549162 997908 549168 997960
rect 549220 997948 549226 997960
rect 551094 997948 551100 997960
rect 549220 997920 551100 997948
rect 549220 997908 549226 997920
rect 551094 997908 551100 997920
rect 551152 997908 551158 997960
rect 621014 997908 621020 997960
rect 621072 997948 621078 997960
rect 625614 997948 625620 997960
rect 621072 997920 625620 997948
rect 621072 997908 621078 997920
rect 625614 997908 625620 997920
rect 625672 997908 625678 997960
rect 246850 997840 246856 997892
rect 246908 997880 246914 997892
rect 249058 997880 249064 997892
rect 246908 997852 249064 997880
rect 246908 997840 246914 997852
rect 249058 997840 249064 997852
rect 249116 997840 249122 997892
rect 254762 997840 254768 997892
rect 254820 997880 254826 997892
rect 256970 997880 256976 997892
rect 254820 997852 256976 997880
rect 254820 997840 254826 997852
rect 256970 997840 256976 997852
rect 257028 997840 257034 997892
rect 195204 997784 195974 997812
rect 195204 997772 195210 997784
rect 200022 997772 200028 997824
rect 200080 997812 200086 997824
rect 201862 997812 201868 997824
rect 200080 997784 201868 997812
rect 200080 997772 200086 997784
rect 201862 997772 201868 997784
rect 201920 997772 201926 997824
rect 202322 997772 202328 997824
rect 202380 997812 202386 997824
rect 204714 997812 204720 997824
rect 202380 997784 204720 997812
rect 202380 997772 202386 997784
rect 204714 997772 204720 997784
rect 204772 997772 204778 997824
rect 260190 997772 260196 997824
rect 260248 997812 260254 997824
rect 260926 997812 260932 997824
rect 260248 997784 260932 997812
rect 260248 997772 260254 997784
rect 260926 997772 260932 997784
rect 260984 997772 260990 997824
rect 298094 997772 298100 997824
rect 298152 997812 298158 997824
rect 302878 997812 302884 997824
rect 298152 997784 302884 997812
rect 298152 997772 298158 997784
rect 302878 997772 302884 997784
rect 302936 997772 302942 997824
rect 303246 997772 303252 997824
rect 303304 997812 303310 997824
rect 305822 997812 305828 997824
rect 303304 997784 305828 997812
rect 303304 997772 303310 997784
rect 305822 997772 305828 997784
rect 305880 997772 305886 997824
rect 522482 997772 522488 997824
rect 522540 997812 522546 997824
rect 524046 997812 524052 997824
rect 522540 997784 524052 997812
rect 522540 997772 522546 997784
rect 524046 997772 524052 997784
rect 524104 997772 524110 997824
rect 547782 997772 547788 997824
rect 547840 997812 547846 997824
rect 550266 997812 550272 997824
rect 547840 997784 550272 997812
rect 547840 997772 547846 997784
rect 550266 997772 550272 997784
rect 550324 997772 550330 997824
rect 551278 997772 551284 997824
rect 551336 997812 551342 997824
rect 552290 997812 552296 997824
rect 551336 997784 552296 997812
rect 551336 997772 551342 997784
rect 552290 997772 552296 997784
rect 552348 997772 552354 997824
rect 591298 997772 591304 997824
rect 591356 997812 591362 997824
rect 625246 997812 625252 997824
rect 591356 997784 625252 997812
rect 591356 997772 591362 997784
rect 625246 997772 625252 997784
rect 625304 997772 625310 997824
rect 92474 997704 92480 997756
rect 92532 997744 92538 997756
rect 106366 997744 106372 997756
rect 92532 997716 106372 997744
rect 92532 997704 92538 997716
rect 106366 997704 106372 997716
rect 106424 997704 106430 997756
rect 144822 997704 144828 997756
rect 144880 997744 144886 997756
rect 153930 997744 153936 997756
rect 144880 997716 153936 997744
rect 144880 997704 144886 997716
rect 153930 997704 153936 997716
rect 153988 997704 153994 997756
rect 246666 997704 246672 997756
rect 246724 997744 246730 997756
rect 254762 997744 254768 997756
rect 246724 997716 254768 997744
rect 246724 997704 246730 997716
rect 254762 997704 254768 997716
rect 254820 997704 254826 997756
rect 362218 997704 362224 997756
rect 362276 997744 362282 997756
rect 372522 997744 372528 997756
rect 362276 997716 372528 997744
rect 362276 997704 362282 997716
rect 372522 997704 372528 997716
rect 372580 997704 372586 997756
rect 431218 997704 431224 997756
rect 431276 997744 431282 997756
rect 439866 997744 439872 997756
rect 431276 997716 439872 997744
rect 431276 997704 431282 997716
rect 439866 997704 439872 997716
rect 439924 997704 439930 997756
rect 500862 997704 500868 997756
rect 500920 997744 500926 997756
rect 516686 997744 516692 997756
rect 500920 997716 516692 997744
rect 500920 997704 500926 997716
rect 516686 997704 516692 997716
rect 516744 997704 516750 997756
rect 164878 997636 164884 997688
rect 164936 997676 164942 997688
rect 170306 997676 170312 997688
rect 164936 997648 170312 997676
rect 164936 997636 164942 997648
rect 170306 997636 170312 997648
rect 170364 997636 170370 997688
rect 551922 997636 551928 997688
rect 551980 997676 551986 997688
rect 621014 997676 621020 997688
rect 551980 997648 621020 997676
rect 551980 997636 551986 997648
rect 621014 997636 621020 997648
rect 621072 997636 621078 997688
rect 359458 997568 359464 997620
rect 359516 997608 359522 997620
rect 372338 997608 372344 997620
rect 359516 997580 372344 997608
rect 359516 997568 359522 997580
rect 372338 997568 372344 997580
rect 372396 997568 372402 997620
rect 425054 997568 425060 997620
rect 425112 997608 425118 997620
rect 439682 997608 439688 997620
rect 425112 997580 439688 997608
rect 425112 997568 425118 997580
rect 439682 997568 439688 997580
rect 439740 997568 439746 997620
rect 514202 997568 514208 997620
rect 514260 997608 514266 997620
rect 516870 997608 516876 997620
rect 514260 997580 516876 997608
rect 514260 997568 514266 997580
rect 516870 997568 516876 997580
rect 516928 997568 516934 997620
rect 558178 997500 558184 997552
rect 558236 997540 558242 997552
rect 590562 997540 590568 997552
rect 558236 997512 590568 997540
rect 558236 997500 558242 997512
rect 590562 997500 590568 997512
rect 590620 997500 590626 997552
rect 574738 997364 574744 997416
rect 574796 997404 574802 997416
rect 591298 997404 591304 997416
rect 574796 997376 591304 997404
rect 574796 997364 574802 997376
rect 591298 997364 591304 997376
rect 591356 997364 591362 997416
rect 144362 997296 144368 997348
rect 144420 997336 144426 997348
rect 149882 997336 149888 997348
rect 144420 997308 149888 997336
rect 144420 997296 144426 997308
rect 149882 997296 149888 997308
rect 149940 997296 149946 997348
rect 551278 997296 551284 997348
rect 551336 997336 551342 997348
rect 572714 997336 572720 997348
rect 551336 997308 572720 997336
rect 551336 997296 551342 997308
rect 572714 997296 572720 997308
rect 572772 997296 572778 997348
rect 200206 997228 200212 997280
rect 200264 997268 200270 997280
rect 203334 997268 203340 997280
rect 200264 997240 203340 997268
rect 200264 997228 200270 997240
rect 203334 997228 203340 997240
rect 203392 997228 203398 997280
rect 319438 997160 319444 997212
rect 319496 997200 319502 997212
rect 332594 997200 332600 997212
rect 319496 997172 332600 997200
rect 319496 997160 319502 997172
rect 332594 997160 332600 997172
rect 332652 997160 332658 997212
rect 556798 997160 556804 997212
rect 556856 997200 556862 997212
rect 570230 997200 570236 997212
rect 556856 997172 570236 997200
rect 556856 997160 556862 997172
rect 570230 997160 570236 997172
rect 570288 997160 570294 997212
rect 573542 997160 573548 997212
rect 573600 997200 573606 997212
rect 622394 997200 622400 997212
rect 573600 997172 622400 997200
rect 573600 997160 573606 997172
rect 622394 997160 622400 997172
rect 622452 997160 622458 997212
rect 318058 997024 318064 997076
rect 318116 997064 318122 997076
rect 349154 997064 349160 997076
rect 318116 997036 349160 997064
rect 318116 997024 318122 997036
rect 349154 997024 349160 997036
rect 349212 997024 349218 997076
rect 363598 997024 363604 997076
rect 363656 997064 363662 997076
rect 372706 997064 372712 997076
rect 363656 997036 372712 997064
rect 363656 997024 363662 997036
rect 372706 997024 372712 997036
rect 372764 997024 372770 997076
rect 437474 997024 437480 997076
rect 437532 997064 437538 997076
rect 448514 997064 448520 997076
rect 437532 997036 448520 997064
rect 437532 997024 437538 997036
rect 448514 997024 448520 997036
rect 448572 997024 448578 997076
rect 457438 997024 457444 997076
rect 457496 997064 457502 997076
rect 471790 997064 471796 997076
rect 457496 997036 471796 997064
rect 457496 997024 457502 997036
rect 471790 997024 471796 997036
rect 471848 997024 471854 997076
rect 567838 997024 567844 997076
rect 567896 997064 567902 997076
rect 618162 997064 618168 997076
rect 567896 997036 618168 997064
rect 567896 997024 567902 997036
rect 618162 997024 618168 997036
rect 618220 997024 618226 997076
rect 106918 996888 106924 996940
rect 106976 996928 106982 996940
rect 111886 996928 111892 996940
rect 106976 996900 111892 996928
rect 106976 996888 106982 996900
rect 111886 996888 111892 996900
rect 111944 996888 111950 996940
rect 566642 996888 566648 996940
rect 566700 996928 566706 996940
rect 590562 996928 590568 996940
rect 566700 996900 590568 996928
rect 566700 996888 566706 996900
rect 590562 996888 590568 996900
rect 590620 996888 590626 996940
rect 571242 996752 571248 996804
rect 571300 996792 571306 996804
rect 591114 996792 591120 996804
rect 571300 996764 591120 996792
rect 571300 996752 571306 996764
rect 591114 996752 591120 996764
rect 591172 996752 591178 996804
rect 421006 996412 421012 996464
rect 421064 996452 421070 996464
rect 425054 996452 425060 996464
rect 421064 996424 425060 996452
rect 421064 996412 421070 996424
rect 425054 996412 425060 996424
rect 425112 996412 425118 996464
rect 366542 996208 366548 996260
rect 366600 996248 366606 996260
rect 375466 996248 375472 996260
rect 366600 996220 375472 996248
rect 366600 996208 366606 996220
rect 375466 996208 375472 996220
rect 375524 996208 375530 996260
rect 504358 996208 504364 996260
rect 504416 996248 504422 996260
rect 510982 996248 510988 996260
rect 504416 996220 510988 996248
rect 504416 996208 504422 996220
rect 510982 996208 510988 996220
rect 511040 996208 511046 996260
rect 516042 996208 516048 996260
rect 516100 996248 516106 996260
rect 523678 996248 523684 996260
rect 516100 996220 523684 996248
rect 516100 996208 516106 996220
rect 523678 996208 523684 996220
rect 523736 996208 523742 996260
rect 109494 996072 109500 996124
rect 109552 996112 109558 996124
rect 158714 996112 158720 996124
rect 109552 996084 158720 996112
rect 109552 996072 109558 996084
rect 158714 996072 158720 996084
rect 158772 996072 158778 996124
rect 159358 996072 159364 996124
rect 159416 996112 159422 996124
rect 208394 996112 208400 996124
rect 159416 996084 208400 996112
rect 159416 996072 159422 996084
rect 208394 996072 208400 996084
rect 208452 996072 208458 996124
rect 229738 996072 229744 996124
rect 229796 996112 229802 996124
rect 262214 996112 262220 996124
rect 229796 996084 262220 996112
rect 229796 996072 229802 996084
rect 262214 996072 262220 996084
rect 262272 996072 262278 996124
rect 262858 996072 262864 996124
rect 262916 996112 262922 996124
rect 313274 996112 313280 996124
rect 262916 996084 313280 996112
rect 262916 996072 262922 996084
rect 313274 996072 313280 996084
rect 313332 996072 313338 996124
rect 364978 996072 364984 996124
rect 365036 996112 365042 996124
rect 432230 996112 432236 996124
rect 365036 996084 432236 996112
rect 365036 996072 365042 996084
rect 432230 996072 432236 996084
rect 432288 996072 432294 996124
rect 471238 996072 471244 996124
rect 471296 996112 471302 996124
rect 507854 996112 507860 996124
rect 471296 996084 507860 996112
rect 471296 996072 471302 996084
rect 507854 996072 507860 996084
rect 507912 996072 507918 996124
rect 509694 996072 509700 996124
rect 509752 996112 509758 996124
rect 560386 996112 560392 996124
rect 509752 996084 560392 996112
rect 509752 996072 509758 996084
rect 560386 996072 560392 996084
rect 560444 996072 560450 996124
rect 572714 996072 572720 996124
rect 572772 996112 572778 996124
rect 625430 996112 625436 996124
rect 572772 996084 625436 996112
rect 572772 996072 572778 996084
rect 625430 996072 625436 996084
rect 625488 996072 625494 996124
rect 126238 995936 126244 995988
rect 126296 995976 126302 995988
rect 160370 995976 160376 995988
rect 126296 995948 160376 995976
rect 126296 995936 126302 995948
rect 160370 995936 160376 995948
rect 160428 995936 160434 995988
rect 162118 995936 162124 995988
rect 162176 995976 162182 995988
rect 210050 995976 210056 995988
rect 162176 995948 210056 995976
rect 162176 995936 162182 995948
rect 210050 995936 210056 995948
rect 210108 995936 210114 995988
rect 213178 995936 213184 995988
rect 213236 995976 213242 995988
rect 261110 995976 261116 995988
rect 213236 995948 261116 995976
rect 213236 995936 213242 995948
rect 261110 995936 261116 995948
rect 261168 995936 261174 995988
rect 264238 995936 264244 995988
rect 264296 995976 264302 995988
rect 281902 995976 281908 995988
rect 264296 995948 281908 995976
rect 264296 995936 264302 995948
rect 281902 995936 281908 995948
rect 281960 995936 281966 995988
rect 298646 995936 298652 995988
rect 298704 995976 298710 995988
rect 314654 995976 314660 995988
rect 298704 995948 314660 995976
rect 298704 995936 298710 995948
rect 314654 995936 314660 995948
rect 314712 995936 314718 995988
rect 365162 995936 365168 995988
rect 365220 995976 365226 995988
rect 432046 995976 432052 995988
rect 365220 995948 432052 995976
rect 365220 995936 365226 995948
rect 432046 995936 432052 995948
rect 432104 995936 432110 995988
rect 434162 995936 434168 995988
rect 434220 995976 434226 995988
rect 510798 995976 510804 995988
rect 434220 995948 510804 995976
rect 434220 995936 434226 995948
rect 510798 995936 510804 995948
rect 510856 995936 510862 995988
rect 511258 995936 511264 995988
rect 511316 995976 511322 995988
rect 563054 995976 563060 995988
rect 511316 995948 563060 995976
rect 511316 995936 511322 995948
rect 563054 995936 563060 995948
rect 563112 995936 563118 995988
rect 284956 995880 292574 995908
rect 124858 995800 124864 995852
rect 124916 995840 124922 995852
rect 160186 995840 160192 995852
rect 124916 995812 160192 995840
rect 124916 995800 124922 995812
rect 160186 995800 160192 995812
rect 160244 995800 160250 995852
rect 175918 995800 175924 995852
rect 175976 995840 175982 995852
rect 211154 995840 211160 995852
rect 175976 995812 211160 995840
rect 175976 995800 175982 995812
rect 211154 995800 211160 995812
rect 211212 995800 211218 995852
rect 228358 995800 228364 995852
rect 228416 995840 228422 995852
rect 263594 995840 263600 995852
rect 228416 995812 263600 995840
rect 228416 995800 228422 995812
rect 263594 995800 263600 995812
rect 263652 995800 263658 995852
rect 278038 995800 278044 995852
rect 278096 995840 278102 995852
rect 284956 995840 284984 995880
rect 278096 995812 284984 995840
rect 292546 995840 292574 995880
rect 316034 995840 316040 995852
rect 292546 995812 316040 995840
rect 278096 995800 278102 995812
rect 316034 995800 316040 995812
rect 316092 995800 316098 995852
rect 366358 995800 366364 995852
rect 366416 995840 366422 995852
rect 433518 995840 433524 995852
rect 366416 995812 433524 995840
rect 366416 995800 366422 995812
rect 433518 995800 433524 995812
rect 433576 995800 433582 995852
rect 433978 995800 433984 995852
rect 434036 995840 434042 995852
rect 504358 995840 504364 995852
rect 434036 995812 504364 995840
rect 434036 995800 434042 995812
rect 504358 995800 504364 995812
rect 504416 995800 504422 995852
rect 510062 995800 510068 995852
rect 510120 995840 510126 995852
rect 554130 995840 554136 995852
rect 510120 995812 554136 995840
rect 510120 995800 510126 995812
rect 554130 995800 554136 995812
rect 554188 995800 554194 995852
rect 618162 995800 618168 995852
rect 618220 995840 618226 995852
rect 625246 995840 625252 995852
rect 618220 995812 625252 995840
rect 618220 995800 618226 995812
rect 625246 995800 625252 995812
rect 625304 995800 625310 995852
rect 143442 995528 143448 995580
rect 143500 995568 143506 995580
rect 146938 995568 146944 995580
rect 143500 995540 146944 995568
rect 143500 995528 143506 995540
rect 146938 995528 146944 995540
rect 146996 995528 147002 995580
rect 195238 995528 195244 995580
rect 195296 995568 195302 995580
rect 204898 995568 204904 995580
rect 195296 995540 204904 995568
rect 195296 995528 195302 995540
rect 204898 995528 204904 995540
rect 204956 995528 204962 995580
rect 298094 995528 298100 995580
rect 298152 995568 298158 995580
rect 310606 995568 310612 995580
rect 298152 995540 310612 995568
rect 298152 995528 298158 995540
rect 310606 995528 310612 995540
rect 310664 995528 310670 995580
rect 324958 995528 324964 995580
rect 325016 995568 325022 995580
rect 364978 995568 364984 995580
rect 325016 995540 364984 995568
rect 325016 995528 325022 995540
rect 364978 995528 364984 995540
rect 365036 995528 365042 995580
rect 375466 995528 375472 995580
rect 375524 995568 375530 995580
rect 375524 995540 379514 995568
rect 375524 995528 375530 995540
rect 111058 995392 111064 995444
rect 111116 995432 111122 995444
rect 144546 995432 144552 995444
rect 111116 995404 144552 995432
rect 111116 995392 111122 995404
rect 144546 995392 144552 995404
rect 144604 995392 144610 995444
rect 152642 995432 152648 995444
rect 145392 995404 152648 995432
rect 89622 995324 89628 995376
rect 89680 995364 89686 995376
rect 92474 995364 92480 995376
rect 89680 995336 92480 995364
rect 89680 995324 89686 995336
rect 92474 995324 92480 995336
rect 92532 995324 92538 995376
rect 142062 995256 142068 995308
rect 142120 995296 142126 995308
rect 145392 995296 145420 995404
rect 152642 995392 152648 995404
rect 152700 995392 152706 995444
rect 211798 995392 211804 995444
rect 211856 995432 211862 995444
rect 260926 995432 260932 995444
rect 211856 995404 260932 995432
rect 211856 995392 211862 995404
rect 260926 995392 260932 995404
rect 260984 995392 260990 995444
rect 281902 995392 281908 995444
rect 281960 995432 281966 995444
rect 298646 995432 298652 995444
rect 281960 995404 292574 995432
rect 281960 995392 281966 995404
rect 194318 995324 194324 995376
rect 194376 995364 194382 995376
rect 195514 995364 195520 995376
rect 194376 995336 195520 995364
rect 194376 995324 194382 995336
rect 195514 995324 195520 995336
rect 195572 995324 195578 995376
rect 292546 995364 292574 995404
rect 295076 995404 298652 995432
rect 294690 995364 294696 995376
rect 292546 995336 294696 995364
rect 294690 995324 294696 995336
rect 294748 995324 294754 995376
rect 142120 995268 145420 995296
rect 142120 995256 142126 995268
rect 146938 995256 146944 995308
rect 146996 995296 147002 995308
rect 152458 995296 152464 995308
rect 146996 995268 152464 995296
rect 146996 995256 147002 995268
rect 152458 995256 152464 995268
rect 152516 995256 152522 995308
rect 242066 995256 242072 995308
rect 242124 995296 242130 995308
rect 246850 995296 246856 995308
rect 242124 995268 246856 995296
rect 242124 995256 242130 995268
rect 246850 995256 246856 995268
rect 246908 995256 246914 995308
rect 280798 995188 280804 995240
rect 280856 995228 280862 995240
rect 295076 995228 295104 995404
rect 298646 995392 298652 995404
rect 298704 995392 298710 995444
rect 295242 995256 295248 995308
rect 295300 995296 295306 995308
rect 298462 995296 298468 995308
rect 295300 995268 298468 995296
rect 295300 995256 295306 995268
rect 298462 995256 298468 995268
rect 298520 995256 298526 995308
rect 379486 995296 379514 995540
rect 383286 995528 383292 995580
rect 383344 995568 383350 995580
rect 385034 995568 385040 995580
rect 383344 995540 385040 995568
rect 383344 995528 383350 995540
rect 385034 995528 385040 995540
rect 385092 995528 385098 995580
rect 440878 995528 440884 995580
rect 440936 995568 440942 995580
rect 472250 995568 472256 995580
rect 440936 995540 472256 995568
rect 440936 995528 440942 995540
rect 472250 995528 472256 995540
rect 472308 995528 472314 995580
rect 472434 995528 472440 995580
rect 472492 995568 472498 995580
rect 473354 995568 473360 995580
rect 472492 995540 473360 995568
rect 472492 995528 472498 995540
rect 473354 995528 473360 995540
rect 473412 995528 473418 995580
rect 524046 995528 524052 995580
rect 524104 995568 524110 995580
rect 524782 995568 524788 995580
rect 524104 995540 524788 995568
rect 524104 995528 524110 995540
rect 524782 995528 524788 995540
rect 524840 995528 524846 995580
rect 625246 995528 625252 995580
rect 625304 995568 625310 995580
rect 625614 995568 625620 995580
rect 625304 995540 625620 995568
rect 625304 995528 625310 995540
rect 625614 995528 625620 995540
rect 625672 995528 625678 995580
rect 625798 995528 625804 995580
rect 625856 995568 625862 995580
rect 626534 995568 626540 995580
rect 625856 995540 626540 995568
rect 625856 995528 625862 995540
rect 626534 995528 626540 995540
rect 626592 995528 626598 995580
rect 381722 995392 381728 995444
rect 381780 995432 381786 995444
rect 388622 995432 388628 995444
rect 381780 995404 388628 995432
rect 381780 995392 381786 995404
rect 388622 995392 388628 995404
rect 388680 995392 388686 995444
rect 432598 995392 432604 995444
rect 432656 995432 432662 995444
rect 506474 995432 506480 995444
rect 432656 995404 506480 995432
rect 432656 995392 432662 995404
rect 506474 995392 506480 995404
rect 506532 995392 506538 995444
rect 523862 995392 523868 995444
rect 523920 995432 523926 995444
rect 525334 995432 525340 995444
rect 523920 995404 525340 995432
rect 523920 995392 523926 995404
rect 525334 995392 525340 995404
rect 525392 995392 525398 995444
rect 529014 995432 529020 995444
rect 525536 995404 529020 995432
rect 400858 995364 400864 995376
rect 389146 995336 400864 995364
rect 389146 995296 389174 995336
rect 400858 995324 400864 995336
rect 400916 995324 400922 995376
rect 379486 995268 389174 995296
rect 523678 995256 523684 995308
rect 523736 995296 523742 995308
rect 525536 995296 525564 995404
rect 529014 995392 529020 995404
rect 529072 995392 529078 995444
rect 560570 995432 560576 995444
rect 538186 995404 560576 995432
rect 523736 995268 525564 995296
rect 523736 995256 523742 995268
rect 305638 995228 305644 995240
rect 280856 995200 295104 995228
rect 302206 995200 305644 995228
rect 280856 995188 280862 995200
rect 77662 995120 77668 995172
rect 77720 995160 77726 995172
rect 97258 995160 97264 995172
rect 77720 995132 97264 995160
rect 77720 995120 77726 995132
rect 97258 995120 97264 995132
rect 97316 995120 97322 995172
rect 137922 995120 137928 995172
rect 137980 995160 137986 995172
rect 144178 995160 144184 995172
rect 137980 995132 144184 995160
rect 137980 995120 137986 995132
rect 144178 995120 144184 995132
rect 144236 995120 144242 995172
rect 242710 995120 242716 995172
rect 242768 995160 242774 995172
rect 253474 995160 253480 995172
rect 242768 995132 253480 995160
rect 242768 995120 242774 995132
rect 253474 995120 253480 995132
rect 253532 995120 253538 995172
rect 296622 995120 296628 995172
rect 296680 995160 296686 995172
rect 302206 995160 302234 995200
rect 305638 995188 305644 995200
rect 305696 995188 305702 995240
rect 489730 995188 489736 995240
rect 489788 995228 489794 995240
rect 489788 995200 489914 995228
rect 489788 995188 489794 995200
rect 296680 995132 302234 995160
rect 296680 995120 296686 995132
rect 377398 995120 377404 995172
rect 377456 995160 377462 995172
rect 384666 995160 384672 995172
rect 377456 995132 384672 995160
rect 377456 995120 377462 995132
rect 384666 995120 384672 995132
rect 384724 995120 384730 995172
rect 294690 995052 294696 995104
rect 294748 995092 294754 995104
rect 296438 995092 296444 995104
rect 294748 995064 296444 995092
rect 294748 995052 294754 995064
rect 296438 995052 296444 995064
rect 296496 995052 296502 995104
rect 77018 994984 77024 995036
rect 77076 995024 77082 995036
rect 102778 995024 102784 995036
rect 77076 994996 102784 995024
rect 77076 994984 77082 994996
rect 102778 994984 102784 994996
rect 102836 994984 102842 995036
rect 181438 994984 181444 995036
rect 181496 995024 181502 995036
rect 207014 995024 207020 995036
rect 181496 994996 207020 995024
rect 181496 994984 181502 994996
rect 207014 994984 207020 994996
rect 207072 994984 207078 995036
rect 232866 994984 232872 995036
rect 232924 995024 232930 995036
rect 258074 995024 258080 995036
rect 232924 994996 258080 995024
rect 232924 994984 232930 994996
rect 258074 994984 258080 994996
rect 258132 994984 258138 995036
rect 358722 994984 358728 995036
rect 358780 995024 358786 995036
rect 398834 995024 398840 995036
rect 358780 994996 398840 995024
rect 358780 994984 358786 994996
rect 398834 994984 398840 994996
rect 398892 994984 398898 995036
rect 129734 994916 129740 994968
rect 129792 994956 129798 994968
rect 155954 994956 155960 994968
rect 129792 994928 155960 994956
rect 129792 994916 129798 994928
rect 155954 994916 155960 994928
rect 156012 994916 156018 994968
rect 282822 994916 282828 994968
rect 282880 994956 282886 994968
rect 311894 994956 311900 994968
rect 282880 994928 311900 994956
rect 282880 994916 282886 994928
rect 311894 994916 311900 994928
rect 311952 994916 311958 994968
rect 422938 994916 422944 994968
rect 422996 994956 423002 994968
rect 489886 994956 489914 995200
rect 522298 995120 522304 995172
rect 522356 995160 522362 995172
rect 538186 995160 538214 995404
rect 560570 995392 560576 995404
rect 560628 995392 560634 995444
rect 622394 995392 622400 995444
rect 622452 995432 622458 995444
rect 622452 995404 640334 995432
rect 622452 995392 622458 995404
rect 640306 995364 640334 995404
rect 640702 995364 640708 995376
rect 640306 995336 640708 995364
rect 640702 995324 640708 995336
rect 640760 995324 640766 995376
rect 571978 995256 571984 995308
rect 572036 995296 572042 995308
rect 625246 995296 625252 995308
rect 572036 995268 625252 995296
rect 572036 995256 572042 995268
rect 625246 995256 625252 995268
rect 625304 995256 625310 995308
rect 625430 995256 625436 995308
rect 625488 995296 625494 995308
rect 631502 995296 631508 995308
rect 625488 995268 631508 995296
rect 625488 995256 625494 995268
rect 631502 995256 631508 995268
rect 631560 995256 631566 995308
rect 522356 995132 538214 995160
rect 522356 995120 522362 995132
rect 569862 995120 569868 995172
rect 569920 995160 569926 995172
rect 569920 995132 629800 995160
rect 569920 995120 569926 995132
rect 629772 995092 629800 995132
rect 630122 995120 630128 995172
rect 630180 995160 630186 995172
rect 633986 995160 633992 995172
rect 630180 995132 633992 995160
rect 630180 995120 630186 995132
rect 633986 995120 633992 995132
rect 634044 995120 634050 995172
rect 629772 995064 629984 995092
rect 499482 994984 499488 995036
rect 499540 995024 499546 995036
rect 530026 995024 530032 995036
rect 499540 994996 530032 995024
rect 499540 994984 499546 994996
rect 530026 994984 530032 994996
rect 530084 994984 530090 995036
rect 555142 994984 555148 995036
rect 555200 995024 555206 995036
rect 625108 995024 625114 995036
rect 555200 994996 625114 995024
rect 555200 994984 555206 994996
rect 625108 994984 625114 994996
rect 625166 994984 625172 995036
rect 625246 994984 625252 995036
rect 625304 995024 625310 995036
rect 629570 995024 629576 995036
rect 625304 994996 629576 995024
rect 625304 994984 625310 994996
rect 629570 994984 629576 994996
rect 629628 994984 629634 995036
rect 629956 995024 629984 995064
rect 635182 995024 635188 995036
rect 629956 994996 635188 995024
rect 635182 994984 635188 994996
rect 635240 994984 635246 995036
rect 422996 994928 489914 994956
rect 422996 994916 423002 994928
rect 78306 994848 78312 994900
rect 78364 994888 78370 994900
rect 101398 994888 101404 994900
rect 78364 994860 101404 994888
rect 78364 994848 78370 994860
rect 101398 994848 101404 994860
rect 101456 994848 101462 994900
rect 180150 994848 180156 994900
rect 180208 994888 180214 994900
rect 209866 994888 209872 994900
rect 180208 994860 209872 994888
rect 180208 994848 180214 994860
rect 209866 994848 209872 994860
rect 209924 994848 209930 994900
rect 232222 994848 232228 994900
rect 232280 994888 232286 994900
rect 242894 994888 242900 994900
rect 232280 994860 242900 994888
rect 232280 994848 232286 994860
rect 242894 994848 242900 994860
rect 242952 994848 242958 994900
rect 244550 994848 244556 994900
rect 244608 994888 244614 994900
rect 259454 994888 259460 994900
rect 244608 994860 259460 994888
rect 244608 994848 244614 994860
rect 259454 994848 259460 994860
rect 259512 994848 259518 994900
rect 372706 994848 372712 994900
rect 372764 994888 372770 994900
rect 396994 994888 397000 994900
rect 372764 994860 397000 994888
rect 372764 994848 372770 994860
rect 396994 994848 397000 994860
rect 397052 994848 397058 994900
rect 502978 994848 502984 994900
rect 503036 994888 503042 994900
rect 538030 994888 538036 994900
rect 503036 994860 538036 994888
rect 503036 994848 503042 994860
rect 538030 994848 538036 994860
rect 538088 994848 538094 994900
rect 573358 994848 573364 994900
rect 573416 994888 573422 994900
rect 639506 994888 639512 994900
rect 573416 994860 639512 994888
rect 573416 994848 573422 994860
rect 639506 994848 639512 994860
rect 639564 994848 639570 994900
rect 128446 994780 128452 994832
rect 128504 994820 128510 994832
rect 154574 994820 154580 994832
rect 128504 994792 154580 994820
rect 128504 994780 128510 994792
rect 154574 994780 154580 994792
rect 154632 994780 154638 994832
rect 284110 994780 284116 994832
rect 284168 994820 284174 994832
rect 298094 994820 298100 994832
rect 284168 994792 298100 994820
rect 284168 994780 284174 994792
rect 298094 994780 298100 994792
rect 298152 994780 298158 994832
rect 448514 994780 448520 994832
rect 448572 994820 448578 994832
rect 448572 994792 484348 994820
rect 448572 994780 448578 994792
rect 81342 994712 81348 994764
rect 81400 994752 81406 994764
rect 98638 994752 98644 994764
rect 81400 994724 98644 994752
rect 81400 994712 81406 994724
rect 98638 994712 98644 994724
rect 98696 994712 98702 994764
rect 180610 994712 180616 994764
rect 180668 994752 180674 994764
rect 202138 994752 202144 994764
rect 180668 994724 202144 994752
rect 180668 994712 180674 994724
rect 202138 994712 202144 994724
rect 202196 994712 202202 994764
rect 235902 994712 235908 994764
rect 235960 994752 235966 994764
rect 242710 994752 242716 994764
rect 235960 994724 242716 994752
rect 235960 994712 235966 994724
rect 242710 994712 242716 994724
rect 242768 994712 242774 994764
rect 243078 994712 243084 994764
rect 243136 994752 243142 994764
rect 255958 994752 255964 994764
rect 243136 994724 255964 994752
rect 243136 994712 243142 994724
rect 255958 994712 255964 994724
rect 256016 994712 256022 994764
rect 356698 994712 356704 994764
rect 356756 994752 356762 994764
rect 378594 994752 378600 994764
rect 356756 994724 378600 994752
rect 356756 994712 356762 994724
rect 378594 994712 378600 994724
rect 378652 994712 378658 994764
rect 393958 994752 393964 994764
rect 378796 994724 393964 994752
rect 129090 994644 129096 994696
rect 129148 994684 129154 994696
rect 151078 994684 151084 994696
rect 129148 994656 151084 994684
rect 129148 994644 129154 994656
rect 151078 994644 151084 994656
rect 151136 994644 151142 994696
rect 285950 994644 285956 994696
rect 286008 994684 286014 994696
rect 308398 994684 308404 994696
rect 286008 994656 308404 994684
rect 286008 994644 286014 994656
rect 308398 994644 308404 994656
rect 308456 994644 308462 994696
rect 90266 994576 90272 994628
rect 90324 994616 90330 994628
rect 93302 994616 93308 994628
rect 90324 994588 93308 994616
rect 90324 994576 90330 994588
rect 93302 994576 93308 994588
rect 93360 994576 93366 994628
rect 195974 994616 195980 994628
rect 180766 994588 195980 994616
rect 135898 994508 135904 994560
rect 135956 994548 135962 994560
rect 142062 994548 142068 994560
rect 135956 994520 142068 994548
rect 135956 994508 135962 994520
rect 142062 994508 142068 994520
rect 142120 994508 142126 994560
rect 180610 994440 180616 994492
rect 180668 994480 180674 994492
rect 180766 994480 180794 994588
rect 195974 994576 195980 994588
rect 196032 994576 196038 994628
rect 231578 994576 231584 994628
rect 231636 994616 231642 994628
rect 231636 994588 243584 994616
rect 231636 994576 231642 994588
rect 180668 994452 180794 994480
rect 180668 994440 180674 994452
rect 183278 994440 183284 994492
rect 183336 994480 183342 994492
rect 195238 994480 195244 994492
rect 183336 994452 195244 994480
rect 183336 994440 183342 994452
rect 195238 994440 195244 994452
rect 195296 994440 195302 994492
rect 234522 994440 234528 994492
rect 234580 994480 234586 994492
rect 243354 994480 243360 994492
rect 234580 994452 243360 994480
rect 234580 994440 234586 994452
rect 243354 994440 243360 994452
rect 243412 994440 243418 994492
rect 243556 994480 243584 994588
rect 243722 994576 243728 994628
rect 243780 994616 243786 994628
rect 253106 994616 253112 994628
rect 243780 994588 253112 994616
rect 243780 994576 243786 994588
rect 253106 994576 253112 994588
rect 253164 994576 253170 994628
rect 372890 994576 372896 994628
rect 372948 994616 372954 994628
rect 378796 994616 378824 994724
rect 393958 994712 393964 994724
rect 394016 994712 394022 994764
rect 459554 994644 459560 994696
rect 459612 994684 459618 994696
rect 484118 994684 484124 994696
rect 459612 994656 484124 994684
rect 459612 994644 459618 994656
rect 484118 994644 484124 994656
rect 484176 994644 484182 994696
rect 484320 994684 484348 994792
rect 486602 994780 486608 994832
rect 486660 994820 486666 994832
rect 489730 994820 489736 994832
rect 486660 994792 489736 994820
rect 486660 994780 486666 994792
rect 489730 994780 489736 994792
rect 489788 994780 489794 994832
rect 505738 994712 505744 994764
rect 505796 994752 505802 994764
rect 533982 994752 533988 994764
rect 505796 994724 533988 994752
rect 505796 994712 505802 994724
rect 533982 994712 533988 994724
rect 534040 994712 534046 994764
rect 539226 994752 539232 994764
rect 538186 994724 539232 994752
rect 487798 994684 487804 994696
rect 484320 994656 487804 994684
rect 487798 994644 487804 994656
rect 487856 994644 487862 994696
rect 397638 994616 397644 994628
rect 372948 994588 378824 994616
rect 379486 994588 397644 994616
rect 372948 994576 372954 994588
rect 283466 994508 283472 994560
rect 283524 994548 283530 994560
rect 296622 994548 296628 994560
rect 283524 994520 296628 994548
rect 283524 994508 283530 994520
rect 296622 994508 296628 994520
rect 296680 994508 296686 994560
rect 257338 994480 257344 994492
rect 243556 994452 257344 994480
rect 257338 994440 257344 994452
rect 257396 994440 257402 994492
rect 378594 994440 378600 994492
rect 378652 994480 378658 994492
rect 379486 994480 379514 994588
rect 397638 994576 397644 994588
rect 397696 994576 397702 994628
rect 504542 994576 504548 994628
rect 504600 994616 504606 994628
rect 538186 994616 538214 994724
rect 539226 994712 539232 994724
rect 539284 994712 539290 994764
rect 569218 994712 569224 994764
rect 569276 994752 569282 994764
rect 639046 994752 639052 994764
rect 569276 994724 639052 994752
rect 569276 994712 569282 994724
rect 639046 994712 639052 994724
rect 639104 994712 639110 994764
rect 504600 994588 538214 994616
rect 504600 994576 504606 994588
rect 625154 994576 625160 994628
rect 625212 994616 625218 994628
rect 630858 994616 630864 994628
rect 625212 994588 630864 994616
rect 625212 994576 625218 994588
rect 630858 994576 630864 994588
rect 630916 994576 630922 994628
rect 468754 994508 468760 994560
rect 468812 994548 468818 994560
rect 482922 994548 482928 994560
rect 468812 994520 482928 994548
rect 468812 994508 468818 994520
rect 482922 994508 482928 994520
rect 482980 994508 482986 994560
rect 565078 994508 565084 994560
rect 565136 994548 565142 994560
rect 592034 994548 592040 994560
rect 565136 994520 592040 994548
rect 565136 994508 565142 994520
rect 592034 994508 592040 994520
rect 592092 994508 592098 994560
rect 378652 994452 379514 994480
rect 378652 994440 378658 994452
rect 132126 994372 132132 994424
rect 132184 994412 132190 994424
rect 143442 994412 143448 994424
rect 132184 994384 143448 994412
rect 132184 994372 132190 994384
rect 143442 994372 143448 994384
rect 143500 994372 143506 994424
rect 472250 994372 472256 994424
rect 472308 994412 472314 994424
rect 485958 994412 485964 994424
rect 472308 994384 485964 994412
rect 472308 994372 472314 994384
rect 485958 994372 485964 994384
rect 486016 994372 486022 994424
rect 549162 994372 549168 994424
rect 549220 994412 549226 994424
rect 667934 994412 667940 994424
rect 549220 994384 667940 994412
rect 549220 994372 549226 994384
rect 667934 994372 667940 994384
rect 667992 994372 667998 994424
rect 235258 994304 235264 994356
rect 235316 994344 235322 994356
rect 243722 994344 243728 994356
rect 235316 994316 243728 994344
rect 235316 994304 235322 994316
rect 243722 994304 243728 994316
rect 243780 994304 243786 994356
rect 88702 994236 88708 994288
rect 88760 994276 88766 994288
rect 121730 994276 121736 994288
rect 88760 994248 121736 994276
rect 88760 994236 88766 994248
rect 121730 994236 121736 994248
rect 121788 994236 121794 994288
rect 140130 994236 140136 994288
rect 140188 994276 140194 994288
rect 186498 994276 186504 994288
rect 140188 994248 186504 994276
rect 140188 994236 140194 994248
rect 186498 994236 186504 994248
rect 186556 994236 186562 994288
rect 207750 994236 207756 994288
rect 207808 994276 207814 994288
rect 213914 994276 213920 994288
rect 207808 994248 213920 994276
rect 207808 994236 207814 994248
rect 213914 994236 213920 994248
rect 213972 994236 213978 994288
rect 294874 994236 294880 994288
rect 294932 994276 294938 994288
rect 381170 994276 381176 994288
rect 294932 994248 381176 994276
rect 294932 994236 294938 994248
rect 381170 994236 381176 994248
rect 381228 994236 381234 994288
rect 425054 994236 425060 994288
rect 425112 994276 425118 994288
rect 446122 994276 446128 994288
rect 425112 994248 446128 994276
rect 425112 994236 425118 994248
rect 446122 994236 446128 994248
rect 446180 994236 446186 994288
rect 547782 994236 547788 994288
rect 547840 994276 547846 994288
rect 666554 994276 666560 994288
rect 547840 994248 666560 994276
rect 547840 994236 547846 994248
rect 666554 994236 666560 994248
rect 666612 994236 666618 994288
rect 243354 994168 243360 994220
rect 243412 994208 243418 994220
rect 244550 994208 244556 994220
rect 243412 994180 244556 994208
rect 243412 994168 243418 994180
rect 244550 994168 244556 994180
rect 244608 994168 244614 994220
rect 265618 994100 265624 994152
rect 265676 994140 265682 994152
rect 267734 994140 267740 994152
rect 265676 994112 267740 994140
rect 265676 994100 265682 994112
rect 267734 994100 267740 994112
rect 267792 994100 267798 994152
rect 568482 994100 568488 994152
rect 568540 994140 568546 994152
rect 635826 994140 635832 994152
rect 568540 994112 635832 994140
rect 568540 994100 568546 994112
rect 635826 994100 635832 994112
rect 635884 994100 635890 994152
rect 496722 993284 496728 993336
rect 496780 993324 496786 993336
rect 666738 993324 666744 993336
rect 496780 993296 666744 993324
rect 496780 993284 496786 993296
rect 666738 993284 666744 993296
rect 666796 993284 666802 993336
rect 351822 993148 351828 993200
rect 351880 993188 351886 993200
rect 667382 993188 667388 993200
rect 351880 993160 667388 993188
rect 351880 993148 351886 993160
rect 667382 993148 667388 993160
rect 667440 993148 667446 993200
rect 51718 993012 51724 993064
rect 51776 993052 51782 993064
rect 107930 993052 107936 993064
rect 51776 993024 107936 993052
rect 51776 993012 51782 993024
rect 107930 993012 107936 993024
rect 107988 993012 107994 993064
rect 148962 993012 148968 993064
rect 149020 993052 149026 993064
rect 652754 993052 652760 993064
rect 149020 993024 652760 993052
rect 149020 993012 149026 993024
rect 652754 993012 652760 993024
rect 652812 993012 652818 993064
rect 46198 992876 46204 992928
rect 46256 992916 46262 992928
rect 107746 992916 107752 992928
rect 46256 992888 107752 992916
rect 46256 992876 46262 992888
rect 107746 992876 107752 992888
rect 107804 992876 107810 992928
rect 147582 992876 147588 992928
rect 147640 992916 147646 992928
rect 652478 992916 652484 992928
rect 147640 992888 652484 992916
rect 147640 992876 147646 992888
rect 652478 992876 652484 992888
rect 652536 992876 652542 992928
rect 512638 991856 512644 991908
rect 512696 991896 512702 991908
rect 527634 991896 527640 991908
rect 512696 991868 527640 991896
rect 512696 991856 512702 991868
rect 527634 991856 527640 991868
rect 527692 991856 527698 991908
rect 563698 991856 563704 991908
rect 563756 991896 563762 991908
rect 576302 991896 576308 991908
rect 563756 991868 576308 991896
rect 563756 991856 563762 991868
rect 576302 991856 576308 991868
rect 576360 991856 576366 991908
rect 266998 991720 267004 991772
rect 267056 991760 267062 991772
rect 284294 991760 284300 991772
rect 267056 991732 284300 991760
rect 267056 991720 267062 991732
rect 284294 991720 284300 991732
rect 284352 991720 284358 991772
rect 367738 991720 367744 991772
rect 367796 991760 367802 991772
rect 415026 991760 415032 991772
rect 367796 991732 415032 991760
rect 367796 991720 367802 991732
rect 415026 991720 415032 991732
rect 415084 991720 415090 991772
rect 419442 991720 419448 991772
rect 419500 991760 419506 991772
rect 666922 991760 666928 991772
rect 419500 991732 666928 991760
rect 419500 991720 419506 991732
rect 666922 991720 666928 991732
rect 666980 991720 666986 991772
rect 73430 991584 73436 991636
rect 73488 991624 73494 991636
rect 112070 991624 112076 991636
rect 73488 991596 112076 991624
rect 73488 991584 73494 991596
rect 112070 991584 112076 991596
rect 112128 991584 112134 991636
rect 198642 991584 198648 991636
rect 198700 991624 198706 991636
rect 650914 991624 650920 991636
rect 198700 991596 650920 991624
rect 198700 991584 198706 991596
rect 650914 991584 650920 991596
rect 650972 991584 650978 991636
rect 50338 991448 50344 991500
rect 50396 991488 50402 991500
rect 110414 991488 110420 991500
rect 50396 991460 110420 991488
rect 50396 991448 50402 991460
rect 110414 991448 110420 991460
rect 110472 991448 110478 991500
rect 138290 991448 138296 991500
rect 138348 991488 138354 991500
rect 162854 991488 162860 991500
rect 138348 991460 162860 991488
rect 138348 991448 138354 991460
rect 162854 991448 162860 991460
rect 162912 991448 162918 991500
rect 200022 991448 200028 991500
rect 200080 991488 200086 991500
rect 651466 991488 651472 991500
rect 200080 991460 651472 991488
rect 200080 991448 200086 991460
rect 651466 991448 651472 991460
rect 651524 991448 651530 991500
rect 562502 990224 562508 990276
rect 562560 990264 562566 990276
rect 672718 990264 672724 990276
rect 562560 990236 672724 990264
rect 562560 990224 562566 990236
rect 672718 990224 672724 990236
rect 672776 990224 672782 990276
rect 48958 990088 48964 990140
rect 49016 990128 49022 990140
rect 109034 990128 109040 990140
rect 49016 990100 109040 990128
rect 49016 990088 49022 990100
rect 109034 990088 109040 990100
rect 109092 990088 109098 990140
rect 249702 990088 249708 990140
rect 249760 990128 249766 990140
rect 650086 990128 650092 990140
rect 249760 990100 650092 990128
rect 249760 990088 249766 990100
rect 650086 990088 650092 990100
rect 650144 990088 650150 990140
rect 422202 988864 422208 988916
rect 422260 988904 422266 988916
rect 668302 988904 668308 988916
rect 422260 988876 668308 988904
rect 422260 988864 422266 988876
rect 668302 988864 668308 988876
rect 668360 988864 668366 988916
rect 250990 988728 250996 988780
rect 251048 988768 251054 988780
rect 650730 988768 650736 988780
rect 251048 988740 650736 988768
rect 251048 988728 251054 988740
rect 650730 988728 650736 988740
rect 650788 988728 650794 988780
rect 562318 987640 562324 987692
rect 562376 987680 562382 987692
rect 658918 987680 658924 987692
rect 562376 987652 658924 987680
rect 562376 987640 562382 987652
rect 658918 987640 658924 987652
rect 658976 987640 658982 987692
rect 354582 987504 354588 987556
rect 354640 987544 354646 987556
rect 668118 987544 668124 987556
rect 354640 987516 668124 987544
rect 354640 987504 354646 987516
rect 668118 987504 668124 987516
rect 668176 987504 668182 987556
rect 96338 987368 96344 987420
rect 96396 987408 96402 987420
rect 651098 987408 651104 987420
rect 96396 987380 651104 987408
rect 96396 987368 96402 987380
rect 651098 987368 651104 987380
rect 651156 987368 651162 987420
rect 203150 986620 203156 986672
rect 203208 986660 203214 986672
rect 207750 986660 207756 986672
rect 203208 986632 207756 986660
rect 203208 986620 203214 986632
rect 207750 986620 207756 986632
rect 207808 986620 207814 986672
rect 217318 986620 217324 986672
rect 217376 986660 217382 986672
rect 219434 986660 219440 986672
rect 217376 986632 219440 986660
rect 217376 986620 217382 986632
rect 219434 986620 219440 986632
rect 219492 986620 219498 986672
rect 566458 986212 566464 986264
rect 566516 986252 566522 986264
rect 608778 986252 608784 986264
rect 566516 986224 608784 986252
rect 566516 986212 566522 986224
rect 608778 986212 608784 986224
rect 608836 986212 608842 986264
rect 370498 986076 370504 986128
rect 370556 986116 370562 986128
rect 397822 986116 397828 986128
rect 370556 986088 397828 986116
rect 370556 986076 370562 986088
rect 397822 986076 397828 986088
rect 397880 986076 397886 986128
rect 465718 986076 465724 986128
rect 465776 986116 465782 986128
rect 495158 986116 495164 986128
rect 465776 986088 495164 986116
rect 465776 986076 465782 986088
rect 495158 986076 495164 986088
rect 495216 986076 495222 986128
rect 515398 986076 515404 986128
rect 515456 986116 515462 986128
rect 543826 986116 543832 986128
rect 515456 986088 543832 986116
rect 515456 986076 515462 986088
rect 543826 986076 543832 986088
rect 543884 986076 543890 986128
rect 559558 986076 559564 986128
rect 559616 986116 559622 986128
rect 559616 986088 567194 986116
rect 559616 986076 559622 986088
rect 89622 985940 89628 985992
rect 89680 985980 89686 985992
rect 106918 985980 106924 985992
rect 89680 985952 106924 985980
rect 89680 985940 89686 985952
rect 106918 985940 106924 985952
rect 106976 985940 106982 985992
rect 215938 985940 215944 985992
rect 215996 985980 216002 985992
rect 235626 985980 235632 985992
rect 215996 985952 235632 985980
rect 215996 985940 216002 985952
rect 235626 985940 235632 985952
rect 235684 985940 235690 985992
rect 279418 985940 279424 985992
rect 279476 985980 279482 985992
rect 300486 985980 300492 985992
rect 279476 985952 300492 985980
rect 279476 985940 279482 985952
rect 300486 985940 300492 985952
rect 300544 985940 300550 985992
rect 369118 985940 369124 985992
rect 369176 985980 369182 985992
rect 414106 985980 414112 985992
rect 369176 985952 414112 985980
rect 369176 985940 369182 985952
rect 414106 985940 414112 985952
rect 414164 985940 414170 985992
rect 415026 985940 415032 985992
rect 415084 985980 415090 985992
rect 430298 985980 430304 985992
rect 415084 985952 430304 985980
rect 415084 985940 415090 985952
rect 430298 985940 430304 985952
rect 430356 985940 430362 985992
rect 436738 985940 436744 985992
rect 436796 985980 436802 985992
rect 478966 985980 478972 985992
rect 436796 985952 478972 985980
rect 436796 985940 436802 985952
rect 478966 985940 478972 985952
rect 479024 985940 479030 985992
rect 514018 985940 514024 985992
rect 514076 985980 514082 985992
rect 560110 985980 560116 985992
rect 514076 985952 560116 985980
rect 514076 985940 514082 985952
rect 560110 985940 560116 985952
rect 560168 985940 560174 985992
rect 567166 985980 567194 986088
rect 570598 986076 570604 986128
rect 570656 986116 570662 986128
rect 624970 986116 624976 986128
rect 570656 986088 624976 986116
rect 570656 986076 570662 986088
rect 624970 986076 624976 986088
rect 625028 986076 625034 986128
rect 669958 985980 669964 985992
rect 567166 985952 669964 985980
rect 669958 985940 669964 985952
rect 670016 985940 670022 985992
rect 560938 985124 560944 985176
rect 560996 985164 561002 985176
rect 671338 985164 671344 985176
rect 560996 985136 671344 985164
rect 560996 985124 561002 985136
rect 671338 985124 671344 985136
rect 671396 985124 671402 985176
rect 498102 984988 498108 985040
rect 498160 985028 498166 985040
rect 667658 985028 667664 985040
rect 498160 985000 667664 985028
rect 498160 984988 498166 985000
rect 667658 984988 667664 985000
rect 667716 984988 667722 985040
rect 331858 984852 331864 984904
rect 331916 984892 331922 984904
rect 664438 984892 664444 984904
rect 331916 984864 664444 984892
rect 331916 984852 331922 984864
rect 664438 984852 664444 984864
rect 664496 984852 664502 984904
rect 332042 984716 332048 984768
rect 332100 984756 332106 984768
rect 665818 984756 665824 984768
rect 332100 984728 665824 984756
rect 332100 984716 332106 984728
rect 665818 984716 665824 984728
rect 665876 984716 665882 984768
rect 96522 984580 96528 984632
rect 96580 984620 96586 984632
rect 651834 984620 651840 984632
rect 96580 984592 651840 984620
rect 96580 984580 96586 984592
rect 651834 984580 651840 984592
rect 651892 984580 651898 984632
rect 55858 975672 55864 975724
rect 55916 975712 55922 975724
rect 62114 975712 62120 975724
rect 55916 975684 62120 975712
rect 55916 975672 55922 975684
rect 62114 975672 62120 975684
rect 62172 975672 62178 975724
rect 651650 975672 651656 975724
rect 651708 975712 651714 975724
rect 661678 975712 661684 975724
rect 651708 975684 661684 975712
rect 651708 975672 651714 975684
rect 661678 975672 661684 975684
rect 661736 975672 661742 975724
rect 42518 969416 42524 969468
rect 42576 969456 42582 969468
rect 55858 969456 55864 969468
rect 42576 969428 55864 969456
rect 42576 969416 42582 969428
rect 55858 969416 55864 969428
rect 55916 969416 55922 969468
rect 42242 966832 42248 966884
rect 42300 966872 42306 966884
rect 42702 966872 42708 966884
rect 42300 966844 42708 966872
rect 42300 966832 42306 966844
rect 42702 966832 42708 966844
rect 42760 966832 42766 966884
rect 673270 966288 673276 966340
rect 673328 966328 673334 966340
rect 675110 966328 675116 966340
rect 673328 966300 675116 966328
rect 673328 966288 673334 966300
rect 675110 966288 675116 966300
rect 675168 966288 675174 966340
rect 42426 964656 42432 964708
rect 42484 964696 42490 964708
rect 42886 964696 42892 964708
rect 42484 964668 42892 964696
rect 42484 964656 42490 964668
rect 42886 964656 42892 964668
rect 42944 964656 42950 964708
rect 42426 963840 42432 963892
rect 42484 963880 42490 963892
rect 44174 963880 44180 963892
rect 42484 963852 44180 963880
rect 42484 963840 42490 963852
rect 44174 963840 44180 963852
rect 44232 963840 44238 963892
rect 42426 963432 42432 963484
rect 42484 963472 42490 963484
rect 43070 963472 43076 963484
rect 42484 963444 43076 963472
rect 42484 963432 42490 963444
rect 43070 963432 43076 963444
rect 43128 963432 43134 963484
rect 42426 961868 42432 961920
rect 42484 961908 42490 961920
rect 44450 961908 44456 961920
rect 42484 961880 44456 961908
rect 42484 961868 42490 961880
rect 44450 961868 44456 961880
rect 44508 961868 44514 961920
rect 47578 961868 47584 961920
rect 47636 961908 47642 961920
rect 62114 961908 62120 961920
rect 47636 961880 62120 961908
rect 47636 961868 47642 961880
rect 62114 961868 62120 961880
rect 62172 961868 62178 961920
rect 651650 961868 651656 961920
rect 651708 961908 651714 961920
rect 663058 961908 663064 961920
rect 651708 961880 663064 961908
rect 651708 961868 651714 961880
rect 663058 961868 663064 961880
rect 663116 961868 663122 961920
rect 674282 961868 674288 961920
rect 674340 961908 674346 961920
rect 675110 961908 675116 961920
rect 674340 961880 675116 961908
rect 674340 961868 674346 961880
rect 675110 961868 675116 961880
rect 675168 961868 675174 961920
rect 42426 959080 42432 959132
rect 42484 959120 42490 959132
rect 43254 959120 43260 959132
rect 42484 959092 43260 959120
rect 42484 959080 42490 959092
rect 43254 959080 43260 959092
rect 43312 959080 43318 959132
rect 42426 958264 42432 958316
rect 42484 958304 42490 958316
rect 44634 958304 44640 958316
rect 42484 958276 44640 958304
rect 42484 958264 42490 958276
rect 44634 958264 44640 958276
rect 44692 958264 44698 958316
rect 674098 957856 674104 957908
rect 674156 957896 674162 957908
rect 675110 957896 675116 957908
rect 674156 957868 675116 957896
rect 674156 957856 674162 957868
rect 675110 957856 675116 957868
rect 675168 957856 675174 957908
rect 660298 957720 660304 957772
rect 660356 957760 660362 957772
rect 660356 957732 675340 957760
rect 660356 957720 660362 957732
rect 675312 957364 675340 957732
rect 675294 957312 675300 957364
rect 675352 957312 675358 957364
rect 673086 956360 673092 956412
rect 673144 956400 673150 956412
rect 675110 956400 675116 956412
rect 673144 956372 675116 956400
rect 673144 956360 673150 956372
rect 675110 956360 675116 956372
rect 675168 956360 675174 956412
rect 37918 952212 37924 952264
rect 37976 952252 37982 952264
rect 41690 952252 41696 952264
rect 37976 952224 41696 952252
rect 37976 952212 37982 952224
rect 41690 952212 41696 952224
rect 41748 952212 41754 952264
rect 675846 949424 675852 949476
rect 675904 949464 675910 949476
rect 678238 949464 678244 949476
rect 675904 949436 678244 949464
rect 675904 949424 675910 949436
rect 678238 949424 678244 949436
rect 678296 949424 678302 949476
rect 675938 948744 675944 948796
rect 675996 948784 676002 948796
rect 682378 948784 682384 948796
rect 675996 948756 682384 948784
rect 675996 948744 676002 948756
rect 682378 948744 682384 948756
rect 682436 948744 682442 948796
rect 651650 948064 651656 948116
rect 651708 948104 651714 948116
rect 671522 948104 671528 948116
rect 651708 948076 671528 948104
rect 651708 948064 651714 948076
rect 671522 948064 671528 948076
rect 671580 948064 671586 948116
rect 43530 945956 43536 946008
rect 43588 945996 43594 946008
rect 62114 945996 62120 946008
rect 43588 945968 62120 945996
rect 43588 945956 43594 945968
rect 62114 945956 62120 945968
rect 62172 945956 62178 946008
rect 663058 941808 663064 941860
rect 663116 941848 663122 941860
rect 675478 941848 675484 941860
rect 663116 941820 675484 941848
rect 663116 941808 663122 941820
rect 675478 941808 675484 941820
rect 675536 941808 675542 941860
rect 41230 941468 41236 941520
rect 41288 941508 41294 941520
rect 41690 941508 41696 941520
rect 41288 941480 41696 941508
rect 41288 941468 41294 941480
rect 41690 941468 41696 941480
rect 41748 941468 41754 941520
rect 43438 941332 43444 941384
rect 43496 941372 43502 941384
rect 48958 941372 48964 941384
rect 43496 941344 48964 941372
rect 43496 941332 43502 941344
rect 48958 941332 48964 941344
rect 49016 941332 49022 941384
rect 43622 941196 43628 941248
rect 43680 941236 43686 941248
rect 50338 941236 50344 941248
rect 43680 941208 50344 941236
rect 43680 941196 43686 941208
rect 50338 941196 50344 941208
rect 50396 941196 50402 941248
rect 41230 940380 41236 940432
rect 41288 940420 41294 940432
rect 41598 940420 41604 940432
rect 41288 940392 41604 940420
rect 41288 940380 41294 940392
rect 41598 940380 41604 940392
rect 41656 940380 41662 940432
rect 41230 939972 41236 940024
rect 41288 940012 41294 940024
rect 41690 940012 41696 940024
rect 41288 939984 41696 940012
rect 41288 939972 41294 939984
rect 41690 939972 41696 939984
rect 41748 939972 41754 940024
rect 43438 939768 43444 939820
rect 43496 939808 43502 939820
rect 51718 939808 51724 939820
rect 43496 939780 51724 939808
rect 43496 939768 43502 939780
rect 51718 939768 51724 939780
rect 51776 939768 51782 939820
rect 671522 938680 671528 938732
rect 671580 938720 671586 938732
rect 675294 938720 675300 938732
rect 671580 938692 675300 938720
rect 671580 938680 671586 938692
rect 675294 938680 675300 938692
rect 675352 938680 675358 938732
rect 41230 938544 41236 938596
rect 41288 938584 41294 938596
rect 41414 938584 41420 938596
rect 41288 938556 41420 938584
rect 41288 938544 41294 938556
rect 41414 938544 41420 938556
rect 41472 938544 41478 938596
rect 672718 938544 672724 938596
rect 672776 938584 672782 938596
rect 675478 938584 675484 938596
rect 672776 938556 675484 938584
rect 672776 938544 672782 938556
rect 675478 938544 675484 938556
rect 675536 938544 675542 938596
rect 41046 938408 41052 938460
rect 41104 938448 41110 938460
rect 41414 938448 41420 938460
rect 41104 938420 41420 938448
rect 41104 938408 41110 938420
rect 41414 938408 41420 938420
rect 41472 938408 41478 938460
rect 661678 938408 661684 938460
rect 661736 938448 661742 938460
rect 675478 938448 675484 938460
rect 661736 938420 675484 938448
rect 661736 938408 661742 938420
rect 675478 938408 675484 938420
rect 675536 938408 675542 938460
rect 672718 937524 672724 937576
rect 672776 937564 672782 937576
rect 675478 937564 675484 937576
rect 672776 937536 675484 937564
rect 672776 937524 672782 937536
rect 675478 937524 675484 937536
rect 675536 937524 675542 937576
rect 671338 937320 671344 937372
rect 671396 937360 671402 937372
rect 675478 937360 675484 937372
rect 671396 937332 675484 937360
rect 671396 937320 671402 937332
rect 675478 937320 675484 937332
rect 675536 937320 675542 937372
rect 658918 937184 658924 937236
rect 658976 937224 658982 937236
rect 675294 937224 675300 937236
rect 658976 937196 675300 937224
rect 658976 937184 658982 937196
rect 675294 937184 675300 937196
rect 675352 937184 675358 937236
rect 672534 937048 672540 937100
rect 672592 937088 672598 937100
rect 674926 937088 674932 937100
rect 672592 937060 674932 937088
rect 672592 937048 672598 937060
rect 674926 937048 674932 937060
rect 674984 937048 674990 937100
rect 44634 936980 44640 937032
rect 44692 937020 44698 937032
rect 62114 937020 62120 937032
rect 44692 936992 62120 937020
rect 44692 936980 44698 936992
rect 62114 936980 62120 936992
rect 62172 936980 62178 937032
rect 651650 936980 651656 937032
rect 651708 937020 651714 937032
rect 660298 937020 660304 937032
rect 651708 936992 660304 937020
rect 651708 936980 651714 936992
rect 660298 936980 660304 936992
rect 660356 936980 660362 937032
rect 669958 935892 669964 935944
rect 670016 935932 670022 935944
rect 675478 935932 675484 935944
rect 670016 935904 675484 935932
rect 670016 935892 670022 935904
rect 675478 935892 675484 935904
rect 675536 935892 675542 935944
rect 670970 935756 670976 935808
rect 671028 935796 671034 935808
rect 675478 935796 675484 935808
rect 671028 935768 675484 935796
rect 671028 935756 671034 935768
rect 675478 935756 675484 935768
rect 675536 935756 675542 935808
rect 671798 935620 671804 935672
rect 671856 935660 671862 935672
rect 675294 935660 675300 935672
rect 671856 935632 675300 935660
rect 671856 935620 671862 935632
rect 675294 935620 675300 935632
rect 675352 935620 675358 935672
rect 673270 933036 673276 933088
rect 673328 933076 673334 933088
rect 675478 933076 675484 933088
rect 673328 933048 675484 933076
rect 673328 933036 673334 933048
rect 675478 933036 675484 933048
rect 675536 933036 675542 933088
rect 42978 932900 42984 932952
rect 43036 932940 43042 932952
rect 54478 932940 54484 932952
rect 43036 932912 54484 932940
rect 43036 932900 43042 932912
rect 54478 932900 54484 932912
rect 54536 932900 54542 932952
rect 672902 932900 672908 932952
rect 672960 932940 672966 932952
rect 675294 932940 675300 932952
rect 672960 932912 675300 932940
rect 672960 932900 672966 932912
rect 675294 932900 675300 932912
rect 675352 932900 675358 932952
rect 42794 931540 42800 931592
rect 42852 931580 42858 931592
rect 53098 931580 53104 931592
rect 42852 931552 53104 931580
rect 42852 931540 42858 931552
rect 53098 931540 53104 931552
rect 53156 931540 53162 931592
rect 674098 931404 674104 931456
rect 674156 931444 674162 931456
rect 675478 931444 675484 931456
rect 674156 931416 675484 931444
rect 674156 931404 674162 931416
rect 675478 931404 675484 931416
rect 675536 931404 675542 931456
rect 673086 930112 673092 930164
rect 673144 930152 673150 930164
rect 675478 930152 675484 930164
rect 673144 930124 675484 930152
rect 673144 930112 673150 930124
rect 675478 930112 675484 930124
rect 675536 930112 675542 930164
rect 678238 930044 678244 930096
rect 678296 930084 678302 930096
rect 683114 930084 683120 930096
rect 678296 930056 683120 930084
rect 678296 930044 678302 930056
rect 683114 930044 683120 930056
rect 683172 930044 683178 930096
rect 673270 928752 673276 928804
rect 673328 928792 673334 928804
rect 675478 928792 675484 928804
rect 673328 928764 675484 928792
rect 673328 928752 673334 928764
rect 675478 928752 675484 928764
rect 675536 928752 675542 928804
rect 670602 927392 670608 927444
rect 670660 927432 670666 927444
rect 675478 927432 675484 927444
rect 670660 927404 675484 927432
rect 670660 927392 670666 927404
rect 675478 927392 675484 927404
rect 675536 927392 675542 927444
rect 47578 923244 47584 923296
rect 47636 923284 47642 923296
rect 62114 923284 62120 923296
rect 47636 923256 62120 923284
rect 47636 923244 47642 923256
rect 62114 923244 62120 923256
rect 62172 923244 62178 923296
rect 651650 921816 651656 921868
rect 651708 921856 651714 921868
rect 663058 921856 663064 921868
rect 651708 921828 663064 921856
rect 651708 921816 651714 921828
rect 663058 921816 663064 921828
rect 663116 921816 663122 921868
rect 50338 909440 50344 909492
rect 50396 909480 50402 909492
rect 62114 909480 62120 909492
rect 50396 909452 62120 909480
rect 50396 909440 50402 909452
rect 62114 909440 62120 909452
rect 62172 909440 62178 909492
rect 651650 909440 651656 909492
rect 651708 909480 651714 909492
rect 671338 909480 671344 909492
rect 651708 909452 671344 909480
rect 651708 909440 651714 909452
rect 671338 909440 671344 909452
rect 671396 909440 671402 909492
rect 46198 896996 46204 897048
rect 46256 897036 46262 897048
rect 62114 897036 62120 897048
rect 46256 897008 62120 897036
rect 46256 896996 46262 897008
rect 62114 896996 62120 897008
rect 62172 896996 62178 897048
rect 651650 895636 651656 895688
rect 651708 895676 651714 895688
rect 664622 895676 664628 895688
rect 651708 895648 664628 895676
rect 651708 895636 651714 895648
rect 664622 895636 664628 895648
rect 664680 895636 664686 895688
rect 42426 884688 42432 884740
rect 42484 884728 42490 884740
rect 62114 884728 62120 884740
rect 42484 884700 62120 884728
rect 42484 884688 42490 884700
rect 62114 884688 62120 884700
rect 62172 884688 62178 884740
rect 651650 881832 651656 881884
rect 651708 881872 651714 881884
rect 671522 881872 671528 881884
rect 651708 881844 671528 881872
rect 651708 881832 651714 881844
rect 671522 881832 671528 881844
rect 671580 881832 671586 881884
rect 670418 879044 670424 879096
rect 670476 879084 670482 879096
rect 675294 879084 675300 879096
rect 670476 879056 675300 879084
rect 670476 879044 670482 879056
rect 675294 879044 675300 879056
rect 675352 879044 675358 879096
rect 43438 870816 43444 870868
rect 43496 870856 43502 870868
rect 62114 870856 62120 870868
rect 43496 870828 62120 870856
rect 43496 870816 43502 870828
rect 62114 870816 62120 870828
rect 62172 870816 62178 870868
rect 651650 869388 651656 869440
rect 651708 869428 651714 869440
rect 658918 869428 658924 869440
rect 651708 869400 658924 869428
rect 651708 869388 651714 869400
rect 658918 869388 658924 869400
rect 658976 869388 658982 869440
rect 671522 868980 671528 869032
rect 671580 869020 671586 869032
rect 675018 869020 675024 869032
rect 671580 868992 675024 869020
rect 671580 868980 671586 868992
rect 675018 868980 675024 868992
rect 675076 868980 675082 869032
rect 673822 868028 673828 868080
rect 673880 868068 673886 868080
rect 675110 868068 675116 868080
rect 673880 868040 675116 868068
rect 673880 868028 673886 868040
rect 675110 868028 675116 868040
rect 675168 868028 675174 868080
rect 671154 866668 671160 866720
rect 671212 866708 671218 866720
rect 675110 866708 675116 866720
rect 671212 866680 675116 866708
rect 671212 866668 671218 866680
rect 675110 866668 675116 866680
rect 675168 866668 675174 866720
rect 674834 865376 674840 865428
rect 674892 865416 674898 865428
rect 674892 865388 675340 865416
rect 674892 865376 674898 865388
rect 670050 865240 670056 865292
rect 670108 865280 670114 865292
rect 674834 865280 674840 865292
rect 670108 865252 674840 865280
rect 670108 865240 670114 865252
rect 674834 865240 674840 865252
rect 674892 865240 674898 865292
rect 675312 865088 675340 865388
rect 675294 865036 675300 865088
rect 675352 865036 675358 865088
rect 51902 858372 51908 858424
rect 51960 858412 51966 858424
rect 62114 858412 62120 858424
rect 51960 858384 62120 858412
rect 51960 858372 51966 858384
rect 62114 858372 62120 858384
rect 62172 858372 62178 858424
rect 651650 855584 651656 855636
rect 651708 855624 651714 855636
rect 659102 855624 659108 855636
rect 651708 855596 659108 855624
rect 651708 855584 651714 855596
rect 659102 855584 659108 855596
rect 659160 855584 659166 855636
rect 44818 844568 44824 844620
rect 44876 844608 44882 844620
rect 62114 844608 62120 844620
rect 44876 844580 62120 844608
rect 44876 844568 44882 844580
rect 62114 844568 62120 844580
rect 62172 844568 62178 844620
rect 651650 841780 651656 841832
rect 651708 841820 651714 841832
rect 661862 841820 661868 841832
rect 651708 841792 661868 841820
rect 651708 841780 651714 841792
rect 661862 841780 661868 841792
rect 661920 841780 661926 841832
rect 55858 832124 55864 832176
rect 55916 832164 55922 832176
rect 62114 832164 62120 832176
rect 55916 832136 62120 832164
rect 55916 832124 55922 832136
rect 62114 832124 62120 832136
rect 62172 832124 62178 832176
rect 651650 829404 651656 829456
rect 651708 829444 651714 829456
rect 660298 829444 660304 829456
rect 651708 829416 660304 829444
rect 651708 829404 651714 829416
rect 660298 829404 660304 829416
rect 660356 829404 660362 829456
rect 51718 818320 51724 818372
rect 51776 818360 51782 818372
rect 62114 818360 62120 818372
rect 51776 818332 62120 818360
rect 51776 818320 51782 818332
rect 62114 818320 62120 818332
rect 62172 818320 62178 818372
rect 35802 817096 35808 817148
rect 35860 817136 35866 817148
rect 40678 817136 40684 817148
rect 35860 817108 40684 817136
rect 35860 817096 35866 817108
rect 40678 817096 40684 817108
rect 40736 817096 40742 817148
rect 35618 816960 35624 817012
rect 35676 817000 35682 817012
rect 40218 817000 40224 817012
rect 35676 816972 40224 817000
rect 35676 816960 35682 816972
rect 40218 816960 40224 816972
rect 40276 816960 40282 817012
rect 35802 816212 35808 816264
rect 35860 816252 35866 816264
rect 39574 816252 39580 816264
rect 35860 816224 39580 816252
rect 35860 816212 35866 816224
rect 39574 816212 39580 816224
rect 39632 816212 39638 816264
rect 35618 815940 35624 815992
rect 35676 815980 35682 815992
rect 41690 815980 41696 815992
rect 35676 815952 41696 815980
rect 35676 815940 35682 815952
rect 41690 815940 41696 815952
rect 41748 815940 41754 815992
rect 35802 815804 35808 815856
rect 35860 815844 35866 815856
rect 41598 815844 41604 815856
rect 35860 815816 41604 815844
rect 35860 815804 35866 815816
rect 41598 815804 41604 815816
rect 41656 815804 41662 815856
rect 35434 815600 35440 815652
rect 35492 815640 35498 815652
rect 41690 815640 41696 815652
rect 35492 815612 41696 815640
rect 35492 815600 35498 815612
rect 41690 815600 41696 815612
rect 41748 815600 41754 815652
rect 42058 815600 42064 815652
rect 42116 815640 42122 815652
rect 50338 815640 50344 815652
rect 42116 815612 50344 815640
rect 42116 815600 42122 815612
rect 50338 815600 50344 815612
rect 50396 815600 50402 815652
rect 651650 815600 651656 815652
rect 651708 815640 651714 815652
rect 661678 815640 661684 815652
rect 651708 815612 661684 815640
rect 651708 815600 651714 815612
rect 661678 815600 661684 815612
rect 661736 815600 661742 815652
rect 35802 814580 35808 814632
rect 35860 814620 35866 814632
rect 35860 814580 35894 814620
rect 35866 814552 35894 814580
rect 39758 814552 39764 814564
rect 35866 814524 39764 814552
rect 39758 814512 39764 814524
rect 39816 814512 39822 814564
rect 35802 814376 35808 814428
rect 35860 814416 35866 814428
rect 41690 814416 41696 814428
rect 35860 814388 41696 814416
rect 35860 814376 35866 814388
rect 41690 814376 41696 814388
rect 41748 814376 41754 814428
rect 42058 814376 42064 814428
rect 42116 814416 42122 814428
rect 42886 814416 42892 814428
rect 42116 814388 42892 814416
rect 42116 814376 42122 814388
rect 42886 814376 42892 814388
rect 42944 814376 42950 814428
rect 35618 814240 35624 814292
rect 35676 814280 35682 814292
rect 41690 814280 41696 814292
rect 35676 814252 41696 814280
rect 35676 814240 35682 814252
rect 41690 814240 41696 814252
rect 41748 814240 41754 814292
rect 42058 814240 42064 814292
rect 42116 814280 42122 814292
rect 44174 814280 44180 814292
rect 42116 814252 44180 814280
rect 42116 814240 42122 814252
rect 44174 814240 44180 814252
rect 44232 814240 44238 814292
rect 41046 812948 41052 813000
rect 41104 812988 41110 813000
rect 41414 812988 41420 813000
rect 41104 812960 41420 812988
rect 41104 812948 41110 812960
rect 41414 812948 41420 812960
rect 41472 812948 41478 813000
rect 41322 811724 41328 811776
rect 41380 811764 41386 811776
rect 41690 811764 41696 811776
rect 41380 811736 41696 811764
rect 41380 811724 41386 811736
rect 41690 811724 41696 811736
rect 41748 811724 41754 811776
rect 40770 810704 40776 810756
rect 40828 810744 40834 810756
rect 41690 810744 41696 810756
rect 40828 810716 41696 810744
rect 40828 810704 40834 810716
rect 41690 810704 41696 810716
rect 41748 810704 41754 810756
rect 42058 810568 42064 810620
rect 42116 810608 42122 810620
rect 42610 810608 42616 810620
rect 42116 810580 42616 810608
rect 42116 810568 42122 810580
rect 42610 810568 42616 810580
rect 42668 810568 42674 810620
rect 41322 807304 41328 807356
rect 41380 807344 41386 807356
rect 41690 807344 41696 807356
rect 41380 807316 41696 807344
rect 41380 807304 41386 807316
rect 41690 807304 41696 807316
rect 41748 807304 41754 807356
rect 42058 807304 42064 807356
rect 42116 807344 42122 807356
rect 48958 807344 48964 807356
rect 42116 807316 48964 807344
rect 42116 807304 42122 807316
rect 48958 807304 48964 807316
rect 49016 807304 49022 807356
rect 50338 805944 50344 805996
rect 50396 805984 50402 805996
rect 62114 805984 62120 805996
rect 50396 805956 62120 805984
rect 50396 805944 50402 805956
rect 62114 805944 62120 805956
rect 62172 805944 62178 805996
rect 651650 803224 651656 803276
rect 651708 803264 651714 803276
rect 663242 803264 663248 803276
rect 651708 803236 663248 803264
rect 651708 803224 651714 803236
rect 663242 803224 663248 803236
rect 663300 803224 663306 803276
rect 32398 802544 32404 802596
rect 32456 802584 32462 802596
rect 41690 802584 41696 802596
rect 32456 802556 41696 802584
rect 32456 802544 32462 802556
rect 41690 802544 41696 802556
rect 41748 802544 41754 802596
rect 31662 802272 31668 802324
rect 31720 802312 31726 802324
rect 39758 802312 39764 802324
rect 31720 802284 39764 802312
rect 31720 802272 31726 802284
rect 39758 802272 39764 802284
rect 39816 802272 39822 802324
rect 36538 801592 36544 801644
rect 36596 801632 36602 801644
rect 40310 801632 40316 801644
rect 36596 801604 40316 801632
rect 36596 801592 36602 801604
rect 40310 801592 40316 801604
rect 40368 801592 40374 801644
rect 33778 801048 33784 801100
rect 33836 801088 33842 801100
rect 40586 801088 40592 801100
rect 33836 801060 40592 801088
rect 33836 801048 33842 801060
rect 40586 801048 40592 801060
rect 40644 801048 40650 801100
rect 43622 799008 43628 799060
rect 43680 799048 43686 799060
rect 47578 799048 47584 799060
rect 43680 799020 47584 799048
rect 43680 799008 43686 799020
rect 47578 799008 47584 799020
rect 47636 799008 47642 799060
rect 42518 798328 42524 798380
rect 42576 798328 42582 798380
rect 42242 798124 42248 798176
rect 42300 798164 42306 798176
rect 42536 798164 42564 798328
rect 42300 798136 42564 798164
rect 42300 798124 42306 798136
rect 44634 796328 44640 796340
rect 42260 796300 44640 796328
rect 42260 795660 42288 796300
rect 44634 796288 44640 796300
rect 44692 796288 44698 796340
rect 42242 795608 42248 795660
rect 42300 795608 42306 795660
rect 47762 793568 47768 793620
rect 47820 793608 47826 793620
rect 62114 793608 62120 793620
rect 47820 793580 62120 793608
rect 47820 793568 47826 793580
rect 62114 793568 62120 793580
rect 62172 793568 62178 793620
rect 651650 789352 651656 789404
rect 651708 789392 651714 789404
rect 660482 789392 660488 789404
rect 651708 789364 660488 789392
rect 651708 789352 651714 789364
rect 660482 789352 660488 789364
rect 660540 789352 660546 789404
rect 669774 789352 669780 789404
rect 669832 789392 669838 789404
rect 674926 789392 674932 789404
rect 669832 789364 674932 789392
rect 669832 789352 669838 789364
rect 674926 789352 674932 789364
rect 674984 789352 674990 789404
rect 674926 788672 674932 788724
rect 674984 788672 674990 788724
rect 674944 788236 674972 788672
rect 675294 788236 675300 788248
rect 674944 788208 675300 788236
rect 675294 788196 675300 788208
rect 675352 788196 675358 788248
rect 670786 787992 670792 788044
rect 670844 788032 670850 788044
rect 675110 788032 675116 788044
rect 670844 788004 675116 788032
rect 670844 787992 670850 788004
rect 675110 787992 675116 788004
rect 675168 787992 675174 788044
rect 672166 786632 672172 786684
rect 672224 786672 672230 786684
rect 675110 786672 675116 786684
rect 672224 786644 675116 786672
rect 672224 786632 672230 786644
rect 675110 786632 675116 786644
rect 675168 786632 675174 786684
rect 674466 783844 674472 783896
rect 674524 783884 674530 783896
rect 675202 783884 675208 783896
rect 674524 783856 675208 783884
rect 674524 783844 674530 783856
rect 675202 783844 675208 783856
rect 675260 783844 675266 783896
rect 670234 783708 670240 783760
rect 670292 783748 670298 783760
rect 675386 783748 675392 783760
rect 670292 783720 675392 783748
rect 670292 783708 670298 783720
rect 675386 783708 675392 783720
rect 675444 783708 675450 783760
rect 674006 782620 674012 782672
rect 674064 782660 674070 782672
rect 675202 782660 675208 782672
rect 674064 782632 675208 782660
rect 674064 782620 674070 782632
rect 675202 782620 675208 782632
rect 675260 782620 675266 782672
rect 669038 782484 669044 782536
rect 669096 782524 669102 782536
rect 675294 782524 675300 782536
rect 669096 782496 675300 782524
rect 669096 782484 669102 782496
rect 675294 782484 675300 782496
rect 675352 782484 675358 782536
rect 56226 780036 56232 780088
rect 56284 780076 56290 780088
rect 62114 780076 62120 780088
rect 56284 780048 62120 780076
rect 56284 780036 56290 780048
rect 62114 780036 62120 780048
rect 62172 780036 62178 780088
rect 674282 779152 674288 779204
rect 674340 779192 674346 779204
rect 675294 779192 675300 779204
rect 674340 779164 675300 779192
rect 674340 779152 674346 779164
rect 675294 779152 675300 779164
rect 675352 779152 675358 779204
rect 660298 778948 660304 779000
rect 660356 778988 660362 779000
rect 675110 778988 675116 779000
rect 660356 778960 675116 778988
rect 660356 778948 660362 778960
rect 675110 778948 675116 778960
rect 675168 778948 675174 779000
rect 674098 778336 674104 778388
rect 674156 778376 674162 778388
rect 675294 778376 675300 778388
rect 674156 778348 675300 778376
rect 674156 778336 674162 778348
rect 675294 778336 675300 778348
rect 675352 778336 675358 778388
rect 671522 776976 671528 777028
rect 671580 777016 671586 777028
rect 675294 777016 675300 777028
rect 671580 776988 675300 777016
rect 671580 776976 671586 776988
rect 675294 776976 675300 776988
rect 675352 776976 675358 777028
rect 651650 775548 651656 775600
rect 651708 775588 651714 775600
rect 663426 775588 663432 775600
rect 651708 775560 663432 775588
rect 651708 775548 651714 775560
rect 663426 775548 663432 775560
rect 663484 775548 663490 775600
rect 674926 775412 674932 775464
rect 674984 775452 674990 775464
rect 675294 775452 675300 775464
rect 674984 775424 675300 775452
rect 674984 775412 674990 775424
rect 675294 775412 675300 775424
rect 675352 775412 675358 775464
rect 35802 774324 35808 774376
rect 35860 774364 35866 774376
rect 40034 774364 40040 774376
rect 35860 774336 40040 774364
rect 35860 774324 35866 774336
rect 40034 774324 40040 774336
rect 40092 774324 40098 774376
rect 35526 773372 35532 773424
rect 35584 773412 35590 773424
rect 40862 773412 40868 773424
rect 35584 773384 40868 773412
rect 35584 773372 35590 773384
rect 40862 773372 40868 773384
rect 40920 773372 40926 773424
rect 35802 773276 35808 773288
rect 35636 773248 35808 773276
rect 35636 773004 35664 773248
rect 35802 773236 35808 773248
rect 35860 773236 35866 773288
rect 35802 773100 35808 773152
rect 35860 773140 35866 773152
rect 41690 773140 41696 773152
rect 35860 773112 41696 773140
rect 35860 773100 35866 773112
rect 41690 773100 41696 773112
rect 41748 773100 41754 773152
rect 42058 773100 42064 773152
rect 42116 773140 42122 773152
rect 44450 773140 44456 773152
rect 42116 773112 44456 773140
rect 42116 773100 42122 773112
rect 44450 773100 44456 773112
rect 44508 773100 44514 773152
rect 41690 773004 41696 773016
rect 35636 772976 41696 773004
rect 41690 772964 41696 772976
rect 41748 772964 41754 773016
rect 42058 772964 42064 773016
rect 42116 773004 42122 773016
rect 55858 773004 55864 773016
rect 42116 772976 55864 773004
rect 42116 772964 42122 772976
rect 55858 772964 55864 772976
rect 55916 772964 55922 773016
rect 35342 772828 35348 772880
rect 35400 772868 35406 772880
rect 51902 772868 51908 772880
rect 35400 772840 41736 772868
rect 35400 772828 35406 772840
rect 41708 772744 41736 772840
rect 42076 772840 51908 772868
rect 42076 772744 42104 772840
rect 51902 772828 51908 772840
rect 51960 772828 51966 772880
rect 41690 772692 41696 772744
rect 41748 772692 41754 772744
rect 42058 772692 42064 772744
rect 42116 772692 42122 772744
rect 675846 772080 675852 772132
rect 675904 772120 675910 772132
rect 683206 772120 683212 772132
rect 675904 772092 683212 772120
rect 675904 772080 675910 772092
rect 683206 772080 683212 772092
rect 683264 772080 683270 772132
rect 35894 772012 35900 772064
rect 35952 772052 35958 772064
rect 39758 772052 39764 772064
rect 35952 772024 39764 772052
rect 35952 772012 35958 772024
rect 39758 772012 39764 772024
rect 39816 772012 39822 772064
rect 35526 771876 35532 771928
rect 35584 771916 35590 771928
rect 39850 771916 39856 771928
rect 35584 771888 39856 771916
rect 35584 771876 35590 771888
rect 39850 771876 39856 771888
rect 39908 771876 39914 771928
rect 35710 771604 35716 771656
rect 35768 771644 35774 771656
rect 35768 771616 35894 771644
rect 35768 771604 35774 771616
rect 35866 771588 35894 771616
rect 35866 771548 35900 771588
rect 35894 771536 35900 771548
rect 35952 771536 35958 771588
rect 35342 771400 35348 771452
rect 35400 771440 35406 771452
rect 39114 771440 39120 771452
rect 35400 771412 39120 771440
rect 35400 771400 35406 771412
rect 39114 771400 39120 771412
rect 39172 771400 39178 771452
rect 675846 771264 675852 771316
rect 675904 771304 675910 771316
rect 680998 771304 681004 771316
rect 675904 771276 681004 771304
rect 675904 771264 675910 771276
rect 680998 771264 681004 771276
rect 681056 771264 681062 771316
rect 35802 770448 35808 770500
rect 35860 770488 35866 770500
rect 41414 770488 41420 770500
rect 35860 770460 41420 770488
rect 35860 770448 35866 770460
rect 41414 770448 41420 770460
rect 41472 770448 41478 770500
rect 41690 770284 41696 770296
rect 41386 770256 41696 770284
rect 35618 770176 35624 770228
rect 35676 770216 35682 770228
rect 41386 770216 41414 770256
rect 41690 770244 41696 770256
rect 41748 770244 41754 770296
rect 42058 770244 42064 770296
rect 42116 770284 42122 770296
rect 43254 770284 43260 770296
rect 42116 770256 43260 770284
rect 42116 770244 42122 770256
rect 43254 770244 43260 770256
rect 43312 770244 43318 770296
rect 35676 770188 41414 770216
rect 35676 770176 35682 770188
rect 35434 770040 35440 770092
rect 35492 770080 35498 770092
rect 41690 770080 41696 770092
rect 35492 770052 41696 770080
rect 35492 770040 35498 770052
rect 41690 770040 41696 770052
rect 41748 770040 41754 770092
rect 42058 770040 42064 770092
rect 42116 770080 42122 770092
rect 44542 770080 44548 770092
rect 42116 770052 44548 770080
rect 42116 770040 42122 770052
rect 44542 770040 44548 770052
rect 44600 770040 44606 770092
rect 35802 768952 35808 769004
rect 35860 768992 35866 769004
rect 39850 768992 39856 769004
rect 35860 768964 39856 768992
rect 35860 768952 35866 768964
rect 39850 768952 39856 768964
rect 39908 768952 39914 769004
rect 35526 768816 35532 768868
rect 35584 768856 35590 768868
rect 39298 768856 39304 768868
rect 35584 768828 39304 768856
rect 35584 768816 35590 768828
rect 39298 768816 39304 768828
rect 39356 768816 39362 768868
rect 35342 768680 35348 768732
rect 35400 768720 35406 768732
rect 40034 768720 40040 768732
rect 35400 768692 40040 768720
rect 35400 768680 35406 768692
rect 40034 768680 40040 768692
rect 40092 768680 40098 768732
rect 35802 767320 35808 767372
rect 35860 767360 35866 767372
rect 36538 767360 36544 767372
rect 35860 767332 36544 767360
rect 35860 767320 35866 767332
rect 36538 767320 36544 767332
rect 36596 767320 36602 767372
rect 43622 767320 43628 767372
rect 43680 767360 43686 767372
rect 62114 767360 62120 767372
rect 43680 767332 62120 767360
rect 43680 767320 43686 767332
rect 62114 767320 62120 767332
rect 62172 767320 62178 767372
rect 35802 766300 35808 766352
rect 35860 766340 35866 766352
rect 35860 766300 35894 766340
rect 35866 766204 35894 766300
rect 40402 766204 40408 766216
rect 35866 766176 40408 766204
rect 40402 766164 40408 766176
rect 40460 766164 40466 766216
rect 41690 766000 41696 766012
rect 41386 765972 41696 766000
rect 35802 765892 35808 765944
rect 35860 765932 35866 765944
rect 41386 765932 41414 765972
rect 41690 765960 41696 765972
rect 41748 765960 41754 766012
rect 35860 765904 41414 765932
rect 35860 765892 35866 765904
rect 42058 765892 42064 765944
rect 42116 765932 42122 765944
rect 45002 765932 45008 765944
rect 42116 765904 45008 765932
rect 42116 765892 42122 765904
rect 45002 765892 45008 765904
rect 45060 765892 45066 765944
rect 40034 765348 40040 765400
rect 40092 765388 40098 765400
rect 41690 765388 41696 765400
rect 40092 765360 41696 765388
rect 40092 765348 40098 765360
rect 41690 765348 41696 765360
rect 41748 765348 41754 765400
rect 673638 765280 673644 765332
rect 673696 765320 673702 765332
rect 674098 765320 674104 765332
rect 673696 765292 674104 765320
rect 673696 765280 673702 765292
rect 674098 765280 674104 765292
rect 674156 765280 674162 765332
rect 35802 764668 35808 764720
rect 35860 764708 35866 764720
rect 40402 764708 40408 764720
rect 35860 764680 40408 764708
rect 35860 764668 35866 764680
rect 40402 764668 40408 764680
rect 40460 764668 40466 764720
rect 35802 763648 35808 763700
rect 35860 763688 35866 763700
rect 37918 763688 37924 763700
rect 35860 763660 37924 763688
rect 35860 763648 35866 763660
rect 37918 763648 37924 763660
rect 37976 763648 37982 763700
rect 35618 763240 35624 763292
rect 35676 763280 35682 763292
rect 41506 763280 41512 763292
rect 35676 763252 41512 763280
rect 35676 763240 35682 763252
rect 41506 763240 41512 763252
rect 41564 763240 41570 763292
rect 651650 763240 651656 763292
rect 651708 763280 651714 763292
rect 651708 763252 654134 763280
rect 651708 763240 651714 763252
rect 654106 763212 654134 763252
rect 660298 763212 660304 763224
rect 654106 763184 660304 763212
rect 660298 763172 660304 763184
rect 660356 763172 660362 763224
rect 35802 761880 35808 761932
rect 35860 761920 35866 761932
rect 40494 761920 40500 761932
rect 35860 761892 40500 761920
rect 35860 761880 35866 761892
rect 40494 761880 40500 761892
rect 40552 761880 40558 761932
rect 673822 761880 673828 761932
rect 673880 761880 673886 761932
rect 673840 761796 673868 761880
rect 673822 761744 673828 761796
rect 673880 761744 673886 761796
rect 671338 761540 671344 761592
rect 671396 761580 671402 761592
rect 675478 761580 675484 761592
rect 671396 761552 675484 761580
rect 671396 761540 671402 761552
rect 675478 761540 675484 761552
rect 675536 761540 675542 761592
rect 673638 761404 673644 761456
rect 673696 761444 673702 761456
rect 674006 761444 674012 761456
rect 673696 761416 674012 761444
rect 673696 761404 673702 761416
rect 674006 761404 674012 761416
rect 674064 761404 674070 761456
rect 664622 760520 664628 760572
rect 664680 760560 664686 760572
rect 675478 760560 675484 760572
rect 664680 760532 675484 760560
rect 664680 760520 664686 760532
rect 675478 760520 675484 760532
rect 675536 760520 675542 760572
rect 663058 760384 663064 760436
rect 663116 760424 663122 760436
rect 675294 760424 675300 760436
rect 663116 760396 675300 760424
rect 663116 760384 663122 760396
rect 675294 760384 675300 760396
rect 675352 760384 675358 760436
rect 672534 760248 672540 760300
rect 672592 760288 672598 760300
rect 675478 760288 675484 760300
rect 672592 760260 675484 760288
rect 672592 760248 672598 760260
rect 675478 760248 675484 760260
rect 675536 760248 675542 760300
rect 671982 759840 671988 759892
rect 672040 759880 672046 759892
rect 675478 759880 675484 759892
rect 672040 759852 675484 759880
rect 672040 759840 672046 759852
rect 675478 759840 675484 759852
rect 675536 759840 675542 759892
rect 672718 759500 672724 759552
rect 672776 759540 672782 759552
rect 675478 759540 675484 759552
rect 672776 759512 675484 759540
rect 672776 759500 672782 759512
rect 675478 759500 675484 759512
rect 675536 759500 675542 759552
rect 36538 759024 36544 759076
rect 36596 759064 36602 759076
rect 41414 759064 41420 759076
rect 36596 759036 41420 759064
rect 36596 759024 36602 759036
rect 41414 759024 41420 759036
rect 41472 759024 41478 759076
rect 672626 759024 672632 759076
rect 672684 759064 672690 759076
rect 675478 759064 675484 759076
rect 672684 759036 675484 759064
rect 672684 759024 672690 759036
rect 675478 759024 675484 759036
rect 675536 759024 675542 759076
rect 670970 758684 670976 758736
rect 671028 758724 671034 758736
rect 675478 758724 675484 758736
rect 671028 758696 675484 758724
rect 671028 758684 671034 758696
rect 675478 758684 675484 758696
rect 675536 758684 675542 758736
rect 671798 758344 671804 758396
rect 671856 758384 671862 758396
rect 675294 758384 675300 758396
rect 671856 758356 675300 758384
rect 671856 758344 671862 758356
rect 675294 758344 675300 758356
rect 675352 758344 675358 758396
rect 35158 758276 35164 758328
rect 35216 758316 35222 758328
rect 40402 758316 40408 758328
rect 35216 758288 40408 758316
rect 35216 758276 35222 758288
rect 40402 758276 40408 758288
rect 40460 758276 40466 758328
rect 671798 758208 671804 758260
rect 671856 758248 671862 758260
rect 675478 758248 675484 758260
rect 671856 758220 675484 758248
rect 671856 758208 671862 758220
rect 675478 758208 675484 758220
rect 675536 758208 675542 758260
rect 37918 757732 37924 757784
rect 37976 757772 37982 757784
rect 41690 757772 41696 757784
rect 37976 757744 41696 757772
rect 37976 757732 37982 757744
rect 41690 757732 41696 757744
rect 41748 757732 41754 757784
rect 671338 757392 671344 757444
rect 671396 757432 671402 757444
rect 675478 757432 675484 757444
rect 671396 757404 675484 757432
rect 671396 757392 671402 757404
rect 675478 757392 675484 757404
rect 675536 757392 675542 757444
rect 670050 755012 670056 755064
rect 670108 755052 670114 755064
rect 675478 755052 675484 755064
rect 670108 755024 675484 755052
rect 670108 755012 670114 755024
rect 675478 755012 675484 755024
rect 675536 755012 675542 755064
rect 43806 754876 43812 754928
rect 43864 754916 43870 754928
rect 45002 754916 45008 754928
rect 43864 754888 45008 754916
rect 43864 754876 43870 754888
rect 45002 754876 45008 754888
rect 45060 754876 45066 754928
rect 670418 754604 670424 754656
rect 670476 754644 670482 754656
rect 675478 754644 675484 754656
rect 670476 754616 675484 754644
rect 670476 754604 670482 754616
rect 675478 754604 675484 754616
rect 675536 754604 675542 754656
rect 42426 754468 42432 754520
rect 42484 754508 42490 754520
rect 45186 754508 45192 754520
rect 42484 754480 45192 754508
rect 42484 754468 42490 754480
rect 45186 754468 45192 754480
rect 45244 754468 45250 754520
rect 50522 753516 50528 753568
rect 50580 753556 50586 753568
rect 62114 753556 62120 753568
rect 50580 753528 62120 753556
rect 50580 753516 50586 753528
rect 62114 753516 62120 753528
rect 62172 753516 62178 753568
rect 671154 753380 671160 753432
rect 671212 753420 671218 753432
rect 675478 753420 675484 753432
rect 671212 753392 675484 753420
rect 671212 753380 671218 753392
rect 675478 753380 675484 753392
rect 675536 753380 675542 753432
rect 673822 752972 673828 753024
rect 673880 753012 673886 753024
rect 675478 753012 675484 753024
rect 673880 752984 675484 753012
rect 673880 752972 673886 752984
rect 675478 752972 675484 752984
rect 675536 752972 675542 753024
rect 672994 752088 673000 752140
rect 673052 752128 673058 752140
rect 673362 752128 673368 752140
rect 673052 752100 673368 752128
rect 673052 752088 673058 752100
rect 673362 752088 673368 752100
rect 673420 752088 673426 752140
rect 672350 751748 672356 751800
rect 672408 751788 672414 751800
rect 675478 751788 675484 751800
rect 672408 751760 675484 751788
rect 672408 751748 672414 751760
rect 675478 751748 675484 751760
rect 675536 751748 675542 751800
rect 672350 751272 672356 751324
rect 672408 751312 672414 751324
rect 675478 751312 675484 751324
rect 672408 751284 675484 751312
rect 672408 751272 672414 751284
rect 675478 751272 675484 751284
rect 675536 751272 675542 751324
rect 675846 751068 675852 751120
rect 675904 751108 675910 751120
rect 683114 751108 683120 751120
rect 675904 751080 683120 751108
rect 675904 751068 675910 751080
rect 683114 751068 683120 751080
rect 683172 751068 683178 751120
rect 669958 750048 669964 750100
rect 670016 750088 670022 750100
rect 675478 750088 675484 750100
rect 670016 750060 675484 750088
rect 670016 750048 670022 750060
rect 675478 750048 675484 750060
rect 675536 750048 675542 750100
rect 652018 749368 652024 749420
rect 652076 749408 652082 749420
rect 659286 749408 659292 749420
rect 652076 749380 659292 749408
rect 652076 749368 652082 749380
rect 659286 749368 659292 749380
rect 659344 749368 659350 749420
rect 673730 748824 673736 748876
rect 673788 748864 673794 748876
rect 674098 748864 674104 748876
rect 673788 748836 674104 748864
rect 673788 748824 673794 748836
rect 674098 748824 674104 748836
rect 674156 748824 674162 748876
rect 673914 748688 673920 748740
rect 673972 748728 673978 748740
rect 673972 748700 674144 748728
rect 673972 748688 673978 748700
rect 42242 748552 42248 748604
rect 42300 748592 42306 748604
rect 43254 748592 43260 748604
rect 42300 748564 43260 748592
rect 42300 748552 42306 748564
rect 43254 748552 43260 748564
rect 43312 748552 43318 748604
rect 674116 748400 674144 748700
rect 674098 748348 674104 748400
rect 674156 748348 674162 748400
rect 42242 747124 42248 747176
rect 42300 747124 42306 747176
rect 42260 746904 42288 747124
rect 42242 746852 42248 746904
rect 42300 746852 42306 746904
rect 42242 745288 42248 745340
rect 42300 745288 42306 745340
rect 42260 745136 42288 745288
rect 669590 745220 669596 745272
rect 669648 745260 669654 745272
rect 675294 745260 675300 745272
rect 669648 745232 675300 745260
rect 669648 745220 669654 745232
rect 675294 745220 675300 745232
rect 675352 745220 675358 745272
rect 42242 745084 42248 745136
rect 42300 745084 42306 745136
rect 669222 743792 669228 743844
rect 669280 743832 669286 743844
rect 669590 743832 669596 743844
rect 669280 743804 669596 743832
rect 669280 743792 669286 743804
rect 669590 743792 669596 743804
rect 669648 743792 669654 743844
rect 666094 742432 666100 742484
rect 666152 742472 666158 742484
rect 675294 742472 675300 742484
rect 666152 742444 675300 742472
rect 666152 742432 666158 742444
rect 675294 742432 675300 742444
rect 675352 742432 675358 742484
rect 674834 741616 674840 741668
rect 674892 741656 674898 741668
rect 675478 741656 675484 741668
rect 674892 741628 675484 741656
rect 674892 741616 674898 741628
rect 675478 741616 675484 741628
rect 675536 741616 675542 741668
rect 56042 741072 56048 741124
rect 56100 741112 56106 741124
rect 62114 741112 62120 741124
rect 56100 741084 62120 741112
rect 56100 741072 56106 741084
rect 62114 741072 62120 741084
rect 62172 741072 62178 741124
rect 672994 738420 673000 738472
rect 673052 738460 673058 738472
rect 675110 738460 675116 738472
rect 673052 738432 675116 738460
rect 673052 738420 673058 738432
rect 675110 738420 675116 738432
rect 675168 738420 675174 738472
rect 651650 735564 651656 735616
rect 651708 735604 651714 735616
rect 664622 735604 664628 735616
rect 651708 735576 664628 735604
rect 651708 735564 651714 735576
rect 664622 735564 664628 735576
rect 664680 735564 664686 735616
rect 663426 734816 663432 734868
rect 663484 734856 663490 734868
rect 663484 734828 663794 734856
rect 663484 734816 663490 734828
rect 663766 734788 663794 734828
rect 663766 734760 669314 734788
rect 669286 734720 669314 734760
rect 675294 734748 675300 734800
rect 675352 734748 675358 734800
rect 675018 734720 675024 734732
rect 669286 734692 675024 734720
rect 675018 734680 675024 734692
rect 675076 734680 675082 734732
rect 675312 734596 675340 734748
rect 675294 734544 675300 734596
rect 675352 734544 675358 734596
rect 42426 731144 42432 731196
rect 42484 731184 42490 731196
rect 56226 731184 56232 731196
rect 42484 731156 56232 731184
rect 42484 731144 42490 731156
rect 56226 731144 56232 731156
rect 56284 731144 56290 731196
rect 41138 730056 41144 730108
rect 41196 730096 41202 730108
rect 41690 730096 41696 730108
rect 41196 730068 41696 730096
rect 41196 730056 41202 730068
rect 41690 730056 41696 730068
rect 41748 730056 41754 730108
rect 42058 730056 42064 730108
rect 42116 730096 42122 730108
rect 50338 730096 50344 730108
rect 42116 730068 50344 730096
rect 42116 730056 42122 730068
rect 50338 730056 50344 730068
rect 50396 730056 50402 730108
rect 675202 728968 675208 729020
rect 675260 728968 675266 729020
rect 675018 728764 675024 728816
rect 675076 728804 675082 728816
rect 675220 728804 675248 728968
rect 675076 728776 675248 728804
rect 675076 728764 675082 728776
rect 674374 728356 674380 728408
rect 674432 728396 674438 728408
rect 675478 728396 675484 728408
rect 674432 728368 675484 728396
rect 674432 728356 674438 728368
rect 675478 728356 675484 728368
rect 675536 728356 675542 728408
rect 41690 727648 41696 727660
rect 41386 727620 41696 727648
rect 41046 727540 41052 727592
rect 41104 727580 41110 727592
rect 41386 727580 41414 727620
rect 41690 727608 41696 727620
rect 41748 727608 41754 727660
rect 42058 727608 42064 727660
rect 42116 727648 42122 727660
rect 42886 727648 42892 727660
rect 42116 727620 42892 727648
rect 42116 727608 42122 727620
rect 42886 727608 42892 727620
rect 42944 727608 42950 727660
rect 41104 727552 41414 727580
rect 41104 727540 41110 727552
rect 41690 727512 41696 727524
rect 41524 727484 41696 727512
rect 41322 727404 41328 727456
rect 41380 727444 41386 727456
rect 41524 727444 41552 727484
rect 41690 727472 41696 727484
rect 41748 727472 41754 727524
rect 42058 727472 42064 727524
rect 42116 727512 42122 727524
rect 44266 727512 44272 727524
rect 42116 727484 44272 727512
rect 42116 727472 42122 727484
rect 44266 727472 44272 727484
rect 44324 727472 44330 727524
rect 41380 727416 41552 727444
rect 41380 727404 41386 727416
rect 40862 727268 40868 727320
rect 40920 727308 40926 727320
rect 41690 727308 41696 727320
rect 40920 727280 41696 727308
rect 40920 727268 40926 727280
rect 41690 727268 41696 727280
rect 41748 727268 41754 727320
rect 42058 727268 42064 727320
rect 42116 727308 42122 727320
rect 44542 727308 44548 727320
rect 42116 727280 44548 727308
rect 42116 727268 42122 727280
rect 44542 727268 44548 727280
rect 44600 727268 44606 727320
rect 51902 727268 51908 727320
rect 51960 727308 51966 727320
rect 62114 727308 62120 727320
rect 51960 727280 62120 727308
rect 51960 727268 51966 727280
rect 62114 727268 62120 727280
rect 62172 727268 62178 727320
rect 676030 726792 676036 726844
rect 676088 726832 676094 726844
rect 683114 726832 683120 726844
rect 676088 726804 683120 726832
rect 676088 726792 676094 726804
rect 683114 726792 683120 726804
rect 683172 726792 683178 726844
rect 675846 726520 675852 726572
rect 675904 726560 675910 726572
rect 683482 726560 683488 726572
rect 675904 726532 683488 726560
rect 675904 726520 675910 726532
rect 683482 726520 683488 726532
rect 683540 726520 683546 726572
rect 41322 726180 41328 726232
rect 41380 726220 41386 726232
rect 41690 726220 41696 726232
rect 41380 726192 41696 726220
rect 41380 726180 41386 726192
rect 41690 726180 41696 726192
rect 41748 726180 41754 726232
rect 42058 726180 42064 726232
rect 42116 726220 42122 726232
rect 42518 726220 42524 726232
rect 42116 726192 42524 726220
rect 42116 726180 42122 726192
rect 42518 726180 42524 726192
rect 42576 726180 42582 726232
rect 41138 726044 41144 726096
rect 41196 726084 41202 726096
rect 41598 726084 41604 726096
rect 41196 726056 41604 726084
rect 41196 726044 41202 726056
rect 41598 726044 41604 726056
rect 41656 726044 41662 726096
rect 651650 723120 651656 723172
rect 651708 723160 651714 723172
rect 659470 723160 659476 723172
rect 651708 723132 659476 723160
rect 651708 723120 651714 723132
rect 659470 723120 659476 723132
rect 659528 723120 659534 723172
rect 31754 720264 31760 720316
rect 31812 720304 31818 720316
rect 40034 720304 40040 720316
rect 31812 720276 40040 720304
rect 31812 720264 31818 720276
rect 40034 720264 40040 720276
rect 40092 720264 40098 720316
rect 675846 719652 675852 719704
rect 675904 719692 675910 719704
rect 683298 719692 683304 719704
rect 675904 719664 683304 719692
rect 675904 719652 675910 719664
rect 683298 719652 683304 719664
rect 683356 719652 683362 719704
rect 43438 719108 43444 719160
rect 43496 719148 43502 719160
rect 55858 719148 55864 719160
rect 43496 719120 55864 719148
rect 43496 719108 43502 719120
rect 55858 719108 55864 719120
rect 55916 719108 55922 719160
rect 659102 716252 659108 716304
rect 659160 716292 659166 716304
rect 675478 716292 675484 716304
rect 659160 716264 675484 716292
rect 659160 716252 659166 716264
rect 675478 716252 675484 716264
rect 675536 716252 675542 716304
rect 672626 715816 672632 715828
rect 672368 715788 672632 715816
rect 35158 715640 35164 715692
rect 35216 715680 35222 715692
rect 39206 715680 39212 715692
rect 35216 715652 39212 715680
rect 35216 715640 35222 715652
rect 39206 715640 39212 715652
rect 39264 715640 39270 715692
rect 672368 715624 672396 715788
rect 672626 715776 672632 715788
rect 672684 715776 672690 715828
rect 672350 715572 672356 715624
rect 672408 715572 672414 715624
rect 37918 715368 37924 715420
rect 37976 715408 37982 715420
rect 41506 715408 41512 715420
rect 37976 715380 41512 715408
rect 37976 715368 37982 715380
rect 41506 715368 41512 715380
rect 41564 715368 41570 715420
rect 671982 715300 671988 715352
rect 672040 715340 672046 715352
rect 674834 715340 674840 715352
rect 672040 715312 674840 715340
rect 672040 715300 672046 715312
rect 674834 715300 674840 715312
rect 674892 715300 674898 715352
rect 33778 715232 33784 715284
rect 33836 715272 33842 715284
rect 41690 715272 41696 715284
rect 33836 715244 41696 715272
rect 33836 715232 33842 715244
rect 41690 715232 41696 715244
rect 41748 715232 41754 715284
rect 661862 715096 661868 715148
rect 661920 715136 661926 715148
rect 675478 715136 675484 715148
rect 661920 715108 675484 715136
rect 661920 715096 661926 715108
rect 675478 715096 675484 715108
rect 675536 715096 675542 715148
rect 670970 714960 670976 715012
rect 671028 715000 671034 715012
rect 671028 714972 675524 715000
rect 671028 714960 671034 714972
rect 675496 714876 675524 714972
rect 50706 714824 50712 714876
rect 50764 714864 50770 714876
rect 62114 714864 62120 714876
rect 50764 714836 62120 714864
rect 50764 714824 50770 714836
rect 62114 714824 62120 714836
rect 62172 714824 62178 714876
rect 658918 714824 658924 714876
rect 658976 714864 658982 714876
rect 675294 714864 675300 714876
rect 658976 714836 675300 714864
rect 658976 714824 658982 714836
rect 675294 714824 675300 714836
rect 675352 714824 675358 714876
rect 675478 714824 675484 714876
rect 675536 714824 675542 714876
rect 672350 714484 672356 714536
rect 672408 714524 672414 714536
rect 675478 714524 675484 714536
rect 672408 714496 675484 714524
rect 672408 714484 672414 714496
rect 675478 714484 675484 714496
rect 675536 714484 675542 714536
rect 40678 714212 40684 714264
rect 40736 714252 40742 714264
rect 41690 714252 41696 714264
rect 40736 714224 41696 714252
rect 40736 714212 40742 714224
rect 41690 714212 41696 714224
rect 41748 714212 41754 714264
rect 42058 714212 42064 714264
rect 42116 714252 42122 714264
rect 42702 714252 42708 714264
rect 42116 714224 42708 714252
rect 42116 714212 42122 714224
rect 42702 714212 42708 714224
rect 42760 714212 42766 714264
rect 671154 714008 671160 714060
rect 671212 714048 671218 714060
rect 675478 714048 675484 714060
rect 671212 714020 675484 714048
rect 671212 714008 671218 714020
rect 675478 714008 675484 714020
rect 675536 714008 675542 714060
rect 671798 713668 671804 713720
rect 671856 713708 671862 713720
rect 675478 713708 675484 713720
rect 671856 713680 675484 713708
rect 671856 713668 671862 713680
rect 675478 713668 675484 713680
rect 675536 713668 675542 713720
rect 676030 713396 676036 713448
rect 676088 713436 676094 713448
rect 677686 713436 677692 713448
rect 676088 713408 677692 713436
rect 676088 713396 676094 713408
rect 677686 713396 677692 713408
rect 677744 713396 677750 713448
rect 671890 713192 671896 713244
rect 671948 713232 671954 713244
rect 675478 713232 675484 713244
rect 671948 713204 675484 713232
rect 671948 713192 671954 713204
rect 675478 713192 675484 713204
rect 675536 713192 675542 713244
rect 671522 712852 671528 712904
rect 671580 712892 671586 712904
rect 675478 712892 675484 712904
rect 671580 712864 675484 712892
rect 671580 712852 671586 712864
rect 675478 712852 675484 712864
rect 675536 712852 675542 712904
rect 671706 712376 671712 712428
rect 671764 712416 671770 712428
rect 675478 712416 675484 712428
rect 671764 712388 675484 712416
rect 671764 712376 671770 712388
rect 675478 712376 675484 712388
rect 675536 712376 675542 712428
rect 51718 712280 51724 712292
rect 51046 712252 51724 712280
rect 51046 712144 51074 712252
rect 51718 712240 51724 712252
rect 51776 712240 51782 712292
rect 42260 712116 51074 712144
rect 42260 711136 42288 712116
rect 672166 712036 672172 712088
rect 672224 712076 672230 712088
rect 675478 712076 675484 712088
rect 672224 712048 675484 712076
rect 672224 712036 672230 712048
rect 675478 712036 675484 712048
rect 675536 712036 675542 712088
rect 670786 711220 670792 711272
rect 670844 711260 670850 711272
rect 675478 711260 675484 711272
rect 670844 711232 675484 711260
rect 670844 711220 670850 711232
rect 675478 711220 675484 711232
rect 675536 711220 675542 711272
rect 42242 711084 42248 711136
rect 42300 711084 42306 711136
rect 673086 709996 673092 710048
rect 673144 710036 673150 710048
rect 675294 710036 675300 710048
rect 673144 710008 675300 710036
rect 673144 709996 673150 710008
rect 675294 709996 675300 710008
rect 675352 709996 675358 710048
rect 669038 709724 669044 709776
rect 669096 709764 669102 709776
rect 675478 709764 675484 709776
rect 669096 709736 675484 709764
rect 669096 709724 669102 709736
rect 675478 709724 675484 709736
rect 675536 709724 675542 709776
rect 669774 709588 669780 709640
rect 669832 709628 669838 709640
rect 675478 709628 675484 709640
rect 669832 709600 675484 709628
rect 669832 709588 669838 709600
rect 675478 709588 675484 709600
rect 675536 709588 675542 709640
rect 651650 709316 651656 709368
rect 651708 709356 651714 709368
rect 663058 709356 663064 709368
rect 651708 709328 663064 709356
rect 651708 709316 651714 709328
rect 663058 709316 663064 709328
rect 663116 709316 663122 709368
rect 670234 708772 670240 708824
rect 670292 708812 670298 708824
rect 675478 708812 675484 708824
rect 670292 708784 675484 708812
rect 670292 708772 670298 708784
rect 675478 708772 675484 708784
rect 675536 708772 675542 708824
rect 671522 708364 671528 708416
rect 671580 708404 671586 708416
rect 675478 708404 675484 708416
rect 671580 708376 675484 708404
rect 671580 708364 671586 708376
rect 675478 708364 675484 708376
rect 675536 708364 675542 708416
rect 674098 707548 674104 707600
rect 674156 707588 674162 707600
rect 675478 707588 675484 707600
rect 674156 707560 675484 707588
rect 674156 707548 674162 707560
rect 675478 707548 675484 707560
rect 675536 707548 675542 707600
rect 42242 706528 42248 706580
rect 42300 706568 42306 706580
rect 43254 706568 43260 706580
rect 42300 706540 43260 706568
rect 42300 706528 42306 706540
rect 43254 706528 43260 706540
rect 43312 706528 43318 706580
rect 672258 706256 672264 706308
rect 672316 706296 672322 706308
rect 675478 706296 675484 706308
rect 672316 706268 675484 706296
rect 672316 706256 672322 706268
rect 675478 706256 675484 706268
rect 675536 706256 675542 706308
rect 675846 705304 675852 705356
rect 675904 705344 675910 705356
rect 683114 705344 683120 705356
rect 675904 705316 683120 705344
rect 675904 705304 675910 705316
rect 683114 705304 683120 705316
rect 683172 705304 683178 705356
rect 670142 705032 670148 705084
rect 670200 705072 670206 705084
rect 675478 705072 675484 705084
rect 670200 705044 675484 705072
rect 670200 705032 670206 705044
rect 675478 705032 675484 705044
rect 675536 705032 675542 705084
rect 42242 704216 42248 704268
rect 42300 704216 42306 704268
rect 42260 704064 42288 704216
rect 42242 704012 42248 704064
rect 42300 704012 42306 704064
rect 42150 702856 42156 702908
rect 42208 702896 42214 702908
rect 42702 702896 42708 702908
rect 42208 702868 42708 702896
rect 42208 702856 42214 702868
rect 42702 702856 42708 702868
rect 42760 702856 42766 702908
rect 51718 701020 51724 701072
rect 51776 701060 51782 701072
rect 62114 701060 62120 701072
rect 51776 701032 62120 701060
rect 51776 701020 51782 701032
rect 62114 701020 62120 701032
rect 62172 701020 62178 701072
rect 42058 700544 42064 700596
rect 42116 700584 42122 700596
rect 42610 700584 42616 700596
rect 42116 700556 42616 700584
rect 42116 700544 42122 700556
rect 42610 700544 42616 700556
rect 42668 700544 42674 700596
rect 672074 698436 672080 698488
rect 672132 698476 672138 698488
rect 675202 698476 675208 698488
rect 672132 698448 675208 698476
rect 672132 698436 672138 698448
rect 675202 698436 675208 698448
rect 675260 698436 675266 698488
rect 673086 697076 673092 697128
rect 673144 697116 673150 697128
rect 675110 697116 675116 697128
rect 673144 697088 675116 697116
rect 673144 697076 673150 697088
rect 675110 697076 675116 697088
rect 675168 697076 675174 697128
rect 651650 696940 651656 696992
rect 651708 696980 651714 696992
rect 661862 696980 661868 696992
rect 651708 696952 661868 696980
rect 651708 696940 651714 696952
rect 661862 696940 661868 696952
rect 661920 696940 661926 696992
rect 674282 694764 674288 694816
rect 674340 694804 674346 694816
rect 675110 694804 675116 694816
rect 674340 694776 675116 694804
rect 674340 694764 674346 694776
rect 675110 694764 675116 694776
rect 675168 694764 675174 694816
rect 674466 694152 674472 694204
rect 674524 694192 674530 694204
rect 675386 694192 675392 694204
rect 674524 694164 675392 694192
rect 674524 694152 674530 694164
rect 675386 694152 675392 694164
rect 675444 694152 675450 694204
rect 666278 692792 666284 692844
rect 666336 692832 666342 692844
rect 675110 692832 675116 692844
rect 666336 692804 675116 692832
rect 666336 692792 666342 692804
rect 675110 692792 675116 692804
rect 675168 692792 675174 692844
rect 659470 689256 659476 689308
rect 659528 689296 659534 689308
rect 674926 689296 674932 689308
rect 659528 689268 674932 689296
rect 659528 689256 659534 689268
rect 674926 689256 674932 689268
rect 674984 689256 674990 689308
rect 674098 689120 674104 689172
rect 674156 689160 674162 689172
rect 675110 689160 675116 689172
rect 674156 689132 675116 689160
rect 674156 689120 674162 689132
rect 675110 689120 675116 689132
rect 675168 689120 675174 689172
rect 43806 688644 43812 688696
rect 43864 688684 43870 688696
rect 62114 688684 62120 688696
rect 43864 688656 62120 688684
rect 43864 688644 43870 688656
rect 62114 688644 62120 688656
rect 62172 688644 62178 688696
rect 42518 687692 42524 687744
rect 42576 687732 42582 687744
rect 50522 687732 50528 687744
rect 42576 687704 50528 687732
rect 42576 687692 42582 687704
rect 50522 687692 50528 687704
rect 50580 687692 50586 687744
rect 43438 687352 43444 687404
rect 43496 687392 43502 687404
rect 51902 687392 51908 687404
rect 43496 687364 51908 687392
rect 43496 687352 43502 687364
rect 51902 687352 51908 687364
rect 51960 687352 51966 687404
rect 40954 687216 40960 687268
rect 41012 687256 41018 687268
rect 41690 687256 41696 687268
rect 41012 687228 41696 687256
rect 41012 687216 41018 687228
rect 41690 687216 41696 687228
rect 41748 687216 41754 687268
rect 42058 687216 42064 687268
rect 42116 687256 42122 687268
rect 56042 687256 56048 687268
rect 42116 687228 56048 687256
rect 42116 687216 42122 687228
rect 56042 687216 56048 687228
rect 56100 687216 56106 687268
rect 672626 687216 672632 687268
rect 672684 687256 672690 687268
rect 675110 687256 675116 687268
rect 672684 687228 675116 687256
rect 672684 687216 672690 687228
rect 675110 687216 675116 687228
rect 675168 687216 675174 687268
rect 41690 686100 41696 686112
rect 41386 686072 41696 686100
rect 41386 686044 41414 686072
rect 41690 686060 41696 686072
rect 41748 686060 41754 686112
rect 42058 686060 42064 686112
rect 42116 686100 42122 686112
rect 45186 686100 45192 686112
rect 42116 686072 45192 686100
rect 42116 686060 42122 686072
rect 45186 686060 45192 686072
rect 45244 686060 45250 686112
rect 41322 685992 41328 686044
rect 41380 686004 41414 686044
rect 41380 685992 41386 686004
rect 41138 685856 41144 685908
rect 41196 685896 41202 685908
rect 41690 685896 41696 685908
rect 41196 685868 41696 685896
rect 41196 685856 41202 685868
rect 41690 685856 41696 685868
rect 41748 685856 41754 685908
rect 42058 685856 42064 685908
rect 42116 685896 42122 685908
rect 45002 685896 45008 685908
rect 42116 685868 45008 685896
rect 42116 685856 42122 685868
rect 45002 685856 45008 685868
rect 45060 685856 45066 685908
rect 669774 685856 669780 685908
rect 669832 685896 669838 685908
rect 674834 685896 674840 685908
rect 669832 685868 674840 685896
rect 669832 685856 669838 685868
rect 674834 685856 674840 685868
rect 674892 685856 674898 685908
rect 40862 684768 40868 684820
rect 40920 684768 40926 684820
rect 40880 684536 40908 684768
rect 41690 684740 41696 684752
rect 41386 684712 41696 684740
rect 41138 684632 41144 684684
rect 41196 684672 41202 684684
rect 41386 684672 41414 684712
rect 41690 684700 41696 684712
rect 41748 684700 41754 684752
rect 42058 684700 42064 684752
rect 42116 684740 42122 684752
rect 43070 684740 43076 684752
rect 42116 684712 43076 684740
rect 42116 684700 42122 684712
rect 43070 684700 43076 684712
rect 43128 684700 43134 684752
rect 41196 684644 41414 684672
rect 41196 684632 41202 684644
rect 41690 684536 41696 684548
rect 40880 684508 41696 684536
rect 41690 684496 41696 684508
rect 41748 684496 41754 684548
rect 42058 684496 42064 684548
rect 42116 684536 42122 684548
rect 44450 684536 44456 684548
rect 42116 684508 44456 684536
rect 42116 684496 42122 684508
rect 44450 684496 44456 684508
rect 44508 684496 44514 684548
rect 41322 683544 41328 683596
rect 41380 683584 41386 683596
rect 41690 683584 41696 683596
rect 41380 683556 41696 683584
rect 41380 683544 41386 683556
rect 41690 683544 41696 683556
rect 41748 683544 41754 683596
rect 42058 683476 42064 683528
rect 42116 683516 42122 683528
rect 42518 683516 42524 683528
rect 42116 683488 42524 683516
rect 42116 683476 42122 683488
rect 42518 683476 42524 683488
rect 42576 683476 42582 683528
rect 42058 683340 42064 683392
rect 42116 683380 42122 683392
rect 42794 683380 42800 683392
rect 42116 683352 42800 683380
rect 42116 683340 42122 683352
rect 42794 683340 42800 683352
rect 42852 683340 42858 683392
rect 40770 683272 40776 683324
rect 40828 683312 40834 683324
rect 41690 683312 41696 683324
rect 40828 683284 41696 683312
rect 40828 683272 40834 683284
rect 41690 683272 41696 683284
rect 41748 683272 41754 683324
rect 41138 683136 41144 683188
rect 41196 683176 41202 683188
rect 41690 683176 41696 683188
rect 41196 683148 41696 683176
rect 41196 683136 41202 683148
rect 41690 683136 41696 683148
rect 41748 683136 41754 683188
rect 42058 683136 42064 683188
rect 42116 683176 42122 683188
rect 42886 683176 42892 683188
rect 42116 683148 42892 683176
rect 42116 683136 42122 683148
rect 42886 683136 42892 683148
rect 42944 683136 42950 683188
rect 651650 683136 651656 683188
rect 651708 683176 651714 683188
rect 658918 683176 658924 683188
rect 651708 683148 658924 683176
rect 651708 683136 651714 683148
rect 658918 683136 658924 683148
rect 658976 683136 658982 683188
rect 41322 682456 41328 682508
rect 41380 682456 41386 682508
rect 41340 682304 41368 682456
rect 675846 682388 675852 682440
rect 675904 682428 675910 682440
rect 683206 682428 683212 682440
rect 675904 682400 683212 682428
rect 675904 682388 675910 682400
rect 683206 682388 683212 682400
rect 683264 682388 683270 682440
rect 41322 682252 41328 682304
rect 41380 682252 41386 682304
rect 676030 682252 676036 682304
rect 676088 682292 676094 682304
rect 683390 682292 683396 682304
rect 676088 682264 683396 682292
rect 676088 682252 676094 682264
rect 683390 682252 683396 682264
rect 683448 682252 683454 682304
rect 42058 676336 42064 676388
rect 42116 676376 42122 676388
rect 50338 676376 50344 676388
rect 42116 676348 50344 676376
rect 42116 676336 42122 676348
rect 50338 676336 50344 676348
rect 50396 676336 50402 676388
rect 42058 675588 42064 675640
rect 42116 675628 42122 675640
rect 42702 675628 42708 675640
rect 42116 675600 42708 675628
rect 42116 675588 42122 675600
rect 42702 675588 42708 675600
rect 42760 675588 42766 675640
rect 34422 675452 34428 675504
rect 34480 675492 34486 675504
rect 39758 675492 39764 675504
rect 34480 675464 39764 675492
rect 34480 675452 34486 675464
rect 39758 675452 39764 675464
rect 39816 675452 39822 675504
rect 47762 674840 47768 674892
rect 47820 674880 47826 674892
rect 62114 674880 62120 674892
rect 47820 674852 62120 674880
rect 47820 674840 47826 674852
rect 62114 674840 62120 674852
rect 62172 674840 62178 674892
rect 31018 672664 31024 672716
rect 31076 672704 31082 672716
rect 40402 672704 40408 672716
rect 31076 672676 40408 672704
rect 31076 672664 31082 672676
rect 40402 672664 40408 672676
rect 40460 672664 40466 672716
rect 36538 672052 36544 672104
rect 36596 672092 36602 672104
rect 41690 672092 41696 672104
rect 36596 672064 41696 672092
rect 36596 672052 36602 672064
rect 41690 672052 41696 672064
rect 41748 672052 41754 672104
rect 675478 671140 675484 671152
rect 663766 671112 675484 671140
rect 663242 670828 663248 670880
rect 663300 670868 663306 670880
rect 663766 670868 663794 671112
rect 675478 671100 675484 671112
rect 675536 671100 675542 671152
rect 663300 670840 663794 670868
rect 663300 670828 663306 670840
rect 661678 670692 661684 670744
rect 661736 670732 661742 670744
rect 675478 670732 675484 670744
rect 661736 670704 675484 670732
rect 661736 670692 661742 670704
rect 675478 670692 675484 670704
rect 675536 670692 675542 670744
rect 674006 670352 674012 670404
rect 674064 670392 674070 670404
rect 675478 670392 675484 670404
rect 674064 670364 675484 670392
rect 674064 670352 674070 670364
rect 675478 670352 675484 670364
rect 675536 670352 675542 670404
rect 670970 669740 670976 669792
rect 671028 669780 671034 669792
rect 675478 669780 675484 669792
rect 671028 669752 675484 669780
rect 671028 669740 671034 669752
rect 675478 669740 675484 669752
rect 675536 669740 675542 669792
rect 671154 669604 671160 669656
rect 671212 669644 671218 669656
rect 675478 669644 675484 669656
rect 671212 669616 675484 669644
rect 671212 669604 671218 669616
rect 675478 669604 675484 669616
rect 675536 669604 675542 669656
rect 660482 669468 660488 669520
rect 660540 669508 660546 669520
rect 674006 669508 674012 669520
rect 660540 669480 674012 669508
rect 660540 669468 660546 669480
rect 674006 669468 674012 669480
rect 674064 669468 674070 669520
rect 651650 669332 651656 669384
rect 651708 669372 651714 669384
rect 662046 669372 662052 669384
rect 651708 669344 662052 669372
rect 651708 669332 651714 669344
rect 662046 669332 662052 669344
rect 662104 669332 662110 669384
rect 671154 669332 671160 669384
rect 671212 669372 671218 669384
rect 674834 669372 674840 669384
rect 671212 669344 674840 669372
rect 671212 669332 671218 669344
rect 674834 669332 674840 669344
rect 674892 669332 674898 669384
rect 671798 668516 671804 668568
rect 671856 668556 671862 668568
rect 675478 668556 675484 668568
rect 671856 668528 675484 668556
rect 671856 668516 671862 668528
rect 675478 668516 675484 668528
rect 675536 668516 675542 668568
rect 671522 667700 671528 667752
rect 671580 667740 671586 667752
rect 675478 667740 675484 667752
rect 671580 667712 675484 667740
rect 671580 667700 671586 667712
rect 675478 667700 675484 667712
rect 675536 667700 675542 667752
rect 671614 667564 671620 667616
rect 671672 667604 671678 667616
rect 674006 667604 674012 667616
rect 671672 667576 674012 667604
rect 671672 667564 671678 667576
rect 674006 667564 674012 667576
rect 674064 667564 674070 667616
rect 670970 667224 670976 667276
rect 671028 667264 671034 667276
rect 675478 667264 675484 667276
rect 671028 667236 675484 667264
rect 671028 667224 671034 667236
rect 675478 667224 675484 667236
rect 675536 667224 675542 667276
rect 42242 667088 42248 667140
rect 42300 667128 42306 667140
rect 43438 667128 43444 667140
rect 42300 667100 43444 667128
rect 42300 667088 42306 667100
rect 43438 667088 43444 667100
rect 43496 667088 43502 667140
rect 43438 666544 43444 666596
rect 43496 666584 43502 666596
rect 45186 666584 45192 666596
rect 43496 666556 45192 666584
rect 43496 666544 43502 666556
rect 45186 666544 45192 666556
rect 45244 666544 45250 666596
rect 669590 666068 669596 666120
rect 669648 666108 669654 666120
rect 675478 666108 675484 666120
rect 669648 666080 675484 666108
rect 669648 666068 669654 666080
rect 675478 666068 675484 666080
rect 675536 666068 675542 666120
rect 666094 665184 666100 665236
rect 666152 665224 666158 665236
rect 675478 665224 675484 665236
rect 666152 665196 675484 665224
rect 666152 665184 666158 665196
rect 675478 665184 675484 665196
rect 675536 665184 675542 665236
rect 42242 664844 42248 664896
rect 42300 664884 42306 664896
rect 43438 664884 43444 664896
rect 42300 664856 43444 664884
rect 42300 664844 42306 664856
rect 43438 664844 43444 664856
rect 43496 664844 43502 664896
rect 672902 664028 672908 664080
rect 672960 664068 672966 664080
rect 674834 664068 674840 664080
rect 672960 664040 674840 664068
rect 672960 664028 672966 664040
rect 674834 664028 674840 664040
rect 674892 664028 674898 664080
rect 669222 663892 669228 663944
rect 669280 663932 669286 663944
rect 675478 663932 675484 663944
rect 669280 663904 675484 663932
rect 669280 663892 669286 663904
rect 675478 663892 675484 663904
rect 675536 663892 675542 663944
rect 668578 663756 668584 663808
rect 668636 663796 668642 663808
rect 675478 663796 675484 663808
rect 668636 663768 675484 663796
rect 668636 663756 668642 663768
rect 675478 663756 675484 663768
rect 675536 663756 675542 663808
rect 42242 663484 42248 663536
rect 42300 663524 42306 663536
rect 42702 663524 42708 663536
rect 42300 663496 42708 663524
rect 42300 663484 42306 663496
rect 42702 663484 42708 663496
rect 42760 663484 42766 663536
rect 673822 663212 673828 663264
rect 673880 663252 673886 663264
rect 675478 663252 675484 663264
rect 673880 663224 675484 663252
rect 673880 663212 673886 663224
rect 675478 663212 675484 663224
rect 675536 663212 675542 663264
rect 42242 662804 42248 662856
rect 42300 662844 42306 662856
rect 43254 662844 43260 662856
rect 42300 662816 43260 662844
rect 42300 662804 42306 662816
rect 43254 662804 43260 662816
rect 43312 662804 43318 662856
rect 670418 662804 670424 662856
rect 670476 662844 670482 662856
rect 675478 662844 675484 662856
rect 670476 662816 675484 662844
rect 670476 662804 670482 662816
rect 675478 662804 675484 662816
rect 675536 662804 675542 662856
rect 43438 662396 43444 662448
rect 43496 662436 43502 662448
rect 62114 662436 62120 662448
rect 43496 662408 62120 662436
rect 43496 662396 43502 662408
rect 62114 662396 62120 662408
rect 62172 662396 62178 662448
rect 671338 661580 671344 661632
rect 671396 661620 671402 661632
rect 675478 661620 675484 661632
rect 671396 661592 675484 661620
rect 671396 661580 671402 661592
rect 675478 661580 675484 661592
rect 675536 661580 675542 661632
rect 671338 661104 671344 661156
rect 671396 661144 671402 661156
rect 675478 661144 675484 661156
rect 671396 661116 675484 661144
rect 671396 661104 671402 661116
rect 675478 661104 675484 661116
rect 675536 661104 675542 661156
rect 670326 659880 670332 659932
rect 670384 659920 670390 659932
rect 675478 659920 675484 659932
rect 670384 659892 675484 659920
rect 670384 659880 670390 659892
rect 675478 659880 675484 659892
rect 675536 659880 675542 659932
rect 675846 659812 675852 659864
rect 675904 659852 675910 659864
rect 683114 659852 683120 659864
rect 675904 659824 683120 659852
rect 675904 659812 675910 659824
rect 683114 659812 683120 659824
rect 683172 659812 683178 659864
rect 42150 657364 42156 657416
rect 42208 657404 42214 657416
rect 42610 657404 42616 657416
rect 42208 657376 42616 657404
rect 42208 657364 42214 657376
rect 42610 657364 42616 657376
rect 42668 657364 42674 657416
rect 651650 656888 651656 656940
rect 651708 656928 651714 656940
rect 661678 656928 661684 656940
rect 651708 656900 661684 656928
rect 651708 656888 651714 656900
rect 661678 656888 661684 656900
rect 661736 656888 661742 656940
rect 665450 654236 665456 654288
rect 665508 654276 665514 654288
rect 675386 654276 675392 654288
rect 665508 654248 675392 654276
rect 665508 654236 665514 654248
rect 675386 654236 675392 654248
rect 675444 654236 675450 654288
rect 672902 651380 672908 651432
rect 672960 651420 672966 651432
rect 675386 651420 675392 651432
rect 672960 651392 675392 651420
rect 672960 651380 672966 651392
rect 675386 651380 675392 651392
rect 675444 651380 675450 651432
rect 669222 650020 669228 650072
rect 669280 650060 669286 650072
rect 674834 650060 674840 650072
rect 669280 650032 674840 650060
rect 669280 650020 669286 650032
rect 674834 650020 674840 650032
rect 674892 650020 674898 650072
rect 671706 649068 671712 649120
rect 671764 649108 671770 649120
rect 675386 649108 675392 649120
rect 671764 649080 675392 649108
rect 671764 649068 671770 649080
rect 675386 649068 675392 649080
rect 675444 649068 675450 649120
rect 674834 648592 674840 648644
rect 674892 648632 674898 648644
rect 675386 648632 675392 648644
rect 674892 648604 675392 648632
rect 674892 648592 674898 648604
rect 675386 648592 675392 648604
rect 675444 648592 675450 648644
rect 51902 647844 51908 647896
rect 51960 647884 51966 647896
rect 62114 647884 62120 647896
rect 51960 647856 62120 647884
rect 51960 647844 51966 647856
rect 62114 647844 62120 647856
rect 62172 647844 62178 647896
rect 665266 647708 665272 647760
rect 665324 647748 665330 647760
rect 670786 647748 670792 647760
rect 665324 647720 670792 647748
rect 665324 647708 665330 647720
rect 670786 647708 670792 647720
rect 670844 647708 670850 647760
rect 35802 644716 35808 644768
rect 35860 644756 35866 644768
rect 38838 644756 38844 644768
rect 35860 644728 38844 644756
rect 35860 644716 35866 644728
rect 38838 644716 38844 644728
rect 38896 644716 38902 644768
rect 35526 644444 35532 644496
rect 35584 644484 35590 644496
rect 41230 644484 41236 644496
rect 35584 644456 41236 644484
rect 35584 644444 35590 644456
rect 41230 644444 41236 644456
rect 41288 644444 41294 644496
rect 662046 643696 662052 643748
rect 662104 643736 662110 643748
rect 662104 643708 663794 643736
rect 662104 643696 662110 643708
rect 663766 643668 663794 643708
rect 670786 643668 670792 643680
rect 663766 643640 670792 643668
rect 670786 643628 670792 643640
rect 670844 643628 670850 643680
rect 35802 643492 35808 643544
rect 35860 643532 35866 643544
rect 40310 643532 40316 643544
rect 35860 643504 40316 643532
rect 35860 643492 35866 643504
rect 40310 643492 40316 643504
rect 40368 643492 40374 643544
rect 41690 643328 41696 643340
rect 41386 643300 41696 643328
rect 35526 643220 35532 643272
rect 35584 643260 35590 643272
rect 41386 643260 41414 643300
rect 41690 643288 41696 643300
rect 41748 643288 41754 643340
rect 42058 643288 42064 643340
rect 42116 643328 42122 643340
rect 44266 643328 44272 643340
rect 42116 643300 44272 643328
rect 42116 643288 42122 643300
rect 44266 643288 44272 643300
rect 44324 643288 44330 643340
rect 35584 643232 41414 643260
rect 35584 643220 35590 643232
rect 35342 643084 35348 643136
rect 35400 643124 35406 643136
rect 41690 643124 41696 643136
rect 35400 643096 41696 643124
rect 35400 643084 35406 643096
rect 41690 643084 41696 643096
rect 41748 643084 41754 643136
rect 42058 643084 42064 643136
rect 42116 643124 42122 643136
rect 51718 643124 51724 643136
rect 42116 643096 51724 643124
rect 42116 643084 42122 643096
rect 51718 643084 51724 643096
rect 51776 643084 51782 643136
rect 651650 643084 651656 643136
rect 651708 643124 651714 643136
rect 664806 643124 664812 643136
rect 651708 643096 664812 643124
rect 651708 643084 651714 643096
rect 664806 643084 664812 643096
rect 664864 643084 664870 643136
rect 39022 642240 39028 642252
rect 38626 642212 39028 642240
rect 35802 642132 35808 642184
rect 35860 642172 35866 642184
rect 38626 642172 38654 642212
rect 39022 642200 39028 642212
rect 39080 642200 39086 642252
rect 35860 642144 38654 642172
rect 35860 642132 35866 642144
rect 39666 641968 39672 641980
rect 36004 641940 39672 641968
rect 35434 641860 35440 641912
rect 35492 641900 35498 641912
rect 36004 641900 36032 641940
rect 39666 641928 39672 641940
rect 39724 641928 39730 641980
rect 35492 641872 36032 641900
rect 35492 641860 35498 641872
rect 670786 641860 670792 641912
rect 670844 641900 670850 641912
rect 675294 641900 675300 641912
rect 670844 641872 675300 641900
rect 670844 641860 670850 641872
rect 675294 641860 675300 641872
rect 675352 641860 675358 641912
rect 35618 641724 35624 641776
rect 35676 641764 35682 641776
rect 39758 641764 39764 641776
rect 35676 641736 39764 641764
rect 35676 641724 35682 641736
rect 39758 641724 39764 641736
rect 39816 641724 39822 641776
rect 666094 641724 666100 641776
rect 666152 641764 666158 641776
rect 670786 641764 670792 641776
rect 666152 641736 670792 641764
rect 666152 641724 666158 641736
rect 670786 641724 670792 641736
rect 670844 641724 670850 641776
rect 42058 640908 42064 640960
rect 42116 640948 42122 640960
rect 42886 640948 42892 640960
rect 42116 640920 42892 640948
rect 42116 640908 42122 640920
rect 42886 640908 42892 640920
rect 42944 640908 42950 640960
rect 35802 640704 35808 640756
rect 35860 640744 35866 640756
rect 39850 640744 39856 640756
rect 35860 640716 39856 640744
rect 35860 640704 35866 640716
rect 39850 640704 39856 640716
rect 39908 640704 39914 640756
rect 35526 640432 35532 640484
rect 35584 640472 35590 640484
rect 41690 640472 41696 640484
rect 35584 640444 41696 640472
rect 35584 640432 35590 640444
rect 41690 640432 41696 640444
rect 41748 640432 41754 640484
rect 35342 640296 35348 640348
rect 35400 640336 35406 640348
rect 41690 640336 41696 640348
rect 35400 640308 41696 640336
rect 35400 640296 35406 640308
rect 41690 640296 41696 640308
rect 41748 640296 41754 640348
rect 42058 640296 42064 640348
rect 42116 640336 42122 640348
rect 43162 640336 43168 640348
rect 42116 640308 43168 640336
rect 42116 640296 42122 640308
rect 43162 640296 43168 640308
rect 43220 640296 43226 640348
rect 670786 640024 670792 640076
rect 670844 640064 670850 640076
rect 675294 640064 675300 640076
rect 670844 640036 675300 640064
rect 670844 640024 670850 640036
rect 675294 640024 675300 640036
rect 675352 640024 675358 640076
rect 35802 639072 35808 639124
rect 35860 639112 35866 639124
rect 40218 639112 40224 639124
rect 35860 639084 40224 639112
rect 35860 639072 35866 639084
rect 40218 639072 40224 639084
rect 40276 639072 40282 639124
rect 673454 639004 673460 639056
rect 673512 639044 673518 639056
rect 675294 639044 675300 639056
rect 673512 639016 675300 639044
rect 673512 639004 673518 639016
rect 675294 639004 675300 639016
rect 675352 639004 675358 639056
rect 35526 638936 35532 638988
rect 35584 638976 35590 638988
rect 40034 638976 40040 638988
rect 35584 638948 40040 638976
rect 35584 638936 35590 638948
rect 40034 638936 40040 638948
rect 40092 638936 40098 638988
rect 34422 638188 34428 638240
rect 34480 638228 34486 638240
rect 41690 638228 41696 638240
rect 34480 638200 41696 638228
rect 34480 638188 34486 638200
rect 41690 638188 41696 638200
rect 41748 638188 41754 638240
rect 42058 638120 42064 638172
rect 42116 638160 42122 638172
rect 42702 638160 42708 638172
rect 42116 638132 42708 638160
rect 42116 638120 42122 638132
rect 42702 638120 42708 638132
rect 42760 638120 42766 638172
rect 35526 637916 35532 637968
rect 35584 637956 35590 637968
rect 41690 637956 41696 637968
rect 35584 637928 41696 637956
rect 35584 637916 35590 637928
rect 41690 637916 41696 637928
rect 41748 637916 41754 637968
rect 42058 637848 42064 637900
rect 42116 637888 42122 637900
rect 43622 637888 43628 637900
rect 42116 637860 43628 637888
rect 42116 637848 42122 637860
rect 43622 637848 43628 637860
rect 43680 637848 43686 637900
rect 35802 637712 35808 637764
rect 35860 637752 35866 637764
rect 41506 637752 41512 637764
rect 35860 637724 41512 637752
rect 35860 637712 35866 637724
rect 41506 637712 41512 637724
rect 41564 637712 41570 637764
rect 675846 637440 675852 637492
rect 675904 637480 675910 637492
rect 679618 637480 679624 637492
rect 675904 637452 679624 637480
rect 675904 637440 675910 637452
rect 679618 637440 679624 637452
rect 679676 637440 679682 637492
rect 674374 636896 674380 636948
rect 674432 636936 674438 636948
rect 674432 636908 674834 636936
rect 674432 636896 674438 636908
rect 674806 636868 674834 636908
rect 675478 636868 675484 636880
rect 674806 636840 675484 636868
rect 675478 636828 675484 636840
rect 675536 636828 675542 636880
rect 35802 636352 35808 636404
rect 35860 636392 35866 636404
rect 41322 636392 41328 636404
rect 35860 636364 41328 636392
rect 35860 636352 35866 636364
rect 41322 636352 41328 636364
rect 41380 636352 41386 636404
rect 49142 636216 49148 636268
rect 49200 636256 49206 636268
rect 62114 636256 62120 636268
rect 49200 636228 62120 636256
rect 49200 636216 49206 636228
rect 62114 636216 62120 636228
rect 62172 636216 62178 636268
rect 675846 636148 675852 636200
rect 675904 636188 675910 636200
rect 682378 636188 682384 636200
rect 675904 636160 682384 636188
rect 675904 636148 675910 636160
rect 682378 636148 682384 636160
rect 682436 636148 682442 636200
rect 35802 635060 35808 635112
rect 35860 635100 35866 635112
rect 39758 635100 39764 635112
rect 35860 635072 39764 635100
rect 35860 635060 35866 635072
rect 39758 635060 39764 635072
rect 39816 635060 39822 635112
rect 35618 634788 35624 634840
rect 35676 634828 35682 634840
rect 39298 634828 39304 634840
rect 35676 634800 39304 634828
rect 35676 634788 35682 634800
rect 39298 634788 39304 634800
rect 39356 634788 39362 634840
rect 35802 633632 35808 633684
rect 35860 633672 35866 633684
rect 41690 633672 41696 633684
rect 35860 633644 41696 633672
rect 35860 633632 35866 633644
rect 41690 633632 41696 633644
rect 41748 633632 41754 633684
rect 42058 633632 42064 633684
rect 42116 633672 42122 633684
rect 51718 633672 51724 633684
rect 42116 633644 51724 633672
rect 42116 633632 42122 633644
rect 51718 633632 51724 633644
rect 51776 633632 51782 633684
rect 35618 633428 35624 633480
rect 35676 633468 35682 633480
rect 41690 633468 41696 633480
rect 35676 633440 41696 633468
rect 35676 633428 35682 633440
rect 41690 633428 41696 633440
rect 41748 633428 41754 633480
rect 42058 633428 42064 633480
rect 42116 633468 42122 633480
rect 50522 633468 50528 633480
rect 42116 633440 50528 633468
rect 42116 633428 42122 633440
rect 50522 633428 50528 633440
rect 50580 633428 50586 633480
rect 33778 630028 33784 630080
rect 33836 630068 33842 630080
rect 41690 630068 41696 630080
rect 33836 630040 41696 630068
rect 33836 630028 33842 630040
rect 41690 630028 41696 630040
rect 41748 630028 41754 630080
rect 42058 629960 42064 630012
rect 42116 630000 42122 630012
rect 42702 630000 42708 630012
rect 42116 629972 42708 630000
rect 42116 629960 42122 629972
rect 42702 629960 42708 629972
rect 42760 629960 42766 630012
rect 32398 629892 32404 629944
rect 32456 629932 32462 629944
rect 41690 629932 41696 629944
rect 32456 629904 41696 629932
rect 32456 629892 32462 629904
rect 41690 629892 41696 629904
rect 41748 629892 41754 629944
rect 652018 629280 652024 629332
rect 652076 629320 652082 629332
rect 659102 629320 659108 629332
rect 652076 629292 659108 629320
rect 652076 629280 652082 629292
rect 659102 629280 659108 629292
rect 659160 629280 659166 629332
rect 50706 626668 50712 626680
rect 42628 626640 50712 626668
rect 42628 626544 42656 626640
rect 50706 626628 50712 626640
rect 50764 626628 50770 626680
rect 42610 626492 42616 626544
rect 42668 626492 42674 626544
rect 659286 625404 659292 625456
rect 659344 625444 659350 625456
rect 675294 625444 675300 625456
rect 659344 625416 675300 625444
rect 659344 625404 659350 625416
rect 675294 625404 675300 625416
rect 675352 625404 675358 625456
rect 664622 625268 664628 625320
rect 664680 625308 664686 625320
rect 675478 625308 675484 625320
rect 664680 625280 675484 625308
rect 664680 625268 664686 625280
rect 675478 625268 675484 625280
rect 675536 625268 675542 625320
rect 660298 625132 660304 625184
rect 660356 625172 660362 625184
rect 675110 625172 675116 625184
rect 660356 625144 675116 625172
rect 660356 625132 660362 625144
rect 675110 625132 675116 625144
rect 675168 625132 675174 625184
rect 671522 624248 671528 624300
rect 671580 624288 671586 624300
rect 675478 624288 675484 624300
rect 671580 624260 675484 624288
rect 671580 624248 671586 624260
rect 675478 624248 675484 624260
rect 675536 624248 675542 624300
rect 671154 624044 671160 624096
rect 671212 624084 671218 624096
rect 675294 624084 675300 624096
rect 671212 624056 675300 624084
rect 671212 624044 671218 624056
rect 675294 624044 675300 624056
rect 675352 624044 675358 624096
rect 671154 623908 671160 623960
rect 671212 623948 671218 623960
rect 675478 623948 675484 623960
rect 671212 623920 675484 623948
rect 671212 623908 671218 623920
rect 675478 623908 675484 623920
rect 675536 623908 675542 623960
rect 43806 623812 43812 623824
rect 42352 623784 43812 623812
rect 42352 623416 42380 623784
rect 43806 623772 43812 623784
rect 43864 623772 43870 623824
rect 47762 623772 47768 623824
rect 47820 623812 47826 623824
rect 62114 623812 62120 623824
rect 47820 623784 62120 623812
rect 47820 623772 47826 623784
rect 62114 623772 62120 623784
rect 62172 623772 62178 623824
rect 670786 623772 670792 623824
rect 670844 623812 670850 623824
rect 675110 623812 675116 623824
rect 670844 623784 675116 623812
rect 670844 623772 670850 623784
rect 675110 623772 675116 623784
rect 675168 623772 675174 623824
rect 42334 623364 42340 623416
rect 42392 623364 42398 623416
rect 671614 622820 671620 622872
rect 671672 622860 671678 622872
rect 675478 622860 675484 622872
rect 671672 622832 675484 622860
rect 671672 622820 671678 622832
rect 675478 622820 675484 622832
rect 675536 622820 675542 622872
rect 671706 622548 671712 622600
rect 671764 622588 671770 622600
rect 675294 622588 675300 622600
rect 671764 622560 675300 622588
rect 671764 622548 671770 622560
rect 675294 622548 675300 622560
rect 675352 622548 675358 622600
rect 45186 622452 45192 622464
rect 42444 622424 45192 622452
rect 42444 622056 42472 622424
rect 45186 622412 45192 622424
rect 45244 622412 45250 622464
rect 670970 622412 670976 622464
rect 671028 622452 671034 622464
rect 675478 622452 675484 622464
rect 671028 622424 675484 622452
rect 671028 622412 671034 622424
rect 675478 622412 675484 622424
rect 675536 622412 675542 622464
rect 42426 622004 42432 622056
rect 42484 622004 42490 622056
rect 671890 621188 671896 621240
rect 671948 621228 671954 621240
rect 675478 621228 675484 621240
rect 671948 621200 675484 621228
rect 671948 621188 671954 621200
rect 675478 621188 675484 621200
rect 675536 621188 675542 621240
rect 671890 620984 671896 621036
rect 671948 621024 671954 621036
rect 675294 621024 675300 621036
rect 671948 620996 675300 621024
rect 671948 620984 671954 620996
rect 675294 620984 675300 620996
rect 675352 620984 675358 621036
rect 669774 619828 669780 619880
rect 669832 619868 669838 619880
rect 675294 619868 675300 619880
rect 669832 619840 675300 619868
rect 669832 619828 669838 619840
rect 675294 619828 675300 619840
rect 675352 619828 675358 619880
rect 666278 619624 666284 619676
rect 666336 619664 666342 619676
rect 675478 619664 675484 619676
rect 666336 619636 675484 619664
rect 666336 619624 666342 619636
rect 675478 619624 675484 619636
rect 675536 619624 675542 619676
rect 673086 619420 673092 619472
rect 673144 619460 673150 619472
rect 675478 619460 675484 619472
rect 673144 619432 675484 619460
rect 673144 619420 673150 619432
rect 675478 619420 675484 619432
rect 675536 619420 675542 619472
rect 42610 618876 42616 618928
rect 42668 618916 42674 618928
rect 43622 618916 43628 618928
rect 42668 618888 43628 618916
rect 42668 618876 42674 618888
rect 43622 618876 43628 618888
rect 43680 618876 43686 618928
rect 672626 618196 672632 618248
rect 672684 618236 672690 618248
rect 675478 618236 675484 618248
rect 672684 618208 675484 618236
rect 672684 618196 672690 618208
rect 675478 618196 675484 618208
rect 675536 618196 675542 618248
rect 651650 616836 651656 616888
rect 651708 616876 651714 616888
rect 660482 616876 660488 616888
rect 651708 616848 660488 616876
rect 651708 616836 651714 616848
rect 660482 616836 660488 616848
rect 660540 616836 660546 616888
rect 671522 616632 671528 616684
rect 671580 616672 671586 616684
rect 671890 616672 671896 616684
rect 671580 616644 671896 616672
rect 671580 616632 671586 616644
rect 671890 616632 671896 616644
rect 671948 616632 671954 616684
rect 671706 616496 671712 616548
rect 671764 616496 671770 616548
rect 671724 616412 671752 616496
rect 671706 616360 671712 616412
rect 671764 616360 671770 616412
rect 670970 616088 670976 616140
rect 671028 616128 671034 616140
rect 675294 616128 675300 616140
rect 671028 616100 675300 616128
rect 671028 616088 671034 616100
rect 675294 616088 675300 616100
rect 675352 616088 675358 616140
rect 668762 615748 668768 615800
rect 668820 615788 668826 615800
rect 675478 615788 675484 615800
rect 668820 615760 675484 615788
rect 668820 615748 668826 615760
rect 675478 615748 675484 615760
rect 675536 615748 675542 615800
rect 42242 615680 42248 615732
rect 42300 615680 42306 615732
rect 42260 615528 42288 615680
rect 675846 615612 675852 615664
rect 675904 615652 675910 615664
rect 683114 615652 683120 615664
rect 675904 615624 683120 615652
rect 675904 615612 675910 615624
rect 683114 615612 683120 615624
rect 683172 615612 683178 615664
rect 42242 615476 42248 615528
rect 42300 615476 42306 615528
rect 663702 614116 663708 614168
rect 663760 614156 663766 614168
rect 675478 614156 675484 614168
rect 663760 614128 675484 614156
rect 663760 614116 663766 614128
rect 675478 614116 675484 614128
rect 675536 614116 675542 614168
rect 42150 613572 42156 613624
rect 42208 613612 42214 613624
rect 44450 613612 44456 613624
rect 42208 613584 44456 613612
rect 42208 613572 42214 613584
rect 44450 613572 44456 613584
rect 44508 613572 44514 613624
rect 668578 610104 668584 610156
rect 668636 610144 668642 610156
rect 671338 610144 671344 610156
rect 668636 610116 671344 610144
rect 668636 610104 668642 610116
rect 671338 610104 671344 610116
rect 671396 610104 671402 610156
rect 666370 609968 666376 610020
rect 666428 610008 666434 610020
rect 675110 610008 675116 610020
rect 666428 609980 675116 610008
rect 666428 609968 666434 609980
rect 675110 609968 675116 609980
rect 675168 609968 675174 610020
rect 43622 609220 43628 609272
rect 43680 609260 43686 609272
rect 62114 609260 62120 609272
rect 43680 609232 62120 609260
rect 43680 609220 43686 609232
rect 62114 609220 62120 609232
rect 62172 609220 62178 609272
rect 673086 607588 673092 607640
rect 673144 607628 673150 607640
rect 675294 607628 675300 607640
rect 673144 607600 675300 607628
rect 673144 607588 673150 607600
rect 675294 607588 675300 607600
rect 675352 607588 675358 607640
rect 672534 605820 672540 605872
rect 672592 605860 672598 605872
rect 675110 605860 675116 605872
rect 672592 605832 675116 605860
rect 672592 605820 672598 605832
rect 675110 605820 675116 605832
rect 675168 605820 675174 605872
rect 674650 603304 674656 603356
rect 674708 603344 674714 603356
rect 675386 603344 675392 603356
rect 674708 603316 675392 603344
rect 674708 603304 674714 603316
rect 675386 603304 675392 603316
rect 675444 603304 675450 603356
rect 669286 603180 674144 603208
rect 652018 603100 652024 603152
rect 652076 603140 652082 603152
rect 660298 603140 660304 603152
rect 652076 603112 660304 603140
rect 652076 603100 652082 603112
rect 660298 603100 660304 603112
rect 660356 603100 660362 603152
rect 665634 603100 665640 603152
rect 665692 603140 665698 603152
rect 669286 603140 669314 603180
rect 665692 603112 669314 603140
rect 665692 603100 665698 603112
rect 674116 603072 674144 603180
rect 675294 603072 675300 603084
rect 674116 603044 675300 603072
rect 675294 603032 675300 603044
rect 675352 603032 675358 603084
rect 35802 601672 35808 601724
rect 35860 601712 35866 601724
rect 41690 601712 41696 601724
rect 35860 601684 41696 601712
rect 35860 601672 35866 601684
rect 41690 601672 41696 601684
rect 41748 601672 41754 601724
rect 42058 601672 42064 601724
rect 42116 601712 42122 601724
rect 49142 601712 49148 601724
rect 42116 601684 49148 601712
rect 42116 601672 42122 601684
rect 49142 601672 49148 601684
rect 49200 601672 49206 601724
rect 674006 601332 674012 601384
rect 674064 601372 674070 601384
rect 674650 601372 674656 601384
rect 674064 601344 674656 601372
rect 674064 601332 674070 601344
rect 674650 601332 674656 601344
rect 674708 601332 674714 601384
rect 42610 600380 42616 600432
rect 42668 600420 42674 600432
rect 42668 600392 51074 600420
rect 42668 600380 42674 600392
rect 51046 600352 51074 600392
rect 51902 600352 51908 600364
rect 51046 600324 51908 600352
rect 51902 600312 51908 600324
rect 51960 600312 51966 600364
rect 660482 599564 660488 599616
rect 660540 599604 660546 599616
rect 660540 599576 663794 599604
rect 660540 599564 660546 599576
rect 663766 599400 663794 599576
rect 674282 599496 674288 599548
rect 674340 599536 674346 599548
rect 675110 599536 675116 599548
rect 674340 599508 675116 599536
rect 674340 599496 674346 599508
rect 675110 599496 675116 599508
rect 675168 599496 675174 599548
rect 675110 599400 675116 599412
rect 663766 599372 675116 599400
rect 675110 599360 675116 599372
rect 675168 599360 675174 599412
rect 41322 598952 41328 599004
rect 41380 598992 41386 599004
rect 41690 598992 41696 599004
rect 41380 598964 41696 598992
rect 41380 598952 41386 598964
rect 41690 598952 41696 598964
rect 41748 598952 41754 599004
rect 42058 598952 42064 599004
rect 42116 598992 42122 599004
rect 44450 598992 44456 599004
rect 42116 598964 44456 598992
rect 42116 598952 42122 598964
rect 44450 598952 44456 598964
rect 44508 598952 44514 599004
rect 668854 598748 668860 598800
rect 668912 598788 668918 598800
rect 668912 598760 669314 598788
rect 668912 598748 668918 598760
rect 669286 598720 669314 598760
rect 675294 598720 675300 598732
rect 669286 598692 675300 598720
rect 675294 598680 675300 598692
rect 675352 598680 675358 598732
rect 41322 597796 41328 597848
rect 41380 597836 41386 597848
rect 41690 597836 41696 597848
rect 41380 597808 41696 597836
rect 41380 597796 41386 597808
rect 41690 597796 41696 597808
rect 41748 597796 41754 597848
rect 42058 597796 42064 597848
rect 42116 597836 42122 597848
rect 42794 597836 42800 597848
rect 42116 597808 42800 597836
rect 42116 597796 42122 597808
rect 42794 597796 42800 597808
rect 42852 597796 42858 597848
rect 41046 597660 41052 597712
rect 41104 597700 41110 597712
rect 41690 597700 41696 597712
rect 41104 597672 41696 597700
rect 41104 597660 41110 597672
rect 41690 597660 41696 597672
rect 41748 597660 41754 597712
rect 42058 597660 42064 597712
rect 42116 597700 42122 597712
rect 42978 597700 42984 597712
rect 42116 597672 42984 597700
rect 42116 597660 42122 597672
rect 42978 597660 42984 597672
rect 43036 597660 43042 597712
rect 40862 597524 40868 597576
rect 40920 597564 40926 597576
rect 41690 597564 41696 597576
rect 40920 597536 41696 597564
rect 40920 597524 40926 597536
rect 41690 597524 41696 597536
rect 41748 597524 41754 597576
rect 42058 597524 42064 597576
rect 42116 597564 42122 597576
rect 43070 597564 43076 597576
rect 42116 597536 43076 597564
rect 42116 597524 42122 597536
rect 43070 597524 43076 597536
rect 43128 597524 43134 597576
rect 49142 597524 49148 597576
rect 49200 597564 49206 597576
rect 62114 597564 62120 597576
rect 49200 597536 62120 597564
rect 49200 597524 49206 597536
rect 62114 597524 62120 597536
rect 62172 597524 62178 597576
rect 674558 597456 674564 597508
rect 674616 597496 674622 597508
rect 675294 597496 675300 597508
rect 674616 597468 675300 597496
rect 674616 597456 674622 597468
rect 675294 597456 675300 597468
rect 675352 597456 675358 597508
rect 41322 596436 41328 596488
rect 41380 596476 41386 596488
rect 41690 596476 41696 596488
rect 41380 596448 41696 596476
rect 41380 596436 41386 596448
rect 41690 596436 41696 596448
rect 41748 596436 41754 596488
rect 41138 596028 41144 596080
rect 41196 596068 41202 596080
rect 41598 596068 41604 596080
rect 41196 596040 41604 596068
rect 41196 596028 41202 596040
rect 41598 596028 41604 596040
rect 41656 596028 41662 596080
rect 41322 594736 41328 594788
rect 41380 594776 41386 594788
rect 41690 594776 41696 594788
rect 41380 594748 41696 594776
rect 41380 594736 41386 594748
rect 41690 594736 41696 594748
rect 41748 594736 41754 594788
rect 40586 593036 40592 593088
rect 40644 593076 40650 593088
rect 41598 593076 41604 593088
rect 40644 593048 41604 593076
rect 40644 593036 40650 593048
rect 41598 593036 41604 593048
rect 41656 593036 41662 593088
rect 40770 592696 40776 592748
rect 40828 592736 40834 592748
rect 41598 592736 41604 592748
rect 40828 592708 41604 592736
rect 40828 592696 40834 592708
rect 41598 592696 41604 592708
rect 41656 592696 41662 592748
rect 673914 591540 673920 591592
rect 673972 591580 673978 591592
rect 675478 591580 675484 591592
rect 673972 591552 675484 591580
rect 673972 591540 673978 591552
rect 675478 591540 675484 591552
rect 675536 591540 675542 591592
rect 675846 591404 675852 591456
rect 675904 591444 675910 591456
rect 683206 591444 683212 591456
rect 675904 591416 683212 591444
rect 675904 591404 675910 591416
rect 683206 591404 683212 591416
rect 683264 591404 683270 591456
rect 675846 591268 675852 591320
rect 675904 591308 675910 591320
rect 683390 591308 683396 591320
rect 675904 591280 683396 591308
rect 675904 591268 675910 591280
rect 683390 591268 683396 591280
rect 683448 591268 683454 591320
rect 43806 590656 43812 590708
rect 43864 590696 43870 590708
rect 56042 590696 56048 590708
rect 43864 590668 56048 590696
rect 43864 590656 43870 590668
rect 56042 590656 56048 590668
rect 56100 590656 56106 590708
rect 651650 590656 651656 590708
rect 651708 590696 651714 590708
rect 663242 590696 663248 590708
rect 651708 590668 663248 590696
rect 651708 590656 651714 590668
rect 663242 590656 663248 590668
rect 663300 590656 663306 590708
rect 33042 586984 33048 587036
rect 33100 587024 33106 587036
rect 40126 587024 40132 587036
rect 33100 586996 40132 587024
rect 33100 586984 33106 586996
rect 40126 586984 40132 586996
rect 40184 586984 40190 587036
rect 35158 585896 35164 585948
rect 35216 585936 35222 585948
rect 41598 585936 41604 585948
rect 35216 585908 41604 585936
rect 35216 585896 35222 585908
rect 41598 585896 41604 585908
rect 41656 585896 41662 585948
rect 31018 585692 31024 585744
rect 31076 585732 31082 585744
rect 41598 585732 41604 585744
rect 31076 585704 41604 585732
rect 31076 585692 31082 585704
rect 41598 585692 41604 585704
rect 41656 585692 41662 585744
rect 39942 585352 39948 585404
rect 40000 585392 40006 585404
rect 41414 585392 41420 585404
rect 40000 585364 41420 585392
rect 40000 585352 40006 585364
rect 41414 585352 41420 585364
rect 41472 585352 41478 585404
rect 36538 585148 36544 585200
rect 36596 585188 36602 585200
rect 39390 585188 39396 585200
rect 36596 585160 39396 585188
rect 36596 585148 36602 585160
rect 39390 585148 39396 585160
rect 39448 585148 39454 585200
rect 42058 584400 42064 584452
rect 42116 584440 42122 584452
rect 42702 584440 42708 584452
rect 42116 584412 42708 584440
rect 42116 584400 42122 584412
rect 42702 584400 42708 584412
rect 42760 584400 42766 584452
rect 51902 583720 51908 583772
rect 51960 583760 51966 583772
rect 62114 583760 62120 583772
rect 51960 583732 62120 583760
rect 51960 583720 51966 583732
rect 62114 583720 62120 583732
rect 62172 583720 62178 583772
rect 661862 581000 661868 581052
rect 661920 581040 661926 581052
rect 675478 581040 675484 581052
rect 661920 581012 675484 581040
rect 661920 581000 661926 581012
rect 675478 581000 675484 581012
rect 675536 581000 675542 581052
rect 42426 580592 42432 580644
rect 42484 580632 42490 580644
rect 44634 580632 44640 580644
rect 42484 580604 44640 580632
rect 42484 580592 42490 580604
rect 44634 580592 44640 580604
rect 44692 580592 44698 580644
rect 670786 579980 670792 580032
rect 670844 580020 670850 580032
rect 674742 580020 674748 580032
rect 670844 579992 674748 580020
rect 670844 579980 670850 579992
rect 674742 579980 674748 579992
rect 674800 579980 674806 580032
rect 663058 579776 663064 579828
rect 663116 579816 663122 579828
rect 675294 579816 675300 579828
rect 663116 579788 675300 579816
rect 663116 579776 663122 579788
rect 675294 579776 675300 579788
rect 675352 579776 675358 579828
rect 658918 579640 658924 579692
rect 658976 579680 658982 579692
rect 675478 579680 675484 579692
rect 658976 579652 675484 579680
rect 658976 579640 658982 579652
rect 675478 579640 675484 579652
rect 675536 579640 675542 579692
rect 671154 579368 671160 579420
rect 671212 579408 671218 579420
rect 675478 579408 675484 579420
rect 671212 579380 675484 579408
rect 671212 579368 671218 579380
rect 675478 579368 675484 579380
rect 675536 579368 675542 579420
rect 671338 579028 671344 579080
rect 671396 579068 671402 579080
rect 675478 579068 675484 579080
rect 671396 579040 675484 579068
rect 671396 579028 671402 579040
rect 675478 579028 675484 579040
rect 675536 579028 675542 579080
rect 42242 578688 42248 578740
rect 42300 578688 42306 578740
rect 42260 578468 42288 578688
rect 672718 578552 672724 578604
rect 672776 578592 672782 578604
rect 675478 578592 675484 578604
rect 672776 578564 675484 578592
rect 672776 578552 672782 578564
rect 675478 578552 675484 578564
rect 675536 578552 675542 578604
rect 42242 578416 42248 578468
rect 42300 578416 42306 578468
rect 672902 578212 672908 578264
rect 672960 578252 672966 578264
rect 675478 578252 675484 578264
rect 672960 578224 675484 578252
rect 672960 578212 672966 578224
rect 675478 578212 675484 578224
rect 675536 578212 675542 578264
rect 671614 578008 671620 578060
rect 671672 578048 671678 578060
rect 675294 578048 675300 578060
rect 671672 578020 675300 578048
rect 671672 578008 671678 578020
rect 675294 578008 675300 578020
rect 675352 578008 675358 578060
rect 671522 577736 671528 577788
rect 671580 577776 671586 577788
rect 675294 577776 675300 577788
rect 671580 577748 675300 577776
rect 671580 577736 671586 577748
rect 675294 577736 675300 577748
rect 675352 577736 675358 577788
rect 673730 577532 673736 577584
rect 673788 577572 673794 577584
rect 674098 577572 674104 577584
rect 673788 577544 674104 577572
rect 673788 577532 673794 577544
rect 674098 577532 674104 577544
rect 674156 577532 674162 577584
rect 671338 577396 671344 577448
rect 671396 577436 671402 577448
rect 675294 577436 675300 577448
rect 671396 577408 675300 577436
rect 671396 577396 671402 577408
rect 675294 577396 675300 577408
rect 675352 577396 675358 577448
rect 671338 576920 671344 576972
rect 671396 576960 671402 576972
rect 675294 576960 675300 576972
rect 671396 576932 675300 576960
rect 671396 576920 671402 576932
rect 675294 576920 675300 576932
rect 675352 576920 675358 576972
rect 651650 576852 651656 576904
rect 651708 576892 651714 576904
rect 664622 576892 664628 576904
rect 651708 576864 664628 576892
rect 651708 576852 651714 576864
rect 664622 576852 664628 576864
rect 664680 576852 664686 576904
rect 675478 574308 675484 574320
rect 669286 574280 675484 574308
rect 665450 574200 665456 574252
rect 665508 574240 665514 574252
rect 669286 574240 669314 574280
rect 675478 574268 675484 574280
rect 675536 574268 675542 574320
rect 665508 574212 669314 574240
rect 665508 574200 665514 574212
rect 665266 574064 665272 574116
rect 665324 574104 665330 574116
rect 675294 574104 675300 574116
rect 665324 574076 675300 574104
rect 665324 574064 665330 574076
rect 675294 574064 675300 574076
rect 675352 574064 675358 574116
rect 671798 573724 671804 573776
rect 671856 573764 671862 573776
rect 675478 573764 675484 573776
rect 671856 573736 675484 573764
rect 671856 573724 671862 573736
rect 675478 573724 675484 573736
rect 675536 573724 675542 573776
rect 669590 572908 669596 572960
rect 669648 572948 669654 572960
rect 675478 572948 675484 572960
rect 669648 572920 675484 572948
rect 669648 572908 669654 572920
rect 675478 572908 675484 572920
rect 675536 572908 675542 572960
rect 674098 572500 674104 572552
rect 674156 572540 674162 572552
rect 675478 572540 675484 572552
rect 674156 572512 675484 572540
rect 674156 572500 674162 572512
rect 675478 572500 675484 572512
rect 675536 572500 675542 572552
rect 43438 571344 43444 571396
rect 43496 571384 43502 571396
rect 62114 571384 62120 571396
rect 43496 571356 62120 571384
rect 43496 571344 43502 571356
rect 62114 571344 62120 571356
rect 62172 571344 62178 571396
rect 669222 571344 669228 571396
rect 669280 571384 669286 571396
rect 675478 571384 675484 571396
rect 669280 571356 675484 571384
rect 669280 571344 669286 571356
rect 675478 571344 675484 571356
rect 675536 571344 675542 571396
rect 42058 570936 42064 570988
rect 42116 570976 42122 570988
rect 42610 570976 42616 570988
rect 42116 570948 42616 570976
rect 42116 570936 42122 570948
rect 42610 570936 42616 570948
rect 42668 570936 42674 570988
rect 671706 570800 671712 570852
rect 671764 570840 671770 570852
rect 675478 570840 675484 570852
rect 671764 570812 675484 570840
rect 671764 570800 671770 570812
rect 675478 570800 675484 570812
rect 675536 570800 675542 570852
rect 666094 570120 666100 570172
rect 666152 570160 666158 570172
rect 675478 570160 675484 570172
rect 666152 570132 675484 570160
rect 666152 570120 666158 570132
rect 675478 570120 675484 570132
rect 675536 570120 675542 570172
rect 675846 570052 675852 570104
rect 675904 570092 675910 570104
rect 683114 570092 683120 570104
rect 675904 570064 683120 570092
rect 675904 570052 675910 570064
rect 683114 570052 683120 570064
rect 683172 570052 683178 570104
rect 670786 569576 670792 569628
rect 670844 569616 670850 569628
rect 675478 569616 675484 569628
rect 670844 569588 675484 569616
rect 670844 569576 670850 569588
rect 675478 569576 675484 569588
rect 675536 569576 675542 569628
rect 671338 565224 671344 565276
rect 671396 565224 671402 565276
rect 671154 565060 671160 565072
rect 670988 565032 671160 565060
rect 670988 564788 671016 565032
rect 671154 565020 671160 565032
rect 671212 565020 671218 565072
rect 671154 564884 671160 564936
rect 671212 564924 671218 564936
rect 671356 564924 671384 565224
rect 671212 564896 671384 564924
rect 671212 564884 671218 564896
rect 671338 564788 671344 564800
rect 670988 564760 671344 564788
rect 671338 564748 671344 564760
rect 671396 564748 671402 564800
rect 665082 564408 665088 564460
rect 665140 564448 665146 564460
rect 675294 564448 675300 564460
rect 665140 564420 675300 564448
rect 665140 564408 665146 564420
rect 675294 564408 675300 564420
rect 675352 564408 675358 564460
rect 651650 563048 651656 563100
rect 651708 563088 651714 563100
rect 658918 563088 658924 563100
rect 651708 563060 658924 563088
rect 651708 563048 651714 563060
rect 658918 563048 658924 563060
rect 658976 563048 658982 563100
rect 673730 561688 673736 561740
rect 673788 561728 673794 561740
rect 675110 561728 675116 561740
rect 673788 561700 675116 561728
rect 673788 561688 673794 561700
rect 675110 561688 675116 561700
rect 675168 561688 675174 561740
rect 666186 560328 666192 560380
rect 666244 560368 666250 560380
rect 675294 560368 675300 560380
rect 666244 560340 675300 560368
rect 666244 560328 666250 560340
rect 675294 560328 675300 560340
rect 675352 560328 675358 560380
rect 41690 557784 41696 557796
rect 41386 557756 41696 557784
rect 41386 557728 41414 557756
rect 41690 557744 41696 557756
rect 41748 557744 41754 557796
rect 42058 557744 42064 557796
rect 42116 557784 42122 557796
rect 49142 557784 49148 557796
rect 42116 557756 49148 557784
rect 42116 557744 42122 557756
rect 49142 557744 49148 557756
rect 49200 557744 49206 557796
rect 41322 557676 41328 557728
rect 41380 557688 41414 557728
rect 41380 557676 41386 557688
rect 674098 557676 674104 557728
rect 674156 557716 674162 557728
rect 675110 557716 675116 557728
rect 674156 557688 675116 557716
rect 674156 557676 674162 557688
rect 675110 557676 675116 557688
rect 675168 557676 675174 557728
rect 43806 557540 43812 557592
rect 43864 557580 43870 557592
rect 51902 557580 51908 557592
rect 43864 557552 51908 557580
rect 43864 557540 43870 557552
rect 51902 557540 51908 557552
rect 51960 557540 51966 557592
rect 54846 557540 54852 557592
rect 54904 557580 54910 557592
rect 62114 557580 62120 557592
rect 54904 557552 62120 557580
rect 54904 557540 54910 557552
rect 62114 557540 62120 557552
rect 62172 557540 62178 557592
rect 666094 557540 666100 557592
rect 666152 557580 666158 557592
rect 675294 557580 675300 557592
rect 666152 557552 675300 557580
rect 666152 557540 666158 557552
rect 675294 557540 675300 557552
rect 675352 557540 675358 557592
rect 42058 555364 42064 555416
rect 42116 555404 42122 555416
rect 43162 555404 43168 555416
rect 42116 555376 43168 555404
rect 42116 555364 42122 555376
rect 43162 555364 43168 555376
rect 43220 555364 43226 555416
rect 41138 555296 41144 555348
rect 41196 555296 41202 555348
rect 41156 555200 41184 555296
rect 41156 555172 41276 555200
rect 41248 555132 41276 555172
rect 41690 555132 41696 555144
rect 41248 555104 41696 555132
rect 41690 555092 41696 555104
rect 41748 555092 41754 555144
rect 41046 554888 41052 554940
rect 41104 554928 41110 554940
rect 41690 554928 41696 554940
rect 41104 554900 41696 554928
rect 41104 554888 41110 554900
rect 41690 554888 41696 554900
rect 41748 554888 41754 554940
rect 42058 554888 42064 554940
rect 42116 554928 42122 554940
rect 42978 554928 42984 554940
rect 42116 554900 42984 554928
rect 42116 554888 42122 554900
rect 42978 554888 42984 554900
rect 43036 554888 43042 554940
rect 40586 554752 40592 554804
rect 40644 554792 40650 554804
rect 41690 554792 41696 554804
rect 40644 554764 41696 554792
rect 40644 554752 40650 554764
rect 41690 554752 41696 554764
rect 41748 554752 41754 554804
rect 42058 554752 42064 554804
rect 42116 554792 42122 554804
rect 44266 554792 44272 554804
rect 42116 554764 44272 554792
rect 42116 554752 42122 554764
rect 44266 554752 44272 554764
rect 44324 554752 44330 554804
rect 669774 554752 669780 554804
rect 669832 554792 669838 554804
rect 675294 554792 675300 554804
rect 669832 554764 675300 554792
rect 669832 554752 669838 554764
rect 675294 554752 675300 554764
rect 675352 554752 675358 554804
rect 674466 554276 674472 554328
rect 674524 554316 674530 554328
rect 675110 554316 675116 554328
rect 674524 554288 675116 554316
rect 674524 554276 674530 554288
rect 675110 554276 675116 554288
rect 675168 554276 675174 554328
rect 658918 554004 658924 554056
rect 658976 554044 658982 554056
rect 675110 554044 675116 554056
rect 658976 554016 675116 554044
rect 658976 554004 658982 554016
rect 675110 554004 675116 554016
rect 675168 554004 675174 554056
rect 671890 553460 671896 553512
rect 671948 553500 671954 553512
rect 675294 553500 675300 553512
rect 671948 553472 675300 553500
rect 671948 553460 671954 553472
rect 675294 553460 675300 553472
rect 675352 553460 675358 553512
rect 651650 550604 651656 550656
rect 651708 550644 651714 550656
rect 659286 550644 659292 550656
rect 651708 550616 659292 550644
rect 651708 550604 651714 550616
rect 659286 550604 659292 550616
rect 659344 550604 659350 550656
rect 664254 550604 664260 550656
rect 664312 550644 664318 550656
rect 675018 550644 675024 550656
rect 664312 550616 675024 550644
rect 664312 550604 664318 550616
rect 675018 550604 675024 550616
rect 675076 550604 675082 550656
rect 40034 550400 40040 550452
rect 40092 550440 40098 550452
rect 41690 550440 41696 550452
rect 40092 550412 41696 550440
rect 40092 550400 40098 550412
rect 41690 550400 41696 550412
rect 41748 550400 41754 550452
rect 42058 550400 42064 550452
rect 42116 550440 42122 550452
rect 42518 550440 42524 550452
rect 42116 550412 42524 550440
rect 42116 550400 42122 550412
rect 42518 550400 42524 550412
rect 42576 550400 42582 550452
rect 45554 548632 45560 548684
rect 45612 548632 45618 548684
rect 45572 548548 45600 548632
rect 45554 548496 45560 548548
rect 45612 548496 45618 548548
rect 42334 547884 42340 547936
rect 42392 547924 42398 547936
rect 53282 547924 53288 547936
rect 42392 547896 53288 547924
rect 42392 547884 42398 547896
rect 53282 547884 53288 547896
rect 53340 547884 53346 547936
rect 31754 547408 31760 547460
rect 31812 547448 31818 547460
rect 38562 547448 38568 547460
rect 31812 547420 38568 547448
rect 31812 547408 31818 547420
rect 38562 547408 38568 547420
rect 38620 547408 38626 547460
rect 675938 547272 675944 547324
rect 675996 547312 676002 547324
rect 678238 547312 678244 547324
rect 675996 547284 678244 547312
rect 675996 547272 676002 547284
rect 678238 547272 678244 547284
rect 678296 547272 678302 547324
rect 676122 547136 676128 547188
rect 676180 547176 676186 547188
rect 683390 547176 683396 547188
rect 676180 547148 683396 547176
rect 676180 547136 676186 547148
rect 683390 547136 683396 547148
rect 683448 547136 683454 547188
rect 43438 546592 43444 546644
rect 43496 546632 43502 546644
rect 49142 546632 49148 546644
rect 43496 546604 49148 546632
rect 43496 546592 43502 546604
rect 49142 546592 49148 546604
rect 49200 546592 49206 546644
rect 675938 545708 675944 545760
rect 675996 545748 676002 545760
rect 683206 545748 683212 545760
rect 675996 545720 683212 545748
rect 675996 545708 676002 545720
rect 683206 545708 683212 545720
rect 683264 545708 683270 545760
rect 43438 545096 43444 545148
rect 43496 545136 43502 545148
rect 62114 545136 62120 545148
rect 43496 545108 62120 545136
rect 43496 545096 43502 545108
rect 62114 545096 62120 545108
rect 62172 545096 62178 545148
rect 29638 544348 29644 544400
rect 29696 544388 29702 544400
rect 41506 544388 41512 544400
rect 29696 544360 41512 544388
rect 29696 544348 29702 544360
rect 41506 544348 41512 544360
rect 41564 544348 41570 544400
rect 38562 542308 38568 542360
rect 38620 542348 38626 542360
rect 41690 542348 41696 542360
rect 38620 542320 41696 542348
rect 38620 542308 38626 542320
rect 41690 542308 41696 542320
rect 41748 542308 41754 542360
rect 652018 536800 652024 536852
rect 652076 536840 652082 536852
rect 660482 536840 660488 536852
rect 652076 536812 660488 536840
rect 652076 536800 652082 536812
rect 660482 536800 660488 536812
rect 660540 536800 660546 536852
rect 42242 536256 42248 536308
rect 42300 536296 42306 536308
rect 45370 536296 45376 536308
rect 42300 536268 45376 536296
rect 42300 536256 42306 536268
rect 45370 536256 45376 536268
rect 45428 536256 45434 536308
rect 664806 535644 664812 535696
rect 664864 535684 664870 535696
rect 675478 535684 675484 535696
rect 664864 535656 675484 535684
rect 664864 535644 664870 535656
rect 675478 535644 675484 535656
rect 675536 535644 675542 535696
rect 661678 535440 661684 535492
rect 661736 535480 661742 535492
rect 675478 535480 675484 535492
rect 661736 535452 675484 535480
rect 661736 535440 661742 535452
rect 675478 535440 675484 535452
rect 675536 535440 675542 535492
rect 672626 534556 672632 534608
rect 672684 534596 672690 534608
rect 674742 534596 674748 534608
rect 672684 534568 674748 534596
rect 672684 534556 672690 534568
rect 674742 534556 674748 534568
rect 674800 534556 674806 534608
rect 675478 534556 675484 534608
rect 675536 534556 675542 534608
rect 671338 534352 671344 534404
rect 671396 534392 671402 534404
rect 675496 534392 675524 534556
rect 671396 534364 675524 534392
rect 671396 534352 671402 534364
rect 659102 534216 659108 534268
rect 659160 534256 659166 534268
rect 674558 534256 674564 534268
rect 659160 534228 674564 534256
rect 659160 534216 659166 534228
rect 674558 534216 674564 534228
rect 674616 534216 674622 534268
rect 42426 534148 42432 534200
rect 42484 534188 42490 534200
rect 45738 534188 45744 534200
rect 42484 534160 45744 534188
rect 42484 534148 42490 534160
rect 45738 534148 45744 534160
rect 45796 534148 45802 534200
rect 672626 534080 672632 534132
rect 672684 534120 672690 534132
rect 675478 534120 675484 534132
rect 672684 534092 675484 534120
rect 672684 534080 672690 534092
rect 675478 534080 675484 534092
rect 675536 534080 675542 534132
rect 42610 533944 42616 533996
rect 42668 533984 42674 533996
rect 43990 533984 43996 533996
rect 42668 533956 43996 533984
rect 42668 533944 42674 533956
rect 43990 533944 43996 533956
rect 44048 533944 44054 533996
rect 671522 532856 671528 532908
rect 671580 532896 671586 532908
rect 675478 532896 675484 532908
rect 671580 532868 675484 532896
rect 671580 532856 671586 532868
rect 675478 532856 675484 532868
rect 675536 532856 675542 532908
rect 673546 531768 673552 531820
rect 673604 531808 673610 531820
rect 675478 531808 675484 531820
rect 673604 531780 675484 531808
rect 673604 531768 673610 531780
rect 675478 531768 675484 531780
rect 675536 531768 675542 531820
rect 672442 531564 672448 531616
rect 672500 531604 672506 531616
rect 675478 531604 675484 531616
rect 672500 531576 675484 531604
rect 672500 531564 672506 531576
rect 675478 531564 675484 531576
rect 675536 531564 675542 531616
rect 671154 531428 671160 531480
rect 671212 531468 671218 531480
rect 673546 531468 673552 531480
rect 671212 531440 673552 531468
rect 671212 531428 671218 531440
rect 673546 531428 673552 531440
rect 673604 531428 673610 531480
rect 45186 531332 45192 531344
rect 42812 531304 45192 531332
rect 42242 530884 42248 530936
rect 42300 530924 42306 530936
rect 42610 530924 42616 530936
rect 42300 530896 42616 530924
rect 42300 530884 42306 530896
rect 42610 530884 42616 530896
rect 42668 530884 42674 530936
rect 42610 530748 42616 530800
rect 42668 530788 42674 530800
rect 42812 530788 42840 531304
rect 45186 531292 45192 531304
rect 45244 531292 45250 531344
rect 672534 531292 672540 531344
rect 672592 531332 672598 531344
rect 674742 531332 674748 531344
rect 672592 531304 674748 531332
rect 672592 531292 672598 531304
rect 674742 531292 674748 531304
rect 674800 531292 674806 531344
rect 42668 530760 42840 530788
rect 42668 530748 42674 530760
rect 42242 530272 42248 530324
rect 42300 530312 42306 530324
rect 42610 530312 42616 530324
rect 42300 530284 42616 530312
rect 42300 530272 42306 530284
rect 42610 530272 42616 530284
rect 42668 530272 42674 530324
rect 673086 530068 673092 530120
rect 673144 530108 673150 530120
rect 675478 530108 675484 530120
rect 673144 530080 675484 530108
rect 673144 530068 673150 530080
rect 675478 530068 675484 530080
rect 675536 530068 675542 530120
rect 665634 529932 665640 529984
rect 665692 529972 665698 529984
rect 675478 529972 675484 529984
rect 665692 529944 675484 529972
rect 665692 529932 665698 529944
rect 675478 529932 675484 529944
rect 675536 529932 675542 529984
rect 669038 529320 669044 529372
rect 669096 529360 669102 529372
rect 675478 529360 675484 529372
rect 669096 529332 675484 529360
rect 669096 529320 669102 529332
rect 675478 529320 675484 529332
rect 675536 529320 675542 529372
rect 42426 529048 42432 529100
rect 42484 529088 42490 529100
rect 43806 529088 43812 529100
rect 42484 529060 43812 529088
rect 42484 529048 42490 529060
rect 43806 529048 43812 529060
rect 43864 529048 43870 529100
rect 666462 528572 666468 528624
rect 666520 528612 666526 528624
rect 675478 528612 675484 528624
rect 666520 528584 675484 528612
rect 666520 528572 666526 528584
rect 675478 528572 675484 528584
rect 675536 528572 675542 528624
rect 673914 528300 673920 528352
rect 673972 528340 673978 528352
rect 675478 528340 675484 528352
rect 673972 528312 675484 528340
rect 673972 528300 673978 528312
rect 675478 528300 675484 528312
rect 675536 528300 675542 528352
rect 674098 528096 674104 528148
rect 674156 528096 674162 528148
rect 674116 527944 674144 528096
rect 674098 527892 674104 527944
rect 674156 527892 674162 527944
rect 673914 527620 673920 527672
rect 673972 527660 673978 527672
rect 675478 527660 675484 527672
rect 673972 527632 675484 527660
rect 673972 527620 673978 527632
rect 675478 527620 675484 527632
rect 675536 527620 675542 527672
rect 668854 525784 668860 525836
rect 668912 525824 668918 525836
rect 675478 525824 675484 525836
rect 668912 525796 675484 525824
rect 668912 525784 668918 525796
rect 675478 525784 675484 525796
rect 675536 525784 675542 525836
rect 678238 525716 678244 525768
rect 678296 525756 678302 525768
rect 683114 525756 683120 525768
rect 678296 525728 683120 525756
rect 678296 525716 678302 525728
rect 683114 525716 683120 525728
rect 683172 525716 683178 525768
rect 671246 524424 671252 524476
rect 671304 524464 671310 524476
rect 675478 524464 675484 524476
rect 671304 524436 675484 524464
rect 671304 524424 671310 524436
rect 675478 524424 675484 524436
rect 675536 524424 675542 524476
rect 42518 523676 42524 523728
rect 42576 523716 42582 523728
rect 62758 523716 62764 523728
rect 42576 523688 62764 523716
rect 42576 523676 42582 523688
rect 62758 523676 62764 523688
rect 62816 523676 62822 523728
rect 651650 522996 651656 523048
rect 651708 523036 651714 523048
rect 661678 523036 661684 523048
rect 651708 523008 661684 523036
rect 651708 522996 651714 523008
rect 661678 522996 661684 523008
rect 661736 522996 661742 523048
rect 42058 518916 42064 518968
rect 42116 518956 42122 518968
rect 62114 518956 62120 518968
rect 42116 518928 62120 518956
rect 42116 518916 42122 518928
rect 62114 518916 62120 518928
rect 62172 518916 62178 518968
rect 651650 510620 651656 510672
rect 651708 510660 651714 510672
rect 659102 510660 659108 510672
rect 651708 510632 659108 510660
rect 651708 510620 651714 510632
rect 659102 510620 659108 510632
rect 659160 510620 659166 510672
rect 52270 506472 52276 506524
rect 52328 506512 52334 506524
rect 62114 506512 62120 506524
rect 52328 506484 62120 506512
rect 52328 506472 52334 506484
rect 62114 506472 62120 506484
rect 62172 506472 62178 506524
rect 676122 503480 676128 503532
rect 676180 503520 676186 503532
rect 679618 503520 679624 503532
rect 676180 503492 679624 503520
rect 676180 503480 676186 503492
rect 679618 503480 679624 503492
rect 679676 503480 679682 503532
rect 651650 496816 651656 496868
rect 651708 496856 651714 496868
rect 661862 496856 661868 496868
rect 651708 496828 661868 496856
rect 651708 496816 651714 496828
rect 661862 496816 661868 496828
rect 661920 496816 661926 496868
rect 43622 491920 43628 491972
rect 43680 491960 43686 491972
rect 62114 491960 62120 491972
rect 43680 491932 62120 491960
rect 43680 491920 43686 491932
rect 62114 491920 62120 491932
rect 62172 491920 62178 491972
rect 664622 491580 664628 491632
rect 664680 491620 664686 491632
rect 675478 491620 675484 491632
rect 664680 491592 675484 491620
rect 664680 491580 664686 491592
rect 675478 491580 675484 491592
rect 675536 491580 675542 491632
rect 663242 491444 663248 491496
rect 663300 491484 663306 491496
rect 674742 491484 674748 491496
rect 663300 491456 674748 491484
rect 663300 491444 663306 491456
rect 674742 491444 674748 491456
rect 674800 491444 674806 491496
rect 660298 491308 660304 491360
rect 660356 491348 660362 491360
rect 675110 491348 675116 491360
rect 660356 491320 675116 491348
rect 660356 491308 660362 491320
rect 675110 491308 675116 491320
rect 675168 491308 675174 491360
rect 672718 490016 672724 490068
rect 672776 490056 672782 490068
rect 675478 490056 675484 490068
rect 672776 490028 675484 490056
rect 672776 490016 672782 490028
rect 675478 490016 675484 490028
rect 675536 490016 675542 490068
rect 672534 487296 672540 487348
rect 672592 487336 672598 487348
rect 675478 487336 675484 487348
rect 672592 487308 675484 487336
rect 672592 487296 672598 487308
rect 675478 487296 675484 487308
rect 675536 487296 675542 487348
rect 666094 485936 666100 485988
rect 666152 485976 666158 485988
rect 675478 485976 675484 485988
rect 666152 485948 675484 485976
rect 666152 485936 666158 485948
rect 675478 485936 675484 485948
rect 675536 485936 675542 485988
rect 665082 485800 665088 485852
rect 665140 485840 665146 485852
rect 675294 485840 675300 485852
rect 665140 485812 675300 485840
rect 665140 485800 665146 485812
rect 675294 485800 675300 485812
rect 675352 485800 675358 485852
rect 673730 485460 673736 485512
rect 673788 485500 673794 485512
rect 674742 485500 674748 485512
rect 673788 485472 674748 485500
rect 673788 485460 673794 485472
rect 674742 485460 674748 485472
rect 674800 485460 674806 485512
rect 664254 484508 664260 484560
rect 664312 484548 664318 484560
rect 675478 484548 675484 484560
rect 664312 484520 675484 484548
rect 664312 484508 664318 484520
rect 675478 484508 675484 484520
rect 675536 484508 675542 484560
rect 651650 484440 651656 484492
rect 651708 484480 651714 484492
rect 651708 484452 654134 484480
rect 651708 484440 651714 484452
rect 654106 484412 654134 484452
rect 664990 484412 664996 484424
rect 654106 484384 664996 484412
rect 664990 484372 664996 484384
rect 665048 484372 665054 484424
rect 669774 483964 669780 484016
rect 669832 484004 669838 484016
rect 675294 484004 675300 484016
rect 669832 483976 675300 484004
rect 669832 483964 669838 483976
rect 675294 483964 675300 483976
rect 675352 483964 675358 484016
rect 672902 483556 672908 483608
rect 672960 483596 672966 483608
rect 675294 483596 675300 483608
rect 672960 483568 675300 483596
rect 672960 483556 672966 483568
rect 675294 483556 675300 483568
rect 675352 483556 675358 483608
rect 666278 483080 666284 483132
rect 666336 483120 666342 483132
rect 675478 483120 675484 483132
rect 666336 483092 675484 483120
rect 666336 483080 666342 483092
rect 675478 483080 675484 483092
rect 675536 483080 675542 483132
rect 671890 482332 671896 482384
rect 671948 482372 671954 482384
rect 675478 482372 675484 482384
rect 671948 482344 675484 482372
rect 671948 482332 671954 482344
rect 675478 482332 675484 482344
rect 675536 482332 675542 482384
rect 673730 481856 673736 481908
rect 673788 481896 673794 481908
rect 675478 481896 675484 481908
rect 673788 481868 675484 481896
rect 673788 481856 673794 481868
rect 675478 481856 675484 481868
rect 675536 481856 675542 481908
rect 671430 480632 671436 480684
rect 671488 480672 671494 480684
rect 675478 480672 675484 480684
rect 671488 480644 675484 480672
rect 671488 480632 671494 480644
rect 675478 480632 675484 480644
rect 675536 480632 675542 480684
rect 47946 480224 47952 480276
rect 48004 480264 48010 480276
rect 62114 480264 62120 480276
rect 48004 480236 62120 480264
rect 48004 480224 48010 480236
rect 62114 480224 62120 480236
rect 62172 480224 62178 480276
rect 668762 474036 668768 474088
rect 668820 474076 668826 474088
rect 671706 474076 671712 474088
rect 668820 474048 671712 474076
rect 668820 474036 668826 474048
rect 671706 474036 671712 474048
rect 671764 474036 671770 474088
rect 651650 470568 651656 470620
rect 651708 470608 651714 470620
rect 663242 470608 663248 470620
rect 651708 470580 663248 470608
rect 651708 470568 651714 470580
rect 663242 470568 663248 470580
rect 663300 470568 663306 470620
rect 49326 466420 49332 466472
rect 49384 466460 49390 466472
rect 62114 466460 62120 466472
rect 49384 466432 62120 466460
rect 49384 466420 49390 466432
rect 62114 466420 62120 466432
rect 62172 466420 62178 466472
rect 651650 456764 651656 456816
rect 651708 456804 651714 456816
rect 663426 456804 663432 456816
rect 651708 456776 663432 456804
rect 651708 456764 651714 456776
rect 663426 456764 663432 456776
rect 663484 456764 663490 456816
rect 46566 446360 46572 446412
rect 46624 446400 46630 446412
rect 62758 446400 62764 446412
rect 46624 446372 62764 446400
rect 46624 446360 46630 446372
rect 62758 446360 62764 446372
rect 62816 446360 62822 446412
rect 651650 444456 651656 444508
rect 651708 444496 651714 444508
rect 651708 444468 654134 444496
rect 651708 444456 651714 444468
rect 654106 444428 654134 444468
rect 660666 444428 660672 444440
rect 654106 444400 660672 444428
rect 660666 444388 660672 444400
rect 660724 444388 660730 444440
rect 43806 433984 43812 434036
rect 43864 434024 43870 434036
rect 62114 434024 62120 434036
rect 43864 433996 62120 434024
rect 43864 433984 43870 433996
rect 62114 433984 62120 433996
rect 62172 433984 62178 434036
rect 652018 430584 652024 430636
rect 652076 430624 652082 430636
rect 658918 430624 658924 430636
rect 652076 430596 658924 430624
rect 652076 430584 652082 430596
rect 658918 430584 658924 430596
rect 658976 430584 658982 430636
rect 41322 429564 41328 429616
rect 41380 429604 41386 429616
rect 41690 429604 41696 429616
rect 41380 429576 41696 429604
rect 41380 429564 41386 429576
rect 41690 429564 41696 429576
rect 41748 429564 41754 429616
rect 41138 429428 41144 429480
rect 41196 429468 41202 429480
rect 41690 429468 41696 429480
rect 41196 429440 41696 429468
rect 41196 429428 41202 429440
rect 41690 429428 41696 429440
rect 41748 429428 41754 429480
rect 42058 429428 42064 429480
rect 42116 429468 42122 429480
rect 43438 429468 43444 429480
rect 42116 429440 43444 429468
rect 42116 429428 42122 429440
rect 43438 429428 43444 429440
rect 43496 429428 43502 429480
rect 41322 429292 41328 429344
rect 41380 429332 41386 429344
rect 41690 429332 41696 429344
rect 41380 429304 41696 429332
rect 41380 429292 41386 429304
rect 41690 429292 41696 429304
rect 41748 429292 41754 429344
rect 42058 429292 42064 429344
rect 42116 429332 42122 429344
rect 43990 429332 43996 429344
rect 42116 429304 43996 429332
rect 42116 429292 42122 429304
rect 43990 429292 43996 429304
rect 44048 429292 44054 429344
rect 40954 429156 40960 429208
rect 41012 429196 41018 429208
rect 41690 429196 41696 429208
rect 41012 429168 41696 429196
rect 41012 429156 41018 429168
rect 41690 429156 41696 429168
rect 41748 429156 41754 429208
rect 42058 429156 42064 429208
rect 42116 429196 42122 429208
rect 44542 429196 44548 429208
rect 42116 429168 44548 429196
rect 42116 429156 42122 429168
rect 44542 429156 44548 429168
rect 44600 429156 44606 429208
rect 56226 427796 56232 427848
rect 56284 427836 56290 427848
rect 62114 427836 62120 427848
rect 56284 427808 62120 427836
rect 56284 427796 56290 427808
rect 62114 427796 62120 427808
rect 62172 427796 62178 427848
rect 41138 426436 41144 426488
rect 41196 426476 41202 426488
rect 41690 426476 41696 426488
rect 41196 426448 41696 426476
rect 41196 426436 41202 426448
rect 41690 426436 41696 426448
rect 41748 426436 41754 426488
rect 42058 426436 42064 426488
rect 42116 426476 42122 426488
rect 44542 426476 44548 426488
rect 42116 426448 44548 426476
rect 42116 426436 42122 426448
rect 44542 426436 44548 426448
rect 44600 426436 44606 426488
rect 45186 419500 45192 419552
rect 45244 419540 45250 419552
rect 51902 419540 51908 419552
rect 45244 419512 51908 419540
rect 45244 419500 45250 419512
rect 51902 419500 51908 419512
rect 51960 419500 51966 419552
rect 42610 418140 42616 418192
rect 42668 418180 42674 418192
rect 54662 418180 54668 418192
rect 42668 418152 54668 418180
rect 42668 418140 42674 418152
rect 54662 418140 54668 418152
rect 54720 418140 54726 418192
rect 651650 416780 651656 416832
rect 651708 416820 651714 416832
rect 660298 416820 660304 416832
rect 651708 416792 660304 416820
rect 651708 416780 651714 416792
rect 660298 416780 660304 416792
rect 660356 416780 660362 416832
rect 45186 415420 45192 415472
rect 45244 415460 45250 415472
rect 62114 415460 62120 415472
rect 45244 415432 62120 415460
rect 45244 415420 45250 415432
rect 62114 415420 62120 415432
rect 62172 415420 62178 415472
rect 42242 409776 42248 409828
rect 42300 409816 42306 409828
rect 43162 409816 43168 409828
rect 42300 409788 43168 409816
rect 42300 409776 42306 409788
rect 43162 409776 43168 409788
rect 43220 409776 43226 409828
rect 42426 408416 42432 408468
rect 42484 408456 42490 408468
rect 54846 408456 54852 408468
rect 42484 408428 54852 408456
rect 42484 408416 42490 408428
rect 54846 408416 54852 408428
rect 54904 408416 54910 408468
rect 42426 408280 42432 408332
rect 42484 408320 42490 408332
rect 44358 408320 44364 408332
rect 42484 408292 44364 408320
rect 42484 408280 42490 408292
rect 44358 408280 44364 408292
rect 44416 408280 44422 408332
rect 42426 407056 42432 407108
rect 42484 407096 42490 407108
rect 45370 407096 45376 407108
rect 42484 407068 45376 407096
rect 42484 407056 42490 407068
rect 45370 407056 45376 407068
rect 45428 407056 45434 407108
rect 651650 404336 651656 404388
rect 651708 404376 651714 404388
rect 664806 404376 664812 404388
rect 651708 404348 664812 404376
rect 651708 404336 651714 404348
rect 664806 404336 664812 404348
rect 664864 404336 664870 404388
rect 42426 404132 42432 404184
rect 42484 404172 42490 404184
rect 45554 404172 45560 404184
rect 42484 404144 45560 404172
rect 42484 404132 42490 404144
rect 45554 404132 45560 404144
rect 45612 404132 45618 404184
rect 667198 403384 667204 403436
rect 667256 403424 667262 403436
rect 675294 403424 675300 403436
rect 667256 403396 675300 403424
rect 667256 403384 667262 403396
rect 675294 403384 675300 403396
rect 675352 403384 675358 403436
rect 659286 403248 659292 403300
rect 659344 403288 659350 403300
rect 659344 403260 668624 403288
rect 659344 403248 659350 403260
rect 660482 403112 660488 403164
rect 660540 403152 660546 403164
rect 667198 403152 667204 403164
rect 660540 403124 667204 403152
rect 660540 403112 660546 403124
rect 667198 403112 667204 403124
rect 667256 403112 667262 403164
rect 668596 403152 668624 403260
rect 675478 403220 675484 403232
rect 669286 403192 675484 403220
rect 669286 403152 669314 403192
rect 675478 403180 675484 403192
rect 675536 403180 675542 403232
rect 668596 403124 669314 403152
rect 661678 402976 661684 403028
rect 661736 403016 661742 403028
rect 675478 403016 675484 403028
rect 661736 402988 675484 403016
rect 661736 402976 661742 402988
rect 675478 402976 675484 402988
rect 675536 402976 675542 403028
rect 42426 402500 42432 402552
rect 42484 402540 42490 402552
rect 43346 402540 43352 402552
rect 42484 402512 43352 402540
rect 42484 402500 42490 402512
rect 43346 402500 43352 402512
rect 43404 402500 43410 402552
rect 50706 401616 50712 401668
rect 50764 401656 50770 401668
rect 62114 401656 62120 401668
rect 50764 401628 62120 401656
rect 50764 401616 50770 401628
rect 62114 401616 62120 401628
rect 62172 401616 62178 401668
rect 673914 401344 673920 401396
rect 673972 401384 673978 401396
rect 675478 401384 675484 401396
rect 673972 401356 675484 401384
rect 673972 401344 673978 401356
rect 675478 401344 675484 401356
rect 675536 401344 675542 401396
rect 672718 400528 672724 400580
rect 672776 400568 672782 400580
rect 675478 400568 675484 400580
rect 672776 400540 675484 400568
rect 672776 400528 672782 400540
rect 675478 400528 675484 400540
rect 675536 400528 675542 400580
rect 673086 399712 673092 399764
rect 673144 399752 673150 399764
rect 675478 399752 675484 399764
rect 673144 399724 675484 399752
rect 673144 399712 673150 399724
rect 675478 399712 675484 399724
rect 675536 399712 675542 399764
rect 42426 397400 42432 397452
rect 42484 397440 42490 397452
rect 46934 397440 46940 397452
rect 42484 397412 46940 397440
rect 42484 397400 42490 397412
rect 46934 397400 46940 397412
rect 46992 397400 46998 397452
rect 671798 396312 671804 396364
rect 671856 396352 671862 396364
rect 675478 396352 675484 396364
rect 671856 396324 675484 396352
rect 671856 396312 671862 396324
rect 675478 396312 675484 396324
rect 675536 396312 675542 396364
rect 672534 396040 672540 396092
rect 672592 396080 672598 396092
rect 675294 396080 675300 396092
rect 672592 396052 675300 396080
rect 672592 396040 672598 396052
rect 675294 396040 675300 396052
rect 675352 396040 675358 396092
rect 673454 394272 673460 394324
rect 673512 394312 673518 394324
rect 675478 394312 675484 394324
rect 673512 394284 675484 394312
rect 673512 394272 673518 394284
rect 675478 394272 675484 394284
rect 675536 394272 675542 394324
rect 672902 393320 672908 393372
rect 672960 393360 672966 393372
rect 675478 393360 675484 393372
rect 672960 393332 675484 393360
rect 672960 393320 672966 393332
rect 675478 393320 675484 393332
rect 675536 393320 675542 393372
rect 671614 391960 671620 392012
rect 671672 392000 671678 392012
rect 675478 392000 675484 392012
rect 671672 391972 675484 392000
rect 671672 391960 671678 391972
rect 675478 391960 675484 391972
rect 675536 391960 675542 392012
rect 651650 390532 651656 390584
rect 651708 390572 651714 390584
rect 663058 390572 663064 390584
rect 651708 390544 663064 390572
rect 651708 390532 651714 390544
rect 663058 390532 663064 390544
rect 663116 390532 663122 390584
rect 48130 389240 48136 389292
rect 48188 389280 48194 389292
rect 62114 389280 62120 389292
rect 48188 389252 62120 389280
rect 48188 389240 48194 389252
rect 62114 389240 62120 389252
rect 62172 389240 62178 389292
rect 35802 387472 35808 387524
rect 35860 387512 35866 387524
rect 39942 387512 39948 387524
rect 35860 387484 39948 387512
rect 35860 387472 35866 387484
rect 39942 387472 39948 387484
rect 40000 387472 40006 387524
rect 35802 386792 35808 386844
rect 35860 386832 35866 386844
rect 40126 386832 40132 386844
rect 35860 386804 40132 386832
rect 35860 386792 35866 386804
rect 40126 386792 40132 386804
rect 40184 386792 40190 386844
rect 35342 386520 35348 386572
rect 35400 386560 35406 386572
rect 40310 386560 40316 386572
rect 35400 386532 40316 386560
rect 35400 386520 35406 386532
rect 40310 386520 40316 386532
rect 40368 386520 40374 386572
rect 42058 386452 42064 386504
rect 42116 386492 42122 386504
rect 49326 386492 49332 386504
rect 42116 386464 49332 386492
rect 42116 386452 42122 386464
rect 49326 386452 49332 386464
rect 49384 386452 49390 386504
rect 35526 386384 35532 386436
rect 35584 386424 35590 386436
rect 41690 386424 41696 386436
rect 35584 386396 41696 386424
rect 35584 386384 35590 386396
rect 41690 386384 41696 386396
rect 41748 386384 41754 386436
rect 35802 385432 35808 385484
rect 35860 385472 35866 385484
rect 39574 385472 39580 385484
rect 35860 385444 39580 385472
rect 35860 385432 35866 385444
rect 39574 385432 39580 385444
rect 39632 385432 39638 385484
rect 41690 385268 41696 385280
rect 41386 385240 41696 385268
rect 35526 385160 35532 385212
rect 35584 385200 35590 385212
rect 41386 385200 41414 385240
rect 41690 385228 41696 385240
rect 41748 385228 41754 385280
rect 42058 385228 42064 385280
rect 42116 385268 42122 385280
rect 42886 385268 42892 385280
rect 42116 385240 42892 385268
rect 42116 385228 42122 385240
rect 42886 385228 42892 385240
rect 42944 385228 42950 385280
rect 35584 385172 41414 385200
rect 35584 385160 35590 385172
rect 35342 385024 35348 385076
rect 35400 385064 35406 385076
rect 41690 385064 41696 385076
rect 35400 385036 41696 385064
rect 35400 385024 35406 385036
rect 41690 385024 41696 385036
rect 41748 385024 41754 385076
rect 42058 385024 42064 385076
rect 42116 385064 42122 385076
rect 43254 385064 43260 385076
rect 42116 385036 43260 385064
rect 42116 385024 42122 385036
rect 43254 385024 43260 385036
rect 43312 385024 43318 385076
rect 35802 384072 35808 384124
rect 35860 384112 35866 384124
rect 39666 384112 39672 384124
rect 35860 384084 39672 384112
rect 35860 384072 35866 384084
rect 39666 384072 39672 384084
rect 39724 384072 39730 384124
rect 42058 383868 42064 383920
rect 42116 383908 42122 383920
rect 44542 383908 44548 383920
rect 42116 383880 44548 383908
rect 42116 383868 42122 383880
rect 44542 383868 44548 383880
rect 44600 383868 44606 383920
rect 35618 383800 35624 383852
rect 35676 383840 35682 383852
rect 41690 383840 41696 383852
rect 35676 383812 41696 383840
rect 35676 383800 35682 383812
rect 41690 383800 41696 383812
rect 41748 383800 41754 383852
rect 35802 383664 35808 383716
rect 35860 383704 35866 383716
rect 41690 383704 41696 383716
rect 35860 383676 41696 383704
rect 35860 383664 35866 383676
rect 41690 383664 41696 383676
rect 41748 383664 41754 383716
rect 42058 383664 42064 383716
rect 42116 383704 42122 383716
rect 44174 383704 44180 383716
rect 42116 383676 44180 383704
rect 42116 383664 42122 383676
rect 44174 383664 44180 383676
rect 44232 383664 44238 383716
rect 35526 382644 35532 382696
rect 35584 382684 35590 382696
rect 40034 382684 40040 382696
rect 35584 382656 40040 382684
rect 35584 382644 35590 382656
rect 40034 382644 40040 382656
rect 40092 382644 40098 382696
rect 35802 382508 35808 382560
rect 35860 382548 35866 382560
rect 41690 382548 41696 382560
rect 35860 382520 41696 382548
rect 35860 382508 35866 382520
rect 41690 382508 41696 382520
rect 41748 382508 41754 382560
rect 35802 382372 35808 382424
rect 35860 382412 35866 382424
rect 40218 382412 40224 382424
rect 35860 382384 40224 382412
rect 35860 382372 35866 382384
rect 40218 382372 40224 382384
rect 40276 382372 40282 382424
rect 671798 382304 671804 382356
rect 671856 382344 671862 382356
rect 675386 382344 675392 382356
rect 671856 382316 675392 382344
rect 671856 382304 671862 382316
rect 675386 382304 675392 382316
rect 675444 382304 675450 382356
rect 35342 382236 35348 382288
rect 35400 382276 35406 382288
rect 41414 382276 41420 382288
rect 35400 382248 41420 382276
rect 35400 382236 35406 382248
rect 41414 382236 41420 382248
rect 41472 382236 41478 382288
rect 674282 382168 674288 382220
rect 674340 382208 674346 382220
rect 675110 382208 675116 382220
rect 674340 382180 675116 382208
rect 674340 382168 674346 382180
rect 675110 382168 675116 382180
rect 675168 382168 675174 382220
rect 35618 381012 35624 381064
rect 35676 381052 35682 381064
rect 40034 381052 40040 381064
rect 35676 381024 40040 381052
rect 35676 381012 35682 381024
rect 40034 381012 40040 381024
rect 40092 381012 40098 381064
rect 35802 380876 35808 380928
rect 35860 380916 35866 380928
rect 39850 380916 39856 380928
rect 35860 380888 39856 380916
rect 35860 380876 35866 380888
rect 39850 380876 39856 380888
rect 39908 380876 39914 380928
rect 35618 379924 35624 379976
rect 35676 379964 35682 379976
rect 41046 379964 41052 379976
rect 35676 379936 41052 379964
rect 35676 379924 35682 379936
rect 41046 379924 41052 379936
rect 41104 379924 41110 379976
rect 35802 379652 35808 379704
rect 35860 379692 35866 379704
rect 39758 379692 39764 379704
rect 35860 379664 39764 379692
rect 35860 379652 35866 379664
rect 39758 379652 39764 379664
rect 39816 379652 39822 379704
rect 35434 379516 35440 379568
rect 35492 379556 35498 379568
rect 41506 379556 41512 379568
rect 35492 379528 41512 379556
rect 35492 379516 35498 379528
rect 41506 379516 41512 379528
rect 41564 379516 41570 379568
rect 35802 378292 35808 378344
rect 35860 378332 35866 378344
rect 39574 378332 39580 378344
rect 35860 378304 39580 378332
rect 35860 378292 35866 378304
rect 39574 378292 39580 378304
rect 39632 378292 39638 378344
rect 651650 378156 651656 378208
rect 651708 378196 651714 378208
rect 661678 378196 661684 378208
rect 651708 378168 661684 378196
rect 651708 378156 651714 378168
rect 661678 378156 661684 378168
rect 661736 378156 661742 378208
rect 673362 377816 673368 377868
rect 673420 377856 673426 377868
rect 675294 377856 675300 377868
rect 673420 377828 675300 377856
rect 673420 377816 673426 377828
rect 675294 377816 675300 377828
rect 675352 377816 675358 377868
rect 35618 377000 35624 377052
rect 35676 377040 35682 377052
rect 35676 377012 38654 377040
rect 35676 377000 35682 377012
rect 38626 376972 38654 377012
rect 41506 376972 41512 376984
rect 38626 376944 41512 376972
rect 41506 376932 41512 376944
rect 41564 376932 41570 376984
rect 42058 376796 42064 376848
rect 42116 376836 42122 376848
rect 42116 376808 51074 376836
rect 42116 376796 42122 376808
rect 35802 376728 35808 376780
rect 35860 376768 35866 376780
rect 41690 376768 41696 376780
rect 35860 376740 41696 376768
rect 35860 376728 35866 376740
rect 41690 376728 41696 376740
rect 41748 376728 41754 376780
rect 51046 376768 51074 376808
rect 53466 376768 53472 376780
rect 51046 376740 53472 376768
rect 53466 376728 53472 376740
rect 53524 376728 53530 376780
rect 672902 376456 672908 376508
rect 672960 376496 672966 376508
rect 675110 376496 675116 376508
rect 672960 376468 675116 376496
rect 672960 376456 672966 376468
rect 675110 376456 675116 376468
rect 675168 376456 675174 376508
rect 28810 375844 28816 375896
rect 28868 375884 28874 375896
rect 33778 375884 33784 375896
rect 28868 375856 33784 375884
rect 28868 375844 28874 375856
rect 33778 375844 33784 375856
rect 33836 375844 33842 375896
rect 35802 375572 35808 375624
rect 35860 375612 35866 375624
rect 41690 375612 41696 375624
rect 35860 375584 41696 375612
rect 35860 375572 35866 375584
rect 41690 375572 41696 375584
rect 41748 375572 41754 375624
rect 42058 375504 42064 375556
rect 42116 375544 42122 375556
rect 52086 375544 52092 375556
rect 42116 375516 52092 375544
rect 42116 375504 42122 375516
rect 52086 375504 52092 375516
rect 52144 375504 52150 375556
rect 49326 375368 49332 375420
rect 49384 375408 49390 375420
rect 62114 375408 62120 375420
rect 49384 375380 62120 375408
rect 49384 375368 49390 375380
rect 62114 375368 62120 375380
rect 62172 375368 62178 375420
rect 674466 375300 674472 375352
rect 674524 375340 674530 375352
rect 675110 375340 675116 375352
rect 674524 375312 675116 375340
rect 674524 375300 674530 375312
rect 675110 375300 675116 375312
rect 675168 375300 675174 375352
rect 33778 373260 33784 373312
rect 33836 373300 33842 373312
rect 41690 373300 41696 373312
rect 33836 373272 41696 373300
rect 33836 373260 33842 373272
rect 41690 373260 41696 373272
rect 41748 373260 41754 373312
rect 32398 371832 32404 371884
rect 32456 371872 32462 371884
rect 41690 371872 41696 371884
rect 32456 371844 41696 371872
rect 32456 371832 32462 371844
rect 41690 371832 41696 371844
rect 41748 371832 41754 371884
rect 42058 371696 42064 371748
rect 42116 371736 42122 371748
rect 42610 371736 42616 371748
rect 42116 371708 42616 371736
rect 42116 371696 42122 371708
rect 42610 371696 42616 371708
rect 42668 371696 42674 371748
rect 651650 364352 651656 364404
rect 651708 364392 651714 364404
rect 664622 364392 664628 364404
rect 651708 364364 664628 364392
rect 651708 364352 651714 364364
rect 664622 364352 664628 364364
rect 664680 364352 664686 364404
rect 42242 364284 42248 364336
rect 42300 364324 42306 364336
rect 52270 364324 52276 364336
rect 42300 364296 52276 364324
rect 42300 364284 42306 364296
rect 52270 364284 52276 364296
rect 52328 364284 52334 364336
rect 42334 364080 42340 364132
rect 42392 364120 42398 364132
rect 43622 364120 43628 364132
rect 42392 364092 43628 364120
rect 42392 364080 42398 364092
rect 43622 364080 43628 364092
rect 43680 364080 43686 364132
rect 42426 360136 42432 360188
rect 42484 360176 42490 360188
rect 44542 360176 44548 360188
rect 42484 360148 44548 360176
rect 42484 360136 42490 360148
rect 44542 360136 44548 360148
rect 44600 360136 44606 360188
rect 42150 359932 42156 359984
rect 42208 359972 42214 359984
rect 43438 359972 43444 359984
rect 42208 359944 43444 359972
rect 42208 359932 42214 359944
rect 43438 359932 43444 359944
rect 43496 359932 43502 359984
rect 664990 357688 664996 357740
rect 665048 357728 665054 357740
rect 675478 357728 675484 357740
rect 665048 357700 675484 357728
rect 665048 357688 665054 357700
rect 675478 357688 675484 357700
rect 675536 357688 675542 357740
rect 661862 357552 661868 357604
rect 661920 357592 661926 357604
rect 675294 357592 675300 357604
rect 661920 357564 675300 357592
rect 661920 357552 661926 357564
rect 675294 357552 675300 357564
rect 675352 357552 675358 357604
rect 659102 357416 659108 357468
rect 659160 357456 659166 357468
rect 675110 357456 675116 357468
rect 659160 357428 675116 357456
rect 659160 357416 659166 357428
rect 675110 357416 675116 357428
rect 675168 357416 675174 357468
rect 673914 357280 673920 357332
rect 673972 357320 673978 357332
rect 674742 357320 674748 357332
rect 673972 357292 674748 357320
rect 673972 357280 673978 357292
rect 674742 357280 674748 357292
rect 674800 357280 674806 357332
rect 673914 357008 673920 357060
rect 673972 357048 673978 357060
rect 675478 357048 675484 357060
rect 673972 357020 675484 357048
rect 673972 357008 673978 357020
rect 675478 357008 675484 357020
rect 675536 357008 675542 357060
rect 42426 355988 42432 356040
rect 42484 356028 42490 356040
rect 45370 356028 45376 356040
rect 42484 356000 45376 356028
rect 42484 355988 42490 356000
rect 45370 355988 45376 356000
rect 45428 355988 45434 356040
rect 672718 355172 672724 355224
rect 672776 355212 672782 355224
rect 675478 355212 675484 355224
rect 672776 355184 675484 355212
rect 672776 355172 672782 355184
rect 675478 355172 675484 355184
rect 675536 355172 675542 355224
rect 673086 354832 673092 354884
rect 673144 354872 673150 354884
rect 675478 354872 675484 354884
rect 673144 354844 675484 354872
rect 673144 354832 673150 354844
rect 675478 354832 675484 354844
rect 675536 354832 675542 354884
rect 673086 354696 673092 354748
rect 673144 354736 673150 354748
rect 675294 354736 675300 354748
rect 673144 354708 675300 354736
rect 673144 354696 673150 354708
rect 675294 354696 675300 354708
rect 675352 354696 675358 354748
rect 673362 353540 673368 353592
rect 673420 353580 673426 353592
rect 675478 353580 675484 353592
rect 673420 353552 675484 353580
rect 673420 353540 673426 353552
rect 675478 353540 675484 353552
rect 675536 353540 675542 353592
rect 672810 353404 672816 353456
rect 672868 353444 672874 353456
rect 675110 353444 675116 353456
rect 672868 353416 675116 353444
rect 672868 353404 672874 353416
rect 675110 353404 675116 353416
rect 675168 353404 675174 353456
rect 669774 353268 669780 353320
rect 669832 353308 669838 353320
rect 675294 353308 675300 353320
rect 669832 353280 675300 353308
rect 669832 353268 669838 353280
rect 675294 353268 675300 353280
rect 675352 353268 675358 353320
rect 671890 351908 671896 351960
rect 671948 351948 671954 351960
rect 675478 351948 675484 351960
rect 671948 351920 675484 351948
rect 671948 351908 671954 351920
rect 675478 351908 675484 351920
rect 675536 351908 675542 351960
rect 669590 350684 669596 350736
rect 669648 350724 669654 350736
rect 675478 350724 675484 350736
rect 669648 350696 675484 350724
rect 669648 350684 669654 350696
rect 675478 350684 675484 350696
rect 675536 350684 675542 350736
rect 651650 350548 651656 350600
rect 651708 350588 651714 350600
rect 661862 350588 661868 350600
rect 651708 350560 661868 350588
rect 651708 350548 651714 350560
rect 661862 350548 661868 350560
rect 661920 350548 661926 350600
rect 671798 350548 671804 350600
rect 671856 350588 671862 350600
rect 675294 350588 675300 350600
rect 671856 350560 675300 350588
rect 671856 350548 671862 350560
rect 675294 350548 675300 350560
rect 675352 350548 675358 350600
rect 673546 349256 673552 349308
rect 673604 349296 673610 349308
rect 675478 349296 675484 349308
rect 673604 349268 675484 349296
rect 673604 349256 673610 349268
rect 675478 349256 675484 349268
rect 675536 349256 675542 349308
rect 672626 348848 672632 348900
rect 672684 348888 672690 348900
rect 675478 348888 675484 348900
rect 672684 348860 675484 348888
rect 672684 348848 672690 348860
rect 675478 348848 675484 348860
rect 675536 348848 675542 348900
rect 45370 347012 45376 347064
rect 45428 347052 45434 347064
rect 62942 347052 62948 347064
rect 45428 347024 62948 347052
rect 45428 347012 45434 347024
rect 62942 347012 62948 347024
rect 63000 347012 63006 347064
rect 675846 346400 675852 346452
rect 675904 346440 675910 346452
rect 683114 346440 683120 346452
rect 675904 346412 683120 346440
rect 675904 346400 675910 346412
rect 683114 346400 683120 346412
rect 683172 346400 683178 346452
rect 671706 344972 671712 345024
rect 671764 345012 671770 345024
rect 675478 345012 675484 345024
rect 671764 344984 675484 345012
rect 671764 344972 671770 344984
rect 675478 344972 675484 344984
rect 675536 344972 675542 345024
rect 35802 344020 35808 344072
rect 35860 344060 35866 344072
rect 39574 344060 39580 344072
rect 35860 344032 39580 344060
rect 35860 344020 35866 344032
rect 39574 344020 39580 344032
rect 39632 344020 39638 344072
rect 40402 343856 40408 343868
rect 36004 343828 40408 343856
rect 35618 343748 35624 343800
rect 35676 343788 35682 343800
rect 36004 343788 36032 343828
rect 40402 343816 40408 343828
rect 40460 343816 40466 343868
rect 35676 343760 36032 343788
rect 35676 343748 35682 343760
rect 35342 343612 35348 343664
rect 35400 343652 35406 343664
rect 41690 343652 41696 343664
rect 35400 343624 41696 343652
rect 35400 343612 35406 343624
rect 41690 343612 41696 343624
rect 41748 343612 41754 343664
rect 42058 343612 42064 343664
rect 42116 343652 42122 343664
rect 56226 343652 56232 343664
rect 42116 343624 56232 343652
rect 42116 343612 42122 343624
rect 56226 343612 56232 343624
rect 56284 343612 56290 343664
rect 35802 342660 35808 342712
rect 35860 342700 35866 342712
rect 39942 342700 39948 342712
rect 35860 342672 39948 342700
rect 35860 342660 35866 342672
rect 39942 342660 39948 342672
rect 40000 342660 40006 342712
rect 39574 342496 39580 342508
rect 36004 342468 39580 342496
rect 35342 342388 35348 342440
rect 35400 342428 35406 342440
rect 36004 342428 36032 342468
rect 39574 342456 39580 342468
rect 39632 342456 39638 342508
rect 35400 342400 36032 342428
rect 35400 342388 35406 342400
rect 35526 342252 35532 342304
rect 35584 342292 35590 342304
rect 40310 342292 40316 342304
rect 35584 342264 40316 342292
rect 35584 342252 35590 342264
rect 40310 342252 40316 342264
rect 40368 342252 40374 342304
rect 35802 341436 35808 341488
rect 35860 341476 35866 341488
rect 39758 341476 39764 341488
rect 35860 341448 39764 341476
rect 35860 341436 35866 341448
rect 39758 341436 39764 341448
rect 39816 341436 39822 341488
rect 40310 341272 40316 341284
rect 36004 341244 40316 341272
rect 35618 341164 35624 341216
rect 35676 341204 35682 341216
rect 36004 341204 36032 341244
rect 40310 341232 40316 341244
rect 40368 341232 40374 341284
rect 35676 341176 36032 341204
rect 35676 341164 35682 341176
rect 35618 341028 35624 341080
rect 35676 341068 35682 341080
rect 41690 341068 41696 341080
rect 35676 341040 41696 341068
rect 35676 341028 35682 341040
rect 41690 341028 41696 341040
rect 41748 341028 41754 341080
rect 42058 341028 42064 341080
rect 42116 341068 42122 341080
rect 45186 341068 45192 341080
rect 42116 341040 45192 341068
rect 42116 341028 42122 341040
rect 45186 341028 45192 341040
rect 45244 341028 45250 341080
rect 35802 340892 35808 340944
rect 35860 340932 35866 340944
rect 41690 340932 41696 340944
rect 35860 340904 41696 340932
rect 35860 340892 35866 340904
rect 41690 340892 41696 340904
rect 41748 340892 41754 340944
rect 42058 340892 42064 340944
rect 42116 340932 42122 340944
rect 44174 340932 44180 340944
rect 42116 340904 44180 340932
rect 42116 340892 42122 340904
rect 44174 340892 44180 340904
rect 44232 340892 44238 340944
rect 673362 340688 673368 340740
rect 673420 340728 673426 340740
rect 675110 340728 675116 340740
rect 673420 340700 675116 340728
rect 673420 340688 673426 340700
rect 675110 340688 675116 340700
rect 675168 340688 675174 340740
rect 35618 339600 35624 339652
rect 35676 339640 35682 339652
rect 39574 339640 39580 339652
rect 35676 339612 39580 339640
rect 35676 339600 35682 339612
rect 39574 339600 39580 339612
rect 39632 339600 39638 339652
rect 35802 338308 35808 338360
rect 35860 338348 35866 338360
rect 41506 338348 41512 338360
rect 35860 338320 41512 338348
rect 35860 338308 35866 338320
rect 41506 338308 41512 338320
rect 41564 338308 41570 338360
rect 35618 338104 35624 338156
rect 35676 338144 35682 338156
rect 41690 338144 41696 338156
rect 35676 338116 41696 338144
rect 35676 338104 35682 338116
rect 41690 338104 41696 338116
rect 41748 338104 41754 338156
rect 42058 338104 42064 338156
rect 42116 338144 42122 338156
rect 47210 338144 47216 338156
rect 42116 338116 47216 338144
rect 42116 338104 42122 338116
rect 47210 338104 47216 338116
rect 47268 338104 47274 338156
rect 651650 338104 651656 338156
rect 651708 338144 651714 338156
rect 667106 338144 667112 338156
rect 651708 338116 667112 338144
rect 651708 338104 651714 338116
rect 667106 338104 667112 338116
rect 667164 338104 667170 338156
rect 673270 337968 673276 338020
rect 673328 338008 673334 338020
rect 675110 338008 675116 338020
rect 673328 337980 675116 338008
rect 673328 337968 673334 337980
rect 675110 337968 675116 337980
rect 675168 337968 675174 338020
rect 35802 337152 35808 337204
rect 35860 337192 35866 337204
rect 40034 337192 40040 337204
rect 35860 337164 40040 337192
rect 35860 337152 35866 337164
rect 40034 337152 40040 337164
rect 40092 337152 40098 337204
rect 41690 336988 41696 337000
rect 41386 336960 41696 336988
rect 35526 336880 35532 336932
rect 35584 336920 35590 336932
rect 41386 336920 41414 336960
rect 41690 336948 41696 336960
rect 41748 336948 41754 337000
rect 42058 336948 42064 337000
rect 42116 336988 42122 337000
rect 43070 336988 43076 337000
rect 42116 336960 43076 336988
rect 42116 336948 42122 336960
rect 43070 336948 43076 336960
rect 43128 336948 43134 337000
rect 35584 336892 41414 336920
rect 35584 336880 35590 336892
rect 35802 336744 35808 336796
rect 35860 336784 35866 336796
rect 41690 336784 41696 336796
rect 35860 336756 41696 336784
rect 35860 336744 35866 336756
rect 41690 336744 41696 336756
rect 41748 336744 41754 336796
rect 42058 336744 42064 336796
rect 42116 336784 42122 336796
rect 43806 336784 43812 336796
rect 42116 336756 43812 336784
rect 42116 336744 42122 336756
rect 43806 336744 43812 336756
rect 43864 336744 43870 336796
rect 46750 336744 46756 336796
rect 46808 336784 46814 336796
rect 62114 336784 62120 336796
rect 46808 336756 62120 336784
rect 46808 336744 46814 336756
rect 62114 336744 62120 336756
rect 62172 336744 62178 336796
rect 674466 336676 674472 336728
rect 674524 336716 674530 336728
rect 675110 336716 675116 336728
rect 674524 336688 675116 336716
rect 674524 336676 674530 336688
rect 675110 336676 675116 336688
rect 675168 336676 675174 336728
rect 35618 335588 35624 335640
rect 35676 335628 35682 335640
rect 40310 335628 40316 335640
rect 35676 335600 40316 335628
rect 35676 335588 35682 335600
rect 40310 335588 40316 335600
rect 40368 335588 40374 335640
rect 669590 335588 669596 335640
rect 669648 335628 669654 335640
rect 674466 335628 674472 335640
rect 669648 335600 674472 335628
rect 669648 335588 669654 335600
rect 674466 335588 674472 335600
rect 674524 335588 674530 335640
rect 673546 335452 673552 335504
rect 673604 335492 673610 335504
rect 675110 335492 675116 335504
rect 673604 335464 675116 335492
rect 673604 335452 673610 335464
rect 675110 335452 675116 335464
rect 675168 335452 675174 335504
rect 35802 335316 35808 335368
rect 35860 335356 35866 335368
rect 39666 335356 39672 335368
rect 35860 335328 39672 335356
rect 35860 335316 35866 335328
rect 39666 335316 39672 335328
rect 39724 335316 39730 335368
rect 674466 335112 674472 335164
rect 674524 335152 674530 335164
rect 674834 335152 674840 335164
rect 674524 335124 674840 335152
rect 674524 335112 674530 335124
rect 674834 335112 674840 335124
rect 674892 335112 674898 335164
rect 35802 334364 35808 334416
rect 35860 334404 35866 334416
rect 40310 334404 40316 334416
rect 35860 334376 40316 334404
rect 35860 334364 35866 334376
rect 40310 334364 40316 334376
rect 40368 334364 40374 334416
rect 36004 334172 38654 334200
rect 35434 334092 35440 334144
rect 35492 334132 35498 334144
rect 36004 334132 36032 334172
rect 35492 334104 36032 334132
rect 38626 334132 38654 334172
rect 39574 334132 39580 334144
rect 38626 334104 39580 334132
rect 35492 334092 35498 334104
rect 39574 334092 39580 334104
rect 39632 334092 39638 334144
rect 42058 334092 42064 334144
rect 42116 334132 42122 334144
rect 42116 334104 51074 334132
rect 42116 334092 42122 334104
rect 35618 333956 35624 334008
rect 35676 333996 35682 334008
rect 41690 333996 41696 334008
rect 35676 333968 41696 333996
rect 35676 333956 35682 333968
rect 41690 333956 41696 333968
rect 41748 333956 41754 334008
rect 51046 333996 51074 334104
rect 54846 333996 54852 334008
rect 51046 333968 54852 333996
rect 54846 333956 54852 333968
rect 54904 333956 54910 334008
rect 671890 333888 671896 333940
rect 671948 333928 671954 333940
rect 675294 333928 675300 333940
rect 671948 333900 675300 333928
rect 671948 333888 671954 333900
rect 675294 333888 675300 333900
rect 675352 333888 675358 333940
rect 35618 332732 35624 332784
rect 35676 332772 35682 332784
rect 39574 332772 39580 332784
rect 35676 332744 39580 332772
rect 35676 332732 35682 332744
rect 39574 332732 39580 332744
rect 39632 332732 39638 332784
rect 35802 332596 35808 332648
rect 35860 332636 35866 332648
rect 41690 332636 41696 332648
rect 35860 332608 41696 332636
rect 35860 332596 35866 332608
rect 41690 332596 41696 332608
rect 41748 332596 41754 332648
rect 42058 332596 42064 332648
rect 42116 332636 42122 332648
rect 56226 332636 56232 332648
rect 42116 332608 56232 332636
rect 42116 332596 42122 332608
rect 56226 332596 56232 332608
rect 56284 332596 56290 332648
rect 672626 332392 672632 332444
rect 672684 332432 672690 332444
rect 675110 332432 675116 332444
rect 672684 332404 675116 332432
rect 672684 332392 672690 332404
rect 675110 332392 675116 332404
rect 675168 332392 675174 332444
rect 42426 327020 42432 327072
rect 42484 327060 42490 327072
rect 43438 327060 43444 327072
rect 42484 327032 43444 327060
rect 42484 327020 42490 327032
rect 43438 327020 43444 327032
rect 43496 327020 43502 327072
rect 42426 325592 42432 325644
rect 42484 325632 42490 325644
rect 45554 325632 45560 325644
rect 42484 325604 45560 325632
rect 42484 325592 42490 325604
rect 45554 325592 45560 325604
rect 45612 325592 45618 325644
rect 669774 325592 669780 325644
rect 669832 325632 669838 325644
rect 674926 325632 674932 325644
rect 669832 325604 674932 325632
rect 669832 325592 669838 325604
rect 674926 325592 674932 325604
rect 674984 325592 674990 325644
rect 669222 325456 669228 325508
rect 669280 325496 669286 325508
rect 675110 325496 675116 325508
rect 669280 325468 675116 325496
rect 669280 325456 669286 325468
rect 675110 325456 675116 325468
rect 675168 325456 675174 325508
rect 651650 324300 651656 324352
rect 651708 324340 651714 324352
rect 673546 324340 673552 324352
rect 651708 324312 673552 324340
rect 651708 324300 651714 324312
rect 673546 324300 673552 324312
rect 673604 324300 673610 324352
rect 42426 324232 42432 324284
rect 42484 324272 42490 324284
rect 46566 324272 46572 324284
rect 42484 324244 46572 324272
rect 42484 324232 42490 324244
rect 46566 324232 46572 324244
rect 46624 324232 46630 324284
rect 49510 322940 49516 322992
rect 49568 322980 49574 322992
rect 62114 322980 62120 322992
rect 49568 322952 62120 322980
rect 49568 322940 49574 322952
rect 62114 322940 62120 322952
rect 62172 322940 62178 322992
rect 42426 321512 42432 321564
rect 42484 321552 42490 321564
rect 43622 321552 43628 321564
rect 42484 321524 43628 321552
rect 42484 321512 42490 321524
rect 43622 321512 43628 321524
rect 43680 321512 43686 321564
rect 42242 321240 42248 321292
rect 42300 321280 42306 321292
rect 44450 321280 44456 321292
rect 42300 321252 44456 321280
rect 42300 321240 42306 321252
rect 44450 321240 44456 321252
rect 44508 321240 44514 321292
rect 42426 320084 42432 320136
rect 42484 320124 42490 320136
rect 44634 320124 44640 320136
rect 42484 320096 44640 320124
rect 42484 320084 42490 320096
rect 44634 320084 44640 320096
rect 44692 320084 44698 320136
rect 42426 318792 42432 318844
rect 42484 318832 42490 318844
rect 47026 318832 47032 318844
rect 42484 318804 47032 318832
rect 42484 318792 42490 318804
rect 47026 318792 47032 318804
rect 47084 318792 47090 318844
rect 43622 318044 43628 318096
rect 43680 318084 43686 318096
rect 62758 318084 62764 318096
rect 43680 318056 62764 318084
rect 43680 318044 43686 318056
rect 62758 318044 62764 318056
rect 62816 318044 62822 318096
rect 42426 317364 42432 317416
rect 42484 317404 42490 317416
rect 43806 317404 43812 317416
rect 42484 317376 43812 317404
rect 42484 317364 42490 317376
rect 43806 317364 43812 317376
rect 43864 317364 43870 317416
rect 42242 317228 42248 317280
rect 42300 317268 42306 317280
rect 43990 317268 43996 317280
rect 42300 317240 43996 317268
rect 42300 317228 42306 317240
rect 43990 317228 43996 317240
rect 44048 317228 44054 317280
rect 42426 315868 42432 315920
rect 42484 315908 42490 315920
rect 43070 315908 43076 315920
rect 42484 315880 43076 315908
rect 42484 315868 42490 315880
rect 43070 315868 43076 315880
rect 43128 315868 43134 315920
rect 666370 313556 666376 313608
rect 666428 313596 666434 313608
rect 666428 313568 673454 313596
rect 666428 313556 666434 313568
rect 663242 313420 663248 313472
rect 663300 313460 663306 313472
rect 673426 313460 673454 313568
rect 675478 313460 675484 313472
rect 663300 313432 668624 313460
rect 673426 313432 675484 313460
rect 663300 313420 663306 313432
rect 663426 313284 663432 313336
rect 663484 313324 663490 313336
rect 666370 313324 666376 313336
rect 663484 313296 666376 313324
rect 663484 313284 663490 313296
rect 666370 313284 666376 313296
rect 666428 313284 666434 313336
rect 668596 313324 668624 313432
rect 675478 313420 675484 313432
rect 675536 313420 675542 313472
rect 675478 313324 675484 313336
rect 668596 313296 675484 313324
rect 675478 313284 675484 313296
rect 675536 313284 675542 313336
rect 673914 312468 673920 312520
rect 673972 312508 673978 312520
rect 675478 312508 675484 312520
rect 673972 312480 675484 312508
rect 673972 312468 673978 312480
rect 675478 312468 675484 312480
rect 675536 312468 675542 312520
rect 660666 311992 660672 312044
rect 660724 312032 660730 312044
rect 675294 312032 675300 312044
rect 660724 312004 675300 312032
rect 660724 311992 660730 312004
rect 675294 311992 675300 312004
rect 675352 311992 675358 312044
rect 666186 311856 666192 311908
rect 666244 311896 666250 311908
rect 675478 311896 675484 311908
rect 666244 311868 675484 311896
rect 666244 311856 666250 311868
rect 675478 311856 675484 311868
rect 675536 311856 675542 311908
rect 673086 310836 673092 310888
rect 673144 310876 673150 310888
rect 675294 310876 675300 310888
rect 673144 310848 675300 310876
rect 673144 310836 673150 310848
rect 675294 310836 675300 310848
rect 675352 310836 675358 310888
rect 43438 310496 43444 310548
rect 43496 310536 43502 310548
rect 62114 310536 62120 310548
rect 43496 310508 62120 310536
rect 43496 310496 43502 310508
rect 62114 310496 62120 310508
rect 62172 310496 62178 310548
rect 666370 310496 666376 310548
rect 666428 310536 666434 310548
rect 675478 310536 675484 310548
rect 666428 310508 675484 310536
rect 666428 310496 666434 310508
rect 675478 310496 675484 310508
rect 675536 310496 675542 310548
rect 42426 310360 42432 310412
rect 42484 310400 42490 310412
rect 47210 310400 47216 310412
rect 42484 310372 47216 310400
rect 42484 310360 42490 310372
rect 47210 310360 47216 310372
rect 47268 310360 47274 310412
rect 672810 310020 672816 310072
rect 672868 310060 672874 310072
rect 675478 310060 675484 310072
rect 672868 310032 675484 310060
rect 672868 310020 672874 310032
rect 675478 310020 675484 310032
rect 675536 310020 675542 310072
rect 664254 309340 664260 309392
rect 664312 309380 664318 309392
rect 675478 309380 675484 309392
rect 664312 309352 675484 309380
rect 664312 309340 664318 309352
rect 675478 309340 675484 309352
rect 675536 309340 675542 309392
rect 665082 309136 665088 309188
rect 665140 309176 665146 309188
rect 675294 309176 675300 309188
rect 665140 309148 675300 309176
rect 665140 309136 665146 309148
rect 675294 309136 675300 309148
rect 675352 309136 675358 309188
rect 673086 305464 673092 305516
rect 673144 305504 673150 305516
rect 675478 305504 675484 305516
rect 673144 305476 675484 305504
rect 673144 305464 673150 305476
rect 675478 305464 675484 305476
rect 675536 305464 675542 305516
rect 673362 303832 673368 303884
rect 673420 303872 673426 303884
rect 675478 303872 675484 303884
rect 673420 303844 675484 303872
rect 673420 303832 673426 303844
rect 675478 303832 675484 303844
rect 675536 303832 675542 303884
rect 672534 303424 672540 303476
rect 672592 303464 672598 303476
rect 675478 303464 675484 303476
rect 672592 303436 675484 303464
rect 672592 303424 672598 303436
rect 675478 303424 675484 303436
rect 675536 303424 675542 303476
rect 680354 302200 680360 302252
rect 680412 302240 680418 302252
rect 683114 302240 683120 302252
rect 680412 302212 683120 302240
rect 680412 302200 680418 302212
rect 683114 302200 683120 302212
rect 683172 302200 683178 302252
rect 43806 301180 43812 301232
rect 43864 301220 43870 301232
rect 49326 301220 49332 301232
rect 43864 301192 49332 301220
rect 43864 301180 43870 301192
rect 49326 301180 49332 301192
rect 49384 301180 49390 301232
rect 669774 300772 669780 300824
rect 669832 300812 669838 300824
rect 675478 300812 675484 300824
rect 669832 300784 675484 300812
rect 669832 300772 669838 300784
rect 675478 300772 675484 300784
rect 675536 300772 675542 300824
rect 674788 298460 674794 298512
rect 674846 298500 674852 298512
rect 675018 298500 675024 298512
rect 674846 298472 675024 298500
rect 674846 298460 674852 298472
rect 675018 298460 675024 298472
rect 675076 298460 675082 298512
rect 41690 298364 41696 298376
rect 41386 298336 41696 298364
rect 40954 298256 40960 298308
rect 41012 298256 41018 298308
rect 41138 298256 41144 298308
rect 41196 298296 41202 298308
rect 41386 298296 41414 298336
rect 41690 298324 41696 298336
rect 41748 298324 41754 298376
rect 42058 298324 42064 298376
rect 42116 298364 42122 298376
rect 42886 298364 42892 298376
rect 42116 298336 42892 298364
rect 42116 298324 42122 298336
rect 42886 298324 42892 298336
rect 42944 298324 42950 298376
rect 41196 298268 41414 298296
rect 41196 298256 41202 298268
rect 40972 298160 41000 298256
rect 42058 298188 42064 298240
rect 42116 298228 42122 298240
rect 45186 298228 45192 298240
rect 42116 298200 45192 298228
rect 42116 298188 42122 298200
rect 45186 298188 45192 298200
rect 45244 298188 45250 298240
rect 41690 298160 41696 298172
rect 40972 298132 41696 298160
rect 41690 298120 41696 298132
rect 41748 298120 41754 298172
rect 47946 298120 47952 298172
rect 48004 298160 48010 298172
rect 62114 298160 62120 298172
rect 48004 298132 62120 298160
rect 48004 298120 48010 298132
rect 62114 298120 62120 298132
rect 62172 298120 62178 298172
rect 672350 297712 672356 297764
rect 672408 297752 672414 297764
rect 672718 297752 672724 297764
rect 672408 297724 672724 297752
rect 672408 297712 672414 297724
rect 672718 297712 672724 297724
rect 672776 297712 672782 297764
rect 675846 297168 675852 297220
rect 675904 297208 675910 297220
rect 680998 297208 681004 297220
rect 675904 297180 681004 297208
rect 675904 297168 675910 297180
rect 680998 297168 681004 297180
rect 681056 297168 681062 297220
rect 40954 296692 40960 296744
rect 41012 296732 41018 296744
rect 41690 296732 41696 296744
rect 41012 296704 41696 296732
rect 41012 296692 41018 296704
rect 41690 296692 41696 296704
rect 41748 296692 41754 296744
rect 42058 296692 42064 296744
rect 42116 296732 42122 296744
rect 45186 296732 45192 296744
rect 42116 296704 45192 296732
rect 42116 296692 42122 296704
rect 45186 296692 45192 296704
rect 45244 296692 45250 296744
rect 675478 296216 675484 296268
rect 675536 296216 675542 296268
rect 675496 295928 675524 296216
rect 675478 295876 675484 295928
rect 675536 295876 675542 295928
rect 40494 292544 40500 292596
rect 40552 292584 40558 292596
rect 41598 292584 41604 292596
rect 40552 292556 41604 292584
rect 40552 292544 40558 292556
rect 41598 292544 41604 292556
rect 41656 292544 41662 292596
rect 674466 292272 674472 292324
rect 674524 292312 674530 292324
rect 675110 292312 675116 292324
rect 674524 292284 675116 292312
rect 674524 292272 674530 292284
rect 675110 292272 675116 292284
rect 675168 292272 675174 292324
rect 42886 289960 42892 290012
rect 42944 290000 42950 290012
rect 64138 290000 64144 290012
rect 42944 289972 64144 290000
rect 42944 289960 42950 289972
rect 64138 289960 64144 289972
rect 64196 289960 64202 290012
rect 41138 289824 41144 289876
rect 41196 289864 41202 289876
rect 41690 289864 41696 289876
rect 41196 289836 41696 289864
rect 41196 289824 41202 289836
rect 41690 289824 41696 289836
rect 41748 289824 41754 289876
rect 42058 289824 42064 289876
rect 42116 289864 42122 289876
rect 61378 289864 61384 289876
rect 42116 289836 61384 289864
rect 42116 289824 42122 289836
rect 61378 289824 61384 289836
rect 61436 289824 61442 289876
rect 672350 289824 672356 289876
rect 672408 289864 672414 289876
rect 672718 289864 672724 289876
rect 672408 289836 672724 289864
rect 672408 289824 672414 289836
rect 672718 289824 672724 289836
rect 672776 289824 672782 289876
rect 40954 289076 40960 289128
rect 41012 289116 41018 289128
rect 41690 289116 41696 289128
rect 41012 289088 41696 289116
rect 41012 289076 41018 289088
rect 41690 289076 41696 289088
rect 41748 289076 41754 289128
rect 35158 284928 35164 284980
rect 35216 284968 35222 284980
rect 41690 284968 41696 284980
rect 35216 284940 41696 284968
rect 35216 284928 35222 284940
rect 41690 284928 41696 284940
rect 41748 284928 41754 284980
rect 651650 284316 651656 284368
rect 651708 284356 651714 284368
rect 662046 284356 662052 284368
rect 651708 284328 662052 284356
rect 651708 284316 651714 284328
rect 662046 284316 662052 284328
rect 662104 284316 662110 284368
rect 42242 280100 42248 280152
rect 42300 280140 42306 280152
rect 43990 280140 43996 280152
rect 42300 280112 43996 280140
rect 42300 280100 42306 280112
rect 43990 280100 43996 280112
rect 44048 280100 44054 280152
rect 406930 278672 406936 278724
rect 406988 278712 406994 278724
rect 499574 278712 499580 278724
rect 406988 278684 499580 278712
rect 406988 278672 406994 278684
rect 499574 278672 499580 278684
rect 499632 278672 499638 278724
rect 42426 278536 42432 278588
rect 42484 278576 42490 278588
rect 50706 278576 50712 278588
rect 42484 278548 50712 278576
rect 42484 278536 42490 278548
rect 50706 278536 50712 278548
rect 50764 278536 50770 278588
rect 467558 278536 467564 278588
rect 467616 278576 467622 278588
rect 476482 278576 476488 278588
rect 467616 278548 476488 278576
rect 467616 278536 467622 278548
rect 476482 278536 476488 278548
rect 476540 278536 476546 278588
rect 482278 278536 482284 278588
rect 482336 278576 482342 278588
rect 590562 278576 590568 278588
rect 482336 278548 590568 278576
rect 482336 278536 482342 278548
rect 590562 278536 590568 278548
rect 590620 278536 590626 278588
rect 42426 278400 42432 278452
rect 42484 278440 42490 278452
rect 44358 278440 44364 278452
rect 42484 278412 44364 278440
rect 42484 278400 42490 278412
rect 44358 278400 44364 278412
rect 44416 278400 44422 278452
rect 64138 278400 64144 278452
rect 64196 278440 64202 278452
rect 661034 278440 661040 278452
rect 64196 278412 661040 278440
rect 64196 278400 64202 278412
rect 661034 278400 661040 278412
rect 661092 278400 661098 278452
rect 61378 278264 61384 278316
rect 61436 278304 61442 278316
rect 659654 278304 659660 278316
rect 61436 278276 659660 278304
rect 61436 278264 61442 278276
rect 659654 278264 659660 278276
rect 659712 278264 659718 278316
rect 53282 278128 53288 278180
rect 53340 278168 53346 278180
rect 654134 278168 654140 278180
rect 53340 278140 654140 278168
rect 53340 278128 53346 278140
rect 654134 278128 654140 278140
rect 654192 278128 654198 278180
rect 56226 277992 56232 278044
rect 56284 278032 56290 278044
rect 658274 278032 658280 278044
rect 56284 278004 658280 278032
rect 56284 277992 56290 278004
rect 658274 277992 658280 278004
rect 658332 277992 658338 278044
rect 437198 277788 437204 277840
rect 437256 277828 437262 277840
rect 546678 277828 546684 277840
rect 437256 277800 546684 277828
rect 437256 277788 437262 277800
rect 546678 277788 546684 277800
rect 546736 277788 546742 277840
rect 421926 277652 421932 277704
rect 421984 277692 421990 277704
rect 524322 277692 524328 277704
rect 421984 277664 524328 277692
rect 421984 277652 421990 277664
rect 524322 277652 524328 277664
rect 524380 277652 524386 277704
rect 413646 277516 413652 277568
rect 413704 277556 413710 277568
rect 510338 277556 510344 277568
rect 413704 277528 510344 277556
rect 413704 277516 413710 277528
rect 510338 277516 510344 277528
rect 510396 277516 510402 277568
rect 475930 277420 475936 277432
rect 473326 277392 475936 277420
rect 466086 277312 466092 277364
rect 466144 277352 466150 277364
rect 471238 277352 471244 277364
rect 466144 277324 471244 277352
rect 466144 277312 466150 277324
rect 471238 277312 471244 277324
rect 471296 277312 471302 277364
rect 471422 277312 471428 277364
rect 471480 277352 471486 277364
rect 473326 277352 473354 277392
rect 475930 277380 475936 277392
rect 475988 277380 475994 277432
rect 476482 277380 476488 277432
rect 476540 277420 476546 277432
rect 596634 277420 596640 277432
rect 476540 277392 596640 277420
rect 476540 277380 476546 277392
rect 596634 277380 596640 277392
rect 596692 277380 596698 277432
rect 471480 277324 473354 277352
rect 471480 277312 471486 277324
rect 475764 277256 483014 277284
rect 442534 277176 442540 277228
rect 442592 277216 442598 277228
rect 475764 277216 475792 277256
rect 442592 277188 475792 277216
rect 482986 277216 483014 277256
rect 557626 277216 557632 277228
rect 482986 277188 557632 277216
rect 442592 277176 442598 277188
rect 557626 277176 557632 277188
rect 557684 277176 557690 277228
rect 409322 277040 409328 277092
rect 409380 277080 409386 277092
rect 475562 277080 475568 277092
rect 409380 277052 475568 277080
rect 409380 277040 409386 277052
rect 475562 277040 475568 277052
rect 475620 277040 475626 277092
rect 476390 277040 476396 277092
rect 476448 277080 476454 277092
rect 502334 277080 502340 277092
rect 476448 277052 502340 277080
rect 476448 277040 476454 277052
rect 502334 277040 502340 277052
rect 502392 277040 502398 277092
rect 502518 277040 502524 277092
rect 502576 277080 502582 277092
rect 509050 277080 509056 277092
rect 502576 277052 509056 277080
rect 502576 277040 502582 277052
rect 509050 277040 509056 277052
rect 509108 277040 509114 277092
rect 509234 277040 509240 277092
rect 509292 277080 509298 277092
rect 511994 277080 512000 277092
rect 509292 277052 512000 277080
rect 509292 277040 509298 277052
rect 511994 277040 512000 277052
rect 512052 277040 512058 277092
rect 512178 277040 512184 277092
rect 512236 277080 512242 277092
rect 571978 277080 571984 277092
rect 512236 277052 571984 277080
rect 512236 277040 512242 277052
rect 571978 277040 571984 277052
rect 572036 277040 572042 277092
rect 587158 277080 587164 277092
rect 576826 277052 587164 277080
rect 380710 276904 380716 276956
rect 380768 276944 380774 276956
rect 457162 276944 457168 276956
rect 380768 276916 457168 276944
rect 380768 276904 380774 276916
rect 457162 276904 457168 276916
rect 457220 276904 457226 276956
rect 471238 276904 471244 276956
rect 471296 276944 471302 276956
rect 475746 276944 475752 276956
rect 471296 276916 475752 276944
rect 471296 276904 471302 276916
rect 475746 276904 475752 276916
rect 475804 276904 475810 276956
rect 476666 276904 476672 276956
rect 476724 276944 476730 276956
rect 576826 276944 576854 277052
rect 587158 277040 587164 277052
rect 587216 277040 587222 277092
rect 476724 276916 576854 276944
rect 476724 276904 476730 276916
rect 581638 276904 581644 276956
rect 581696 276944 581702 276956
rect 606110 276944 606116 276956
rect 581696 276916 606116 276944
rect 581696 276904 581702 276916
rect 606110 276904 606116 276916
rect 606168 276904 606174 276956
rect 387334 276768 387340 276820
rect 387392 276808 387398 276820
rect 467834 276808 467840 276820
rect 387392 276780 467840 276808
rect 387392 276768 387398 276780
rect 467834 276768 467840 276780
rect 467892 276768 467898 276820
rect 469030 276768 469036 276820
rect 469088 276808 469094 276820
rect 471422 276808 471428 276820
rect 469088 276780 471428 276808
rect 469088 276768 469094 276780
rect 471422 276768 471428 276780
rect 471480 276768 471486 276820
rect 472894 276768 472900 276820
rect 472952 276808 472958 276820
rect 475746 276808 475752 276820
rect 472952 276780 475752 276808
rect 472952 276768 472958 276780
rect 475746 276768 475752 276780
rect 475804 276768 475810 276820
rect 475930 276768 475936 276820
rect 475988 276808 475994 276820
rect 599026 276808 599032 276820
rect 475988 276780 599032 276808
rect 475988 276768 475994 276780
rect 599026 276768 599032 276780
rect 599084 276768 599090 276820
rect 43806 276632 43812 276684
rect 43864 276672 43870 276684
rect 509050 276672 509056 276684
rect 43864 276644 509056 276672
rect 43864 276632 43870 276644
rect 509050 276632 509056 276644
rect 509108 276632 509114 276684
rect 509234 276632 509240 276684
rect 509292 276672 509298 276684
rect 659838 276672 659844 276684
rect 509292 276644 659844 276672
rect 509292 276632 509298 276644
rect 659838 276632 659844 276644
rect 659896 276632 659902 276684
rect 446306 276496 446312 276548
rect 446364 276536 446370 276548
rect 451274 276536 451280 276548
rect 446364 276508 451280 276536
rect 446364 276496 446370 276508
rect 451274 276496 451280 276508
rect 451332 276496 451338 276548
rect 456978 276496 456984 276548
rect 457036 276536 457042 276548
rect 570690 276536 570696 276548
rect 457036 276508 570696 276536
rect 457036 276496 457042 276508
rect 570690 276496 570696 276508
rect 570748 276496 570754 276548
rect 571978 276496 571984 276548
rect 572036 276536 572042 276548
rect 581638 276536 581644 276548
rect 572036 276508 581644 276536
rect 572036 276496 572042 276508
rect 581638 276496 581644 276508
rect 581696 276496 581702 276548
rect 420362 276360 420368 276412
rect 420420 276400 420426 276412
rect 521010 276400 521016 276412
rect 420420 276372 521016 276400
rect 420420 276360 420426 276372
rect 521010 276360 521016 276372
rect 521068 276360 521074 276412
rect 446950 276224 446956 276276
rect 447008 276264 447014 276276
rect 531222 276264 531228 276276
rect 447008 276236 531228 276264
rect 447008 276224 447014 276236
rect 531222 276224 531228 276236
rect 531280 276224 531286 276276
rect 402790 276088 402796 276140
rect 402848 276128 402854 276140
rect 485728 276128 485734 276140
rect 402848 276100 485734 276128
rect 402848 276088 402854 276100
rect 485728 276088 485734 276100
rect 485786 276088 485792 276140
rect 485866 276088 485872 276140
rect 485924 276128 485930 276140
rect 499390 276128 499396 276140
rect 485924 276100 499396 276128
rect 485924 276088 485930 276100
rect 499390 276088 499396 276100
rect 499448 276088 499454 276140
rect 499528 276088 499534 276140
rect 499586 276128 499592 276140
rect 499586 276100 622440 276128
rect 499586 276088 499592 276100
rect 110782 275952 110788 276004
rect 110840 275992 110846 276004
rect 156414 275992 156420 276004
rect 110840 275964 156420 275992
rect 110840 275952 110846 275964
rect 156414 275952 156420 275964
rect 156472 275952 156478 276004
rect 171042 275952 171048 276004
rect 171100 275992 171106 276004
rect 175642 275992 175648 276004
rect 171100 275964 175648 275992
rect 171100 275952 171106 275964
rect 175642 275952 175648 275964
rect 175700 275952 175706 276004
rect 175826 275952 175832 276004
rect 175884 275992 175890 276004
rect 177390 275992 177396 276004
rect 175884 275964 177396 275992
rect 175884 275952 175890 275964
rect 177390 275952 177396 275964
rect 177448 275952 177454 276004
rect 344002 275952 344008 276004
rect 344060 275992 344066 276004
rect 354306 275992 354312 276004
rect 344060 275964 354312 275992
rect 344060 275952 344066 275964
rect 354306 275952 354312 275964
rect 354364 275952 354370 276004
rect 356974 275952 356980 276004
rect 357032 275992 357038 276004
rect 388622 275992 388628 276004
rect 357032 275964 388628 275992
rect 357032 275952 357038 275964
rect 388622 275952 388628 275964
rect 388680 275952 388686 276004
rect 388990 275952 388996 276004
rect 389048 275992 389054 276004
rect 418154 275992 418160 276004
rect 389048 275964 418160 275992
rect 389048 275952 389054 275964
rect 418154 275952 418160 275964
rect 418212 275952 418218 276004
rect 418338 275952 418344 276004
rect 418396 275992 418402 276004
rect 427630 275992 427636 276004
rect 418396 275964 427636 275992
rect 418396 275952 418402 275964
rect 427630 275952 427636 275964
rect 427688 275952 427694 276004
rect 436738 275992 436744 276004
rect 427832 275964 436744 275992
rect 217134 275884 217140 275936
rect 217192 275924 217198 275936
rect 218514 275924 218520 275936
rect 217192 275896 218520 275924
rect 217192 275884 217198 275896
rect 218514 275884 218520 275896
rect 218572 275884 218578 275936
rect 103698 275816 103704 275868
rect 103756 275856 103762 275868
rect 160646 275856 160652 275868
rect 103756 275828 160652 275856
rect 103756 275816 103762 275828
rect 160646 275816 160652 275828
rect 160704 275816 160710 275868
rect 174630 275816 174636 275868
rect 174688 275856 174694 275868
rect 197538 275856 197544 275868
rect 174688 275828 197544 275856
rect 174688 275816 174694 275828
rect 197538 275816 197544 275828
rect 197596 275816 197602 275868
rect 316770 275816 316776 275868
rect 316828 275856 316834 275868
rect 327074 275856 327080 275868
rect 316828 275828 327080 275856
rect 316828 275816 316834 275828
rect 327074 275816 327080 275828
rect 327132 275816 327138 275868
rect 331214 275816 331220 275868
rect 331272 275856 331278 275868
rect 340138 275856 340144 275868
rect 331272 275828 340144 275856
rect 331272 275816 331278 275828
rect 340138 275816 340144 275828
rect 340196 275816 340202 275868
rect 343818 275816 343824 275868
rect 343876 275856 343882 275868
rect 370866 275856 370872 275868
rect 343876 275828 370872 275856
rect 343876 275816 343882 275828
rect 370866 275816 370872 275828
rect 370924 275816 370930 275868
rect 371050 275816 371056 275868
rect 371108 275856 371114 275868
rect 407482 275856 407488 275868
rect 371108 275828 407488 275856
rect 371108 275816 371114 275828
rect 407482 275816 407488 275828
rect 407540 275816 407546 275868
rect 410058 275816 410064 275868
rect 410116 275856 410122 275868
rect 421650 275856 421656 275868
rect 410116 275828 421656 275856
rect 410116 275816 410122 275828
rect 421650 275816 421656 275828
rect 421708 275816 421714 275868
rect 426066 275816 426072 275868
rect 426124 275856 426130 275868
rect 427832 275856 427860 275964
rect 436738 275952 436744 275964
rect 436796 275952 436802 276004
rect 436922 275952 436928 276004
rect 436980 275992 436986 276004
rect 471238 275992 471244 276004
rect 436980 275964 471244 275992
rect 436980 275952 436986 275964
rect 471238 275952 471244 275964
rect 471296 275952 471302 276004
rect 471422 275952 471428 276004
rect 471480 275992 471486 276004
rect 473722 275992 473728 276004
rect 471480 275964 473728 275992
rect 471480 275952 471486 275964
rect 473722 275952 473728 275964
rect 473780 275952 473786 276004
rect 473906 275952 473912 276004
rect 473964 275992 473970 276004
rect 477218 275992 477224 276004
rect 473964 275964 477224 275992
rect 473964 275952 473970 275964
rect 477218 275952 477224 275964
rect 477276 275952 477282 276004
rect 477402 275952 477408 276004
rect 477460 275992 477466 276004
rect 485222 275992 485228 276004
rect 477460 275964 485228 275992
rect 477460 275952 477466 275964
rect 485222 275952 485228 275964
rect 485280 275952 485286 276004
rect 487890 275992 487896 276004
rect 485746 275964 487896 275992
rect 426124 275828 427860 275856
rect 426124 275816 426130 275828
rect 427998 275816 428004 275868
rect 428056 275856 428062 275868
rect 465534 275856 465540 275868
rect 428056 275828 465540 275856
rect 428056 275816 428062 275828
rect 465534 275816 465540 275828
rect 465592 275816 465598 275868
rect 465718 275816 465724 275868
rect 465776 275856 465782 275868
rect 470870 275856 470876 275868
rect 465776 275828 470876 275856
rect 465776 275816 465782 275828
rect 470870 275816 470876 275828
rect 470928 275816 470934 275868
rect 471054 275816 471060 275868
rect 471112 275856 471118 275868
rect 480806 275856 480812 275868
rect 471112 275828 480812 275856
rect 471112 275816 471118 275828
rect 480806 275816 480812 275828
rect 480864 275816 480870 275868
rect 480990 275816 480996 275868
rect 481048 275856 481054 275868
rect 484302 275856 484308 275868
rect 481048 275828 484308 275856
rect 481048 275816 481054 275828
rect 484302 275816 484308 275828
rect 484360 275816 484366 275868
rect 484486 275816 484492 275868
rect 484544 275856 484550 275868
rect 485746 275856 485774 275964
rect 487890 275952 487896 275964
rect 487948 275952 487954 276004
rect 490558 275952 490564 276004
rect 490616 275992 490622 276004
rect 498562 275992 498568 276004
rect 490616 275964 498568 275992
rect 490616 275952 490622 275964
rect 498562 275952 498568 275964
rect 498620 275952 498626 276004
rect 498746 275952 498752 276004
rect 498804 275992 498810 276004
rect 501782 275992 501788 276004
rect 498804 275964 501788 275992
rect 498804 275952 498810 275964
rect 501782 275952 501788 275964
rect 501840 275952 501846 276004
rect 501966 275952 501972 276004
rect 502024 275992 502030 276004
rect 511534 275992 511540 276004
rect 502024 275964 511540 275992
rect 502024 275952 502030 275964
rect 511534 275952 511540 275964
rect 511592 275952 511598 276004
rect 561030 275952 561036 276004
rect 561088 275992 561094 276004
rect 565906 275992 565912 276004
rect 561088 275964 565912 275992
rect 561088 275952 561094 275964
rect 565906 275952 565912 275964
rect 565964 275952 565970 276004
rect 622412 275992 622440 276100
rect 635642 275992 635648 276004
rect 622412 275964 635648 275992
rect 635642 275952 635648 275964
rect 635700 275952 635706 276004
rect 484544 275828 485774 275856
rect 484544 275816 484550 275828
rect 485866 275816 485872 275868
rect 485924 275856 485930 275868
rect 611998 275856 612004 275868
rect 485924 275828 612004 275856
rect 485924 275816 485930 275828
rect 611998 275816 612004 275828
rect 612056 275816 612062 275868
rect 96614 275680 96620 275732
rect 96672 275720 96678 275732
rect 153838 275720 153844 275732
rect 96672 275692 153844 275720
rect 96672 275680 96678 275692
rect 153838 275680 153844 275692
rect 153896 275680 153902 275732
rect 160462 275680 160468 275732
rect 160520 275720 160526 275732
rect 174446 275720 174452 275732
rect 160520 275692 174452 275720
rect 160520 275680 160526 275692
rect 174446 275680 174452 275692
rect 174504 275680 174510 275732
rect 181714 275680 181720 275732
rect 181772 275720 181778 275732
rect 207014 275720 207020 275732
rect 181772 275692 207020 275720
rect 181772 275680 181778 275692
rect 207014 275680 207020 275692
rect 207072 275680 207078 275732
rect 298002 275680 298008 275732
rect 298060 275720 298066 275732
rect 298060 275692 302556 275720
rect 298060 275680 298066 275692
rect 85942 275544 85948 275596
rect 86000 275584 86006 275596
rect 149054 275584 149060 275596
rect 86000 275556 149060 275584
rect 86000 275544 86006 275556
rect 149054 275544 149060 275556
rect 149112 275544 149118 275596
rect 153286 275544 153292 275596
rect 153344 275584 153350 275596
rect 185762 275584 185768 275596
rect 153344 275556 185768 275584
rect 153344 275544 153350 275556
rect 185762 275544 185768 275556
rect 185820 275544 185826 275596
rect 199470 275544 199476 275596
rect 199528 275584 199534 275596
rect 210970 275584 210976 275596
rect 199528 275556 210976 275584
rect 199528 275544 199534 275556
rect 210970 275544 210976 275556
rect 211028 275544 211034 275596
rect 218330 275544 218336 275596
rect 218388 275584 218394 275596
rect 218388 275556 219434 275584
rect 218388 275544 218394 275556
rect 68186 275408 68192 275460
rect 68244 275448 68250 275460
rect 135254 275448 135260 275460
rect 68244 275420 135260 275448
rect 68244 275408 68250 275420
rect 135254 275408 135260 275420
rect 135312 275408 135318 275460
rect 156874 275408 156880 275460
rect 156932 275448 156938 275460
rect 166166 275448 166172 275460
rect 156932 275420 166172 275448
rect 156932 275408 156938 275420
rect 166166 275408 166172 275420
rect 166224 275408 166230 275460
rect 167546 275408 167552 275460
rect 167604 275448 167610 275460
rect 200022 275448 200028 275460
rect 167604 275420 200028 275448
rect 167604 275408 167610 275420
rect 200022 275408 200028 275420
rect 200080 275408 200086 275460
rect 207750 275408 207756 275460
rect 207808 275448 207814 275460
rect 216674 275448 216680 275460
rect 207808 275420 216680 275448
rect 207808 275408 207814 275420
rect 216674 275408 216680 275420
rect 216732 275408 216738 275460
rect 219406 275448 219434 275556
rect 221918 275544 221924 275596
rect 221976 275584 221982 275596
rect 228450 275584 228456 275596
rect 221976 275556 228456 275584
rect 221976 275544 221982 275556
rect 228450 275544 228456 275556
rect 228508 275544 228514 275596
rect 282914 275544 282920 275596
rect 282972 275584 282978 275596
rect 285766 275584 285772 275596
rect 282972 275556 285772 275584
rect 282972 275544 282978 275556
rect 285766 275544 285772 275556
rect 285824 275544 285830 275596
rect 299014 275544 299020 275596
rect 299072 275584 299078 275596
rect 302326 275584 302332 275596
rect 299072 275556 302332 275584
rect 299072 275544 299078 275556
rect 302326 275544 302332 275556
rect 302384 275544 302390 275596
rect 302528 275584 302556 275692
rect 305086 275680 305092 275732
rect 305144 275720 305150 275732
rect 316494 275720 316500 275732
rect 305144 275692 316500 275720
rect 305144 275680 305150 275692
rect 316494 275680 316500 275692
rect 316552 275680 316558 275732
rect 317322 275680 317328 275732
rect 317380 275720 317386 275732
rect 329466 275720 329472 275732
rect 317380 275692 329472 275720
rect 317380 275680 317386 275692
rect 329466 275680 329472 275692
rect 329524 275680 329530 275732
rect 374362 275720 374368 275732
rect 329760 275692 374368 275720
rect 311710 275584 311716 275596
rect 302528 275556 311716 275584
rect 311710 275544 311716 275556
rect 311768 275544 311774 275596
rect 313274 275544 313280 275596
rect 313332 275584 313338 275596
rect 325970 275584 325976 275596
rect 313332 275556 325976 275584
rect 313332 275544 313338 275556
rect 325970 275544 325976 275556
rect 326028 275544 326034 275596
rect 329190 275544 329196 275596
rect 329248 275584 329254 275596
rect 329760 275584 329788 275692
rect 374362 275680 374368 275692
rect 374420 275680 374426 275732
rect 380894 275680 380900 275732
rect 380952 275720 380958 275732
rect 411070 275720 411076 275732
rect 380952 275692 411076 275720
rect 380952 275680 380958 275692
rect 411070 275680 411076 275692
rect 411128 275680 411134 275732
rect 414198 275680 414204 275732
rect 414256 275720 414262 275732
rect 508682 275720 508688 275732
rect 414256 275692 508688 275720
rect 414256 275680 414262 275692
rect 508682 275680 508688 275692
rect 508740 275680 508746 275732
rect 511350 275680 511356 275732
rect 511408 275720 511414 275732
rect 633342 275720 633348 275732
rect 511408 275692 633348 275720
rect 511408 275680 511414 275692
rect 633342 275680 633348 275692
rect 633400 275680 633406 275732
rect 329248 275556 329788 275584
rect 329248 275544 329254 275556
rect 333606 275544 333612 275596
rect 333664 275584 333670 275596
rect 381538 275584 381544 275596
rect 333664 275556 381544 275584
rect 333664 275544 333670 275556
rect 381538 275544 381544 275556
rect 381596 275544 381602 275596
rect 394602 275544 394608 275596
rect 394660 275584 394666 275596
rect 470502 275584 470508 275596
rect 394660 275556 470508 275584
rect 394660 275544 394666 275556
rect 470502 275544 470508 275556
rect 470560 275544 470566 275596
rect 471238 275544 471244 275596
rect 471296 275584 471302 275596
rect 471296 275556 485084 275584
rect 471296 275544 471302 275556
rect 222838 275448 222844 275460
rect 219406 275420 222844 275448
rect 222838 275408 222844 275420
rect 222896 275408 222902 275460
rect 236086 275408 236092 275460
rect 236144 275448 236150 275460
rect 242250 275448 242256 275460
rect 236144 275420 242256 275448
rect 236144 275408 236150 275420
rect 242250 275408 242256 275420
rect 242308 275408 242314 275460
rect 285858 275408 285864 275460
rect 285916 275448 285922 275460
rect 303430 275448 303436 275460
rect 285916 275420 303436 275448
rect 285916 275408 285922 275420
rect 303430 275408 303436 275420
rect 303488 275408 303494 275460
rect 318794 275448 318800 275460
rect 303632 275420 318800 275448
rect 70578 275272 70584 275324
rect 70636 275312 70642 275324
rect 139762 275312 139768 275324
rect 70636 275284 139768 275312
rect 70636 275272 70642 275284
rect 139762 275272 139768 275284
rect 139820 275272 139826 275324
rect 149790 275272 149796 275324
rect 149848 275312 149854 275324
rect 184750 275312 184756 275324
rect 149848 275284 184756 275312
rect 149848 275272 149854 275284
rect 184750 275272 184756 275284
rect 184808 275272 184814 275324
rect 188798 275272 188804 275324
rect 188856 275312 188862 275324
rect 188856 275284 200114 275312
rect 188856 275272 188862 275284
rect 107194 275136 107200 275188
rect 107252 275176 107258 275188
rect 151170 275176 151176 275188
rect 107252 275148 151176 275176
rect 107252 275136 107258 275148
rect 151170 275136 151176 275148
rect 151228 275136 151234 275188
rect 152182 275136 152188 275188
rect 152240 275176 152246 275188
rect 162578 275176 162584 275188
rect 152240 275148 162584 275176
rect 152240 275136 152246 275148
rect 162578 275136 162584 275148
rect 162636 275136 162642 275188
rect 200086 275108 200114 275284
rect 227806 275272 227812 275324
rect 227864 275312 227870 275324
rect 237374 275312 237380 275324
rect 227864 275284 237380 275312
rect 227864 275272 227870 275284
rect 237374 275272 237380 275284
rect 237432 275272 237438 275324
rect 238478 275272 238484 275324
rect 238536 275312 238542 275324
rect 243722 275312 243728 275324
rect 238536 275284 243728 275312
rect 238536 275272 238542 275284
rect 243722 275272 243728 275284
rect 243780 275272 243786 275324
rect 265894 275272 265900 275324
rect 265952 275312 265958 275324
rect 271506 275312 271512 275324
rect 265952 275284 271512 275312
rect 265952 275272 265958 275284
rect 271506 275272 271512 275284
rect 271564 275272 271570 275324
rect 278406 275272 278412 275324
rect 278464 275312 278470 275324
rect 292850 275312 292856 275324
rect 278464 275284 292856 275312
rect 278464 275272 278470 275284
rect 292850 275272 292856 275284
rect 292908 275272 292914 275324
rect 302234 275272 302240 275324
rect 302292 275312 302298 275324
rect 303632 275312 303660 275420
rect 318794 275408 318800 275420
rect 318852 275408 318858 275460
rect 320082 275408 320088 275460
rect 320140 275448 320146 275460
rect 336550 275448 336556 275460
rect 320140 275420 336556 275448
rect 320140 275408 320146 275420
rect 336550 275408 336556 275420
rect 336608 275408 336614 275460
rect 340230 275408 340236 275460
rect 340288 275448 340294 275460
rect 392118 275448 392124 275460
rect 340288 275420 392124 275448
rect 340288 275408 340294 275420
rect 392118 275408 392124 275420
rect 392176 275408 392182 275460
rect 392302 275408 392308 275460
rect 392360 275448 392366 275460
rect 396902 275448 396908 275460
rect 392360 275420 396908 275448
rect 392360 275408 392366 275420
rect 396902 275408 396908 275420
rect 396960 275408 396966 275460
rect 397086 275408 397092 275460
rect 397144 275448 397150 275460
rect 471054 275448 471060 275460
rect 397144 275420 471060 275448
rect 397144 275408 397150 275420
rect 471054 275408 471060 275420
rect 471112 275408 471118 275460
rect 471238 275408 471244 275460
rect 471296 275448 471302 275460
rect 484854 275448 484860 275460
rect 471296 275420 484860 275448
rect 471296 275408 471302 275420
rect 484854 275408 484860 275420
rect 484912 275408 484918 275460
rect 485056 275448 485084 275556
rect 485222 275544 485228 275596
rect 485280 275584 485286 275596
rect 490558 275584 490564 275596
rect 485280 275556 490564 275584
rect 485280 275544 485286 275556
rect 490558 275544 490564 275556
rect 490616 275544 490622 275596
rect 490742 275544 490748 275596
rect 490800 275584 490806 275596
rect 494974 275584 494980 275596
rect 490800 275556 494980 275584
rect 490800 275544 490806 275556
rect 494974 275544 494980 275556
rect 495032 275544 495038 275596
rect 495158 275544 495164 275596
rect 495216 275584 495222 275596
rect 604914 275584 604920 275596
rect 495216 275556 604920 275584
rect 495216 275544 495222 275556
rect 604914 275544 604920 275556
rect 604972 275544 604978 275596
rect 499390 275448 499396 275460
rect 485056 275420 499396 275448
rect 499390 275408 499396 275420
rect 499448 275408 499454 275460
rect 616782 275448 616788 275460
rect 499546 275420 616788 275448
rect 322382 275312 322388 275324
rect 302292 275284 303660 275312
rect 306346 275284 322388 275312
rect 302292 275272 302298 275284
rect 211246 275204 211252 275256
rect 211304 275244 211310 275256
rect 212442 275244 212448 275256
rect 211304 275216 212448 275244
rect 211304 275204 211310 275216
rect 212442 275204 212448 275216
rect 212500 275204 212506 275256
rect 245562 275136 245568 275188
rect 245620 275176 245626 275188
rect 246298 275176 246304 275188
rect 245620 275148 246304 275176
rect 245620 275136 245626 275148
rect 246298 275136 246304 275148
rect 246356 275136 246362 275188
rect 301498 275136 301504 275188
rect 301556 275176 301562 275188
rect 306346 275176 306374 275284
rect 322382 275272 322388 275284
rect 322440 275272 322446 275324
rect 322566 275272 322572 275324
rect 322624 275312 322630 275324
rect 333054 275312 333060 275324
rect 322624 275284 333060 275312
rect 322624 275272 322630 275284
rect 333054 275272 333060 275284
rect 333112 275272 333118 275324
rect 342254 275272 342260 275324
rect 342312 275312 342318 275324
rect 350718 275312 350724 275324
rect 342312 275284 350724 275312
rect 342312 275272 342318 275284
rect 350718 275272 350724 275284
rect 350776 275272 350782 275324
rect 350902 275272 350908 275324
rect 350960 275312 350966 275324
rect 399202 275312 399208 275324
rect 350960 275284 399208 275312
rect 350960 275272 350966 275284
rect 399202 275272 399208 275284
rect 399260 275272 399266 275324
rect 399846 275272 399852 275324
rect 399904 275312 399910 275324
rect 484486 275312 484492 275324
rect 399904 275284 484492 275312
rect 399904 275272 399910 275284
rect 484486 275272 484492 275284
rect 484544 275272 484550 275324
rect 487338 275312 487344 275324
rect 484964 275284 487344 275312
rect 301556 275148 306374 275176
rect 301556 275136 301562 275148
rect 336458 275136 336464 275188
rect 336516 275176 336522 275188
rect 343634 275176 343640 275188
rect 336516 275148 343640 275176
rect 336516 275136 336522 275148
rect 343634 275136 343640 275148
rect 343692 275136 343698 275188
rect 350534 275136 350540 275188
rect 350592 275176 350598 275188
rect 357894 275176 357900 275188
rect 350592 275148 357900 275176
rect 350592 275136 350598 275148
rect 357894 275136 357900 275148
rect 357952 275136 357958 275188
rect 365622 275136 365628 275188
rect 365680 275176 365686 275188
rect 375558 275176 375564 275188
rect 365680 275148 375564 275176
rect 365680 275136 365686 275148
rect 375558 275136 375564 275148
rect 375616 275136 375622 275188
rect 376018 275136 376024 275188
rect 376076 275176 376082 275188
rect 403986 275176 403992 275188
rect 376076 275148 403992 275176
rect 376076 275136 376082 275148
rect 403986 275136 403992 275148
rect 404044 275136 404050 275188
rect 404262 275136 404268 275188
rect 404320 275176 404326 275188
rect 425238 275176 425244 275188
rect 404320 275148 425244 275176
rect 404320 275136 404326 275148
rect 425238 275136 425244 275148
rect 425296 275136 425302 275188
rect 425422 275136 425428 275188
rect 425480 275176 425486 275188
rect 427998 275176 428004 275188
rect 425480 275148 428004 275176
rect 425480 275136 425486 275148
rect 427998 275136 428004 275148
rect 428056 275136 428062 275188
rect 430574 275136 430580 275188
rect 430632 275176 430638 275188
rect 436554 275176 436560 275188
rect 430632 275148 436560 275176
rect 430632 275136 430638 275148
rect 436554 275136 436560 275148
rect 436612 275136 436618 275188
rect 436738 275136 436744 275188
rect 436796 275176 436802 275188
rect 465718 275176 465724 275188
rect 436796 275148 465724 275176
rect 436796 275136 436802 275148
rect 465718 275136 465724 275148
rect 465776 275136 465782 275188
rect 465902 275136 465908 275188
rect 465960 275176 465966 275188
rect 466408 275176 466414 275188
rect 465960 275148 466414 275176
rect 465960 275136 465966 275148
rect 466408 275136 466414 275148
rect 466466 275136 466472 275188
rect 466546 275136 466552 275188
rect 466604 275176 466610 275188
rect 484964 275176 484992 275284
rect 487338 275272 487344 275284
rect 487396 275272 487402 275324
rect 487522 275272 487528 275324
rect 487580 275312 487586 275324
rect 491478 275312 491484 275324
rect 487580 275284 491484 275312
rect 487580 275272 487586 275284
rect 491478 275272 491484 275284
rect 491536 275272 491542 275324
rect 491662 275272 491668 275324
rect 491720 275312 491726 275324
rect 498746 275312 498752 275324
rect 491720 275284 498752 275312
rect 491720 275272 491726 275284
rect 498746 275272 498752 275284
rect 498804 275272 498810 275324
rect 498930 275272 498936 275324
rect 498988 275312 498994 275324
rect 499546 275312 499574 275420
rect 616782 275408 616788 275420
rect 616840 275408 616846 275460
rect 498988 275284 499574 275312
rect 498988 275272 498994 275284
rect 499666 275272 499672 275324
rect 499724 275312 499730 275324
rect 640426 275312 640432 275324
rect 499724 275284 640432 275312
rect 499724 275272 499730 275284
rect 640426 275272 640432 275284
rect 640484 275272 640490 275324
rect 466604 275148 484992 275176
rect 466604 275136 466610 275148
rect 485222 275136 485228 275188
rect 485280 275176 485286 275188
rect 485280 275148 523724 275176
rect 485280 275136 485286 275148
rect 213914 275108 213920 275120
rect 200086 275080 213920 275108
rect 213914 275068 213920 275080
rect 213972 275068 213978 275120
rect 122806 275012 142568 275040
rect 81250 274932 81256 274984
rect 81308 274972 81314 274984
rect 86218 274972 86224 274984
rect 81308 274944 86224 274972
rect 81308 274932 81314 274944
rect 86218 274932 86224 274944
rect 86276 274932 86282 274984
rect 116670 274864 116676 274916
rect 116728 274904 116734 274916
rect 122806 274904 122834 275012
rect 116728 274876 122834 274904
rect 116728 274864 116734 274876
rect 135622 274864 135628 274916
rect 135680 274904 135686 274916
rect 142540 274904 142568 275012
rect 142706 275000 142712 275052
rect 142764 275040 142770 275052
rect 169754 275040 169760 275052
rect 142764 275012 169760 275040
rect 142764 275000 142770 275012
rect 169754 275000 169760 275012
rect 169812 275000 169818 275052
rect 249058 275000 249064 275052
rect 249116 275040 249122 275052
rect 250346 275040 250352 275052
rect 249116 275012 250352 275040
rect 249116 275000 249122 275012
rect 250346 275000 250352 275012
rect 250404 275000 250410 275052
rect 347038 275000 347044 275052
rect 347096 275040 347102 275052
rect 350902 275040 350908 275052
rect 347096 275012 350908 275040
rect 347096 275000 347102 275012
rect 350902 275000 350908 275012
rect 350960 275000 350966 275052
rect 375282 275000 375288 275052
rect 375340 275040 375346 275052
rect 375340 275012 379376 275040
rect 375340 275000 375346 275012
rect 178126 274932 178132 274984
rect 178184 274972 178190 274984
rect 180058 274972 180064 274984
rect 178184 274944 180064 274972
rect 178184 274932 178190 274944
rect 180058 274932 180064 274944
rect 180116 274932 180122 274984
rect 214834 274932 214840 274984
rect 214892 274972 214898 274984
rect 221458 274972 221464 274984
rect 214892 274944 221464 274972
rect 214892 274932 214898 274944
rect 221458 274932 221464 274944
rect 221516 274932 221522 274984
rect 365254 274932 365260 274984
rect 365312 274972 365318 274984
rect 369670 274972 369676 274984
rect 365312 274944 369676 274972
rect 365312 274932 365318 274944
rect 369670 274932 369676 274944
rect 369728 274932 369734 274984
rect 142982 274904 142988 274916
rect 135680 274876 142154 274904
rect 142540 274876 142988 274904
rect 135680 274864 135686 274876
rect 140314 274728 140320 274780
rect 140372 274768 140378 274780
rect 140774 274768 140780 274780
rect 140372 274740 140780 274768
rect 140372 274728 140378 274740
rect 140774 274728 140780 274740
rect 140832 274728 140838 274780
rect 142126 274768 142154 274876
rect 142982 274864 142988 274876
rect 143040 274864 143046 274916
rect 150986 274864 150992 274916
rect 151044 274904 151050 274916
rect 152642 274904 152648 274916
rect 151044 274876 152648 274904
rect 151044 274864 151050 274876
rect 152642 274864 152648 274876
rect 152700 274864 152706 274916
rect 374546 274864 374552 274916
rect 374604 274904 374610 274916
rect 379146 274904 379152 274916
rect 374604 274876 379152 274904
rect 374604 274864 374610 274876
rect 379146 274864 379152 274876
rect 379204 274864 379210 274916
rect 379348 274904 379376 275012
rect 382366 275000 382372 275052
rect 382424 275040 382430 275052
rect 408678 275040 408684 275052
rect 382424 275012 408684 275040
rect 382424 275000 382430 275012
rect 408678 275000 408684 275012
rect 408736 275000 408742 275052
rect 408862 275000 408868 275052
rect 408920 275040 408926 275052
rect 412450 275040 412456 275052
rect 408920 275012 412456 275040
rect 408920 275000 408926 275012
rect 412450 275000 412456 275012
rect 412508 275000 412514 275052
rect 414014 275000 414020 275052
rect 414072 275040 414078 275052
rect 415762 275040 415768 275052
rect 414072 275012 415768 275040
rect 414072 275000 414078 275012
rect 415762 275000 415768 275012
rect 415820 275000 415826 275052
rect 422110 275000 422116 275052
rect 422168 275040 422174 275052
rect 523402 275040 523408 275052
rect 422168 275012 523408 275040
rect 422168 275000 422174 275012
rect 523402 275000 523408 275012
rect 523460 275000 523466 275052
rect 523696 275040 523724 275148
rect 523862 275136 523868 275188
rect 523920 275176 523926 275188
rect 537570 275176 537576 275188
rect 523920 275148 537576 275176
rect 523920 275136 523926 275148
rect 537570 275136 537576 275148
rect 537628 275136 537634 275188
rect 537754 275136 537760 275188
rect 537812 275176 537818 275188
rect 552934 275176 552940 275188
rect 537812 275148 552940 275176
rect 537812 275136 537818 275148
rect 552934 275136 552940 275148
rect 552992 275136 552998 275188
rect 556154 275136 556160 275188
rect 556212 275176 556218 275188
rect 561214 275176 561220 275188
rect 556212 275148 561220 275176
rect 556212 275136 556218 275148
rect 561214 275136 561220 275148
rect 561272 275136 561278 275188
rect 530486 275040 530492 275052
rect 523696 275012 530492 275040
rect 530486 275000 530492 275012
rect 530544 275000 530550 275052
rect 549346 275040 549352 275052
rect 531056 275012 549352 275040
rect 393314 274904 393320 274916
rect 379348 274876 393320 274904
rect 393314 274864 393320 274876
rect 393372 274864 393378 274916
rect 397362 274864 397368 274916
rect 397420 274904 397426 274916
rect 414566 274904 414572 274916
rect 397420 274876 414572 274904
rect 397420 274864 397426 274876
rect 414566 274864 414572 274876
rect 414624 274864 414630 274916
rect 418062 274864 418068 274916
rect 418120 274904 418126 274916
rect 516226 274904 516232 274916
rect 418120 274876 516232 274904
rect 418120 274864 418126 274876
rect 516226 274864 516232 274876
rect 516284 274864 516290 274916
rect 523862 274904 523868 274916
rect 518866 274876 523868 274904
rect 186406 274796 186412 274848
rect 186464 274836 186470 274848
rect 188430 274836 188436 274848
rect 186464 274808 188436 274836
rect 186464 274796 186470 274808
rect 188430 274796 188436 274808
rect 188488 274796 188494 274848
rect 358722 274796 358728 274848
rect 358780 274836 358786 274848
rect 364978 274836 364984 274848
rect 358780 274808 364984 274836
rect 358780 274796 358786 274808
rect 364978 274796 364984 274808
rect 365036 274796 365042 274848
rect 156598 274768 156604 274780
rect 142126 274740 156604 274768
rect 156598 274728 156604 274740
rect 156656 274728 156662 274780
rect 378778 274728 378784 274780
rect 378836 274768 378842 274780
rect 386230 274768 386236 274780
rect 378836 274740 386236 274768
rect 378836 274728 378842 274740
rect 386230 274728 386236 274740
rect 386288 274728 386294 274780
rect 408494 274728 408500 274780
rect 408552 274768 408558 274780
rect 412266 274768 412272 274780
rect 408552 274740 412272 274768
rect 408552 274728 408558 274740
rect 412266 274728 412272 274740
rect 412324 274728 412330 274780
rect 412450 274728 412456 274780
rect 412508 274768 412514 274780
rect 491662 274768 491668 274780
rect 412508 274740 491668 274768
rect 412508 274728 412514 274740
rect 491662 274728 491668 274740
rect 491720 274728 491726 274780
rect 491846 274728 491852 274780
rect 491904 274768 491910 274780
rect 494146 274768 494152 274780
rect 491904 274740 494152 274768
rect 491904 274728 491910 274740
rect 494146 274728 494152 274740
rect 494204 274728 494210 274780
rect 494330 274728 494336 274780
rect 494388 274768 494394 274780
rect 499390 274768 499396 274780
rect 494388 274740 499396 274768
rect 494388 274728 494394 274740
rect 499390 274728 499396 274740
rect 499448 274728 499454 274780
rect 500126 274728 500132 274780
rect 500184 274768 500190 274780
rect 518866 274768 518894 274876
rect 523862 274864 523868 274876
rect 523920 274864 523926 274916
rect 500184 274740 518894 274768
rect 500184 274728 500190 274740
rect 523678 274728 523684 274780
rect 523736 274768 523742 274780
rect 531056 274768 531084 275012
rect 549346 275000 549352 275012
rect 549404 275000 549410 275052
rect 563054 275000 563060 275052
rect 563112 275040 563118 275052
rect 577774 275040 577780 275052
rect 563112 275012 577780 275040
rect 563112 275000 563118 275012
rect 577774 275000 577780 275012
rect 577832 275000 577838 275052
rect 531222 274864 531228 274916
rect 531280 274904 531286 274916
rect 563514 274904 563520 274916
rect 531280 274876 563520 274904
rect 531280 274864 531286 274876
rect 563514 274864 563520 274876
rect 563572 274864 563578 274916
rect 523736 274740 531084 274768
rect 523736 274728 523742 274740
rect 552658 274728 552664 274780
rect 552716 274768 552722 274780
rect 556430 274768 556436 274780
rect 552716 274740 556436 274768
rect 552716 274728 552722 274740
rect 556430 274728 556436 274740
rect 556488 274728 556494 274780
rect 619450 274728 619456 274780
rect 619508 274768 619514 274780
rect 623866 274768 623872 274780
rect 619508 274740 623872 274768
rect 619508 274728 619514 274740
rect 623866 274728 623872 274740
rect 623924 274728 623930 274780
rect 89530 274660 89536 274712
rect 89588 274700 89594 274712
rect 92474 274700 92480 274712
rect 89588 274672 92480 274700
rect 89588 274660 89594 274672
rect 92474 274660 92480 274672
rect 92532 274660 92538 274712
rect 161566 274660 161572 274712
rect 161624 274700 161630 274712
rect 163682 274700 163688 274712
rect 161624 274672 163688 274700
rect 161624 274660 161630 274672
rect 163682 274660 163688 274672
rect 163740 274660 163746 274712
rect 163958 274660 163964 274712
rect 164016 274700 164022 274712
rect 167822 274700 167828 274712
rect 164016 274672 167828 274700
rect 164016 274660 164022 274672
rect 167822 274660 167828 274672
rect 167880 274660 167886 274712
rect 185210 274660 185216 274712
rect 185268 274700 185274 274712
rect 186958 274700 186964 274712
rect 185268 274672 186964 274700
rect 185268 274660 185274 274672
rect 186958 274660 186964 274672
rect 187016 274660 187022 274712
rect 241974 274660 241980 274712
rect 242032 274700 242038 274712
rect 246022 274700 246028 274712
rect 242032 274672 246028 274700
rect 242032 274660 242038 274672
rect 246022 274660 246028 274672
rect 246080 274660 246086 274712
rect 246758 274660 246764 274712
rect 246816 274700 246822 274712
rect 248874 274700 248880 274712
rect 246816 274672 248880 274700
rect 246816 274660 246822 274672
rect 248874 274660 248880 274672
rect 248932 274660 248938 274712
rect 271138 274660 271144 274712
rect 271196 274700 271202 274712
rect 276290 274700 276296 274712
rect 271196 274672 276296 274700
rect 271196 274660 271202 274672
rect 276290 274660 276296 274672
rect 276348 274660 276354 274712
rect 276658 274660 276664 274712
rect 276716 274700 276722 274712
rect 278682 274700 278688 274712
rect 276716 274672 278688 274700
rect 276716 274660 276722 274672
rect 278682 274660 278688 274672
rect 278740 274660 278746 274712
rect 280706 274660 280712 274712
rect 280764 274700 280770 274712
rect 283374 274700 283380 274712
rect 280764 274672 283380 274700
rect 280764 274660 280770 274672
rect 283374 274660 283380 274672
rect 283432 274660 283438 274712
rect 293218 274660 293224 274712
rect 293276 274700 293282 274712
rect 294046 274700 294052 274712
rect 293276 274672 294052 274700
rect 293276 274660 293282 274672
rect 294046 274660 294052 274672
rect 294104 274660 294110 274712
rect 295518 274660 295524 274712
rect 295576 274700 295582 274712
rect 298738 274700 298744 274712
rect 295576 274672 298744 274700
rect 295576 274660 295582 274672
rect 298738 274660 298744 274672
rect 298796 274660 298802 274712
rect 339218 274660 339224 274712
rect 339276 274700 339282 274712
rect 344830 274700 344836 274712
rect 339276 274672 344836 274700
rect 339276 274660 339282 274672
rect 344830 274660 344836 274672
rect 344888 274660 344894 274712
rect 355686 274660 355692 274712
rect 355744 274700 355750 274712
rect 356698 274700 356704 274712
rect 355744 274672 356704 274700
rect 355744 274660 355750 274672
rect 356698 274660 356704 274672
rect 356756 274660 356762 274712
rect 643738 274660 643744 274712
rect 643796 274700 643802 274712
rect 645118 274700 645124 274712
rect 643796 274672 645124 274700
rect 643796 274660 643802 274672
rect 645118 274660 645124 274672
rect 645176 274660 645182 274712
rect 119338 274632 119344 274644
rect 103486 274604 119344 274632
rect 93026 274456 93032 274508
rect 93084 274496 93090 274508
rect 103486 274496 103514 274604
rect 119338 274592 119344 274604
rect 119396 274592 119402 274644
rect 120258 274592 120264 274644
rect 120316 274632 120322 274644
rect 161428 274632 161434 274644
rect 120316 274604 161434 274632
rect 120316 274592 120322 274604
rect 161428 274592 161434 274604
rect 161486 274592 161492 274644
rect 359458 274592 359464 274644
rect 359516 274632 359522 274644
rect 400398 274632 400404 274644
rect 359516 274604 400404 274632
rect 359516 274592 359522 274604
rect 400398 274592 400404 274604
rect 400456 274592 400462 274644
rect 401318 274592 401324 274644
rect 401376 274632 401382 274644
rect 489822 274632 489828 274644
rect 401376 274604 489828 274632
rect 401376 274592 401382 274604
rect 489822 274592 489828 274604
rect 489880 274592 489886 274644
rect 490006 274592 490012 274644
rect 490064 274632 490070 274644
rect 495250 274632 495256 274644
rect 490064 274604 495256 274632
rect 490064 274592 490070 274604
rect 495250 274592 495256 274604
rect 495308 274592 495314 274644
rect 495388 274592 495394 274644
rect 495446 274632 495452 274644
rect 496998 274632 497004 274644
rect 495446 274604 497004 274632
rect 495446 274592 495452 274604
rect 496998 274592 497004 274604
rect 497056 274592 497062 274644
rect 497182 274592 497188 274644
rect 497240 274632 497246 274644
rect 621474 274632 621480 274644
rect 497240 274604 621480 274632
rect 497240 274592 497246 274604
rect 621474 274592 621480 274604
rect 621532 274592 621538 274644
rect 93084 274468 103514 274496
rect 93084 274456 93090 274468
rect 119062 274456 119068 274508
rect 119120 274496 119126 274508
rect 168466 274496 168472 274508
rect 119120 274468 168472 274496
rect 119120 274456 119126 274468
rect 168466 274456 168472 274468
rect 168524 274456 168530 274508
rect 169754 274456 169760 274508
rect 169812 274496 169818 274508
rect 184934 274496 184940 274508
rect 169812 274468 184940 274496
rect 169812 274456 169818 274468
rect 184934 274456 184940 274468
rect 184992 274456 184998 274508
rect 306190 274456 306196 274508
rect 306248 274496 306254 274508
rect 320082 274496 320088 274508
rect 306248 274468 320088 274496
rect 306248 274456 306254 274468
rect 320082 274456 320088 274468
rect 320140 274456 320146 274508
rect 329650 274456 329656 274508
rect 329708 274496 329714 274508
rect 365622 274496 365628 274508
rect 329708 274468 365628 274496
rect 329708 274456 329714 274468
rect 365622 274456 365628 274468
rect 365680 274456 365686 274508
rect 366358 274456 366364 274508
rect 366416 274496 366422 274508
rect 366416 274468 383654 274496
rect 366416 274456 366422 274468
rect 111978 274320 111984 274372
rect 112036 274360 112042 274372
rect 164234 274360 164240 274372
rect 112036 274332 164240 274360
rect 112036 274320 112042 274332
rect 164234 274320 164240 274332
rect 164292 274320 164298 274372
rect 177390 274320 177396 274372
rect 177448 274360 177454 274372
rect 204254 274360 204260 274372
rect 177448 274332 204260 274360
rect 177448 274320 177454 274332
rect 204254 274320 204260 274332
rect 204312 274320 204318 274372
rect 299198 274320 299204 274372
rect 299256 274360 299262 274372
rect 313274 274360 313280 274372
rect 299256 274332 313280 274360
rect 299256 274320 299262 274332
rect 313274 274320 313280 274332
rect 313332 274320 313338 274372
rect 322750 274320 322756 274372
rect 322808 274360 322814 274372
rect 358722 274360 358728 274372
rect 322808 274332 358728 274360
rect 322808 274320 322814 274332
rect 358722 274320 358728 274332
rect 358780 274320 358786 274372
rect 358906 274320 358912 274372
rect 358964 274360 358970 274372
rect 368014 274360 368020 274372
rect 358964 274332 368020 274360
rect 358964 274320 358970 274332
rect 368014 274320 368020 274332
rect 368072 274320 368078 274372
rect 102502 274184 102508 274236
rect 102560 274224 102566 274236
rect 159082 274224 159088 274236
rect 102560 274196 159088 274224
rect 102560 274184 102566 274196
rect 159082 274184 159088 274196
rect 159140 274184 159146 274236
rect 166350 274184 166356 274236
rect 166408 274224 166414 274236
rect 198918 274224 198924 274236
rect 166408 274196 198924 274224
rect 166408 274184 166414 274196
rect 198918 274184 198924 274196
rect 198976 274184 198982 274236
rect 200574 274184 200580 274236
rect 200632 274224 200638 274236
rect 213178 274224 213184 274236
rect 200632 274196 213184 274224
rect 200632 274184 200638 274196
rect 213178 274184 213184 274196
rect 213236 274184 213242 274236
rect 274358 274184 274364 274236
rect 274416 274224 274422 274236
rect 286870 274224 286876 274236
rect 274416 274196 286876 274224
rect 274416 274184 274422 274196
rect 286870 274184 286876 274196
rect 286928 274184 286934 274236
rect 290458 274184 290464 274236
rect 290516 274224 290522 274236
rect 305822 274224 305828 274236
rect 290516 274196 305828 274224
rect 290516 274184 290522 274196
rect 305822 274184 305828 274196
rect 305880 274184 305886 274236
rect 310054 274184 310060 274236
rect 310112 274224 310118 274236
rect 336458 274224 336464 274236
rect 310112 274196 336464 274224
rect 310112 274184 310118 274196
rect 336458 274184 336464 274196
rect 336516 274184 336522 274236
rect 378778 274224 378784 274236
rect 344986 274196 378784 274224
rect 234890 274116 234896 274168
rect 234948 274156 234954 274168
rect 239490 274156 239496 274168
rect 234948 274128 239496 274156
rect 234948 274116 234954 274128
rect 239490 274116 239496 274128
rect 239548 274116 239554 274168
rect 77662 274048 77668 274100
rect 77720 274088 77726 274100
rect 143626 274088 143632 274100
rect 77720 274060 143632 274088
rect 77720 274048 77726 274060
rect 143626 274048 143632 274060
rect 143684 274048 143690 274100
rect 158070 274048 158076 274100
rect 158128 274088 158134 274100
rect 193214 274088 193220 274100
rect 158128 274060 193220 274088
rect 158128 274048 158134 274060
rect 193214 274048 193220 274060
rect 193272 274048 193278 274100
rect 198274 274048 198280 274100
rect 198332 274088 198338 274100
rect 217962 274088 217968 274100
rect 198332 274060 217968 274088
rect 198332 274048 198338 274060
rect 217962 274048 217968 274060
rect 218020 274048 218026 274100
rect 283926 274048 283932 274100
rect 283984 274088 283990 274100
rect 299014 274088 299020 274100
rect 283984 274060 299020 274088
rect 283984 274048 283990 274060
rect 299014 274048 299020 274060
rect 299072 274048 299078 274100
rect 307570 274048 307576 274100
rect 307628 274088 307634 274100
rect 331214 274088 331220 274100
rect 307628 274060 331220 274088
rect 307628 274048 307634 274060
rect 331214 274048 331220 274060
rect 331272 274048 331278 274100
rect 336550 274048 336556 274100
rect 336608 274088 336614 274100
rect 344986 274088 345014 274196
rect 378778 274184 378784 274196
rect 378836 274184 378842 274236
rect 336608 274060 345014 274088
rect 336608 274048 336614 274060
rect 353938 274048 353944 274100
rect 353996 274088 354002 274100
rect 382642 274088 382648 274100
rect 353996 274060 382648 274088
rect 353996 274048 354002 274060
rect 382642 274048 382648 274060
rect 382700 274048 382706 274100
rect 383626 274088 383654 274468
rect 390278 274456 390284 274508
rect 390336 274496 390342 274508
rect 466408 274496 466414 274508
rect 390336 274468 466414 274496
rect 390336 274456 390342 274468
rect 466408 274456 466414 274468
rect 466466 274456 466472 274508
rect 466546 274456 466552 274508
rect 466604 274496 466610 274508
rect 471054 274496 471060 274508
rect 466604 274468 471060 274496
rect 466604 274456 466610 274468
rect 471054 274456 471060 274468
rect 471112 274456 471118 274508
rect 471238 274456 471244 274508
rect 471296 274496 471302 274508
rect 479610 274496 479616 274508
rect 471296 274468 479616 274496
rect 471296 274456 471302 274468
rect 479610 274456 479616 274468
rect 479668 274456 479674 274508
rect 480346 274456 480352 274508
rect 480404 274496 480410 274508
rect 610802 274496 610808 274508
rect 480404 274468 610808 274496
rect 480404 274456 480410 274468
rect 610802 274456 610808 274468
rect 610860 274456 610866 274508
rect 393222 274320 393228 274372
rect 393280 274360 393286 274372
rect 476206 274360 476212 274372
rect 393280 274332 476212 274360
rect 393280 274320 393286 274332
rect 476206 274320 476212 274332
rect 476264 274320 476270 274372
rect 478598 274320 478604 274372
rect 478656 274360 478662 274372
rect 614390 274360 614396 274372
rect 478656 274332 614396 274360
rect 478656 274320 478662 274332
rect 614390 274320 614396 274332
rect 614448 274320 614454 274372
rect 394326 274184 394332 274236
rect 394384 274224 394390 274236
rect 471238 274224 471244 274236
rect 394384 274196 471244 274224
rect 394384 274184 394390 274196
rect 471238 274184 471244 274196
rect 471296 274184 471302 274236
rect 471422 274184 471428 274236
rect 471480 274224 471486 274236
rect 484854 274224 484860 274236
rect 471480 274196 484860 274224
rect 471480 274184 471486 274196
rect 484854 274184 484860 274196
rect 484912 274184 484918 274236
rect 485222 274184 485228 274236
rect 485280 274224 485286 274236
rect 485280 274196 486096 274224
rect 485280 274184 485286 274196
rect 395706 274088 395712 274100
rect 383626 274060 395712 274088
rect 395706 274048 395712 274060
rect 395764 274048 395770 274100
rect 397178 274048 397184 274100
rect 397236 274088 397242 274100
rect 483198 274088 483204 274100
rect 397236 274060 483204 274088
rect 397236 274048 397242 274060
rect 483198 274048 483204 274060
rect 483256 274048 483262 274100
rect 486068 274088 486096 274196
rect 486418 274184 486424 274236
rect 486476 274224 486482 274236
rect 617978 274224 617984 274236
rect 486476 274196 617984 274224
rect 486476 274184 486482 274196
rect 617978 274184 617984 274196
rect 618036 274184 618042 274236
rect 625062 274088 625068 274100
rect 486068 274060 625068 274088
rect 625062 274048 625068 274060
rect 625120 274048 625126 274100
rect 72970 273912 72976 273964
rect 73028 273952 73034 273964
rect 140958 273952 140964 273964
rect 73028 273924 140964 273952
rect 73028 273912 73034 273924
rect 140958 273912 140964 273924
rect 141016 273912 141022 273964
rect 141786 273912 141792 273964
rect 141844 273952 141850 273964
rect 183738 273952 183744 273964
rect 141844 273924 183744 273952
rect 141844 273912 141850 273924
rect 183738 273912 183744 273924
rect 183796 273912 183802 273964
rect 184474 273912 184480 273964
rect 184532 273952 184538 273964
rect 206278 273952 206284 273964
rect 184532 273924 206284 273952
rect 184532 273912 184538 273924
rect 206278 273912 206284 273924
rect 206336 273912 206342 273964
rect 206554 273912 206560 273964
rect 206612 273952 206618 273964
rect 223850 273952 223856 273964
rect 206612 273924 223856 273952
rect 206612 273912 206618 273924
rect 223850 273912 223856 273924
rect 223908 273912 223914 273964
rect 224218 273912 224224 273964
rect 224276 273952 224282 273964
rect 234890 273952 234896 273964
rect 224276 273924 234896 273952
rect 224276 273912 224282 273924
rect 234890 273912 234896 273924
rect 234948 273912 234954 273964
rect 279878 273912 279884 273964
rect 279936 273952 279942 273964
rect 295150 273952 295156 273964
rect 279936 273924 295156 273952
rect 279936 273912 279942 273924
rect 295150 273912 295156 273924
rect 295208 273912 295214 273964
rect 314102 273952 314108 273964
rect 296686 273924 314108 273952
rect 130838 273776 130844 273828
rect 130896 273816 130902 273828
rect 176746 273816 176752 273828
rect 130896 273788 176752 273816
rect 130896 273776 130902 273788
rect 176746 273776 176752 273788
rect 176804 273776 176810 273828
rect 294598 273776 294604 273828
rect 294656 273816 294662 273828
rect 296686 273816 296714 273924
rect 314102 273912 314108 273924
rect 314160 273912 314166 273964
rect 314470 273912 314476 273964
rect 314528 273952 314534 273964
rect 342254 273952 342260 273964
rect 314528 273924 342260 273952
rect 314528 273912 314534 273924
rect 342254 273912 342260 273924
rect 342312 273912 342318 273964
rect 351178 273912 351184 273964
rect 351236 273952 351242 273964
rect 359458 273952 359464 273964
rect 351236 273924 359464 273952
rect 351236 273912 351242 273924
rect 359458 273912 359464 273924
rect 359516 273912 359522 273964
rect 368014 273912 368020 273964
rect 368072 273952 368078 273964
rect 389726 273952 389732 273964
rect 368072 273924 389732 273952
rect 368072 273912 368078 273924
rect 389726 273912 389732 273924
rect 389784 273912 389790 273964
rect 391842 273912 391848 273964
rect 391900 273952 391906 273964
rect 394602 273952 394608 273964
rect 391900 273924 394608 273952
rect 391900 273912 391906 273924
rect 394602 273912 394608 273924
rect 394660 273912 394666 273964
rect 396718 273912 396724 273964
rect 396776 273952 396782 273964
rect 435174 273952 435180 273964
rect 396776 273924 435180 273952
rect 396776 273912 396782 273924
rect 435174 273912 435180 273924
rect 435232 273912 435238 273964
rect 435358 273912 435364 273964
rect 435416 273952 435422 273964
rect 451228 273952 451234 273964
rect 435416 273924 451234 273952
rect 435416 273912 435422 273924
rect 451228 273912 451234 273924
rect 451286 273912 451292 273964
rect 451366 273912 451372 273964
rect 451424 273952 451430 273964
rect 561030 273952 561036 273964
rect 451424 273924 561036 273952
rect 451424 273912 451430 273924
rect 561030 273912 561036 273924
rect 561088 273912 561094 273964
rect 632698 273912 632704 273964
rect 632756 273952 632762 273964
rect 643922 273952 643928 273964
rect 632756 273924 643928 273952
rect 632756 273912 632762 273924
rect 643922 273912 643928 273924
rect 643980 273912 643986 273964
rect 294656 273788 296714 273816
rect 294656 273776 294662 273788
rect 318702 273776 318708 273828
rect 318760 273816 318766 273828
rect 350534 273816 350540 273828
rect 318760 273788 350540 273816
rect 318760 273776 318766 273788
rect 350534 273776 350540 273788
rect 350592 273776 350598 273828
rect 354214 273776 354220 273828
rect 354272 273816 354278 273828
rect 397362 273816 397368 273828
rect 354272 273788 397368 273816
rect 354272 273776 354278 273788
rect 397362 273776 397368 273788
rect 397420 273776 397426 273828
rect 398742 273776 398748 273828
rect 398800 273816 398806 273828
rect 484302 273816 484308 273828
rect 398800 273788 484308 273816
rect 398800 273776 398806 273788
rect 484302 273776 484308 273788
rect 484360 273776 484366 273828
rect 484854 273776 484860 273828
rect 484912 273816 484918 273828
rect 484912 273788 488028 273816
rect 484912 273776 484918 273788
rect 488000 273748 488028 273788
rect 488718 273776 488724 273828
rect 488776 273816 488782 273828
rect 628558 273816 628564 273828
rect 488776 273788 628564 273816
rect 488776 273776 488782 273788
rect 628558 273776 628564 273788
rect 628616 273776 628622 273828
rect 488000 273720 488304 273748
rect 124950 273640 124956 273692
rect 125008 273680 125014 273692
rect 157978 273680 157984 273692
rect 125008 273652 157984 273680
rect 125008 273640 125014 273652
rect 157978 273640 157984 273652
rect 158036 273640 158042 273692
rect 161474 273640 161480 273692
rect 161532 273680 161538 273692
rect 169938 273680 169944 273692
rect 161532 273652 169944 273680
rect 161532 273640 161538 273652
rect 169938 273640 169944 273652
rect 169996 273640 170002 273692
rect 361206 273640 361212 273692
rect 361264 273680 361270 273692
rect 404262 273680 404268 273692
rect 361264 273652 404268 273680
rect 361264 273640 361270 273652
rect 404262 273640 404268 273652
rect 404320 273640 404326 273692
rect 405550 273640 405556 273692
rect 405608 273680 405614 273692
rect 486878 273680 486884 273692
rect 405608 273652 486884 273680
rect 405608 273640 405614 273652
rect 486878 273640 486884 273652
rect 486936 273640 486942 273692
rect 488276 273680 488304 273720
rect 543458 273680 543464 273692
rect 488276 273652 543464 273680
rect 543458 273640 543464 273652
rect 543516 273640 543522 273692
rect 332502 273504 332508 273556
rect 332560 273544 332566 273556
rect 374546 273544 374552 273556
rect 332560 273516 374552 273544
rect 332560 273504 332566 273516
rect 374546 273504 374552 273516
rect 374604 273504 374610 273556
rect 378778 273504 378784 273556
rect 378836 273544 378842 273556
rect 420546 273544 420552 273556
rect 378836 273516 420552 273544
rect 378836 273504 378842 273516
rect 420546 273504 420552 273516
rect 420604 273504 420610 273556
rect 426250 273504 426256 273556
rect 426308 273544 426314 273556
rect 529290 273544 529296 273556
rect 426308 273516 529296 273544
rect 426308 273504 426314 273516
rect 529290 273504 529296 273516
rect 529348 273504 529354 273556
rect 343542 273368 343548 273420
rect 343600 273408 343606 273420
rect 392302 273408 392308 273420
rect 343600 273380 392308 273408
rect 343600 273368 343606 273380
rect 392302 273368 392308 273380
rect 392360 273368 392366 273420
rect 416130 273368 416136 273420
rect 416188 273408 416194 273420
rect 515122 273408 515128 273420
rect 416188 273380 515128 273408
rect 416188 273368 416194 273380
rect 515122 273368 515128 273380
rect 515180 273368 515186 273420
rect 395430 273300 395436 273352
rect 395488 273340 395494 273352
rect 396902 273340 396908 273352
rect 395488 273312 396908 273340
rect 395488 273300 395494 273312
rect 396902 273300 396908 273312
rect 396960 273300 396966 273352
rect 358170 273232 358176 273284
rect 358228 273272 358234 273284
rect 358722 273272 358728 273284
rect 358228 273244 358728 273272
rect 358228 273232 358234 273244
rect 358722 273232 358728 273244
rect 358780 273232 358786 273284
rect 451090 273232 451096 273284
rect 451148 273272 451154 273284
rect 451228 273272 451234 273284
rect 451148 273244 451234 273272
rect 451148 273232 451154 273244
rect 451228 273232 451234 273244
rect 451286 273232 451292 273284
rect 451366 273232 451372 273284
rect 451424 273272 451430 273284
rect 460750 273272 460756 273284
rect 451424 273244 460756 273272
rect 451424 273232 451430 273244
rect 460750 273232 460756 273244
rect 460808 273232 460814 273284
rect 42426 273164 42432 273216
rect 42484 273204 42490 273216
rect 43070 273204 43076 273216
rect 42484 273176 43076 273204
rect 42484 273164 42490 273176
rect 43070 273164 43076 273176
rect 43128 273164 43134 273216
rect 127342 273164 127348 273216
rect 127400 273204 127406 273216
rect 174262 273204 174268 273216
rect 127400 273176 174268 273204
rect 127400 273164 127406 273176
rect 174262 273164 174268 273176
rect 174320 273164 174326 273216
rect 326890 273164 326896 273216
rect 326948 273204 326954 273216
rect 343818 273204 343824 273216
rect 326948 273176 343824 273204
rect 326948 273164 326954 273176
rect 343818 273164 343824 273176
rect 343876 273164 343882 273216
rect 364334 273164 364340 273216
rect 364392 273204 364398 273216
rect 430758 273204 430764 273216
rect 364392 273176 430764 273204
rect 364392 273164 364398 273176
rect 430758 273164 430764 273176
rect 430816 273164 430822 273216
rect 430942 273164 430948 273216
rect 431000 273204 431006 273216
rect 431000 273176 437152 273204
rect 431000 273164 431006 273176
rect 121362 273028 121368 273080
rect 121420 273068 121426 273080
rect 171594 273068 171600 273080
rect 121420 273040 171600 273068
rect 121420 273028 121426 273040
rect 171594 273028 171600 273040
rect 171652 273028 171658 273080
rect 174446 273028 174452 273080
rect 174504 273068 174510 273080
rect 196158 273068 196164 273080
rect 174504 273040 196164 273068
rect 174504 273028 174510 273040
rect 196158 273028 196164 273040
rect 196216 273028 196222 273080
rect 295150 273028 295156 273080
rect 295208 273068 295214 273080
rect 302234 273068 302240 273080
rect 295208 273040 302240 273068
rect 295208 273028 295214 273040
rect 302234 273028 302240 273040
rect 302292 273028 302298 273080
rect 317138 273028 317144 273080
rect 317196 273068 317202 273080
rect 344002 273068 344008 273080
rect 317196 273040 344008 273068
rect 317196 273028 317202 273040
rect 344002 273028 344008 273040
rect 344060 273028 344066 273080
rect 357986 273028 357992 273080
rect 358044 273068 358050 273080
rect 361390 273068 361396 273080
rect 358044 273040 361396 273068
rect 358044 273028 358050 273040
rect 361390 273028 361396 273040
rect 361448 273028 361454 273080
rect 368842 273028 368848 273080
rect 368900 273068 368906 273080
rect 436922 273068 436928 273080
rect 368900 273040 436928 273068
rect 368900 273028 368906 273040
rect 436922 273028 436928 273040
rect 436980 273028 436986 273080
rect 437124 273068 437152 273176
rect 437428 273164 437434 273216
rect 437486 273204 437492 273216
rect 445478 273204 445484 273216
rect 437486 273176 445484 273204
rect 437486 273164 437492 273176
rect 445478 273164 445484 273176
rect 445536 273164 445542 273216
rect 447686 273204 447692 273216
rect 445680 273176 447692 273204
rect 441614 273068 441620 273080
rect 437124 273040 441620 273068
rect 441614 273028 441620 273040
rect 441672 273028 441678 273080
rect 442074 273028 442080 273080
rect 442132 273068 442138 273080
rect 445680 273068 445708 273176
rect 447686 273164 447692 273176
rect 447744 273164 447750 273216
rect 460934 273164 460940 273216
rect 460992 273204 460998 273216
rect 568298 273204 568304 273216
rect 460992 273176 568304 273204
rect 460992 273164 460998 273176
rect 568298 273164 568304 273176
rect 568356 273164 568362 273216
rect 456766 273108 459692 273136
rect 442132 273040 445708 273068
rect 442132 273028 442138 273040
rect 446122 273028 446128 273080
rect 446180 273068 446186 273080
rect 456766 273068 456794 273108
rect 446180 273040 456794 273068
rect 459664 273068 459692 273108
rect 555234 273068 555240 273080
rect 459664 273040 555240 273068
rect 446180 273028 446186 273040
rect 555234 273028 555240 273040
rect 555292 273028 555298 273080
rect 572162 273028 572168 273080
rect 572220 273068 572226 273080
rect 608502 273068 608508 273080
rect 572220 273040 608508 273068
rect 572220 273028 572226 273040
rect 608502 273028 608508 273040
rect 608560 273028 608566 273080
rect 71774 272892 71780 272944
rect 71832 272932 71838 272944
rect 109678 272932 109684 272944
rect 71832 272904 109684 272932
rect 71832 272892 71838 272904
rect 109678 272892 109684 272904
rect 109736 272892 109742 272944
rect 109954 272892 109960 272944
rect 110012 272932 110018 272944
rect 163314 272932 163320 272944
rect 110012 272904 163320 272932
rect 110012 272892 110018 272904
rect 163314 272892 163320 272904
rect 163372 272892 163378 272944
rect 180794 272892 180800 272944
rect 180852 272932 180858 272944
rect 207474 272932 207480 272944
rect 180852 272904 207480 272932
rect 180852 272892 180858 272904
rect 207474 272892 207480 272904
rect 207532 272892 207538 272944
rect 302878 272892 302884 272944
rect 302936 272932 302942 272944
rect 317690 272932 317696 272944
rect 302936 272904 317696 272932
rect 302936 272892 302942 272904
rect 317690 272892 317696 272904
rect 317748 272892 317754 272944
rect 325510 272892 325516 272944
rect 325568 272932 325574 272944
rect 368474 272932 368480 272944
rect 325568 272904 368480 272932
rect 325568 272892 325574 272904
rect 368474 272892 368480 272904
rect 368532 272892 368538 272944
rect 381354 272892 381360 272944
rect 381412 272932 381418 272944
rect 384482 272932 384488 272944
rect 381412 272904 384488 272932
rect 381412 272892 381418 272904
rect 384482 272892 384488 272904
rect 384540 272892 384546 272944
rect 387794 272892 387800 272944
rect 387852 272932 387858 272944
rect 387852 272904 447272 272932
rect 387852 272892 387858 272904
rect 97718 272756 97724 272808
rect 97776 272796 97782 272808
rect 155402 272796 155408 272808
rect 97776 272768 155408 272796
rect 97776 272756 97782 272768
rect 155402 272756 155408 272768
rect 155460 272756 155466 272808
rect 168650 272756 168656 272808
rect 168708 272796 168714 272808
rect 198734 272796 198740 272808
rect 168708 272768 198740 272796
rect 168708 272756 168714 272768
rect 198734 272756 198740 272768
rect 198792 272756 198798 272808
rect 210602 272796 210608 272808
rect 200086 272768 210608 272796
rect 91830 272620 91836 272672
rect 91888 272660 91894 272672
rect 152366 272660 152372 272672
rect 91888 272632 152372 272660
rect 91888 272620 91894 272632
rect 152366 272620 152372 272632
rect 152424 272620 152430 272672
rect 159266 272620 159272 272672
rect 159324 272660 159330 272672
rect 194778 272660 194784 272672
rect 159324 272632 194784 272660
rect 159324 272620 159330 272632
rect 194778 272620 194784 272632
rect 194836 272620 194842 272672
rect 195698 272620 195704 272672
rect 195756 272660 195762 272672
rect 200086 272660 200114 272768
rect 210602 272756 210608 272768
rect 210660 272756 210666 272808
rect 300670 272756 300676 272808
rect 300728 272796 300734 272808
rect 317322 272796 317328 272808
rect 300728 272768 317328 272796
rect 300728 272756 300734 272768
rect 317322 272756 317328 272768
rect 317380 272756 317386 272808
rect 321462 272756 321468 272808
rect 321520 272796 321526 272808
rect 357986 272796 357992 272808
rect 321520 272768 357992 272796
rect 321520 272756 321526 272768
rect 357986 272756 357992 272768
rect 358044 272756 358050 272808
rect 359458 272756 359464 272808
rect 359516 272796 359522 272808
rect 365254 272796 365260 272808
rect 359516 272768 365260 272796
rect 359516 272756 359522 272768
rect 365254 272756 365260 272768
rect 365312 272756 365318 272808
rect 376570 272756 376576 272808
rect 376628 272796 376634 272808
rect 446306 272796 446312 272808
rect 376628 272768 446312 272796
rect 376628 272756 376634 272768
rect 446306 272756 446312 272768
rect 446364 272756 446370 272808
rect 447244 272796 447272 272904
rect 447410 272892 447416 272944
rect 447468 272932 447474 272944
rect 451090 272932 451096 272944
rect 447468 272904 451096 272932
rect 447468 272892 447474 272904
rect 451090 272892 451096 272904
rect 451148 272892 451154 272944
rect 451918 272892 451924 272944
rect 451976 272932 451982 272944
rect 456610 272932 456616 272944
rect 451976 272904 456616 272932
rect 451976 272892 451982 272904
rect 456610 272892 456616 272904
rect 456668 272892 456674 272944
rect 575382 272932 575388 272944
rect 457272 272904 575388 272932
rect 452102 272796 452108 272808
rect 447244 272768 452108 272796
rect 452102 272756 452108 272768
rect 452160 272756 452166 272808
rect 453850 272756 453856 272808
rect 453908 272796 453914 272808
rect 457272 272796 457300 272904
rect 575382 272892 575388 272904
rect 575440 272892 575446 272944
rect 453908 272768 457300 272796
rect 453908 272756 453914 272768
rect 457438 272756 457444 272808
rect 457496 272796 457502 272808
rect 571794 272796 571800 272808
rect 457496 272768 571800 272796
rect 457496 272756 457502 272768
rect 571794 272756 571800 272768
rect 571852 272756 571858 272808
rect 578878 272756 578884 272808
rect 578936 272796 578942 272808
rect 636838 272796 636844 272808
rect 578936 272768 636844 272796
rect 578936 272756 578942 272768
rect 636838 272756 636844 272768
rect 636896 272756 636902 272808
rect 195756 272632 200114 272660
rect 195756 272620 195762 272632
rect 210050 272620 210056 272672
rect 210108 272660 210114 272672
rect 226426 272660 226432 272672
rect 210108 272632 226432 272660
rect 210108 272620 210114 272632
rect 226426 272620 226432 272632
rect 226484 272620 226490 272672
rect 289078 272620 289084 272672
rect 289136 272660 289142 272672
rect 299934 272660 299940 272672
rect 289136 272632 299940 272660
rect 289136 272620 289142 272632
rect 299934 272620 299940 272632
rect 299992 272620 299998 272672
rect 300118 272620 300124 272672
rect 300176 272660 300182 272672
rect 319622 272660 319628 272672
rect 300176 272632 319628 272660
rect 300176 272620 300182 272632
rect 319622 272620 319628 272632
rect 319680 272620 319686 272672
rect 333238 272620 333244 272672
rect 333296 272660 333302 272672
rect 377950 272660 377956 272672
rect 333296 272632 377956 272660
rect 333296 272620 333302 272632
rect 377950 272620 377956 272632
rect 378008 272620 378014 272672
rect 378134 272620 378140 272672
rect 378192 272660 378198 272672
rect 378192 272632 384344 272660
rect 378192 272620 378198 272632
rect 239674 272552 239680 272604
rect 239732 272592 239738 272604
rect 244550 272592 244556 272604
rect 239732 272564 244556 272592
rect 239732 272552 239738 272564
rect 244550 272552 244556 272564
rect 244608 272552 244614 272604
rect 74074 272484 74080 272536
rect 74132 272524 74138 272536
rect 142154 272524 142160 272536
rect 74132 272496 142160 272524
rect 74132 272484 74138 272496
rect 142154 272484 142160 272496
rect 142212 272484 142218 272536
rect 154482 272484 154488 272536
rect 154540 272524 154546 272536
rect 190730 272524 190736 272536
rect 154540 272496 190736 272524
rect 154540 272484 154546 272496
rect 190730 272484 190736 272496
rect 190788 272484 190794 272536
rect 197078 272484 197084 272536
rect 197136 272524 197142 272536
rect 197136 272496 200114 272524
rect 197136 272484 197142 272496
rect 137922 272348 137928 272400
rect 137980 272388 137986 272400
rect 181162 272388 181168 272400
rect 137980 272360 181168 272388
rect 137980 272348 137986 272360
rect 181162 272348 181168 272360
rect 181220 272348 181226 272400
rect 200086 272388 200114 272496
rect 218514 272484 218520 272536
rect 218572 272524 218578 272536
rect 230566 272524 230572 272536
rect 218572 272496 230572 272524
rect 218572 272484 218578 272496
rect 230566 272484 230572 272496
rect 230624 272484 230630 272536
rect 231394 272484 231400 272536
rect 231452 272524 231458 272536
rect 239306 272524 239312 272536
rect 231452 272496 239312 272524
rect 231452 272484 231458 272496
rect 239306 272484 239312 272496
rect 239364 272484 239370 272536
rect 271690 272484 271696 272536
rect 271748 272524 271754 272536
rect 280982 272524 280988 272536
rect 271748 272496 280988 272524
rect 271748 272484 271754 272496
rect 280982 272484 280988 272496
rect 281040 272484 281046 272536
rect 282178 272484 282184 272536
rect 282236 272524 282242 272536
rect 297542 272524 297548 272536
rect 282236 272496 297548 272524
rect 282236 272484 282242 272496
rect 297542 272484 297548 272496
rect 297600 272484 297606 272536
rect 303430 272484 303436 272536
rect 303488 272524 303494 272536
rect 322566 272524 322572 272536
rect 303488 272496 322572 272524
rect 303488 272484 303494 272496
rect 322566 272484 322572 272496
rect 322624 272484 322630 272536
rect 326706 272484 326712 272536
rect 326764 272524 326770 272536
rect 326764 272496 335354 272524
rect 326764 272484 326770 272496
rect 218238 272388 218244 272400
rect 200086 272360 218244 272388
rect 218238 272348 218244 272360
rect 218296 272348 218302 272400
rect 280982 272348 280988 272400
rect 281040 272388 281046 272400
rect 289262 272388 289268 272400
rect 281040 272360 289268 272388
rect 281040 272348 281046 272360
rect 289262 272348 289268 272360
rect 289320 272348 289326 272400
rect 335326 272388 335354 272496
rect 345658 272484 345664 272536
rect 345716 272524 345722 272536
rect 372062 272524 372068 272536
rect 345716 272496 372068 272524
rect 345716 272484 345722 272496
rect 372062 272484 372068 272496
rect 372120 272484 372126 272536
rect 374454 272484 374460 272536
rect 374512 272524 374518 272536
rect 380894 272524 380900 272536
rect 374512 272496 380900 272524
rect 374512 272484 374518 272496
rect 380894 272484 380900 272496
rect 380952 272484 380958 272536
rect 384316 272524 384344 272632
rect 384482 272620 384488 272672
rect 384540 272660 384546 272672
rect 458358 272660 458364 272672
rect 384540 272632 458364 272660
rect 384540 272620 384546 272632
rect 458358 272620 458364 272632
rect 458416 272620 458422 272672
rect 460474 272620 460480 272672
rect 460532 272660 460538 272672
rect 466270 272660 466276 272672
rect 460532 272632 466276 272660
rect 460532 272620 460538 272632
rect 466270 272620 466276 272632
rect 466328 272620 466334 272672
rect 466454 272620 466460 272672
rect 466512 272660 466518 272672
rect 582466 272660 582472 272672
rect 466512 272632 582472 272660
rect 466512 272620 466518 272632
rect 582466 272620 582472 272632
rect 582524 272620 582530 272672
rect 442074 272524 442080 272536
rect 384316 272496 442080 272524
rect 442074 272484 442080 272496
rect 442132 272484 442138 272536
rect 442276 272496 447180 272524
rect 359458 272388 359464 272400
rect 335326 272360 359464 272388
rect 359458 272348 359464 272360
rect 359516 272348 359522 272400
rect 361850 272348 361856 272400
rect 361908 272388 361914 272400
rect 417234 272388 417240 272400
rect 361908 272360 417240 272388
rect 361908 272348 361914 272360
rect 417234 272348 417240 272360
rect 417292 272348 417298 272400
rect 442276 272388 442304 272496
rect 447152 272456 447180 272496
rect 447410 272484 447416 272536
rect 447468 272524 447474 272536
rect 455874 272524 455880 272536
rect 447468 272496 455880 272524
rect 447468 272484 447474 272496
rect 455874 272484 455880 272496
rect 455932 272484 455938 272536
rect 456058 272484 456064 272536
rect 456116 272524 456122 272536
rect 456116 272496 567194 272524
rect 456116 272484 456122 272496
rect 447152 272428 447272 272456
rect 417436 272360 442304 272388
rect 113174 272212 113180 272264
rect 113232 272252 113238 272264
rect 142798 272252 142804 272264
rect 113232 272224 142804 272252
rect 113232 272212 113238 272224
rect 142798 272212 142804 272224
rect 142856 272212 142862 272264
rect 142982 272212 142988 272264
rect 143040 272252 143046 272264
rect 167454 272252 167460 272264
rect 143040 272224 167460 272252
rect 143040 272212 143046 272224
rect 167454 272212 167460 272224
rect 167512 272212 167518 272264
rect 348418 272212 348424 272264
rect 348476 272252 348482 272264
rect 374638 272252 374644 272264
rect 348476 272224 374644 272252
rect 348476 272212 348482 272224
rect 374638 272212 374644 272224
rect 374696 272212 374702 272264
rect 374822 272212 374828 272264
rect 374880 272252 374886 272264
rect 378134 272252 378140 272264
rect 374880 272224 378140 272252
rect 374880 272212 374886 272224
rect 378134 272212 378140 272224
rect 378192 272212 378198 272264
rect 379146 272212 379152 272264
rect 379204 272252 379210 272264
rect 417436 272252 417464 272360
rect 442718 272348 442724 272400
rect 442776 272388 442782 272400
rect 446766 272388 446772 272400
rect 442776 272360 446772 272388
rect 442776 272348 442782 272360
rect 446766 272348 446772 272360
rect 446824 272348 446830 272400
rect 447244 272388 447272 272428
rect 454218 272388 454224 272400
rect 447244 272360 454224 272388
rect 454218 272348 454224 272360
rect 454276 272348 454282 272400
rect 454402 272348 454408 272400
rect 454460 272388 454466 272400
rect 564710 272388 564716 272400
rect 454460 272360 564716 272388
rect 454460 272348 454466 272360
rect 564710 272348 564716 272360
rect 564768 272348 564774 272400
rect 567166 272388 567194 272496
rect 571978 272484 571984 272536
rect 572036 272524 572042 272536
rect 585594 272524 585600 272536
rect 572036 272496 585600 272524
rect 572036 272484 572042 272496
rect 585594 272484 585600 272496
rect 585652 272484 585658 272536
rect 585778 272484 585784 272536
rect 585836 272524 585842 272536
rect 622670 272524 622676 272536
rect 585836 272496 622676 272524
rect 585836 272484 585842 272496
rect 622670 272484 622676 272496
rect 622728 272484 622734 272536
rect 578510 272388 578516 272400
rect 567166 272360 578516 272388
rect 578510 272348 578516 272360
rect 578568 272348 578574 272400
rect 485728 272252 485734 272264
rect 379204 272224 417464 272252
rect 417528 272224 485734 272252
rect 379204 272212 379210 272224
rect 340690 272076 340696 272128
rect 340748 272116 340754 272128
rect 375282 272116 375288 272128
rect 340748 272088 375288 272116
rect 340748 272076 340754 272088
rect 375282 272076 375288 272088
rect 375340 272076 375346 272128
rect 376754 272076 376760 272128
rect 376812 272116 376818 272128
rect 409874 272116 409880 272128
rect 376812 272088 409880 272116
rect 376812 272076 376818 272088
rect 409874 272076 409880 272088
rect 409932 272076 409938 272128
rect 412266 272076 412272 272128
rect 412324 272116 412330 272128
rect 417528 272116 417556 272224
rect 485728 272212 485734 272224
rect 485786 272212 485792 272264
rect 485866 272212 485872 272264
rect 485924 272252 485930 272264
rect 571978 272252 571984 272264
rect 485924 272224 571984 272252
rect 485924 272212 485930 272224
rect 571978 272212 571984 272224
rect 572036 272212 572042 272264
rect 412324 272088 417556 272116
rect 412324 272076 412330 272088
rect 417694 272076 417700 272128
rect 417752 272116 417758 272128
rect 418338 272116 418344 272128
rect 417752 272088 418344 272116
rect 417752 272076 417758 272088
rect 418338 272076 418344 272088
rect 418396 272076 418402 272128
rect 427768 272116 427774 272128
rect 422956 272088 427774 272116
rect 351730 271940 351736 271992
rect 351788 271980 351794 271992
rect 374454 271980 374460 271992
rect 351788 271952 374460 271980
rect 351788 271940 351794 271952
rect 374454 271940 374460 271952
rect 374512 271940 374518 271992
rect 374638 271940 374644 271992
rect 374696 271980 374702 271992
rect 385034 271980 385040 271992
rect 374696 271952 385040 271980
rect 374696 271940 374702 271952
rect 385034 271940 385040 271952
rect 385092 271940 385098 271992
rect 410702 271940 410708 271992
rect 410760 271980 410766 271992
rect 422956 271980 422984 272088
rect 427768 272076 427774 272088
rect 427826 272076 427832 272128
rect 427906 272076 427912 272128
rect 427964 272116 427970 272128
rect 442718 272116 442724 272128
rect 427964 272088 442724 272116
rect 427964 272076 427970 272088
rect 442718 272076 442724 272088
rect 442776 272076 442782 272128
rect 443362 272076 443368 272128
rect 443420 272116 443426 272128
rect 446122 272116 446128 272128
rect 443420 272088 446128 272116
rect 443420 272076 443426 272088
rect 446122 272076 446128 272088
rect 446180 272076 446186 272128
rect 451274 272076 451280 272128
rect 451332 272116 451338 272128
rect 556154 272116 556160 272128
rect 451332 272088 556160 272116
rect 451332 272076 451338 272088
rect 556154 272076 556160 272088
rect 556212 272076 556218 272128
rect 410760 271952 422984 271980
rect 410760 271940 410766 271952
rect 423490 271940 423496 271992
rect 423548 271980 423554 271992
rect 427078 271980 427084 271992
rect 423548 271952 427084 271980
rect 423548 271940 423554 271952
rect 427078 271940 427084 271952
rect 427136 271940 427142 271992
rect 427262 271940 427268 271992
rect 427320 271980 427326 271992
rect 532786 271980 532792 271992
rect 427320 271952 532792 271980
rect 427320 271940 427326 271952
rect 532786 271940 532792 271952
rect 532844 271940 532850 271992
rect 101306 271804 101312 271856
rect 101364 271844 101370 271856
rect 157610 271844 157616 271856
rect 101364 271816 157616 271844
rect 101364 271804 101370 271816
rect 157610 271804 157616 271816
rect 157668 271804 157674 271856
rect 165154 271804 165160 271856
rect 165212 271844 165218 271856
rect 197354 271844 197360 271856
rect 165212 271816 197360 271844
rect 165212 271804 165218 271816
rect 197354 271804 197360 271816
rect 197412 271804 197418 271856
rect 297358 271804 297364 271856
rect 297416 271844 297422 271856
rect 309410 271844 309416 271856
rect 297416 271816 309416 271844
rect 297416 271804 297422 271816
rect 309410 271804 309416 271816
rect 309468 271804 309474 271856
rect 312538 271804 312544 271856
rect 312596 271844 312602 271856
rect 338574 271844 338580 271856
rect 312596 271816 338580 271844
rect 312596 271804 312602 271816
rect 338574 271804 338580 271816
rect 338632 271804 338638 271856
rect 338942 271804 338948 271856
rect 339000 271844 339006 271856
rect 363782 271844 363788 271856
rect 339000 271816 363788 271844
rect 339000 271804 339006 271816
rect 363782 271804 363788 271816
rect 363840 271804 363846 271856
rect 364812 271816 428412 271844
rect 263410 271736 263416 271788
rect 263468 271776 263474 271788
rect 269206 271776 269212 271788
rect 263468 271748 269212 271776
rect 263468 271736 263474 271748
rect 269206 271736 269212 271748
rect 269264 271736 269270 271788
rect 88610 271668 88616 271720
rect 88668 271708 88674 271720
rect 145558 271708 145564 271720
rect 88668 271680 145564 271708
rect 88668 271668 88674 271680
rect 145558 271668 145564 271680
rect 145616 271668 145622 271720
rect 179322 271668 179328 271720
rect 179380 271708 179386 271720
rect 204898 271708 204904 271720
rect 179380 271680 204904 271708
rect 179380 271668 179386 271680
rect 204898 271668 204904 271680
rect 204956 271668 204962 271720
rect 296622 271668 296628 271720
rect 296680 271708 296686 271720
rect 301498 271708 301504 271720
rect 296680 271680 301504 271708
rect 296680 271668 296686 271680
rect 301498 271668 301504 271680
rect 301556 271668 301562 271720
rect 304902 271668 304908 271720
rect 304960 271708 304966 271720
rect 334158 271708 334164 271720
rect 304960 271680 334164 271708
rect 304960 271668 304966 271680
rect 334158 271668 334164 271680
rect 334216 271668 334222 271720
rect 338022 271668 338028 271720
rect 338080 271708 338086 271720
rect 356974 271708 356980 271720
rect 338080 271680 356980 271708
rect 338080 271668 338086 271680
rect 356974 271668 356980 271680
rect 357032 271668 357038 271720
rect 363690 271668 363696 271720
rect 363748 271708 363754 271720
rect 364812 271708 364840 271816
rect 422754 271708 422760 271720
rect 363748 271680 364840 271708
rect 364904 271680 422760 271708
rect 363748 271668 363754 271680
rect 98914 271532 98920 271584
rect 98972 271572 98978 271584
rect 156230 271572 156236 271584
rect 98972 271544 156236 271572
rect 98972 271532 98978 271544
rect 156230 271532 156236 271544
rect 156288 271532 156294 271584
rect 170122 271532 170128 271584
rect 170180 271572 170186 271584
rect 201034 271572 201040 271584
rect 170180 271544 201040 271572
rect 170180 271532 170186 271544
rect 201034 271532 201040 271544
rect 201092 271532 201098 271584
rect 213638 271532 213644 271584
rect 213696 271572 213702 271584
rect 228266 271572 228272 271584
rect 213696 271544 228272 271572
rect 213696 271532 213702 271544
rect 228266 271532 228272 271544
rect 228324 271532 228330 271584
rect 229002 271532 229008 271584
rect 229060 271572 229066 271584
rect 237834 271572 237840 271584
rect 229060 271544 237840 271572
rect 229060 271532 229066 271544
rect 237834 271532 237840 271544
rect 237892 271532 237898 271584
rect 289630 271532 289636 271584
rect 289688 271572 289694 271584
rect 298002 271572 298008 271584
rect 289688 271544 298008 271572
rect 289688 271532 289694 271544
rect 298002 271532 298008 271544
rect 298060 271532 298066 271584
rect 309042 271532 309048 271584
rect 309100 271572 309106 271584
rect 342438 271572 342444 271584
rect 309100 271544 342444 271572
rect 309100 271532 309106 271544
rect 342438 271532 342444 271544
rect 342496 271532 342502 271584
rect 345842 271532 345848 271584
rect 345900 271572 345906 271584
rect 362586 271572 362592 271584
rect 345900 271544 362592 271572
rect 345900 271532 345906 271544
rect 362586 271532 362592 271544
rect 362644 271532 362650 271584
rect 92474 271396 92480 271448
rect 92532 271436 92538 271448
rect 150434 271436 150440 271448
rect 92532 271408 150440 271436
rect 92532 271396 92538 271408
rect 150434 271396 150440 271408
rect 150492 271396 150498 271448
rect 156598 271396 156604 271448
rect 156656 271436 156662 271448
rect 180794 271436 180800 271448
rect 156656 271408 180800 271436
rect 156656 271396 156662 271408
rect 180794 271396 180800 271408
rect 180852 271396 180858 271448
rect 201770 271396 201776 271448
rect 201828 271436 201834 271448
rect 220998 271436 221004 271448
rect 201828 271408 221004 271436
rect 201828 271396 201834 271408
rect 220998 271396 221004 271408
rect 221056 271396 221062 271448
rect 233694 271396 233700 271448
rect 233752 271436 233758 271448
rect 240778 271436 240784 271448
rect 233752 271408 240784 271436
rect 233752 271396 233758 271408
rect 240778 271396 240784 271408
rect 240836 271396 240842 271448
rect 268838 271396 268844 271448
rect 268896 271436 268902 271448
rect 277486 271436 277492 271448
rect 268896 271408 277492 271436
rect 268896 271396 268902 271408
rect 277486 271396 277492 271408
rect 277544 271396 277550 271448
rect 285582 271396 285588 271448
rect 285640 271436 285646 271448
rect 304626 271436 304632 271448
rect 285640 271408 304632 271436
rect 285640 271396 285646 271408
rect 304626 271396 304632 271408
rect 304684 271396 304690 271448
rect 311710 271396 311716 271448
rect 311768 271436 311774 271448
rect 347222 271436 347228 271448
rect 311768 271408 347228 271436
rect 311768 271396 311774 271408
rect 347222 271396 347228 271408
rect 347280 271396 347286 271448
rect 361482 271396 361488 271448
rect 361540 271436 361546 271448
rect 364904 271436 364932 271680
rect 422754 271668 422760 271680
rect 422812 271668 422818 271720
rect 428182 271708 428188 271720
rect 422956 271680 428188 271708
rect 365530 271532 365536 271584
rect 365588 271572 365594 271584
rect 422956 271572 422984 271680
rect 428182 271668 428188 271680
rect 428240 271668 428246 271720
rect 428384 271708 428412 271816
rect 428550 271804 428556 271856
rect 428608 271844 428614 271856
rect 440602 271844 440608 271856
rect 428608 271816 440608 271844
rect 428608 271804 428614 271816
rect 440602 271804 440608 271816
rect 440660 271804 440666 271856
rect 440970 271804 440976 271856
rect 441028 271844 441034 271856
rect 444558 271844 444564 271856
rect 441028 271816 444564 271844
rect 441028 271804 441034 271816
rect 444558 271804 444564 271816
rect 444616 271804 444622 271856
rect 444742 271804 444748 271856
rect 444800 271844 444806 271856
rect 551738 271844 551744 271856
rect 444800 271816 551744 271844
rect 444800 271804 444806 271816
rect 551738 271804 551744 271816
rect 551796 271804 551802 271856
rect 551922 271804 551928 271856
rect 551980 271844 551986 271856
rect 553854 271844 553860 271856
rect 551980 271816 553860 271844
rect 551980 271804 551986 271816
rect 553854 271804 553860 271816
rect 553912 271804 553918 271856
rect 429194 271708 429200 271720
rect 428384 271680 429200 271708
rect 429194 271668 429200 271680
rect 429252 271668 429258 271720
rect 429378 271668 429384 271720
rect 429436 271708 429442 271720
rect 433334 271708 433340 271720
rect 429436 271680 433340 271708
rect 429436 271668 429442 271680
rect 433334 271668 433340 271680
rect 433392 271668 433398 271720
rect 433518 271668 433524 271720
rect 433576 271708 433582 271720
rect 535178 271708 535184 271720
rect 433576 271680 535184 271708
rect 433576 271668 433582 271680
rect 535178 271668 535184 271680
rect 535236 271668 535242 271720
rect 542998 271668 543004 271720
rect 543056 271708 543062 271720
rect 543056 271680 552704 271708
rect 543056 271668 543062 271680
rect 365588 271544 422984 271572
rect 365588 271532 365594 271544
rect 423122 271532 423128 271584
rect 423180 271572 423186 271584
rect 432598 271572 432604 271584
rect 423180 271544 432604 271572
rect 423180 271532 423186 271544
rect 432598 271532 432604 271544
rect 432656 271532 432662 271584
rect 432782 271532 432788 271584
rect 432840 271572 432846 271584
rect 442258 271572 442264 271584
rect 432840 271544 442264 271572
rect 432840 271532 432846 271544
rect 442258 271532 442264 271544
rect 442316 271532 442322 271584
rect 442718 271532 442724 271584
rect 442776 271572 442782 271584
rect 551922 271572 551928 271584
rect 442776 271544 551928 271572
rect 442776 271532 442782 271544
rect 551922 271532 551928 271544
rect 551980 271532 551986 271584
rect 552676 271572 552704 271680
rect 554038 271668 554044 271720
rect 554096 271708 554102 271720
rect 615586 271708 615592 271720
rect 554096 271680 615592 271708
rect 554096 271668 554102 271680
rect 615586 271668 615592 271680
rect 615644 271668 615650 271720
rect 562318 271572 562324 271584
rect 552676 271544 562324 271572
rect 562318 271532 562324 271544
rect 562376 271532 562382 271584
rect 361540 271408 364932 271436
rect 361540 271396 361546 271408
rect 383194 271396 383200 271448
rect 383252 271436 383258 271448
rect 456794 271436 456800 271448
rect 383252 271408 456800 271436
rect 383252 271396 383258 271408
rect 456794 271396 456800 271408
rect 456852 271396 456858 271448
rect 457438 271396 457444 271448
rect 457496 271436 457502 271448
rect 457496 271408 461716 271436
rect 457496 271396 457502 271408
rect 84746 271260 84752 271312
rect 84804 271300 84810 271312
rect 147674 271300 147680 271312
rect 84804 271272 147680 271300
rect 84804 271260 84810 271272
rect 147674 271260 147680 271272
rect 147732 271260 147738 271312
rect 155678 271260 155684 271312
rect 155736 271300 155742 271312
rect 192386 271300 192392 271312
rect 155736 271272 192392 271300
rect 155736 271260 155742 271272
rect 192386 271260 192392 271272
rect 192444 271260 192450 271312
rect 193490 271260 193496 271312
rect 193548 271300 193554 271312
rect 215754 271300 215760 271312
rect 193548 271272 215760 271300
rect 193548 271260 193554 271272
rect 215754 271260 215760 271272
rect 215812 271260 215818 271312
rect 223114 271260 223120 271312
rect 223172 271300 223178 271312
rect 234154 271300 234160 271312
rect 223172 271272 234160 271300
rect 223172 271260 223178 271272
rect 234154 271260 234160 271272
rect 234212 271260 234218 271312
rect 273070 271260 273076 271312
rect 273128 271300 273134 271312
rect 284570 271300 284576 271312
rect 273128 271272 284576 271300
rect 273128 271260 273134 271272
rect 284570 271260 284576 271272
rect 284628 271260 284634 271312
rect 291838 271260 291844 271312
rect 291896 271300 291902 271312
rect 310514 271300 310520 271312
rect 291896 271272 310520 271300
rect 291896 271260 291902 271272
rect 310514 271260 310520 271272
rect 310572 271260 310578 271312
rect 315942 271260 315948 271312
rect 316000 271300 316006 271312
rect 353110 271300 353116 271312
rect 316000 271272 353116 271300
rect 316000 271260 316006 271272
rect 353110 271260 353116 271272
rect 353168 271260 353174 271312
rect 360194 271300 360200 271312
rect 354646 271272 360200 271300
rect 65886 271124 65892 271176
rect 65944 271164 65950 271176
rect 136634 271164 136640 271176
rect 65944 271136 136640 271164
rect 65944 271124 65950 271136
rect 136634 271124 136640 271136
rect 136692 271124 136698 271176
rect 139118 271124 139124 271176
rect 139176 271164 139182 271176
rect 140038 271164 140044 271176
rect 139176 271136 140044 271164
rect 139176 271124 139182 271136
rect 140038 271124 140044 271136
rect 140096 271124 140102 271176
rect 145006 271124 145012 271176
rect 145064 271164 145070 271176
rect 185578 271164 185584 271176
rect 145064 271136 185584 271164
rect 145064 271124 145070 271136
rect 185578 271124 185584 271136
rect 185636 271124 185642 271176
rect 192202 271124 192208 271176
rect 192260 271164 192266 271176
rect 215294 271164 215300 271176
rect 192260 271136 215300 271164
rect 192260 271124 192266 271136
rect 215294 271124 215300 271136
rect 215352 271124 215358 271176
rect 215938 271124 215944 271176
rect 215996 271164 216002 271176
rect 229738 271164 229744 271176
rect 215996 271136 229744 271164
rect 215996 271124 216002 271136
rect 229738 271124 229744 271136
rect 229796 271124 229802 271176
rect 277302 271124 277308 271176
rect 277360 271164 277366 271176
rect 291654 271164 291660 271176
rect 277360 271136 291660 271164
rect 277360 271124 277366 271136
rect 291654 271124 291660 271136
rect 291712 271124 291718 271176
rect 292390 271124 292396 271176
rect 292448 271164 292454 271176
rect 315298 271164 315304 271176
rect 292448 271136 315304 271164
rect 292448 271124 292454 271136
rect 315298 271124 315304 271136
rect 315356 271124 315362 271176
rect 322198 271124 322204 271176
rect 322256 271164 322262 271176
rect 354646 271164 354674 271272
rect 360194 271260 360200 271272
rect 360252 271260 360258 271312
rect 369946 271260 369952 271312
rect 370004 271300 370010 271312
rect 428550 271300 428556 271312
rect 370004 271272 428556 271300
rect 370004 271260 370010 271272
rect 428550 271260 428556 271272
rect 428608 271260 428614 271312
rect 432598 271260 432604 271312
rect 432656 271300 432662 271312
rect 440970 271300 440976 271312
rect 432656 271272 440976 271300
rect 432656 271260 432662 271272
rect 440970 271260 440976 271272
rect 441028 271260 441034 271312
rect 442258 271260 442264 271312
rect 442316 271300 442322 271312
rect 461688 271300 461716 271408
rect 461854 271396 461860 271448
rect 461912 271436 461918 271448
rect 465166 271436 465172 271448
rect 461912 271408 465172 271436
rect 461912 271396 461918 271408
rect 465166 271396 465172 271408
rect 465224 271396 465230 271448
rect 465626 271396 465632 271448
rect 465684 271436 465690 271448
rect 466408 271436 466414 271448
rect 465684 271408 466414 271436
rect 465684 271396 465690 271408
rect 466408 271396 466414 271408
rect 466466 271396 466472 271448
rect 466546 271396 466552 271448
rect 466604 271436 466610 271448
rect 580074 271436 580080 271448
rect 466604 271408 580080 271436
rect 466604 271396 466610 271408
rect 580074 271396 580080 271408
rect 580132 271396 580138 271448
rect 562134 271300 562140 271312
rect 442316 271272 461624 271300
rect 461688 271272 562140 271300
rect 442316 271260 442322 271272
rect 382366 271164 382372 271176
rect 322256 271136 354674 271164
rect 359476 271136 382372 271164
rect 322256 271124 322262 271136
rect 114278 270988 114284 271040
rect 114336 271028 114342 271040
rect 164878 271028 164884 271040
rect 114336 271000 164884 271028
rect 114336 270988 114342 271000
rect 164878 270988 164884 271000
rect 164936 270988 164942 271040
rect 185762 270988 185768 271040
rect 185820 271028 185826 271040
rect 192202 271028 192208 271040
rect 185820 271000 192208 271028
rect 185820 270988 185826 271000
rect 192202 270988 192208 271000
rect 192260 270988 192266 271040
rect 319438 270988 319444 271040
rect 319496 271028 319502 271040
rect 346026 271028 346032 271040
rect 319496 271000 346032 271028
rect 319496 270988 319502 271000
rect 346026 270988 346032 271000
rect 346084 270988 346090 271040
rect 350442 270988 350448 271040
rect 350500 271028 350506 271040
rect 359476 271028 359504 271136
rect 382366 271124 382372 271136
rect 382424 271124 382430 271176
rect 389818 271124 389824 271176
rect 389876 271164 389882 271176
rect 456794 271164 456800 271176
rect 389876 271136 456800 271164
rect 389876 271124 389882 271136
rect 456794 271124 456800 271136
rect 456852 271124 456858 271176
rect 456978 271124 456984 271176
rect 457036 271164 457042 271176
rect 461394 271164 461400 271176
rect 457036 271136 461400 271164
rect 457036 271124 457042 271136
rect 461394 271124 461400 271136
rect 461452 271124 461458 271176
rect 461596 271164 461624 271272
rect 562134 271260 562140 271272
rect 562192 271260 562198 271312
rect 562318 271260 562324 271312
rect 562376 271300 562382 271312
rect 594334 271300 594340 271312
rect 562376 271272 594340 271300
rect 562376 271260 562382 271272
rect 594334 271260 594340 271272
rect 594392 271260 594398 271312
rect 485728 271164 485734 271176
rect 461596 271136 485734 271164
rect 485728 271124 485734 271136
rect 485786 271124 485792 271176
rect 485866 271124 485872 271176
rect 485924 271164 485930 271176
rect 495434 271164 495440 271176
rect 485924 271136 495440 271164
rect 485924 271124 485930 271136
rect 495434 271124 495440 271136
rect 495492 271124 495498 271176
rect 495618 271124 495624 271176
rect 495676 271164 495682 271176
rect 495676 271136 495940 271164
rect 495676 271124 495682 271136
rect 350500 271000 359504 271028
rect 350500 270988 350506 271000
rect 360102 270988 360108 271040
rect 360160 271028 360166 271040
rect 422478 271028 422484 271040
rect 360160 271000 422484 271028
rect 360160 270988 360166 271000
rect 422478 270988 422484 271000
rect 422536 270988 422542 271040
rect 432782 271028 432788 271040
rect 422956 271000 432788 271028
rect 123754 270852 123760 270904
rect 123812 270892 123818 270904
rect 172698 270892 172704 270904
rect 123812 270864 172704 270892
rect 123812 270852 123818 270864
rect 172698 270852 172704 270864
rect 172756 270852 172762 270904
rect 334618 270852 334624 270904
rect 334676 270892 334682 270904
rect 349614 270892 349620 270904
rect 334676 270864 349620 270892
rect 334676 270852 334682 270864
rect 349614 270852 349620 270864
rect 349672 270852 349678 270904
rect 357158 270852 357164 270904
rect 357216 270892 357222 270904
rect 412588 270892 412594 270904
rect 357216 270864 412594 270892
rect 357216 270852 357222 270864
rect 412588 270852 412594 270864
rect 412646 270852 412652 270904
rect 412726 270852 412732 270904
rect 412784 270892 412790 270904
rect 414014 270892 414020 270904
rect 412784 270864 414020 270892
rect 412784 270852 412790 270864
rect 414014 270852 414020 270864
rect 414072 270852 414078 270904
rect 414658 270852 414664 270904
rect 414716 270892 414722 270904
rect 417234 270892 417240 270904
rect 414716 270864 417240 270892
rect 414716 270852 414722 270864
rect 417234 270852 417240 270864
rect 417292 270852 417298 270904
rect 422956 270892 422984 271000
rect 432782 270988 432788 271000
rect 432840 270988 432846 271040
rect 432966 270988 432972 271040
rect 433024 271028 433030 271040
rect 495618 271028 495624 271040
rect 433024 271000 495624 271028
rect 433024 270988 433030 271000
rect 495618 270988 495624 271000
rect 495676 270988 495682 271040
rect 495912 271028 495940 271136
rect 496538 271124 496544 271176
rect 496596 271164 496602 271176
rect 639230 271164 639236 271176
rect 496596 271136 639236 271164
rect 496596 271124 496602 271136
rect 639230 271124 639236 271136
rect 639288 271124 639294 271176
rect 538398 271028 538404 271040
rect 495912 271000 538404 271028
rect 538398 270988 538404 271000
rect 538456 270988 538462 271040
rect 538858 270988 538864 271040
rect 538916 271028 538922 271040
rect 597830 271028 597836 271040
rect 538916 271000 597836 271028
rect 538916 270988 538922 271000
rect 597830 270988 597836 271000
rect 597888 270988 597894 271040
rect 417436 270864 422984 270892
rect 134426 270716 134432 270768
rect 134484 270756 134490 270768
rect 178954 270756 178960 270768
rect 134484 270728 178960 270756
rect 134484 270716 134490 270728
rect 178954 270716 178960 270728
rect 179012 270716 179018 270768
rect 342530 270716 342536 270768
rect 342588 270756 342594 270768
rect 348142 270756 348148 270768
rect 342588 270728 348148 270756
rect 342588 270716 342594 270728
rect 348142 270716 348148 270728
rect 348200 270716 348206 270768
rect 354490 270716 354496 270768
rect 354548 270756 354554 270768
rect 412082 270756 412088 270768
rect 354548 270728 412088 270756
rect 354548 270716 354554 270728
rect 412082 270716 412088 270728
rect 412140 270716 412146 270768
rect 412450 270716 412456 270768
rect 412508 270756 412514 270768
rect 417436 270756 417464 270864
rect 423306 270852 423312 270904
rect 423364 270892 423370 270904
rect 426434 270892 426440 270904
rect 423364 270864 426440 270892
rect 423364 270852 423370 270864
rect 426434 270852 426440 270864
rect 426492 270852 426498 270904
rect 495066 270892 495072 270904
rect 426636 270864 495072 270892
rect 412508 270728 417464 270756
rect 412508 270716 412514 270728
rect 418246 270716 418252 270768
rect 418304 270756 418310 270768
rect 423122 270756 423128 270768
rect 418304 270728 423128 270756
rect 418304 270716 418310 270728
rect 423122 270716 423128 270728
rect 423180 270716 423186 270768
rect 423306 270716 423312 270768
rect 423364 270756 423370 270768
rect 426636 270756 426664 270864
rect 495066 270852 495072 270864
rect 495124 270852 495130 270904
rect 495802 270852 495808 270904
rect 495860 270892 495866 270904
rect 513834 270892 513840 270904
rect 495860 270864 513840 270892
rect 495860 270852 495866 270864
rect 513834 270852 513840 270864
rect 513892 270852 513898 270904
rect 514018 270852 514024 270904
rect 514076 270892 514082 270904
rect 542998 270892 543004 270904
rect 514076 270864 543004 270892
rect 514076 270852 514082 270864
rect 542998 270852 543004 270864
rect 543056 270852 543062 270904
rect 423364 270728 426664 270756
rect 423364 270716 423370 270728
rect 426986 270716 426992 270768
rect 427044 270756 427050 270768
rect 495066 270756 495072 270768
rect 427044 270728 495072 270756
rect 427044 270716 427050 270728
rect 495066 270716 495072 270728
rect 495124 270716 495130 270768
rect 531590 270756 531596 270768
rect 496096 270728 531596 270756
rect 136818 270580 136824 270632
rect 136876 270620 136882 270632
rect 174630 270620 174636 270632
rect 136876 270592 174636 270620
rect 136876 270580 136882 270592
rect 174630 270580 174636 270592
rect 174688 270580 174694 270632
rect 176764 270592 177896 270620
rect 108942 270444 108948 270496
rect 109000 270484 109006 270496
rect 162394 270484 162400 270496
rect 109000 270456 162400 270484
rect 109000 270444 109006 270456
rect 162394 270444 162400 270456
rect 162452 270444 162458 270496
rect 173802 270444 173808 270496
rect 173860 270484 173866 270496
rect 176764 270484 176792 270592
rect 173860 270456 176792 270484
rect 173860 270444 173866 270456
rect 176930 270444 176936 270496
rect 176988 270484 176994 270496
rect 177868 270484 177896 270592
rect 353202 270580 353208 270632
rect 353260 270620 353266 270632
rect 403986 270620 403992 270632
rect 353260 270592 403992 270620
rect 353260 270580 353266 270592
rect 403986 270580 403992 270592
rect 404044 270580 404050 270632
rect 404170 270580 404176 270632
rect 404228 270620 404234 270632
rect 409506 270620 409512 270632
rect 404228 270592 409512 270620
rect 404228 270580 404234 270592
rect 409506 270580 409512 270592
rect 409564 270580 409570 270632
rect 409690 270580 409696 270632
rect 409748 270620 409754 270632
rect 495434 270620 495440 270632
rect 409748 270592 495440 270620
rect 409748 270580 409754 270592
rect 495434 270580 495440 270592
rect 495492 270580 495498 270632
rect 495894 270580 495900 270632
rect 495952 270620 495958 270632
rect 496096 270620 496124 270728
rect 531590 270716 531596 270728
rect 531648 270716 531654 270768
rect 495952 270592 496124 270620
rect 495952 270580 495958 270592
rect 496354 270580 496360 270632
rect 496412 270620 496418 270632
rect 514018 270620 514024 270632
rect 496412 270592 514024 270620
rect 496412 270580 496418 270592
rect 514018 270580 514024 270592
rect 514076 270580 514082 270632
rect 514202 270580 514208 270632
rect 514260 270620 514266 270632
rect 518618 270620 518624 270632
rect 514260 270592 518624 270620
rect 514260 270580 514266 270592
rect 518618 270580 518624 270592
rect 518676 270580 518682 270632
rect 203610 270484 203616 270496
rect 176988 270456 177804 270484
rect 177868 270456 203616 270484
rect 176988 270444 176994 270456
rect 78858 270308 78864 270360
rect 78916 270348 78922 270360
rect 132586 270348 132592 270360
rect 78916 270320 132592 270348
rect 78916 270308 78922 270320
rect 132586 270308 132592 270320
rect 132644 270308 132650 270360
rect 133782 270308 133788 270360
rect 133840 270348 133846 270360
rect 177574 270348 177580 270360
rect 133840 270320 177580 270348
rect 133840 270308 133846 270320
rect 177574 270308 177580 270320
rect 177632 270308 177638 270360
rect 177776 270348 177804 270456
rect 203610 270444 203616 270456
rect 203668 270444 203674 270496
rect 207014 270444 207020 270496
rect 207072 270484 207078 270496
rect 209498 270484 209504 270496
rect 207072 270456 209504 270484
rect 207072 270444 207078 270456
rect 209498 270444 209504 270456
rect 209556 270444 209562 270496
rect 216674 270444 216680 270496
rect 216732 270484 216738 270496
rect 224954 270484 224960 270496
rect 216732 270456 224960 270484
rect 216732 270444 216738 270456
rect 224954 270444 224960 270456
rect 225012 270444 225018 270496
rect 244366 270444 244372 270496
rect 244424 270484 244430 270496
rect 247770 270484 247776 270496
rect 244424 270456 247776 270484
rect 244424 270444 244430 270456
rect 247770 270444 247776 270456
rect 247828 270444 247834 270496
rect 250162 270444 250168 270496
rect 250220 270484 250226 270496
rect 251450 270484 251456 270496
rect 250220 270456 251456 270484
rect 250220 270444 250226 270456
rect 251450 270444 251456 270456
rect 251508 270444 251514 270496
rect 258810 270444 258816 270496
rect 258868 270484 258874 270496
rect 261294 270484 261300 270496
rect 258868 270456 261300 270484
rect 258868 270444 258874 270456
rect 261294 270444 261300 270456
rect 261352 270444 261358 270496
rect 292666 270444 292672 270496
rect 292724 270484 292730 270496
rect 305086 270484 305092 270496
rect 292724 270456 305092 270484
rect 292724 270444 292730 270456
rect 305086 270444 305092 270456
rect 305144 270444 305150 270496
rect 323578 270444 323584 270496
rect 323636 270484 323642 270496
rect 365806 270484 365812 270496
rect 323636 270456 365812 270484
rect 323636 270444 323642 270456
rect 365806 270444 365812 270456
rect 365864 270444 365870 270496
rect 367738 270444 367744 270496
rect 367796 270484 367802 270496
rect 436094 270484 436100 270496
rect 367796 270456 436100 270484
rect 367796 270444 367802 270456
rect 436094 270444 436100 270456
rect 436152 270444 436158 270496
rect 438394 270444 438400 270496
rect 438452 270484 438458 270496
rect 542998 270484 543004 270496
rect 438452 270456 543004 270484
rect 438452 270444 438458 270456
rect 542998 270444 543004 270456
rect 543056 270444 543062 270496
rect 543182 270444 543188 270496
rect 543240 270484 543246 270496
rect 557810 270484 557816 270496
rect 543240 270456 557816 270484
rect 543240 270444 543246 270456
rect 557810 270444 557816 270456
rect 557868 270444 557874 270496
rect 205818 270348 205824 270360
rect 177776 270320 205824 270348
rect 205818 270308 205824 270320
rect 205876 270308 205882 270360
rect 212258 270308 212264 270360
rect 212316 270348 212322 270360
rect 219434 270348 219440 270360
rect 212316 270320 219440 270348
rect 212316 270308 212322 270320
rect 219434 270308 219440 270320
rect 219492 270308 219498 270360
rect 243170 270308 243176 270360
rect 243228 270348 243234 270360
rect 247034 270348 247040 270360
rect 243228 270320 247040 270348
rect 243228 270308 243234 270320
rect 247034 270308 247040 270320
rect 247092 270308 247098 270360
rect 261018 270308 261024 270360
rect 261076 270348 261082 270360
rect 264974 270348 264980 270360
rect 261076 270320 264980 270348
rect 261076 270308 261082 270320
rect 264974 270308 264980 270320
rect 265032 270308 265038 270360
rect 301958 270308 301964 270360
rect 302016 270348 302022 270360
rect 320266 270348 320272 270360
rect 302016 270320 320272 270348
rect 302016 270308 302022 270320
rect 320266 270308 320272 270320
rect 320324 270308 320330 270360
rect 334986 270308 334992 270360
rect 335044 270348 335050 270360
rect 383654 270348 383660 270360
rect 335044 270320 383660 270348
rect 335044 270308 335050 270320
rect 383654 270308 383660 270320
rect 383712 270308 383718 270360
rect 383838 270308 383844 270360
rect 383896 270348 383902 270360
rect 386414 270348 386420 270360
rect 383896 270320 386420 270348
rect 383896 270308 383902 270320
rect 386414 270308 386420 270320
rect 386472 270308 386478 270360
rect 386598 270308 386604 270360
rect 386656 270348 386662 270360
rect 456610 270348 456616 270360
rect 386656 270320 456616 270348
rect 386656 270308 386662 270320
rect 456610 270308 456616 270320
rect 456668 270308 456674 270360
rect 456748 270308 456754 270360
rect 456806 270348 456812 270360
rect 475930 270348 475936 270360
rect 456806 270320 475936 270348
rect 456806 270308 456812 270320
rect 475930 270308 475936 270320
rect 475988 270308 475994 270360
rect 476482 270308 476488 270360
rect 476540 270348 476546 270360
rect 599394 270348 599400 270360
rect 476540 270320 599400 270348
rect 476540 270308 476546 270320
rect 599394 270308 599400 270320
rect 599452 270308 599458 270360
rect 94222 270172 94228 270224
rect 94280 270212 94286 270224
rect 153562 270212 153568 270224
rect 94280 270184 153568 270212
rect 94280 270172 94286 270184
rect 153562 270172 153568 270184
rect 153620 270172 153626 270224
rect 163682 270172 163688 270224
rect 163740 270212 163746 270224
rect 195514 270212 195520 270224
rect 163740 270184 195520 270212
rect 163740 270172 163746 270184
rect 195514 270172 195520 270184
rect 195572 270172 195578 270224
rect 197538 270172 197544 270224
rect 197596 270212 197602 270224
rect 205082 270212 205088 270224
rect 197596 270184 205088 270212
rect 197596 270172 197602 270184
rect 205082 270172 205088 270184
rect 205140 270172 205146 270224
rect 205542 270172 205548 270224
rect 205600 270212 205606 270224
rect 223482 270212 223488 270224
rect 205600 270184 223488 270212
rect 205600 270172 205606 270184
rect 223482 270172 223488 270184
rect 223540 270172 223546 270224
rect 290826 270172 290832 270224
rect 290884 270212 290890 270224
rect 311894 270212 311900 270224
rect 290884 270184 311900 270212
rect 290884 270172 290890 270184
rect 311894 270172 311900 270184
rect 311952 270172 311958 270224
rect 312814 270172 312820 270224
rect 312872 270212 312878 270224
rect 331398 270212 331404 270224
rect 312872 270184 331404 270212
rect 312872 270172 312878 270184
rect 331398 270172 331404 270184
rect 331456 270172 331462 270224
rect 346394 270172 346400 270224
rect 346452 270212 346458 270224
rect 393498 270212 393504 270224
rect 346452 270184 393504 270212
rect 346452 270172 346458 270184
rect 393498 270172 393504 270184
rect 393556 270172 393562 270224
rect 393866 270172 393872 270224
rect 393924 270212 393930 270224
rect 393924 270184 398328 270212
rect 393924 270172 393930 270184
rect 67542 270036 67548 270088
rect 67600 270076 67606 270088
rect 78214 270076 78220 270088
rect 67600 270048 78220 270076
rect 67600 270036 67606 270048
rect 78214 270036 78220 270048
rect 78272 270036 78278 270088
rect 80054 270036 80060 270088
rect 80112 270076 80118 270088
rect 144454 270076 144460 270088
rect 80112 270048 144460 270076
rect 80112 270036 80118 270048
rect 144454 270036 144460 270048
rect 144512 270036 144518 270088
rect 152642 270036 152648 270088
rect 152700 270076 152706 270088
rect 188890 270076 188896 270088
rect 152700 270048 188896 270076
rect 152700 270036 152706 270048
rect 188890 270036 188896 270048
rect 188948 270036 188954 270088
rect 202966 270036 202972 270088
rect 203024 270076 203030 270088
rect 222010 270076 222016 270088
rect 203024 270048 222016 270076
rect 203024 270036 203030 270048
rect 222010 270036 222016 270048
rect 222068 270036 222074 270088
rect 226610 270036 226616 270088
rect 226668 270076 226674 270088
rect 236730 270076 236736 270088
rect 226668 270048 236736 270076
rect 226668 270036 226674 270048
rect 236730 270036 236736 270048
rect 236788 270036 236794 270088
rect 266170 270036 266176 270088
rect 266228 270076 266234 270088
rect 273254 270076 273260 270088
rect 266228 270048 273260 270076
rect 266228 270036 266234 270048
rect 273254 270036 273260 270048
rect 273312 270036 273318 270088
rect 276474 270036 276480 270088
rect 276532 270076 276538 270088
rect 289814 270076 289820 270088
rect 276532 270048 289820 270076
rect 276532 270036 276538 270048
rect 289814 270036 289820 270048
rect 289872 270036 289878 270088
rect 301222 270036 301228 270088
rect 301280 270076 301286 270088
rect 324314 270076 324320 270088
rect 301280 270048 324320 270076
rect 301280 270036 301286 270048
rect 324314 270036 324320 270048
rect 324372 270036 324378 270088
rect 337194 270036 337200 270088
rect 337252 270076 337258 270088
rect 383838 270076 383844 270088
rect 337252 270048 383844 270076
rect 337252 270036 337258 270048
rect 383838 270036 383844 270048
rect 383896 270036 383902 270088
rect 384114 270036 384120 270088
rect 384172 270076 384178 270088
rect 393682 270076 393688 270088
rect 384172 270048 393688 270076
rect 384172 270036 384178 270048
rect 393682 270036 393688 270048
rect 393740 270036 393746 270088
rect 395982 270036 395988 270088
rect 396040 270076 396046 270088
rect 398300 270076 398328 270184
rect 398466 270172 398472 270224
rect 398524 270212 398530 270224
rect 401870 270212 401876 270224
rect 398524 270184 401876 270212
rect 398524 270172 398530 270184
rect 401870 270172 401876 270184
rect 401928 270172 401934 270224
rect 402238 270172 402244 270224
rect 402296 270212 402302 270224
rect 412588 270212 412594 270224
rect 402296 270184 412594 270212
rect 402296 270172 402302 270184
rect 412588 270172 412594 270184
rect 412646 270172 412652 270224
rect 412726 270172 412732 270224
rect 412784 270212 412790 270224
rect 475746 270212 475752 270224
rect 412784 270184 475752 270212
rect 412784 270172 412790 270184
rect 475746 270172 475752 270184
rect 475804 270172 475810 270224
rect 476206 270172 476212 270224
rect 476264 270212 476270 270224
rect 490282 270212 490288 270224
rect 476264 270184 490288 270212
rect 476264 270172 476270 270184
rect 490282 270172 490288 270184
rect 490340 270172 490346 270224
rect 500218 270212 500224 270224
rect 490576 270184 500224 270212
rect 490576 270144 490604 270184
rect 500218 270172 500224 270184
rect 500276 270172 500282 270224
rect 500402 270172 500408 270224
rect 500460 270212 500466 270224
rect 501966 270212 501972 270224
rect 500460 270184 501972 270212
rect 500460 270172 500466 270184
rect 501966 270172 501972 270184
rect 502024 270172 502030 270224
rect 502150 270172 502156 270224
rect 502208 270212 502214 270224
rect 633618 270212 633624 270224
rect 502208 270184 633624 270212
rect 502208 270172 502214 270184
rect 633618 270172 633624 270184
rect 633676 270172 633682 270224
rect 490484 270116 490604 270144
rect 475746 270076 475752 270088
rect 396040 270048 398236 270076
rect 398300 270048 475752 270076
rect 396040 270036 396046 270048
rect 75822 269900 75828 269952
rect 75880 269940 75886 269952
rect 141786 269940 141792 269952
rect 75880 269912 141792 269940
rect 75880 269900 75886 269912
rect 141786 269900 141792 269912
rect 141844 269900 141850 269952
rect 143902 269900 143908 269952
rect 143960 269940 143966 269952
rect 184474 269940 184480 269952
rect 143960 269912 184480 269940
rect 143960 269900 143966 269912
rect 184474 269900 184480 269912
rect 184532 269900 184538 269952
rect 184750 269900 184756 269952
rect 184808 269940 184814 269952
rect 189626 269940 189632 269952
rect 184808 269912 189632 269940
rect 184808 269900 184814 269912
rect 189626 269900 189632 269912
rect 189684 269900 189690 269952
rect 194594 269900 194600 269952
rect 194652 269940 194658 269952
rect 216858 269940 216864 269952
rect 194652 269912 216864 269940
rect 194652 269900 194658 269912
rect 216858 269900 216864 269912
rect 216916 269900 216922 269952
rect 221458 269900 221464 269952
rect 221516 269940 221522 269952
rect 229370 269940 229376 269952
rect 221516 269912 229376 269940
rect 221516 269900 221522 269912
rect 229370 269900 229376 269912
rect 229428 269900 229434 269952
rect 230382 269900 230388 269952
rect 230440 269940 230446 269952
rect 238938 269940 238944 269952
rect 230440 269912 238944 269940
rect 230440 269900 230446 269912
rect 238938 269900 238944 269912
rect 238996 269900 239002 269952
rect 266906 269900 266912 269952
rect 266964 269940 266970 269952
rect 274634 269940 274640 269952
rect 266964 269912 274640 269940
rect 266964 269900 266970 269912
rect 274634 269900 274640 269912
rect 274692 269900 274698 269952
rect 275002 269900 275008 269952
rect 275060 269940 275066 269952
rect 287054 269940 287060 269952
rect 275060 269912 287060 269940
rect 275060 269900 275066 269912
rect 287054 269900 287060 269912
rect 287112 269900 287118 269952
rect 287514 269900 287520 269952
rect 287572 269940 287578 269952
rect 307754 269940 307760 269952
rect 287572 269912 307760 269940
rect 287572 269900 287578 269912
rect 307754 269900 307760 269912
rect 307812 269900 307818 269952
rect 310330 269900 310336 269952
rect 310388 269940 310394 269952
rect 339218 269940 339224 269952
rect 310388 269912 339224 269940
rect 310388 269900 310394 269912
rect 339218 269900 339224 269912
rect 339276 269900 339282 269952
rect 339402 269900 339408 269952
rect 339460 269940 339466 269952
rect 390554 269940 390560 269952
rect 339460 269912 390560 269940
rect 339460 269900 339466 269912
rect 390554 269900 390560 269912
rect 390612 269900 390618 269952
rect 390738 269900 390744 269952
rect 390796 269940 390802 269952
rect 398208 269940 398236 270048
rect 475746 270036 475752 270048
rect 475804 270036 475810 270088
rect 475930 270036 475936 270088
rect 475988 270076 475994 270088
rect 490484 270076 490512 270116
rect 619450 270076 619456 270088
rect 475988 270048 490512 270076
rect 490668 270048 619456 270076
rect 475988 270036 475994 270048
rect 490668 270008 490696 270048
rect 619450 270036 619456 270048
rect 619508 270036 619514 270088
rect 490576 269980 490696 270008
rect 481634 269940 481640 269952
rect 390796 269912 398144 269940
rect 398208 269912 481640 269940
rect 390796 269900 390802 269912
rect 69382 269764 69388 269816
rect 69440 269804 69446 269816
rect 138842 269804 138848 269816
rect 69440 269776 138848 269804
rect 69440 269764 69446 269776
rect 138842 269764 138848 269776
rect 138900 269764 138906 269816
rect 140774 269764 140780 269816
rect 140832 269804 140838 269816
rect 182266 269804 182272 269816
rect 140832 269776 182272 269804
rect 140832 269764 140838 269776
rect 182266 269764 182272 269776
rect 182324 269764 182330 269816
rect 191742 269764 191748 269816
rect 191800 269804 191806 269816
rect 214650 269804 214656 269816
rect 191800 269776 214656 269804
rect 191800 269764 191806 269776
rect 214650 269764 214656 269776
rect 214708 269764 214714 269816
rect 219618 269764 219624 269816
rect 219676 269804 219682 269816
rect 232314 269804 232320 269816
rect 219676 269776 232320 269804
rect 219676 269764 219682 269776
rect 232314 269764 232320 269776
rect 232372 269764 232378 269816
rect 237190 269764 237196 269816
rect 237248 269804 237254 269816
rect 243354 269804 243360 269816
rect 237248 269776 243360 269804
rect 237248 269764 237254 269776
rect 243354 269764 243360 269776
rect 243412 269764 243418 269816
rect 261754 269764 261760 269816
rect 261812 269804 261818 269816
rect 263594 269804 263600 269816
rect 261812 269776 263600 269804
rect 261812 269764 261818 269776
rect 263594 269764 263600 269776
rect 263652 269764 263658 269816
rect 265434 269764 265440 269816
rect 265492 269804 265498 269816
rect 271874 269804 271880 269816
rect 265492 269776 271880 269804
rect 265492 269764 265498 269776
rect 271874 269764 271880 269776
rect 271932 269764 271938 269816
rect 283098 269764 283104 269816
rect 283156 269804 283162 269816
rect 300854 269804 300860 269816
rect 283156 269776 300860 269804
rect 283156 269764 283162 269776
rect 300854 269764 300860 269776
rect 300912 269764 300918 269816
rect 305546 269764 305552 269816
rect 305604 269804 305610 269816
rect 335354 269804 335360 269816
rect 305604 269776 335360 269804
rect 305604 269764 305610 269776
rect 335354 269764 335360 269776
rect 335412 269764 335418 269816
rect 341242 269764 341248 269816
rect 341300 269804 341306 269816
rect 384114 269804 384120 269816
rect 341300 269776 384120 269804
rect 341300 269764 341306 269776
rect 384114 269764 384120 269776
rect 384172 269764 384178 269816
rect 397546 269804 397552 269816
rect 384316 269776 397552 269804
rect 122742 269628 122748 269680
rect 122800 269668 122806 269680
rect 171226 269668 171232 269680
rect 122800 269640 171232 269668
rect 122800 269628 122806 269640
rect 171226 269628 171232 269640
rect 171284 269628 171290 269680
rect 172422 269628 172428 269680
rect 172480 269668 172486 269680
rect 202138 269668 202144 269680
rect 172480 269640 202144 269668
rect 172480 269628 172486 269640
rect 202138 269628 202144 269640
rect 202196 269628 202202 269680
rect 271874 269628 271880 269680
rect 271932 269668 271938 269680
rect 281534 269668 281540 269680
rect 271932 269640 281540 269668
rect 271932 269628 271938 269640
rect 281534 269628 281540 269640
rect 281592 269628 281598 269680
rect 311526 269628 311532 269680
rect 311584 269668 311590 269680
rect 327258 269668 327264 269680
rect 311584 269640 327264 269668
rect 311584 269628 311590 269640
rect 327258 269628 327264 269640
rect 327316 269628 327322 269680
rect 332318 269628 332324 269680
rect 332376 269668 332382 269680
rect 332376 269640 374684 269668
rect 332376 269628 332382 269640
rect 84102 269492 84108 269544
rect 84160 269532 84166 269544
rect 126698 269532 126704 269544
rect 84160 269504 126704 269532
rect 84160 269492 84166 269504
rect 126698 269492 126704 269504
rect 126756 269492 126762 269544
rect 126882 269492 126888 269544
rect 126940 269532 126946 269544
rect 173434 269532 173440 269544
rect 126940 269504 173440 269532
rect 126940 269492 126946 269504
rect 173434 269492 173440 269504
rect 173492 269492 173498 269544
rect 183462 269492 183468 269544
rect 183520 269532 183526 269544
rect 194502 269532 194508 269544
rect 183520 269504 194508 269532
rect 183520 269492 183526 269504
rect 194502 269492 194508 269504
rect 194560 269492 194566 269544
rect 259638 269492 259644 269544
rect 259696 269532 259702 269544
rect 260834 269532 260840 269544
rect 259696 269504 260840 269532
rect 259696 269492 259702 269504
rect 260834 269492 260840 269504
rect 260892 269492 260898 269544
rect 330202 269492 330208 269544
rect 330260 269532 330266 269544
rect 374454 269532 374460 269544
rect 330260 269504 374460 269532
rect 330260 269492 330266 269504
rect 374454 269492 374460 269504
rect 374512 269492 374518 269544
rect 374656 269532 374684 269640
rect 374822 269628 374828 269680
rect 374880 269668 374886 269680
rect 384316 269668 384344 269776
rect 397546 269764 397552 269776
rect 397604 269764 397610 269816
rect 398116 269804 398144 269912
rect 481634 269900 481640 269912
rect 481692 269900 481698 269952
rect 484302 269900 484308 269952
rect 484360 269940 484366 269952
rect 484360 269912 484900 269940
rect 484360 269900 484366 269912
rect 407942 269804 407948 269816
rect 398116 269776 407948 269804
rect 407942 269764 407948 269776
rect 408000 269764 408006 269816
rect 408126 269764 408132 269816
rect 408184 269804 408190 269816
rect 484670 269804 484676 269816
rect 408184 269776 484676 269804
rect 408184 269764 408190 269776
rect 484670 269764 484676 269776
rect 484728 269764 484734 269816
rect 484872 269804 484900 269912
rect 485038 269900 485044 269952
rect 485096 269940 485102 269952
rect 490190 269940 490196 269952
rect 485096 269912 490196 269940
rect 485096 269900 485102 269912
rect 490190 269900 490196 269912
rect 490248 269900 490254 269952
rect 490576 269804 490604 269980
rect 490834 269900 490840 269952
rect 490892 269940 490898 269952
rect 495250 269940 495256 269952
rect 490892 269912 495256 269940
rect 490892 269900 490898 269912
rect 495250 269900 495256 269912
rect 495308 269900 495314 269952
rect 626534 269940 626540 269952
rect 495406 269912 626540 269940
rect 484872 269776 490604 269804
rect 490834 269764 490840 269816
rect 490892 269804 490898 269816
rect 491386 269804 491392 269816
rect 490892 269776 491392 269804
rect 490892 269764 490898 269776
rect 491386 269764 491392 269776
rect 491444 269764 491450 269816
rect 491570 269764 491576 269816
rect 491628 269804 491634 269816
rect 495406 269804 495434 269912
rect 626534 269900 626540 269912
rect 626592 269900 626598 269952
rect 491628 269776 495434 269804
rect 491628 269764 491634 269776
rect 495526 269764 495532 269816
rect 495584 269804 495590 269816
rect 637574 269804 637580 269816
rect 495584 269776 637580 269804
rect 495584 269764 495590 269776
rect 637574 269764 637580 269776
rect 637632 269764 637638 269816
rect 638310 269764 638316 269816
rect 638368 269804 638374 269816
rect 647234 269804 647240 269816
rect 638368 269776 647240 269804
rect 638368 269764 638374 269776
rect 647234 269764 647240 269776
rect 647292 269764 647298 269816
rect 374880 269640 384344 269668
rect 374880 269628 374886 269640
rect 384482 269628 384488 269680
rect 384540 269668 384546 269680
rect 412726 269668 412732 269680
rect 384540 269640 412732 269668
rect 384540 269628 384546 269640
rect 412726 269628 412732 269640
rect 412784 269628 412790 269680
rect 413094 269628 413100 269680
rect 413152 269668 413158 269680
rect 427814 269668 427820 269680
rect 413152 269640 427820 269668
rect 413152 269628 413158 269640
rect 427814 269628 427820 269640
rect 427872 269628 427878 269680
rect 427998 269628 428004 269680
rect 428056 269668 428062 269680
rect 527174 269668 527180 269680
rect 428056 269640 527180 269668
rect 428056 269628 428062 269640
rect 527174 269628 527180 269640
rect 527232 269628 527238 269680
rect 542998 269628 543004 269680
rect 543056 269668 543062 269680
rect 549898 269668 549904 269680
rect 543056 269640 549904 269668
rect 543056 269628 543062 269640
rect 549898 269628 549904 269640
rect 549956 269628 549962 269680
rect 379514 269532 379520 269544
rect 374656 269504 379520 269532
rect 379514 269492 379520 269504
rect 379572 269492 379578 269544
rect 379698 269492 379704 269544
rect 379756 269532 379762 269544
rect 379756 269504 407804 269532
rect 379756 269492 379762 269504
rect 129366 269356 129372 269408
rect 129424 269396 129430 269408
rect 175642 269396 175648 269408
rect 129424 269368 175648 269396
rect 129424 269356 129430 269368
rect 175642 269356 175648 269368
rect 175700 269356 175706 269408
rect 327994 269356 328000 269408
rect 328052 269396 328058 269408
rect 328052 269368 354674 269396
rect 328052 269356 328058 269368
rect 264698 269288 264704 269340
rect 264756 269328 264762 269340
rect 265894 269328 265900 269340
rect 264756 269300 265900 269328
rect 264756 269288 264762 269300
rect 265894 269288 265900 269300
rect 265952 269288 265958 269340
rect 128538 269220 128544 269272
rect 128596 269260 128602 269272
rect 162946 269260 162952 269272
rect 128596 269232 162952 269260
rect 128596 269220 128602 269232
rect 162946 269220 162952 269232
rect 163004 269220 163010 269272
rect 354646 269260 354674 269368
rect 365714 269356 365720 269408
rect 365772 269396 365778 269408
rect 374822 269396 374828 269408
rect 365772 269368 374828 269396
rect 365772 269356 365778 269368
rect 374822 269356 374828 269368
rect 374880 269356 374886 269408
rect 375006 269356 375012 269408
rect 375064 269396 375070 269408
rect 393406 269396 393412 269408
rect 375064 269368 393412 269396
rect 375064 269356 375070 269368
rect 393406 269356 393412 269368
rect 393464 269356 393470 269408
rect 393590 269356 393596 269408
rect 393648 269396 393654 269408
rect 398282 269396 398288 269408
rect 393648 269368 398288 269396
rect 393648 269356 393654 269368
rect 398282 269356 398288 269368
rect 398340 269356 398346 269408
rect 398466 269356 398472 269408
rect 398524 269396 398530 269408
rect 407776 269396 407804 269504
rect 407942 269492 407948 269544
rect 408000 269532 408006 269544
rect 422570 269532 422576 269544
rect 408000 269504 422576 269532
rect 408000 269492 408006 269504
rect 422570 269492 422576 269504
rect 422628 269492 422634 269544
rect 500034 269532 500040 269544
rect 422956 269504 500040 269532
rect 422956 269464 422984 269504
rect 500034 269492 500040 269504
rect 500092 269492 500098 269544
rect 500218 269492 500224 269544
rect 500276 269532 500282 269544
rect 543182 269532 543188 269544
rect 500276 269504 543188 269532
rect 500276 269492 500282 269504
rect 543182 269492 543188 269504
rect 543240 269492 543246 269544
rect 422772 269436 422984 269464
rect 412910 269396 412916 269408
rect 398524 269368 407712 269396
rect 407776 269368 412916 269396
rect 398524 269356 398530 269368
rect 354646 269232 369854 269260
rect 248322 269084 248328 269136
rect 248380 269124 248386 269136
rect 249978 269124 249984 269136
rect 248380 269096 249984 269124
rect 248380 269084 248386 269096
rect 249978 269084 249984 269096
rect 250036 269084 250042 269136
rect 274634 269084 274640 269136
rect 274692 269124 274698 269136
rect 278958 269124 278964 269136
rect 274692 269096 278964 269124
rect 274692 269084 274698 269096
rect 278958 269084 278964 269096
rect 279016 269084 279022 269136
rect 369826 269124 369854 269232
rect 372522 269220 372528 269272
rect 372580 269260 372586 269272
rect 406102 269260 406108 269272
rect 372580 269232 406108 269260
rect 372580 269220 372586 269232
rect 406102 269220 406108 269232
rect 406160 269220 406166 269272
rect 407684 269260 407712 269368
rect 412910 269356 412916 269368
rect 412968 269356 412974 269408
rect 413094 269356 413100 269408
rect 413152 269396 413158 269408
rect 413922 269396 413928 269408
rect 413152 269368 413928 269396
rect 413152 269356 413158 269368
rect 413922 269356 413928 269368
rect 413980 269356 413986 269408
rect 414106 269356 414112 269408
rect 414164 269396 414170 269408
rect 422772 269396 422800 269436
rect 414164 269368 422800 269396
rect 414164 269356 414170 269368
rect 423122 269356 423128 269408
rect 423180 269396 423186 269408
rect 423674 269396 423680 269408
rect 423180 269368 423680 269396
rect 423180 269356 423186 269368
rect 423674 269356 423680 269368
rect 423732 269356 423738 269408
rect 424410 269356 424416 269408
rect 424468 269396 424474 269408
rect 427630 269396 427636 269408
rect 424468 269368 427636 269396
rect 424468 269356 424474 269368
rect 427630 269356 427636 269368
rect 427688 269356 427694 269408
rect 427814 269356 427820 269408
rect 427872 269396 427878 269408
rect 521654 269396 521660 269408
rect 427872 269368 521660 269396
rect 427872 269356 427878 269368
rect 521654 269356 521660 269368
rect 521712 269356 521718 269408
rect 408126 269260 408132 269272
rect 407684 269232 408132 269260
rect 408126 269220 408132 269232
rect 408184 269220 408190 269272
rect 408310 269220 408316 269272
rect 408368 269260 408374 269272
rect 412450 269260 412456 269272
rect 408368 269232 412456 269260
rect 408368 269220 408374 269232
rect 412450 269220 412456 269232
rect 412508 269220 412514 269272
rect 412726 269220 412732 269272
rect 412784 269260 412790 269272
rect 416406 269260 416412 269272
rect 412784 269232 416412 269260
rect 412784 269220 412790 269232
rect 416406 269220 416412 269232
rect 416464 269220 416470 269272
rect 513374 269260 513380 269272
rect 418126 269232 513380 269260
rect 416682 269152 416688 269204
rect 416740 269192 416746 269204
rect 418126 269192 418154 269232
rect 513374 269220 513380 269232
rect 513432 269220 513438 269272
rect 416740 269164 418154 269192
rect 416740 269152 416746 269164
rect 372706 269124 372712 269136
rect 369826 269096 372712 269124
rect 372706 269084 372712 269096
rect 372764 269084 372770 269136
rect 373902 269084 373908 269136
rect 373960 269124 373966 269136
rect 375006 269124 375012 269136
rect 373960 269096 375012 269124
rect 373960 269084 373966 269096
rect 375006 269084 375012 269096
rect 375064 269084 375070 269136
rect 376938 269124 376944 269136
rect 375208 269096 376944 269124
rect 42334 269016 42340 269068
rect 42392 269056 42398 269068
rect 45554 269056 45560 269068
rect 42392 269028 45560 269056
rect 42392 269016 42398 269028
rect 45554 269016 45560 269028
rect 45612 269016 45618 269068
rect 118602 269016 118608 269068
rect 118660 269056 118666 269068
rect 169754 269056 169760 269068
rect 118660 269028 169760 269056
rect 118660 269016 118666 269028
rect 169754 269016 169760 269028
rect 169812 269016 169818 269068
rect 225414 269016 225420 269068
rect 225472 269056 225478 269068
rect 227622 269056 227628 269068
rect 225472 269028 227628 269056
rect 225472 269016 225478 269028
rect 227622 269016 227628 269028
rect 227680 269016 227686 269068
rect 324314 269016 324320 269068
rect 324372 269056 324378 269068
rect 336734 269056 336740 269068
rect 324372 269028 336740 269056
rect 324372 269016 324378 269028
rect 336734 269016 336740 269028
rect 336792 269016 336798 269068
rect 338482 269016 338488 269068
rect 338540 269056 338546 269068
rect 359090 269056 359096 269068
rect 338540 269028 359096 269056
rect 338540 269016 338546 269028
rect 359090 269016 359096 269028
rect 359148 269016 359154 269068
rect 269114 268948 269120 269000
rect 269172 268988 269178 269000
rect 276658 268988 276664 269000
rect 269172 268960 276664 268988
rect 269172 268948 269178 268960
rect 276658 268948 276664 268960
rect 276716 268948 276722 269000
rect 374454 268948 374460 269000
rect 374512 268988 374518 269000
rect 375208 268988 375236 269096
rect 376938 269084 376944 269096
rect 376996 269084 377002 269136
rect 378042 269016 378048 269068
rect 378100 269056 378106 269068
rect 384298 269056 384304 269068
rect 378100 269028 384304 269056
rect 378100 269016 378106 269028
rect 384298 269016 384304 269028
rect 384356 269016 384362 269068
rect 384482 269016 384488 269068
rect 384540 269056 384546 269068
rect 398098 269056 398104 269068
rect 384540 269028 398104 269056
rect 384540 269016 384546 269028
rect 398098 269016 398104 269028
rect 398156 269016 398162 269068
rect 398282 269016 398288 269068
rect 398340 269056 398346 269068
rect 466270 269056 466276 269068
rect 398340 269028 466276 269056
rect 398340 269016 398346 269028
rect 466270 269016 466276 269028
rect 466328 269016 466334 269068
rect 466454 269016 466460 269068
rect 466512 269056 466518 269068
rect 468110 269056 468116 269068
rect 466512 269028 468116 269056
rect 466512 269016 466518 269028
rect 468110 269016 468116 269028
rect 468168 269016 468174 269068
rect 471238 269016 471244 269068
rect 471296 269056 471302 269068
rect 587894 269056 587900 269068
rect 471296 269028 587900 269056
rect 471296 269016 471302 269028
rect 587894 269016 587900 269028
rect 587952 269016 587958 269068
rect 374512 268960 375236 268988
rect 374512 268948 374518 268960
rect 104894 268880 104900 268932
rect 104952 268920 104958 268932
rect 160186 268920 160192 268932
rect 104952 268892 160192 268920
rect 104952 268880 104958 268892
rect 160186 268880 160192 268892
rect 160244 268880 160250 268932
rect 187510 268880 187516 268932
rect 187568 268920 187574 268932
rect 208486 268920 208492 268932
rect 187568 268892 208492 268920
rect 187568 268880 187574 268892
rect 208486 268880 208492 268892
rect 208544 268880 208550 268932
rect 304166 268880 304172 268932
rect 304224 268920 304230 268932
rect 329834 268920 329840 268932
rect 304224 268892 329840 268920
rect 304224 268880 304230 268892
rect 329834 268880 329840 268892
rect 329892 268880 329898 268932
rect 347406 268880 347412 268932
rect 347464 268920 347470 268932
rect 347464 268892 369854 268920
rect 347464 268880 347470 268892
rect 77202 268744 77208 268796
rect 77260 268784 77266 268796
rect 104894 268784 104900 268796
rect 77260 268756 104900 268784
rect 77260 268744 77266 268756
rect 104894 268744 104900 268756
rect 104952 268744 104958 268796
rect 106274 268744 106280 268796
rect 106332 268784 106338 268796
rect 161658 268784 161664 268796
rect 106332 268756 161664 268784
rect 106332 268744 106338 268756
rect 161658 268744 161664 268756
rect 161716 268744 161722 268796
rect 166166 268744 166172 268796
rect 166224 268784 166230 268796
rect 194042 268784 194048 268796
rect 166224 268756 194048 268784
rect 166224 268744 166230 268756
rect 194042 268744 194048 268756
rect 194100 268744 194106 268796
rect 203886 268744 203892 268796
rect 203944 268784 203950 268796
rect 211154 268784 211160 268796
rect 203944 268756 211160 268784
rect 203944 268744 203950 268756
rect 211154 268744 211160 268756
rect 211212 268744 211218 268796
rect 284570 268744 284576 268796
rect 284628 268784 284634 268796
rect 285858 268784 285864 268796
rect 284628 268756 285864 268784
rect 284628 268744 284634 268756
rect 285858 268744 285864 268756
rect 285916 268744 285922 268796
rect 314746 268744 314752 268796
rect 314804 268784 314810 268796
rect 352098 268784 352104 268796
rect 314804 268756 352104 268784
rect 314804 268744 314810 268756
rect 352098 268744 352104 268756
rect 352156 268744 352162 268796
rect 369826 268784 369854 268892
rect 375834 268880 375840 268932
rect 375892 268920 375898 268932
rect 449894 268920 449900 268932
rect 375892 268892 449900 268920
rect 375892 268880 375898 268892
rect 449894 268880 449900 268892
rect 449952 268880 449958 268932
rect 455322 268880 455328 268932
rect 455380 268920 455386 268932
rect 461394 268920 461400 268932
rect 455380 268892 461400 268920
rect 455380 268880 455386 268892
rect 461394 268880 461400 268892
rect 461452 268880 461458 268932
rect 462498 268880 462504 268932
rect 462556 268920 462562 268932
rect 580994 268920 581000 268932
rect 462556 268892 581000 268920
rect 462556 268880 462562 268892
rect 580994 268880 581000 268892
rect 581052 268880 581058 268932
rect 376018 268784 376024 268796
rect 369826 268756 376024 268784
rect 376018 268744 376024 268756
rect 376076 268744 376082 268796
rect 384298 268744 384304 268796
rect 384356 268784 384362 268796
rect 440418 268784 440424 268796
rect 384356 268756 440424 268784
rect 384356 268744 384362 268756
rect 440418 268744 440424 268756
rect 440476 268744 440482 268796
rect 460106 268784 460112 268796
rect 440620 268756 460112 268784
rect 95418 268608 95424 268660
rect 95476 268648 95482 268660
rect 155034 268648 155040 268660
rect 95476 268620 155040 268648
rect 95476 268608 95482 268620
rect 155034 268608 155040 268620
rect 155092 268608 155098 268660
rect 162578 268608 162584 268660
rect 162636 268648 162642 268660
rect 190086 268648 190092 268660
rect 162636 268620 190092 268648
rect 162636 268608 162642 268620
rect 190086 268608 190092 268620
rect 190144 268608 190150 268660
rect 190362 268608 190368 268660
rect 190420 268648 190426 268660
rect 204070 268648 204076 268660
rect 190420 268620 204076 268648
rect 190420 268608 190426 268620
rect 204070 268608 204076 268620
rect 204128 268608 204134 268660
rect 285766 268608 285772 268660
rect 285824 268648 285830 268660
rect 295334 268648 295340 268660
rect 285824 268620 295340 268648
rect 285824 268608 285830 268620
rect 295334 268608 295340 268620
rect 295392 268608 295398 268660
rect 299290 268608 299296 268660
rect 299348 268648 299354 268660
rect 316770 268648 316776 268660
rect 299348 268620 316776 268648
rect 299348 268608 299354 268620
rect 316770 268608 316776 268620
rect 316828 268608 316834 268660
rect 317690 268608 317696 268660
rect 317748 268648 317754 268660
rect 355686 268648 355692 268660
rect 317748 268620 355692 268648
rect 317748 268608 317754 268620
rect 355686 268608 355692 268620
rect 355744 268608 355750 268660
rect 369210 268608 369216 268660
rect 369268 268648 369274 268660
rect 437290 268648 437296 268660
rect 369268 268620 437296 268648
rect 369268 268608 369274 268620
rect 437290 268608 437296 268620
rect 437348 268608 437354 268660
rect 437428 268608 437434 268660
rect 437486 268648 437492 268660
rect 440620 268648 440648 268756
rect 460106 268744 460112 268756
rect 460164 268744 460170 268796
rect 583846 268784 583852 268796
rect 461780 268756 583852 268784
rect 456426 268648 456432 268660
rect 437486 268620 440648 268648
rect 440712 268620 456432 268648
rect 437486 268608 437492 268620
rect 87138 268472 87144 268524
rect 87196 268512 87202 268524
rect 149882 268512 149888 268524
rect 87196 268484 149888 268512
rect 87196 268472 87202 268484
rect 149882 268472 149888 268484
rect 149940 268472 149946 268524
rect 162762 268472 162768 268524
rect 162820 268512 162826 268524
rect 196986 268512 196992 268524
rect 162820 268484 196992 268512
rect 162820 268472 162826 268484
rect 196986 268472 196992 268484
rect 197044 268472 197050 268524
rect 208854 268472 208860 268524
rect 208912 268512 208918 268524
rect 225690 268512 225696 268524
rect 208912 268484 225696 268512
rect 208912 268472 208918 268484
rect 225690 268472 225696 268484
rect 225748 268472 225754 268524
rect 281626 268472 281632 268524
rect 281684 268512 281690 268524
rect 295518 268512 295524 268524
rect 281684 268484 295524 268512
rect 281684 268472 281690 268484
rect 295518 268472 295524 268484
rect 295576 268472 295582 268524
rect 297082 268472 297088 268524
rect 297140 268512 297146 268524
rect 322934 268512 322940 268524
rect 297140 268484 322940 268512
rect 297140 268472 297146 268484
rect 322934 268472 322940 268484
rect 322992 268472 322998 268524
rect 329466 268472 329472 268524
rect 329524 268512 329530 268524
rect 340874 268512 340880 268524
rect 329524 268484 340880 268512
rect 329524 268472 329530 268484
rect 340874 268472 340880 268484
rect 340932 268472 340938 268524
rect 349338 268472 349344 268524
rect 349396 268512 349402 268524
rect 371050 268512 371056 268524
rect 349396 268484 371056 268512
rect 349396 268472 349402 268484
rect 371050 268472 371056 268484
rect 371108 268472 371114 268524
rect 371418 268472 371424 268524
rect 371476 268512 371482 268524
rect 432598 268512 432604 268524
rect 371476 268484 432604 268512
rect 371476 268472 371482 268484
rect 432598 268472 432604 268484
rect 432656 268472 432662 268524
rect 434714 268472 434720 268524
rect 434772 268512 434778 268524
rect 440712 268512 440740 268620
rect 456426 268608 456432 268620
rect 456484 268608 456490 268660
rect 460290 268608 460296 268660
rect 460348 268648 460354 268660
rect 461780 268648 461808 268756
rect 583846 268744 583852 268756
rect 583904 268744 583910 268796
rect 460348 268620 461808 268648
rect 460348 268608 460354 268620
rect 461946 268608 461952 268660
rect 462004 268648 462010 268660
rect 462004 268620 466684 268648
rect 462004 268608 462010 268620
rect 434772 268484 440740 268512
rect 434772 268472 434778 268484
rect 440878 268472 440884 268524
rect 440936 268512 440942 268524
rect 442810 268512 442816 268524
rect 440936 268484 442816 268512
rect 440936 268472 440942 268484
rect 442810 268472 442816 268484
rect 442868 268472 442874 268524
rect 442994 268472 443000 268524
rect 443052 268512 443058 268524
rect 456426 268512 456432 268524
rect 443052 268484 456432 268512
rect 443052 268472 443058 268484
rect 456426 268472 456432 268484
rect 456484 268472 456490 268524
rect 456978 268472 456984 268524
rect 457036 268512 457042 268524
rect 466408 268512 466414 268524
rect 457036 268484 466414 268512
rect 457036 268472 457042 268484
rect 466408 268472 466414 268484
rect 466466 268472 466472 268524
rect 466656 268512 466684 268620
rect 467098 268608 467104 268660
rect 467156 268648 467162 268660
rect 594794 268648 594800 268660
rect 467156 268620 594800 268648
rect 467156 268608 467162 268620
rect 594794 268608 594800 268620
rect 594852 268608 594858 268660
rect 594978 268608 594984 268660
rect 595036 268648 595042 268660
rect 645854 268648 645860 268660
rect 595036 268620 645860 268648
rect 595036 268608 595042 268620
rect 645854 268608 645860 268620
rect 645912 268608 645918 268660
rect 471238 268512 471244 268524
rect 466656 268484 471244 268512
rect 471238 268472 471244 268484
rect 471296 268472 471302 268524
rect 471422 268472 471428 268524
rect 471480 268512 471486 268524
rect 474734 268512 474740 268524
rect 471480 268484 474740 268512
rect 471480 268472 471486 268484
rect 474734 268472 474740 268484
rect 474792 268472 474798 268524
rect 475194 268472 475200 268524
rect 475252 268512 475258 268524
rect 608686 268512 608692 268524
rect 475252 268484 608692 268512
rect 475252 268472 475258 268484
rect 608686 268472 608692 268484
rect 608744 268472 608750 268524
rect 669314 268472 669320 268524
rect 669372 268512 669378 268524
rect 675478 268512 675484 268524
rect 669372 268484 675484 268512
rect 669372 268472 669378 268484
rect 675478 268472 675484 268484
rect 675536 268472 675542 268524
rect 82722 268336 82728 268388
rect 82780 268376 82786 268388
rect 146938 268376 146944 268388
rect 82780 268348 146944 268376
rect 82780 268336 82786 268348
rect 146938 268336 146944 268348
rect 146996 268336 147002 268388
rect 148870 268336 148876 268388
rect 148928 268376 148934 268388
rect 188154 268376 188160 268388
rect 148928 268348 188160 268376
rect 148928 268336 148934 268348
rect 188154 268336 188160 268348
rect 188212 268336 188218 268388
rect 188430 268336 188436 268388
rect 188488 268376 188494 268388
rect 188488 268348 200114 268376
rect 188488 268336 188494 268348
rect 115750 268200 115756 268252
rect 115808 268240 115814 268252
rect 166810 268240 166816 268252
rect 115808 268212 166816 268240
rect 115808 268200 115814 268212
rect 166810 268200 166816 268212
rect 166868 268200 166874 268252
rect 200086 268240 200114 268348
rect 210970 268336 210976 268388
rect 211028 268376 211034 268388
rect 219802 268376 219808 268388
rect 211028 268348 219808 268376
rect 211028 268336 211034 268348
rect 219802 268336 219808 268348
rect 219860 268336 219866 268388
rect 220722 268336 220728 268388
rect 220780 268376 220786 268388
rect 230750 268376 230756 268388
rect 220780 268348 230756 268376
rect 220780 268336 220786 268348
rect 230750 268336 230756 268348
rect 230808 268336 230814 268388
rect 273530 268336 273536 268388
rect 273588 268376 273594 268388
rect 282914 268376 282920 268388
rect 273588 268348 282920 268376
rect 273588 268336 273594 268348
rect 282914 268336 282920 268348
rect 282972 268336 282978 268388
rect 286778 268336 286784 268388
rect 286836 268376 286842 268388
rect 306374 268376 306380 268388
rect 286836 268348 306380 268376
rect 286836 268336 286842 268348
rect 306374 268336 306380 268348
rect 306432 268336 306438 268388
rect 316954 268336 316960 268388
rect 317012 268376 317018 268388
rect 354674 268376 354680 268388
rect 317012 268348 354680 268376
rect 317012 268336 317018 268348
rect 354674 268336 354680 268348
rect 354732 268336 354738 268388
rect 358538 268336 358544 268388
rect 358596 268376 358602 268388
rect 407390 268376 407396 268388
rect 358596 268348 407396 268376
rect 358596 268336 358602 268348
rect 407390 268336 407396 268348
rect 407448 268336 407454 268388
rect 417418 268376 417424 268388
rect 407776 268348 417424 268376
rect 210970 268240 210976 268252
rect 200086 268212 210976 268240
rect 210970 268200 210976 268212
rect 211028 268200 211034 268252
rect 324682 268200 324688 268252
rect 324740 268240 324746 268252
rect 367094 268240 367100 268252
rect 324740 268212 367100 268240
rect 324740 268200 324746 268212
rect 367094 268200 367100 268212
rect 367152 268200 367158 268252
rect 382458 268200 382464 268252
rect 382516 268240 382522 268252
rect 384482 268240 384488 268252
rect 382516 268212 384488 268240
rect 382516 268200 382522 268212
rect 384482 268200 384488 268212
rect 384540 268200 384546 268252
rect 387610 268200 387616 268252
rect 387668 268240 387674 268252
rect 397914 268240 397920 268252
rect 387668 268212 397920 268240
rect 387668 268200 387674 268212
rect 397914 268200 397920 268212
rect 397972 268200 397978 268252
rect 398098 268200 398104 268252
rect 398156 268240 398162 268252
rect 407776 268240 407804 268348
rect 417418 268336 417424 268348
rect 417476 268336 417482 268388
rect 417602 268336 417608 268388
rect 417660 268376 417666 268388
rect 456610 268376 456616 268388
rect 417660 268348 456616 268376
rect 417660 268336 417666 268348
rect 456610 268336 456616 268348
rect 456668 268336 456674 268388
rect 456794 268336 456800 268388
rect 456852 268376 456858 268388
rect 495066 268376 495072 268388
rect 456852 268348 495072 268376
rect 456852 268336 456858 268348
rect 495066 268336 495072 268348
rect 495124 268336 495130 268388
rect 495526 268336 495532 268388
rect 495584 268376 495590 268388
rect 504910 268376 504916 268388
rect 495584 268348 504916 268376
rect 495584 268336 495590 268348
rect 504910 268336 504916 268348
rect 504968 268336 504974 268388
rect 505048 268336 505054 268388
rect 505106 268376 505112 268388
rect 607214 268376 607220 268388
rect 505106 268348 607220 268376
rect 505106 268336 505112 268348
rect 607214 268336 607220 268348
rect 607272 268336 607278 268388
rect 675478 268308 675484 268320
rect 669286 268280 675484 268308
rect 398156 268212 407804 268240
rect 398156 268200 398162 268212
rect 407942 268200 407948 268252
rect 408000 268240 408006 268252
rect 446766 268240 446772 268252
rect 408000 268212 446772 268240
rect 408000 268200 408006 268212
rect 446766 268200 446772 268212
rect 446824 268200 446830 268252
rect 452378 268200 452384 268252
rect 452436 268240 452442 268252
rect 456610 268240 456616 268252
rect 452436 268212 456616 268240
rect 452436 268200 452442 268212
rect 456610 268200 456616 268212
rect 456668 268200 456674 268252
rect 461578 268200 461584 268252
rect 461636 268240 461642 268252
rect 480898 268240 480904 268252
rect 461636 268212 480904 268240
rect 461636 268200 461642 268212
rect 480898 268200 480904 268212
rect 480956 268200 480962 268252
rect 481082 268200 481088 268252
rect 481140 268240 481146 268252
rect 484854 268240 484860 268252
rect 481140 268212 484860 268240
rect 481140 268200 481146 268212
rect 484854 268200 484860 268212
rect 484912 268200 484918 268252
rect 485682 268200 485688 268252
rect 485740 268240 485746 268252
rect 485866 268240 485872 268252
rect 485740 268212 485872 268240
rect 485740 268200 485746 268212
rect 485866 268200 485872 268212
rect 485924 268200 485930 268252
rect 486050 268200 486056 268252
rect 486108 268240 486114 268252
rect 572714 268240 572720 268252
rect 486108 268212 572720 268240
rect 486108 268200 486114 268212
rect 572714 268200 572720 268212
rect 572772 268200 572778 268252
rect 135254 268064 135260 268116
rect 135312 268104 135318 268116
rect 138106 268104 138112 268116
rect 135312 268076 138112 268104
rect 135312 268064 135318 268076
rect 138106 268064 138112 268076
rect 138164 268064 138170 268116
rect 147490 268064 147496 268116
rect 147548 268104 147554 268116
rect 186682 268104 186688 268116
rect 147548 268076 186688 268104
rect 147548 268064 147554 268076
rect 186682 268064 186688 268076
rect 186740 268064 186746 268116
rect 365346 268064 365352 268116
rect 365404 268104 365410 268116
rect 432046 268104 432052 268116
rect 365404 268076 432052 268104
rect 365404 268064 365410 268076
rect 432046 268064 432052 268076
rect 432104 268064 432110 268116
rect 432598 268064 432604 268116
rect 432656 268104 432662 268116
rect 440234 268104 440240 268116
rect 432656 268076 440240 268104
rect 432656 268064 432662 268076
rect 440234 268064 440240 268076
rect 440292 268064 440298 268116
rect 440418 268064 440424 268116
rect 440476 268104 440482 268116
rect 452654 268104 452660 268116
rect 440476 268076 452660 268104
rect 440476 268064 440482 268076
rect 452654 268064 452660 268076
rect 452712 268064 452718 268116
rect 457530 268064 457536 268116
rect 457588 268104 457594 268116
rect 461026 268104 461032 268116
rect 457588 268076 461032 268104
rect 457588 268064 457594 268076
rect 461026 268064 461032 268076
rect 461084 268064 461090 268116
rect 461394 268064 461400 268116
rect 461452 268104 461458 268116
rect 484670 268104 484676 268116
rect 461452 268076 484676 268104
rect 461452 268064 461458 268076
rect 484670 268064 484676 268076
rect 484728 268064 484734 268116
rect 486418 268064 486424 268116
rect 486476 268104 486482 268116
rect 563054 268104 563060 268116
rect 486476 268076 563060 268104
rect 486476 268064 486482 268076
rect 563054 268064 563060 268076
rect 563112 268064 563118 268116
rect 658918 267996 658924 268048
rect 658976 268036 658982 268048
rect 669286 268036 669314 268280
rect 675478 268268 675484 268280
rect 675536 268268 675542 268320
rect 658976 268008 669314 268036
rect 658976 267996 658982 268008
rect 354674 267928 354680 267980
rect 354732 267968 354738 267980
rect 354732 267940 393314 267968
rect 354732 267928 354738 267940
rect 143442 267832 143448 267844
rect 142632 267804 143448 267832
rect 137554 267764 137560 267776
rect 135732 267736 137560 267764
rect 42518 267656 42524 267708
rect 42576 267696 42582 267708
rect 45922 267696 45928 267708
rect 42576 267668 45928 267696
rect 42576 267656 42582 267668
rect 45922 267656 45928 267668
rect 45980 267656 45986 267708
rect 104894 267656 104900 267708
rect 104952 267696 104958 267708
rect 135732 267696 135760 267736
rect 137554 267724 137560 267736
rect 137612 267724 137618 267776
rect 104952 267668 135760 267696
rect 104952 267656 104958 267668
rect 140038 267656 140044 267708
rect 140096 267696 140102 267708
rect 142632 267696 142660 267804
rect 143442 267792 143448 267804
rect 143500 267792 143506 267844
rect 355962 267792 355968 267844
rect 356020 267832 356026 267844
rect 388990 267832 388996 267844
rect 356020 267804 388996 267832
rect 356020 267792 356026 267804
rect 388990 267792 388996 267804
rect 389048 267792 389054 267844
rect 393286 267832 393314 267940
rect 402606 267928 402612 267980
rect 402664 267968 402670 267980
rect 407942 267968 407948 267980
rect 402664 267940 407948 267968
rect 402664 267928 402670 267940
rect 407942 267928 407948 267940
rect 408000 267928 408006 267980
rect 411162 267928 411168 267980
rect 411220 267968 411226 267980
rect 411220 267940 417280 267968
rect 411220 267928 411226 267940
rect 404446 267832 404452 267844
rect 393286 267804 404452 267832
rect 404446 267792 404452 267804
rect 404504 267792 404510 267844
rect 407390 267792 407396 267844
rect 407448 267832 407454 267844
rect 410058 267832 410064 267844
rect 407448 267804 410064 267832
rect 407448 267792 407454 267804
rect 410058 267792 410064 267804
rect 410116 267792 410122 267844
rect 410242 267792 410248 267844
rect 410300 267832 410306 267844
rect 415302 267832 415308 267844
rect 410300 267804 410932 267832
rect 410300 267792 410306 267804
rect 263962 267724 263968 267776
rect 264020 267764 264026 267776
rect 269574 267764 269580 267776
rect 264020 267736 269580 267764
rect 264020 267724 264026 267736
rect 269574 267724 269580 267736
rect 269632 267724 269638 267776
rect 344186 267724 344192 267776
rect 344244 267764 344250 267776
rect 347038 267764 347044 267776
rect 344244 267736 347044 267764
rect 344244 267724 344250 267736
rect 347038 267724 347044 267736
rect 347096 267724 347102 267776
rect 140096 267668 142660 267696
rect 140096 267656 140102 267668
rect 142798 267656 142804 267708
rect 142856 267696 142862 267708
rect 166074 267696 166080 267708
rect 142856 267668 166080 267696
rect 142856 267656 142862 267668
rect 166074 267656 166080 267668
rect 166132 267656 166138 267708
rect 213178 267656 213184 267708
rect 213236 267696 213242 267708
rect 220538 267696 220544 267708
rect 213236 267668 220544 267696
rect 213236 267656 213242 267668
rect 220538 267656 220544 267668
rect 220596 267656 220602 267708
rect 288250 267656 288256 267708
rect 288308 267696 288314 267708
rect 297358 267696 297364 267708
rect 288308 267668 297364 267696
rect 288308 267656 288314 267668
rect 297358 267656 297364 267668
rect 297416 267656 297422 267708
rect 305914 267656 305920 267708
rect 305972 267696 305978 267708
rect 324314 267696 324320 267708
rect 305972 267668 324320 267696
rect 305972 267656 305978 267668
rect 324314 267656 324320 267668
rect 324372 267656 324378 267708
rect 349816 267668 364656 267696
rect 343358 267588 343364 267640
rect 343416 267628 343422 267640
rect 349816 267628 349844 267668
rect 343416 267600 349844 267628
rect 343416 267588 343422 267600
rect 132402 267520 132408 267572
rect 132460 267560 132466 267572
rect 178586 267560 178592 267572
rect 132460 267532 178592 267560
rect 132460 267520 132466 267532
rect 178586 267520 178592 267532
rect 178644 267520 178650 267572
rect 180058 267520 180064 267572
rect 180116 267560 180122 267572
rect 207290 267560 207296 267572
rect 180116 267532 207296 267560
rect 180116 267520 180122 267532
rect 207290 267520 207296 267532
rect 207348 267520 207354 267572
rect 286042 267520 286048 267572
rect 286100 267560 286106 267572
rect 290458 267560 290464 267572
rect 286100 267532 290464 267560
rect 286100 267520 286106 267532
rect 290458 267520 290464 267532
rect 290516 267520 290522 267572
rect 294874 267520 294880 267572
rect 294932 267560 294938 267572
rect 300118 267560 300124 267572
rect 294932 267532 300124 267560
rect 294932 267520 294938 267532
rect 300118 267520 300124 267532
rect 300176 267520 300182 267572
rect 319162 267520 319168 267572
rect 319220 267560 319226 267572
rect 338482 267560 338488 267572
rect 319220 267532 338488 267560
rect 319220 267520 319226 267532
rect 338482 267520 338488 267532
rect 338540 267520 338546 267572
rect 350258 267520 350264 267572
rect 350316 267560 350322 267572
rect 364150 267560 364156 267572
rect 350316 267532 364156 267560
rect 350316 267520 350322 267532
rect 364150 267520 364156 267532
rect 364208 267520 364214 267572
rect 364628 267560 364656 267668
rect 364794 267656 364800 267708
rect 364852 267696 364858 267708
rect 372522 267696 372528 267708
rect 364852 267668 372528 267696
rect 364852 267656 364858 267668
rect 372522 267656 372528 267668
rect 372580 267656 372586 267708
rect 372890 267656 372896 267708
rect 372948 267696 372954 267708
rect 372948 267668 374868 267696
rect 372948 267656 372954 267668
rect 365714 267560 365720 267572
rect 364628 267532 365720 267560
rect 365714 267520 365720 267532
rect 365772 267520 365778 267572
rect 366266 267520 366272 267572
rect 366324 267560 366330 267572
rect 374454 267560 374460 267572
rect 366324 267532 374460 267560
rect 366324 267520 366330 267532
rect 374454 267520 374460 267532
rect 374512 267520 374518 267572
rect 374840 267560 374868 267668
rect 375006 267656 375012 267708
rect 375064 267696 375070 267708
rect 410702 267696 410708 267708
rect 375064 267668 410708 267696
rect 375064 267656 375070 267668
rect 410702 267656 410708 267668
rect 410760 267656 410766 267708
rect 410904 267696 410932 267804
rect 414676 267804 415308 267832
rect 414676 267696 414704 267804
rect 415302 267792 415308 267804
rect 415360 267792 415366 267844
rect 417252 267832 417280 267940
rect 417418 267928 417424 267980
rect 417476 267968 417482 267980
rect 427630 267968 427636 267980
rect 417476 267940 427636 267968
rect 417476 267928 417482 267940
rect 427630 267928 427636 267940
rect 427688 267928 427694 267980
rect 427814 267928 427820 267980
rect 427872 267968 427878 267980
rect 437290 267968 437296 267980
rect 427872 267940 437296 267968
rect 427872 267928 427878 267940
rect 437290 267928 437296 267940
rect 437348 267928 437354 267980
rect 437428 267928 437434 267980
rect 437486 267968 437492 267980
rect 541342 267968 541348 267980
rect 437486 267940 541348 267968
rect 437486 267928 437492 267940
rect 541342 267928 541348 267940
rect 541400 267928 541406 267980
rect 660298 267860 660304 267912
rect 660356 267900 660362 267912
rect 669314 267900 669320 267912
rect 660356 267872 669320 267900
rect 660356 267860 660362 267872
rect 669314 267860 669320 267872
rect 669372 267860 669378 267912
rect 417602 267832 417608 267844
rect 417252 267804 417608 267832
rect 417602 267792 417608 267804
rect 417660 267792 417666 267844
rect 417786 267792 417792 267844
rect 417844 267832 417850 267844
rect 422294 267832 422300 267844
rect 417844 267804 422300 267832
rect 417844 267792 417850 267804
rect 422294 267792 422300 267804
rect 422352 267792 422358 267844
rect 422938 267792 422944 267844
rect 422996 267832 423002 267844
rect 475746 267832 475752 267844
rect 422996 267804 475752 267832
rect 422996 267792 423002 267804
rect 475746 267792 475752 267804
rect 475804 267792 475810 267844
rect 476206 267792 476212 267844
rect 476264 267832 476270 267844
rect 480714 267832 480720 267844
rect 476264 267804 480720 267832
rect 476264 267792 476270 267804
rect 480714 267792 480720 267804
rect 480772 267792 480778 267844
rect 480898 267792 480904 267844
rect 480956 267832 480962 267844
rect 485038 267832 485044 267844
rect 480956 267804 485044 267832
rect 480956 267792 480962 267804
rect 485038 267792 485044 267804
rect 485096 267792 485102 267844
rect 486234 267792 486240 267844
rect 486292 267832 486298 267844
rect 494514 267832 494520 267844
rect 486292 267804 494520 267832
rect 486292 267792 486298 267804
rect 494514 267792 494520 267804
rect 494572 267792 494578 267844
rect 524690 267832 524696 267844
rect 494716 267804 524696 267832
rect 410904 267668 414704 267696
rect 415302 267656 415308 267708
rect 415360 267696 415366 267708
rect 417878 267696 417884 267708
rect 415360 267668 417884 267696
rect 415360 267656 415366 267668
rect 417878 267656 417884 267668
rect 417936 267656 417942 267708
rect 418338 267656 418344 267708
rect 418396 267696 418402 267708
rect 490190 267696 490196 267708
rect 418396 267668 490196 267696
rect 418396 267656 418402 267668
rect 490190 267656 490196 267668
rect 490248 267656 490254 267708
rect 491386 267656 491392 267708
rect 491444 267696 491450 267708
rect 492582 267696 492588 267708
rect 491444 267668 492588 267696
rect 491444 267656 491450 267668
rect 492582 267656 492588 267668
rect 492640 267656 492646 267708
rect 492766 267656 492772 267708
rect 492824 267696 492830 267708
rect 494716 267696 494744 267804
rect 524690 267792 524696 267804
rect 524748 267792 524754 267844
rect 675478 267832 675484 267844
rect 669516 267804 675484 267832
rect 664806 267724 664812 267776
rect 664864 267764 664870 267776
rect 664864 267736 669360 267764
rect 664864 267724 664870 267736
rect 492824 267668 494744 267696
rect 492824 267656 492830 267668
rect 494882 267656 494888 267708
rect 494940 267696 494946 267708
rect 525978 267696 525984 267708
rect 494940 267668 525984 267696
rect 494940 267656 494946 267668
rect 525978 267656 525984 267668
rect 526036 267656 526042 267708
rect 669332 267696 669360 267736
rect 669516 267696 669544 267804
rect 675478 267792 675484 267804
rect 675536 267792 675542 267844
rect 669332 267668 669544 267696
rect 411990 267560 411996 267572
rect 374840 267532 411996 267560
rect 411990 267520 411996 267532
rect 412048 267520 412054 267572
rect 412174 267520 412180 267572
rect 412232 267560 412238 267572
rect 412588 267560 412594 267572
rect 412232 267532 412594 267560
rect 412232 267520 412238 267532
rect 412588 267520 412594 267532
rect 412646 267520 412652 267572
rect 412726 267520 412732 267572
rect 412784 267560 412790 267572
rect 414658 267560 414664 267572
rect 412784 267532 414664 267560
rect 412784 267520 412790 267532
rect 414658 267520 414664 267532
rect 414716 267520 414722 267572
rect 415302 267520 415308 267572
rect 415360 267560 415366 267572
rect 415360 267532 421328 267560
rect 415360 267520 415366 267532
rect 100662 267384 100668 267436
rect 100720 267424 100726 267436
rect 158714 267424 158720 267436
rect 100720 267396 158720 267424
rect 100720 267384 100726 267396
rect 158714 267384 158720 267396
rect 158772 267384 158778 267436
rect 162946 267384 162952 267436
rect 163004 267424 163010 267436
rect 163004 267396 174400 267424
rect 163004 267384 163010 267396
rect 78214 267248 78220 267300
rect 78272 267288 78278 267300
rect 137370 267288 137376 267300
rect 78272 267260 137376 267288
rect 78272 267248 78278 267260
rect 137370 267248 137376 267260
rect 137428 267248 137434 267300
rect 137554 267248 137560 267300
rect 137612 267288 137618 267300
rect 143258 267288 143264 267300
rect 137612 267260 143264 267288
rect 137612 267248 137618 267260
rect 143258 267248 143264 267260
rect 143316 267248 143322 267300
rect 143442 267248 143448 267300
rect 143500 267288 143506 267300
rect 173894 267288 173900 267300
rect 143500 267260 173900 267288
rect 143500 267248 143506 267260
rect 173894 267248 173900 267260
rect 173952 267248 173958 267300
rect 174372 267288 174400 267396
rect 175918 267384 175924 267436
rect 175976 267424 175982 267436
rect 202874 267424 202880 267436
rect 175976 267396 202880 267424
rect 175976 267384 175982 267396
rect 202874 267384 202880 267396
rect 202932 267384 202938 267436
rect 204070 267384 204076 267436
rect 204128 267424 204134 267436
rect 213178 267424 213184 267436
rect 204128 267396 213184 267424
rect 204128 267384 204134 267396
rect 213178 267384 213184 267396
rect 213236 267384 213242 267436
rect 222838 267384 222844 267436
rect 222896 267424 222902 267436
rect 231578 267424 231584 267436
rect 222896 267396 231584 267424
rect 222896 267384 222902 267396
rect 231578 267384 231584 267396
rect 231636 267384 231642 267436
rect 295610 267384 295616 267436
rect 295668 267424 295674 267436
rect 301958 267424 301964 267436
rect 295668 267396 301964 267424
rect 295668 267384 295674 267396
rect 301958 267384 301964 267396
rect 302016 267384 302022 267436
rect 308122 267384 308128 267436
rect 308180 267424 308186 267436
rect 329466 267424 329472 267436
rect 308180 267396 329472 267424
rect 308180 267384 308186 267396
rect 329466 267384 329472 267396
rect 329524 267384 329530 267436
rect 345842 267424 345848 267436
rect 335326 267396 345848 267424
rect 176378 267288 176384 267300
rect 174372 267260 176384 267288
rect 176378 267248 176384 267260
rect 176436 267248 176442 267300
rect 187418 267288 187424 267300
rect 180766 267260 187424 267288
rect 86218 267112 86224 267164
rect 86276 267152 86282 267164
rect 145926 267152 145932 267164
rect 86276 267124 145932 267152
rect 86276 267112 86282 267124
rect 145926 267112 145932 267124
rect 145984 267112 145990 267164
rect 146202 267112 146208 267164
rect 146260 267152 146266 267164
rect 180766 267152 180794 267260
rect 187418 267248 187424 267260
rect 187476 267248 187482 267300
rect 194502 267248 194508 267300
rect 194560 267288 194566 267300
rect 208762 267288 208768 267300
rect 194560 267260 208768 267288
rect 194560 267248 194566 267260
rect 208762 267248 208768 267260
rect 208820 267248 208826 267300
rect 228450 267248 228456 267300
rect 228508 267288 228514 267300
rect 233786 267288 233792 267300
rect 228508 267260 233792 267288
rect 228508 267248 228514 267260
rect 233786 267248 233792 267260
rect 233844 267248 233850 267300
rect 262858 267248 262864 267300
rect 262916 267288 262922 267300
rect 267918 267288 267924 267300
rect 262916 267260 267924 267288
rect 262916 267248 262922 267260
rect 267918 267248 267924 267260
rect 267976 267248 267982 267300
rect 275738 267248 275744 267300
rect 275796 267288 275802 267300
rect 280982 267288 280988 267300
rect 275796 267260 280988 267288
rect 275796 267248 275802 267260
rect 280982 267248 280988 267260
rect 281040 267248 281046 267300
rect 282362 267248 282368 267300
rect 282420 267288 282426 267300
rect 289078 267288 289084 267300
rect 282420 267260 289084 267288
rect 282420 267248 282426 267260
rect 289078 267248 289084 267260
rect 289136 267248 289142 267300
rect 302878 267288 302884 267300
rect 296686 267260 302884 267288
rect 257338 267180 257344 267232
rect 257396 267220 257402 267232
rect 259454 267220 259460 267232
rect 257396 267192 259460 267220
rect 257396 267180 257402 267192
rect 259454 267180 259460 267192
rect 259512 267180 259518 267232
rect 146260 267124 180794 267152
rect 146260 267112 146266 267124
rect 186958 267112 186964 267164
rect 187016 267152 187022 267164
rect 187016 267124 200114 267152
rect 187016 267112 187022 267124
rect 91002 266976 91008 267028
rect 91060 267016 91066 267028
rect 152090 267016 152096 267028
rect 91060 266988 152096 267016
rect 91060 266976 91066 266988
rect 152090 266976 152096 266988
rect 152148 266976 152154 267028
rect 156506 266976 156512 267028
rect 156564 267016 156570 267028
rect 165338 267016 165344 267028
rect 156564 266988 165344 267016
rect 156564 266976 156570 266988
rect 165338 266976 165344 266988
rect 165396 266976 165402 267028
rect 167914 266976 167920 267028
rect 167972 267016 167978 267028
rect 198458 267016 198464 267028
rect 167972 266988 198464 267016
rect 167972 266976 167978 266988
rect 198458 266976 198464 266988
rect 198516 266976 198522 267028
rect 200086 267016 200114 267124
rect 211154 267112 211160 267164
rect 211212 267152 211218 267164
rect 222746 267152 222752 267164
rect 211212 267124 222752 267152
rect 211212 267112 211218 267124
rect 222746 267112 222752 267124
rect 222804 267112 222810 267164
rect 233234 267112 233240 267164
rect 233292 267152 233298 267164
rect 240410 267152 240416 267164
rect 233292 267124 240416 267152
rect 233292 267112 233298 267124
rect 240410 267112 240416 267124
rect 240468 267112 240474 267164
rect 267642 267112 267648 267164
rect 267700 267152 267706 267164
rect 271138 267152 271144 267164
rect 267700 267124 271144 267152
rect 267700 267112 267706 267124
rect 271138 267112 271144 267124
rect 271196 267112 271202 267164
rect 272058 267112 272064 267164
rect 272116 267152 272122 267164
rect 280706 267152 280712 267164
rect 272116 267124 280712 267152
rect 272116 267112 272122 267124
rect 280706 267112 280712 267124
rect 280764 267112 280770 267164
rect 293402 267112 293408 267164
rect 293460 267152 293466 267164
rect 296686 267152 296714 267260
rect 302878 267248 302884 267260
rect 302936 267248 302942 267300
rect 306650 267248 306656 267300
rect 306708 267288 306714 267300
rect 312538 267288 312544 267300
rect 306708 267260 312544 267288
rect 306708 267248 306714 267260
rect 312538 267248 312544 267260
rect 312596 267248 312602 267300
rect 334618 267288 334624 267300
rect 316006 267260 334624 267288
rect 293460 267124 296714 267152
rect 293460 267112 293466 267124
rect 302234 267112 302240 267164
rect 302292 267152 302298 267164
rect 312814 267152 312820 267164
rect 302292 267124 312820 267152
rect 302292 267112 302298 267124
rect 312814 267112 312820 267124
rect 312872 267112 312878 267164
rect 313274 267112 313280 267164
rect 313332 267152 313338 267164
rect 316006 267152 316034 267260
rect 334618 267248 334624 267260
rect 334676 267248 334682 267300
rect 313332 267124 316034 267152
rect 313332 267112 313338 267124
rect 330478 267112 330484 267164
rect 330536 267152 330542 267164
rect 335326 267152 335354 267396
rect 345842 267384 345848 267396
rect 345900 267384 345906 267436
rect 347682 267384 347688 267436
rect 347740 267424 347746 267436
rect 353938 267424 353944 267436
rect 347740 267396 353944 267424
rect 347740 267384 347746 267396
rect 353938 267384 353944 267396
rect 353996 267384 354002 267436
rect 364978 267424 364984 267436
rect 354646 267396 364984 267424
rect 335722 267248 335728 267300
rect 335780 267288 335786 267300
rect 348418 267288 348424 267300
rect 335780 267260 348424 267288
rect 335780 267248 335786 267260
rect 348418 267248 348424 267260
rect 348476 267248 348482 267300
rect 350074 267248 350080 267300
rect 350132 267288 350138 267300
rect 354646 267288 354674 267396
rect 364978 267384 364984 267396
rect 365036 267384 365042 267436
rect 365162 267384 365168 267436
rect 365220 267424 365226 267436
rect 370498 267424 370504 267436
rect 365220 267396 370504 267424
rect 365220 267384 365226 267396
rect 370498 267384 370504 267396
rect 370556 267384 370562 267436
rect 370682 267384 370688 267436
rect 370740 267424 370746 267436
rect 374822 267424 374828 267436
rect 370740 267396 374828 267424
rect 370740 267384 370746 267396
rect 374822 267384 374828 267396
rect 374880 267384 374886 267436
rect 376754 267424 376760 267436
rect 375024 267396 376760 267424
rect 350132 267260 354674 267288
rect 350132 267248 350138 267260
rect 355226 267248 355232 267300
rect 355284 267288 355290 267300
rect 363230 267288 363236 267300
rect 355284 267260 363236 267288
rect 355284 267248 355290 267260
rect 363230 267248 363236 267260
rect 363288 267248 363294 267300
rect 375024 267288 375052 267396
rect 376754 267384 376760 267396
rect 376812 267384 376818 267436
rect 384298 267424 384304 267436
rect 377048 267396 384304 267424
rect 363432 267260 375052 267288
rect 330536 267124 335354 267152
rect 330536 267112 330542 267124
rect 341978 267112 341984 267164
rect 342036 267152 342042 267164
rect 350258 267152 350264 267164
rect 342036 267124 350264 267152
rect 342036 267112 342042 267124
rect 350258 267112 350264 267124
rect 350316 267112 350322 267164
rect 350810 267112 350816 267164
rect 350868 267152 350874 267164
rect 363432 267152 363460 267260
rect 375466 267248 375472 267300
rect 375524 267288 375530 267300
rect 377048 267288 377076 267396
rect 384298 267384 384304 267396
rect 384356 267384 384362 267436
rect 384482 267384 384488 267436
rect 384540 267424 384546 267436
rect 384540 267396 389174 267424
rect 384540 267384 384546 267396
rect 375524 267260 377076 267288
rect 375524 267248 375530 267260
rect 379514 267248 379520 267300
rect 379572 267288 379578 267300
rect 383654 267288 383660 267300
rect 379572 267260 383660 267288
rect 379572 267248 379578 267260
rect 383654 267248 383660 267260
rect 383712 267248 383718 267300
rect 383930 267248 383936 267300
rect 383988 267288 383994 267300
rect 388990 267288 388996 267300
rect 383988 267260 388996 267288
rect 383988 267248 383994 267260
rect 388990 267248 388996 267260
rect 389048 267248 389054 267300
rect 389146 267288 389174 267396
rect 392026 267384 392032 267436
rect 392084 267424 392090 267436
rect 393222 267424 393228 267436
rect 392084 267396 393228 267424
rect 392084 267384 392090 267396
rect 393222 267384 393228 267396
rect 393280 267384 393286 267436
rect 393406 267384 393412 267436
rect 393464 267424 393470 267436
rect 421098 267424 421104 267436
rect 393464 267396 421104 267424
rect 393464 267384 393470 267396
rect 421098 267384 421104 267396
rect 421156 267384 421162 267436
rect 421300 267424 421328 267532
rect 421466 267520 421472 267572
rect 421524 267560 421530 267572
rect 422110 267560 422116 267572
rect 421524 267532 422116 267560
rect 421524 267520 421530 267532
rect 422110 267520 422116 267532
rect 422168 267520 422174 267572
rect 422294 267520 422300 267572
rect 422352 267560 422358 267572
rect 423490 267560 423496 267572
rect 422352 267532 423496 267560
rect 422352 267520 422358 267532
rect 423490 267520 423496 267532
rect 423548 267520 423554 267572
rect 423674 267520 423680 267572
rect 423732 267560 423738 267572
rect 424962 267560 424968 267572
rect 423732 267532 424968 267560
rect 423732 267520 423738 267532
rect 424962 267520 424968 267532
rect 425020 267520 425026 267572
rect 425146 267520 425152 267572
rect 425204 267560 425210 267572
rect 426250 267560 426256 267572
rect 425204 267532 426256 267560
rect 425204 267520 425210 267532
rect 426250 267520 426256 267532
rect 426308 267520 426314 267572
rect 426434 267520 426440 267572
rect 426492 267560 426498 267572
rect 427768 267560 427774 267572
rect 426492 267532 427774 267560
rect 426492 267520 426498 267532
rect 427768 267520 427774 267532
rect 427826 267520 427832 267572
rect 427906 267520 427912 267572
rect 427964 267560 427970 267572
rect 427964 267532 466454 267560
rect 427964 267520 427970 267532
rect 442258 267424 442264 267436
rect 421300 267396 442264 267424
rect 442258 267384 442264 267396
rect 442316 267384 442322 267436
rect 442718 267384 442724 267436
rect 442776 267424 442782 267436
rect 446582 267424 446588 267436
rect 442776 267396 446588 267424
rect 442776 267384 442782 267396
rect 446582 267384 446588 267396
rect 446640 267384 446646 267436
rect 447226 267384 447232 267436
rect 447284 267424 447290 267436
rect 461578 267424 461584 267436
rect 447284 267396 461584 267424
rect 447284 267384 447290 267396
rect 461578 267384 461584 267396
rect 461636 267384 461642 267436
rect 461762 267384 461768 267436
rect 461820 267424 461826 267436
rect 466086 267424 466092 267436
rect 461820 267396 466092 267424
rect 461820 267384 461826 267396
rect 466086 267384 466092 267396
rect 466144 267384 466150 267436
rect 466426 267424 466454 267532
rect 467834 267520 467840 267572
rect 467892 267560 467898 267572
rect 475746 267560 475752 267572
rect 467892 267532 475752 267560
rect 467892 267520 467898 267532
rect 475746 267520 475752 267532
rect 475804 267520 475810 267572
rect 476114 267520 476120 267572
rect 476172 267560 476178 267572
rect 538858 267560 538864 267572
rect 476172 267532 538864 267560
rect 476172 267520 476178 267532
rect 538858 267520 538864 267532
rect 538916 267520 538922 267572
rect 466426 267396 477356 267424
rect 415486 267288 415492 267300
rect 389146 267260 415492 267288
rect 415486 267248 415492 267260
rect 415544 267248 415550 267300
rect 446766 267288 446772 267300
rect 415872 267260 446772 267288
rect 350868 267124 363460 267152
rect 350868 267112 350874 267124
rect 364978 267112 364984 267164
rect 365036 267152 365042 267164
rect 373902 267152 373908 267164
rect 365036 267124 373908 267152
rect 365036 267112 365042 267124
rect 373902 267112 373908 267124
rect 373960 267112 373966 267164
rect 374454 267112 374460 267164
rect 374512 267152 374518 267164
rect 402238 267152 402244 267164
rect 374512 267124 402244 267152
rect 374512 267112 374518 267124
rect 402238 267112 402244 267124
rect 402296 267112 402302 267164
rect 402974 267112 402980 267164
rect 403032 267152 403038 267164
rect 415872 267152 415900 267260
rect 446766 267248 446772 267260
rect 446824 267248 446830 267300
rect 447410 267248 447416 267300
rect 447468 267288 447474 267300
rect 477126 267288 477132 267300
rect 447468 267260 477132 267288
rect 447468 267248 447474 267260
rect 477126 267248 477132 267260
rect 477184 267248 477190 267300
rect 477328 267288 477356 267396
rect 480346 267384 480352 267436
rect 480404 267424 480410 267436
rect 481450 267424 481456 267436
rect 480404 267396 481456 267424
rect 480404 267384 480410 267396
rect 481450 267384 481456 267396
rect 481508 267384 481514 267436
rect 481634 267384 481640 267436
rect 481692 267424 481698 267436
rect 490558 267424 490564 267436
rect 481692 267396 490564 267424
rect 481692 267384 481698 267396
rect 490558 267384 490564 267396
rect 490616 267384 490622 267436
rect 490834 267384 490840 267436
rect 490892 267424 490898 267436
rect 572162 267424 572168 267436
rect 490892 267396 572168 267424
rect 490892 267384 490898 267396
rect 572162 267384 572168 267396
rect 572220 267384 572226 267436
rect 490558 267288 490564 267300
rect 477328 267260 490564 267288
rect 490558 267248 490564 267260
rect 490616 267248 490622 267300
rect 490834 267248 490840 267300
rect 490892 267288 490898 267300
rect 494882 267288 494888 267300
rect 490892 267260 494888 267288
rect 490892 267248 490898 267260
rect 494882 267248 494888 267260
rect 494940 267248 494946 267300
rect 495406 267260 496400 267288
rect 403032 267124 415900 267152
rect 403032 267112 403038 267124
rect 416314 267112 416320 267164
rect 416372 267152 416378 267164
rect 426434 267152 426440 267164
rect 416372 267124 426440 267152
rect 416372 267112 416378 267124
rect 426434 267112 426440 267124
rect 426492 267112 426498 267164
rect 426618 267112 426624 267164
rect 426676 267152 426682 267164
rect 426676 267124 430896 267152
rect 426676 267112 426682 267124
rect 430868 267084 430896 267124
rect 431218 267112 431224 267164
rect 431276 267152 431282 267164
rect 434714 267152 434720 267164
rect 431276 267124 434720 267152
rect 431276 267112 431282 267124
rect 434714 267112 434720 267124
rect 434772 267112 434778 267164
rect 436186 267112 436192 267164
rect 436244 267152 436250 267164
rect 437106 267152 437112 267164
rect 436244 267124 437112 267152
rect 436244 267112 436250 267124
rect 437106 267112 437112 267124
rect 437164 267112 437170 267164
rect 437290 267112 437296 267164
rect 437348 267152 437354 267164
rect 442074 267152 442080 267164
rect 437348 267124 442080 267152
rect 437348 267112 437354 267124
rect 442074 267112 442080 267124
rect 442132 267112 442138 267164
rect 442258 267112 442264 267164
rect 442316 267152 442322 267164
rect 442316 267124 446996 267152
rect 442316 267112 442322 267124
rect 430868 267056 431080 267084
rect 211706 267016 211712 267028
rect 200086 266988 211712 267016
rect 211706 266976 211712 266988
rect 211764 266976 211770 267028
rect 212442 266976 212448 267028
rect 212500 267016 212506 267028
rect 227162 267016 227168 267028
rect 212500 266988 227168 267016
rect 212500 266976 212506 266988
rect 227162 266976 227168 266988
rect 227220 266976 227226 267028
rect 227622 266976 227628 267028
rect 227680 267016 227686 267028
rect 235994 267016 236000 267028
rect 227680 266988 236000 267016
rect 227680 266976 227686 266988
rect 235994 266976 236000 266988
rect 236052 266976 236058 267028
rect 278682 266976 278688 267028
rect 278740 267016 278746 267028
rect 293218 267016 293224 267028
rect 278740 266988 293224 267016
rect 278740 266976 278746 266988
rect 293218 266976 293224 266988
rect 293276 266976 293282 267028
rect 300026 266976 300032 267028
rect 300084 267016 300090 267028
rect 311526 267016 311532 267028
rect 300084 266988 311532 267016
rect 300084 266976 300090 266988
rect 311526 266976 311532 266988
rect 311584 266976 311590 267028
rect 312538 266976 312544 267028
rect 312596 267016 312602 267028
rect 342530 267016 342536 267028
rect 312596 266988 342536 267016
rect 312596 266976 312602 266988
rect 342530 266976 342536 266988
rect 342588 266976 342594 267028
rect 344922 266976 344928 267028
rect 344980 267016 344986 267028
rect 351178 267016 351184 267028
rect 344980 266988 351184 267016
rect 344980 266976 344986 266988
rect 351178 266976 351184 266988
rect 351236 266976 351242 267028
rect 353018 266976 353024 267028
rect 353076 267016 353082 267028
rect 379698 267016 379704 267028
rect 353076 266988 379704 267016
rect 353076 266976 353082 266988
rect 379698 266976 379704 266988
rect 379756 266976 379762 267028
rect 379882 266976 379888 267028
rect 379940 267016 379946 267028
rect 384482 267016 384488 267028
rect 379940 266988 384488 267016
rect 379940 266976 379946 266988
rect 384482 266976 384488 266988
rect 384540 266976 384546 267028
rect 384666 266976 384672 267028
rect 384724 267016 384730 267028
rect 387794 267016 387800 267028
rect 384724 266988 387800 267016
rect 384724 266976 384730 266988
rect 387794 266976 387800 266988
rect 387852 266976 387858 267028
rect 388346 266976 388352 267028
rect 388404 267016 388410 267028
rect 393130 267016 393136 267028
rect 388404 266988 393136 267016
rect 388404 266976 388410 266988
rect 393130 266976 393136 266988
rect 393188 266976 393194 267028
rect 393314 266976 393320 267028
rect 393372 267016 393378 267028
rect 430666 267016 430672 267028
rect 393372 266988 430672 267016
rect 393372 266976 393378 266988
rect 430666 266976 430672 266988
rect 430724 266976 430730 267028
rect 431052 267016 431080 267056
rect 436738 267016 436744 267028
rect 431052 266988 436744 267016
rect 436738 266976 436744 266988
rect 436796 266976 436802 267028
rect 437106 266976 437112 267028
rect 437164 267016 437170 267028
rect 446766 267016 446772 267028
rect 437164 266988 446772 267016
rect 437164 266976 437170 266988
rect 446766 266976 446772 266988
rect 446824 266976 446830 267028
rect 446968 267016 446996 267124
rect 451918 267112 451924 267164
rect 451976 267152 451982 267164
rect 466408 267152 466414 267164
rect 451976 267124 466414 267152
rect 451976 267112 451982 267124
rect 466408 267112 466414 267124
rect 466466 267112 466472 267164
rect 466546 267112 466552 267164
rect 466604 267152 466610 267164
rect 475746 267152 475752 267164
rect 466604 267124 475752 267152
rect 466604 267112 466610 267124
rect 475746 267112 475752 267124
rect 475804 267112 475810 267164
rect 476086 267124 490052 267152
rect 461394 267016 461400 267028
rect 446968 266988 461400 267016
rect 461394 266976 461400 266988
rect 461452 266976 461458 267028
rect 461578 266976 461584 267028
rect 461636 267016 461642 267028
rect 476086 267016 476114 267124
rect 490024 267084 490052 267124
rect 490834 267112 490840 267164
rect 490892 267152 490898 267164
rect 495406 267152 495434 267260
rect 490892 267124 495434 267152
rect 496372 267152 496400 267260
rect 496538 267248 496544 267300
rect 496596 267288 496602 267300
rect 504910 267288 504916 267300
rect 496596 267260 504916 267288
rect 496596 267248 496602 267260
rect 504910 267248 504916 267260
rect 504968 267248 504974 267300
rect 505048 267248 505054 267300
rect 505106 267288 505112 267300
rect 550358 267288 550364 267300
rect 505106 267260 550364 267288
rect 505106 267248 505112 267260
rect 550358 267248 550364 267260
rect 550416 267248 550422 267300
rect 497458 267152 497464 267164
rect 496372 267124 497464 267152
rect 490892 267112 490898 267124
rect 497458 267112 497464 267124
rect 497516 267112 497522 267164
rect 498746 267112 498752 267164
rect 498804 267152 498810 267164
rect 638310 267152 638316 267164
rect 498804 267124 504772 267152
rect 498804 267112 498810 267124
rect 490558 267084 490564 267096
rect 490024 267056 490564 267084
rect 490558 267044 490564 267056
rect 490616 267044 490622 267096
rect 504744 267084 504772 267124
rect 504928 267124 638316 267152
rect 504928 267084 504956 267124
rect 638310 267112 638316 267124
rect 638368 267112 638374 267164
rect 504744 267056 504956 267084
rect 461636 266988 476114 267016
rect 461636 266976 461642 266988
rect 476390 266976 476396 267028
rect 476448 267016 476454 267028
rect 476942 267016 476948 267028
rect 476448 266988 476948 267016
rect 476448 266976 476454 266988
rect 476942 266976 476948 266988
rect 477000 266976 477006 267028
rect 477126 266976 477132 267028
rect 477184 267016 477190 267028
rect 487522 267016 487528 267028
rect 477184 266988 487528 267016
rect 477184 266976 477190 266988
rect 487522 266976 487528 266988
rect 487580 266976 487586 267028
rect 487706 266976 487712 267028
rect 487764 267016 487770 267028
rect 489822 267016 489828 267028
rect 487764 266988 489828 267016
rect 487764 266976 487770 266988
rect 489822 266976 489828 266988
rect 489880 266976 489886 267028
rect 504542 267016 504548 267028
rect 490944 266988 504548 267016
rect 490944 266948 490972 266988
rect 504542 266976 504548 266988
rect 504600 266976 504606 267028
rect 505186 266976 505192 267028
rect 505244 267016 505250 267028
rect 632698 267016 632704 267028
rect 505244 266988 632704 267016
rect 505244 266976 505250 266988
rect 632698 266976 632704 266988
rect 632756 266976 632762 267028
rect 490760 266920 490972 266948
rect 119338 266840 119344 266892
rect 119396 266880 119402 266892
rect 119396 266852 142154 266880
rect 119396 266840 119402 266852
rect 109678 266704 109684 266756
rect 109736 266744 109742 266756
rect 140314 266744 140320 266756
rect 109736 266716 140320 266744
rect 109736 266704 109742 266716
rect 140314 266704 140320 266716
rect 140372 266704 140378 266756
rect 142126 266744 142154 266852
rect 145558 266840 145564 266892
rect 145616 266880 145622 266892
rect 151354 266880 151360 266892
rect 145616 266852 151360 266880
rect 145616 266840 145622 266852
rect 151354 266840 151360 266852
rect 151412 266840 151418 266892
rect 157978 266840 157984 266892
rect 158036 266880 158042 266892
rect 174170 266880 174176 266892
rect 158036 266852 174176 266880
rect 158036 266840 158042 266852
rect 174170 266840 174176 266852
rect 174228 266840 174234 266892
rect 256510 266840 256516 266892
rect 256568 266880 256574 266892
rect 258074 266880 258080 266892
rect 256568 266852 258080 266880
rect 256568 266840 256574 266852
rect 258074 266840 258080 266852
rect 258132 266840 258138 266892
rect 311066 266840 311072 266892
rect 311124 266880 311130 266892
rect 319438 266880 319444 266892
rect 311124 266852 319444 266880
rect 311124 266840 311130 266852
rect 319438 266840 319444 266852
rect 319496 266840 319502 266892
rect 321278 266840 321284 266892
rect 321336 266880 321342 266892
rect 330478 266880 330484 266892
rect 321336 266852 330484 266880
rect 321336 266840 321342 266852
rect 330478 266840 330484 266852
rect 330536 266840 330542 266892
rect 330680 266852 333468 266880
rect 154298 266744 154304 266756
rect 142126 266716 154304 266744
rect 154298 266704 154304 266716
rect 154356 266704 154362 266756
rect 173894 266704 173900 266756
rect 173952 266744 173958 266756
rect 183002 266744 183008 266756
rect 173952 266716 183008 266744
rect 173952 266704 173958 266716
rect 183002 266704 183008 266716
rect 183060 266704 183066 266756
rect 206278 266704 206284 266756
rect 206336 266744 206342 266756
rect 210234 266744 210240 266756
rect 206336 266716 210240 266744
rect 206336 266704 206342 266716
rect 210234 266704 210240 266716
rect 210292 266704 210298 266756
rect 327258 266704 327264 266756
rect 327316 266744 327322 266756
rect 330680 266744 330708 266852
rect 327316 266716 330708 266744
rect 327316 266704 327322 266716
rect 330938 266704 330944 266756
rect 330996 266744 331002 266756
rect 333238 266744 333244 266756
rect 330996 266716 333244 266744
rect 330996 266704 331002 266716
rect 333238 266704 333244 266716
rect 333296 266704 333302 266756
rect 126698 266568 126704 266620
rect 126756 266608 126762 266620
rect 148410 266608 148416 266620
rect 126756 266580 148416 266608
rect 126756 266568 126762 266580
rect 148410 266568 148416 266580
rect 148468 266568 148474 266620
rect 151170 266568 151176 266620
rect 151228 266608 151234 266620
rect 163130 266608 163136 266620
rect 151228 266580 163136 266608
rect 151228 266568 151234 266580
rect 163130 266568 163136 266580
rect 163188 266568 163194 266620
rect 210602 266568 210608 266620
rect 210660 266608 210666 266620
rect 217594 266608 217600 266620
rect 210660 266580 217600 266608
rect 210660 266568 210666 266580
rect 217594 266568 217600 266580
rect 217652 266568 217658 266620
rect 246298 266568 246304 266620
rect 246356 266608 246362 266620
rect 248506 266608 248512 266620
rect 246356 266580 248512 266608
rect 246356 266568 246362 266580
rect 248506 266568 248512 266580
rect 248564 266568 248570 266620
rect 325786 266568 325792 266620
rect 325844 266608 325850 266620
rect 326706 266608 326712 266620
rect 325844 266580 326712 266608
rect 325844 266568 325850 266580
rect 326706 266568 326712 266580
rect 326764 266568 326770 266620
rect 331674 266568 331680 266620
rect 331732 266608 331738 266620
rect 332502 266608 332508 266620
rect 331732 266580 332508 266608
rect 331732 266568 331738 266580
rect 332502 266568 332508 266580
rect 332560 266568 332566 266620
rect 333440 266608 333468 266852
rect 333882 266840 333888 266892
rect 333940 266880 333946 266892
rect 347682 266880 347688 266892
rect 333940 266852 347688 266880
rect 333940 266840 333946 266852
rect 347682 266840 347688 266852
rect 347740 266840 347746 266892
rect 347866 266840 347872 266892
rect 347924 266880 347930 266892
rect 353570 266880 353576 266892
rect 347924 266852 353576 266880
rect 347924 266840 347930 266852
rect 353570 266840 353576 266852
rect 353628 266840 353634 266892
rect 359642 266840 359648 266892
rect 359700 266880 359706 266892
rect 390738 266880 390744 266892
rect 359700 266852 390744 266880
rect 359700 266840 359706 266852
rect 390738 266840 390744 266852
rect 390796 266840 390802 266892
rect 391290 266840 391296 266892
rect 391348 266880 391354 266892
rect 392210 266880 392216 266892
rect 391348 266852 392216 266880
rect 391348 266840 391354 266852
rect 392210 266840 392216 266852
rect 392268 266840 392274 266892
rect 392762 266840 392768 266892
rect 392820 266880 392826 266892
rect 466270 266880 466276 266892
rect 392820 266852 437244 266880
rect 392820 266840 392826 266852
rect 437216 266812 437244 266852
rect 437400 266852 466276 266880
rect 437400 266812 437428 266852
rect 466270 266840 466276 266852
rect 466328 266840 466334 266892
rect 490760 266880 490788 266920
rect 466426 266852 490788 266880
rect 437216 266784 437428 266812
rect 338298 266704 338304 266756
rect 338356 266744 338362 266756
rect 358170 266744 358176 266756
rect 338356 266716 358176 266744
rect 338356 266704 338362 266716
rect 358170 266704 358176 266716
rect 358228 266704 358234 266756
rect 365162 266744 365168 266756
rect 358740 266716 365168 266744
rect 345658 266608 345664 266620
rect 333440 266580 345664 266608
rect 345658 266568 345664 266580
rect 345716 266568 345722 266620
rect 353570 266568 353576 266620
rect 353628 266608 353634 266620
rect 354674 266608 354680 266620
rect 353628 266580 354680 266608
rect 353628 266568 353634 266580
rect 354674 266568 354680 266580
rect 354732 266568 354738 266620
rect 357434 266568 357440 266620
rect 357492 266608 357498 266620
rect 358740 266608 358768 266716
rect 365162 266704 365168 266716
rect 365220 266704 365226 266756
rect 367002 266704 367008 266756
rect 367060 266744 367066 266756
rect 396718 266744 396724 266756
rect 367060 266716 396724 266744
rect 367060 266704 367066 266716
rect 396718 266704 396724 266716
rect 396776 266704 396782 266756
rect 397178 266704 397184 266756
rect 397236 266744 397242 266756
rect 402790 266744 402796 266756
rect 397236 266716 402796 266744
rect 397236 266704 397242 266716
rect 402790 266704 402796 266716
rect 402848 266704 402854 266756
rect 403066 266704 403072 266756
rect 403124 266744 403130 266756
rect 404170 266744 404176 266756
rect 403124 266716 404176 266744
rect 403124 266704 403130 266716
rect 404170 266704 404176 266716
rect 404228 266704 404234 266756
rect 406010 266704 406016 266756
rect 406068 266744 406074 266756
rect 410242 266744 410248 266756
rect 406068 266716 410248 266744
rect 406068 266704 406074 266716
rect 410242 266704 410248 266716
rect 410300 266704 410306 266756
rect 410426 266704 410432 266756
rect 410484 266744 410490 266756
rect 412082 266744 412088 266756
rect 410484 266716 412088 266744
rect 410484 266704 410490 266716
rect 412082 266704 412088 266716
rect 412140 266704 412146 266756
rect 412450 266704 412456 266756
rect 412508 266744 412514 266756
rect 415302 266744 415308 266756
rect 412508 266716 415308 266744
rect 412508 266704 412514 266716
rect 415302 266704 415308 266716
rect 415360 266704 415366 266756
rect 415578 266704 415584 266756
rect 415636 266744 415642 266756
rect 416682 266744 416688 266756
rect 415636 266716 416688 266744
rect 415636 266704 415642 266716
rect 416682 266704 416688 266716
rect 416740 266704 416746 266756
rect 418246 266704 418252 266756
rect 418304 266744 418310 266756
rect 426618 266744 426624 266756
rect 418304 266716 426624 266744
rect 418304 266704 418310 266716
rect 426618 266704 426624 266716
rect 426676 266704 426682 266756
rect 436554 266744 436560 266756
rect 427786 266716 436560 266744
rect 357492 266580 358768 266608
rect 357492 266568 357498 266580
rect 358906 266568 358912 266620
rect 358964 266608 358970 266620
rect 360102 266608 360108 266620
rect 358964 266580 360108 266608
rect 358964 266568 358970 266580
rect 360102 266568 360108 266580
rect 360160 266568 360166 266620
rect 360378 266568 360384 266620
rect 360436 266608 360442 266620
rect 361206 266608 361212 266620
rect 360436 266580 361212 266608
rect 360436 266568 360442 266580
rect 361206 266568 361212 266580
rect 361264 266568 361270 266620
rect 363230 266568 363236 266620
rect 363288 266608 363294 266620
rect 382182 266608 382188 266620
rect 363288 266580 382188 266608
rect 363288 266568 363294 266580
rect 382182 266568 382188 266580
rect 382240 266568 382246 266620
rect 384942 266608 384948 266620
rect 382384 266580 384948 266608
rect 241330 266500 241336 266552
rect 241388 266540 241394 266552
rect 245562 266540 245568 266552
rect 241388 266512 245568 266540
rect 241388 266500 241394 266512
rect 245562 266500 245568 266512
rect 245620 266500 245626 266552
rect 259914 266500 259920 266552
rect 259972 266540 259978 266552
rect 262582 266540 262588 266552
rect 259972 266512 262588 266540
rect 259972 266500 259978 266512
rect 262582 266500 262588 266512
rect 262640 266500 262646 266552
rect 269850 266500 269856 266552
rect 269908 266540 269914 266552
rect 274634 266540 274640 266552
rect 269908 266512 274640 266540
rect 269908 266500 269914 266512
rect 274634 266500 274640 266512
rect 274692 266500 274698 266552
rect 280154 266500 280160 266552
rect 280212 266540 280218 266552
rect 285766 266540 285772 266552
rect 280212 266512 285772 266540
rect 280212 266500 280218 266512
rect 285766 266500 285772 266512
rect 285824 266500 285830 266552
rect 291194 266500 291200 266552
rect 291252 266540 291258 266552
rect 294598 266540 294604 266552
rect 291252 266512 294604 266540
rect 291252 266500 291258 266512
rect 294598 266500 294604 266512
rect 294656 266500 294662 266552
rect 301498 266500 301504 266552
rect 301556 266540 301562 266552
rect 304166 266540 304172 266552
rect 301556 266512 304172 266540
rect 301556 266500 301562 266512
rect 304166 266500 304172 266512
rect 304224 266500 304230 266552
rect 304442 266500 304448 266552
rect 304500 266540 304506 266552
rect 305546 266540 305552 266552
rect 304500 266512 305552 266540
rect 304500 266500 304506 266512
rect 305546 266500 305552 266512
rect 305604 266500 305610 266552
rect 319898 266500 319904 266552
rect 319956 266540 319962 266552
rect 322198 266540 322204 266552
rect 319956 266512 322204 266540
rect 319956 266500 319962 266512
rect 322198 266500 322204 266512
rect 322256 266500 322262 266552
rect 348602 266500 348608 266552
rect 348660 266540 348666 266552
rect 348660 266512 353432 266540
rect 348660 266500 348666 266512
rect 132586 266432 132592 266484
rect 132644 266472 132650 266484
rect 145466 266472 145472 266484
rect 132644 266444 145472 266472
rect 132644 266432 132650 266444
rect 145466 266432 145472 266444
rect 145524 266432 145530 266484
rect 208486 266432 208492 266484
rect 208544 266472 208550 266484
rect 212442 266472 212448 266484
rect 208544 266444 212448 266472
rect 208544 266432 208550 266444
rect 212442 266432 212448 266444
rect 212500 266432 212506 266484
rect 322474 266432 322480 266484
rect 322532 266472 322538 266484
rect 338942 266472 338948 266484
rect 322532 266444 338948 266472
rect 322532 266432 322538 266444
rect 338942 266432 338948 266444
rect 339000 266432 339006 266484
rect 353404 266472 353432 266512
rect 364794 266472 364800 266484
rect 353404 266444 364800 266472
rect 364794 266432 364800 266444
rect 364852 266432 364858 266484
rect 370498 266432 370504 266484
rect 370556 266472 370562 266484
rect 378778 266472 378784 266484
rect 370556 266444 378784 266472
rect 370556 266432 370562 266444
rect 378778 266432 378784 266444
rect 378836 266432 378842 266484
rect 381722 266432 381728 266484
rect 381780 266472 381786 266484
rect 382384 266472 382412 266580
rect 384942 266568 384948 266580
rect 385000 266568 385006 266620
rect 385402 266568 385408 266620
rect 385460 266608 385466 266620
rect 389818 266608 389824 266620
rect 385460 266580 389824 266608
rect 385460 266568 385466 266580
rect 389818 266568 389824 266580
rect 389876 266568 389882 266620
rect 390554 266568 390560 266620
rect 390612 266608 390618 266620
rect 391842 266608 391848 266620
rect 390612 266580 391848 266608
rect 390612 266568 390618 266580
rect 391842 266568 391848 266580
rect 391900 266568 391906 266620
rect 392210 266568 392216 266620
rect 392268 266608 392274 266620
rect 427786 266608 427814 266716
rect 436554 266704 436560 266716
rect 436612 266704 436618 266756
rect 437934 266704 437940 266756
rect 437992 266744 437998 266756
rect 451918 266744 451924 266756
rect 437992 266716 451924 266744
rect 437992 266704 437998 266716
rect 451918 266704 451924 266716
rect 451976 266704 451982 266756
rect 452102 266704 452108 266756
rect 452160 266744 452166 266756
rect 454586 266744 454592 266756
rect 452160 266716 454592 266744
rect 452160 266704 452166 266716
rect 454586 266704 454592 266716
rect 454644 266704 454650 266756
rect 454770 266704 454776 266756
rect 454828 266744 454834 266756
rect 466426 266744 466454 266852
rect 491202 266840 491208 266892
rect 491260 266880 491266 266892
rect 629294 266880 629300 266892
rect 491260 266852 629300 266880
rect 491260 266840 491266 266852
rect 629294 266840 629300 266852
rect 629352 266840 629358 266892
rect 666186 266772 666192 266824
rect 666244 266812 666250 266824
rect 675478 266812 675484 266824
rect 666244 266784 675484 266812
rect 666244 266772 666250 266784
rect 675478 266772 675484 266784
rect 675536 266772 675542 266824
rect 454828 266716 466454 266744
rect 454828 266704 454834 266716
rect 466730 266704 466736 266756
rect 466788 266744 466794 266756
rect 469858 266744 469864 266756
rect 466788 266716 469864 266744
rect 466788 266704 466794 266716
rect 469858 266704 469864 266716
rect 469916 266704 469922 266756
rect 470042 266704 470048 266756
rect 470100 266744 470106 266756
rect 504726 266744 504732 266756
rect 470100 266716 504732 266744
rect 470100 266704 470106 266716
rect 504726 266704 504732 266716
rect 504784 266704 504790 266756
rect 504910 266704 504916 266756
rect 504968 266744 504974 266756
rect 543734 266744 543740 266756
rect 504968 266716 543740 266744
rect 504968 266704 504974 266716
rect 543734 266704 543740 266716
rect 543792 266704 543798 266756
rect 550358 266704 550364 266756
rect 550416 266744 550422 266756
rect 594978 266744 594984 266756
rect 550416 266716 594984 266744
rect 550416 266704 550422 266716
rect 594978 266704 594984 266716
rect 595036 266704 595042 266756
rect 392268 266580 427814 266608
rect 392268 266568 392274 266580
rect 427906 266568 427912 266620
rect 427964 266608 427970 266620
rect 437106 266608 437112 266620
rect 427964 266580 437112 266608
rect 427964 266568 427970 266580
rect 437106 266568 437112 266580
rect 437164 266568 437170 266620
rect 466546 266608 466552 266620
rect 437400 266580 466552 266608
rect 381780 266444 382412 266472
rect 381780 266432 381786 266444
rect 384298 266432 384304 266484
rect 384356 266472 384362 266484
rect 401134 266472 401140 266484
rect 384356 266444 401140 266472
rect 384356 266432 384362 266444
rect 401134 266432 401140 266444
rect 401192 266432 401198 266484
rect 401594 266432 401600 266484
rect 401652 266472 401658 266484
rect 402606 266472 402612 266484
rect 401652 266444 402612 266472
rect 401652 266432 401658 266444
rect 402606 266432 402612 266444
rect 402664 266432 402670 266484
rect 402790 266432 402796 266484
rect 402848 266472 402854 266484
rect 437400 266472 437428 266580
rect 466546 266568 466552 266580
rect 466604 266568 466610 266620
rect 466914 266568 466920 266620
rect 466972 266608 466978 266620
rect 476022 266608 476028 266620
rect 466972 266580 476028 266608
rect 466972 266568 466978 266580
rect 476022 266568 476028 266580
rect 476080 266568 476086 266620
rect 476206 266568 476212 266620
rect 476264 266608 476270 266620
rect 481634 266608 481640 266620
rect 476264 266580 481640 266608
rect 476264 266568 476270 266580
rect 481634 266568 481640 266580
rect 481692 266568 481698 266620
rect 482554 266568 482560 266620
rect 482612 266608 482618 266620
rect 485590 266608 485596 266620
rect 482612 266580 485596 266608
rect 482612 266568 482618 266580
rect 485590 266568 485596 266580
rect 485648 266568 485654 266620
rect 485774 266568 485780 266620
rect 485832 266608 485838 266620
rect 554038 266608 554044 266620
rect 485832 266580 554044 266608
rect 485832 266568 485838 266580
rect 554038 266568 554044 266580
rect 554096 266568 554102 266620
rect 675478 266608 675484 266620
rect 669286 266580 675484 266608
rect 666370 266500 666376 266552
rect 666428 266540 666434 266552
rect 669286 266540 669314 266580
rect 675478 266568 675484 266580
rect 675536 266568 675542 266620
rect 666428 266512 669314 266540
rect 666428 266500 666434 266512
rect 402848 266444 437428 266472
rect 402848 266432 402854 266444
rect 437750 266432 437756 266484
rect 437808 266472 437814 266484
rect 437808 266444 441936 266472
rect 437808 266432 437814 266444
rect 153838 266364 153844 266416
rect 153896 266404 153902 266416
rect 156138 266404 156144 266416
rect 153896 266376 156144 266404
rect 153896 266364 153902 266376
rect 156138 266364 156144 266376
rect 156196 266364 156202 266416
rect 164878 266364 164884 266416
rect 164936 266404 164942 266416
rect 167546 266404 167552 266416
rect 164936 266376 167552 266404
rect 164936 266364 164942 266376
rect 167546 266364 167552 266376
rect 167604 266364 167610 266416
rect 174722 266364 174728 266416
rect 174780 266404 174786 266416
rect 180058 266404 180064 266416
rect 174780 266376 180064 266404
rect 174780 266364 174786 266376
rect 180058 266364 180064 266376
rect 180116 266364 180122 266416
rect 204898 266364 204904 266416
rect 204956 266404 204962 266416
rect 206554 266404 206560 266416
rect 204956 266376 206560 266404
rect 204956 266364 204962 266376
rect 206554 266364 206560 266376
rect 206612 266364 206618 266416
rect 219434 266364 219440 266416
rect 219492 266404 219498 266416
rect 227898 266404 227904 266416
rect 219492 266376 227904 266404
rect 219492 266364 219498 266376
rect 227898 266364 227904 266376
rect 227956 266364 227962 266416
rect 230750 266364 230756 266416
rect 230808 266404 230814 266416
rect 233050 266404 233056 266416
rect 230808 266376 233056 266404
rect 230808 266364 230814 266376
rect 233050 266364 233056 266376
rect 233108 266364 233114 266416
rect 239490 266364 239496 266416
rect 239548 266404 239554 266416
rect 241882 266404 241888 266416
rect 239548 266376 241888 266404
rect 239548 266364 239554 266376
rect 241882 266364 241888 266376
rect 241940 266364 241946 266416
rect 251174 266364 251180 266416
rect 251232 266404 251238 266416
rect 252186 266404 252192 266416
rect 251232 266376 252192 266404
rect 251232 266364 251238 266376
rect 252186 266364 252192 266376
rect 252244 266364 252250 266416
rect 255866 266364 255872 266416
rect 255924 266404 255930 266416
rect 256694 266404 256700 266416
rect 255924 266376 256700 266404
rect 255924 266364 255930 266376
rect 256694 266364 256700 266376
rect 256752 266364 256758 266416
rect 258074 266364 258080 266416
rect 258132 266404 258138 266416
rect 259638 266404 259644 266416
rect 258132 266376 259644 266404
rect 258132 266364 258138 266376
rect 259638 266364 259644 266376
rect 259696 266364 259702 266416
rect 260282 266364 260288 266416
rect 260340 266404 260346 266416
rect 261754 266404 261760 266416
rect 260340 266376 261760 266404
rect 260340 266364 260346 266376
rect 261754 266364 261760 266376
rect 261812 266364 261818 266416
rect 262122 266364 262128 266416
rect 262180 266404 262186 266416
rect 266354 266404 266360 266416
rect 262180 266376 266360 266404
rect 262180 266364 262186 266376
rect 266354 266364 266360 266376
rect 266412 266364 266418 266416
rect 270586 266364 270592 266416
rect 270644 266404 270650 266416
rect 271598 266404 271604 266416
rect 270644 266376 271604 266404
rect 270644 266364 270650 266376
rect 271598 266364 271604 266376
rect 271656 266364 271662 266416
rect 280890 266364 280896 266416
rect 280948 266404 280954 266416
rect 282178 266404 282184 266416
rect 280948 266376 282184 266404
rect 280948 266364 280954 266376
rect 282178 266364 282184 266376
rect 282236 266364 282242 266416
rect 288986 266364 288992 266416
rect 289044 266404 289050 266416
rect 291838 266404 291844 266416
rect 289044 266376 291844 266404
rect 289044 266364 289050 266376
rect 291838 266364 291844 266376
rect 291896 266364 291902 266416
rect 294138 266364 294144 266416
rect 294196 266404 294202 266416
rect 295150 266404 295156 266416
rect 294196 266376 295156 266404
rect 294196 266364 294202 266376
rect 295150 266364 295156 266376
rect 295208 266364 295214 266416
rect 297818 266364 297824 266416
rect 297876 266404 297882 266416
rect 301222 266404 301228 266416
rect 297876 266376 301228 266404
rect 297876 266364 297882 266376
rect 301222 266364 301228 266376
rect 301280 266364 301286 266416
rect 303706 266364 303712 266416
rect 303764 266404 303770 266416
rect 304902 266404 304908 266416
rect 303764 266376 304908 266404
rect 303764 266364 303770 266376
rect 304902 266364 304908 266376
rect 304960 266364 304966 266416
rect 305178 266364 305184 266416
rect 305236 266404 305242 266416
rect 306190 266404 306196 266416
rect 305236 266376 306196 266404
rect 305236 266364 305242 266376
rect 306190 266364 306196 266376
rect 306248 266364 306254 266416
rect 316218 266364 316224 266416
rect 316276 266404 316282 266416
rect 317138 266404 317144 266416
rect 316276 266376 317144 266404
rect 316276 266364 316282 266376
rect 317138 266364 317144 266376
rect 317196 266364 317202 266416
rect 320634 266364 320640 266416
rect 320692 266404 320698 266416
rect 321462 266404 321468 266416
rect 320692 266376 321468 266404
rect 320692 266364 320698 266376
rect 321462 266364 321468 266376
rect 321520 266364 321526 266416
rect 342714 266364 342720 266416
rect 342772 266404 342778 266416
rect 343542 266404 343548 266416
rect 342772 266376 343548 266404
rect 342772 266364 342778 266376
rect 343542 266364 343548 266376
rect 343600 266364 343606 266416
rect 346394 266364 346400 266416
rect 346452 266404 346458 266416
rect 350074 266404 350080 266416
rect 346452 266376 350080 266404
rect 346452 266364 346458 266376
rect 350074 266364 350080 266376
rect 350132 266364 350138 266416
rect 352282 266364 352288 266416
rect 352340 266404 352346 266416
rect 353202 266404 353208 266416
rect 352340 266376 353208 266404
rect 352340 266364 352346 266376
rect 353202 266364 353208 266376
rect 353260 266364 353266 266416
rect 372154 266296 372160 266348
rect 372212 266336 372218 266348
rect 432598 266336 432604 266348
rect 372212 266308 432604 266336
rect 372212 266296 372218 266308
rect 432598 266296 432604 266308
rect 432656 266296 432662 266348
rect 441706 266336 441712 266348
rect 437446 266308 441712 266336
rect 373626 266160 373632 266212
rect 373684 266200 373690 266212
rect 437446 266200 437474 266308
rect 441706 266296 441712 266308
rect 441764 266296 441770 266348
rect 441908 266336 441936 266444
rect 442074 266432 442080 266484
rect 442132 266472 442138 266484
rect 532970 266472 532976 266484
rect 442132 266444 532976 266472
rect 442132 266432 442138 266444
rect 532970 266432 532976 266444
rect 533028 266432 533034 266484
rect 664806 266364 664812 266416
rect 664864 266404 664870 266416
rect 675294 266404 675300 266416
rect 664864 266376 675300 266404
rect 664864 266364 664870 266376
rect 675294 266364 675300 266376
rect 675352 266364 675358 266416
rect 442718 266336 442724 266348
rect 441908 266308 442724 266336
rect 442718 266296 442724 266308
rect 442776 266296 442782 266348
rect 442902 266296 442908 266348
rect 442960 266336 442966 266348
rect 445938 266336 445944 266348
rect 442960 266308 445944 266336
rect 442960 266296 442966 266308
rect 445938 266296 445944 266308
rect 445996 266296 446002 266348
rect 450538 266296 450544 266348
rect 450596 266336 450602 266348
rect 452102 266336 452108 266348
rect 450596 266308 452108 266336
rect 450596 266296 450602 266308
rect 452102 266296 452108 266308
rect 452160 266296 452166 266348
rect 566274 266336 566280 266348
rect 452304 266308 566280 266336
rect 443178 266200 443184 266212
rect 373684 266172 437474 266200
rect 440344 266172 443184 266200
rect 373684 266160 373690 266172
rect 404170 266024 404176 266076
rect 404228 266064 404234 266076
rect 412450 266064 412456 266076
rect 404228 266036 412456 266064
rect 404228 266024 404234 266036
rect 412450 266024 412456 266036
rect 412508 266024 412514 266076
rect 432598 266024 432604 266076
rect 432656 266064 432662 266076
rect 440344 266064 440372 266172
rect 443178 266160 443184 266172
rect 443236 266160 443242 266212
rect 443914 266160 443920 266212
rect 443972 266200 443978 266212
rect 448514 266200 448520 266212
rect 443972 266172 448520 266200
rect 443972 266160 443978 266172
rect 448514 266160 448520 266172
rect 448572 266160 448578 266212
rect 448698 266160 448704 266212
rect 448756 266200 448762 266212
rect 452304 266200 452332 266308
rect 566274 266296 566280 266308
rect 566332 266296 566338 266348
rect 448756 266172 452332 266200
rect 448756 266160 448762 266172
rect 454586 266160 454592 266212
rect 454644 266200 454650 266212
rect 575750 266200 575756 266212
rect 454644 266172 575756 266200
rect 454644 266160 454650 266172
rect 575750 266160 575756 266172
rect 575808 266160 575814 266212
rect 432656 266036 440372 266064
rect 432656 266024 432662 266036
rect 442258 266024 442264 266076
rect 442316 266064 442322 266076
rect 461578 266064 461584 266076
rect 442316 266036 461584 266064
rect 442316 266024 442322 266036
rect 461578 266024 461584 266036
rect 461636 266024 461642 266076
rect 462130 266024 462136 266076
rect 462188 266064 462194 266076
rect 463970 266064 463976 266076
rect 462188 266036 463976 266064
rect 462188 266024 462194 266036
rect 463970 266024 463976 266036
rect 464028 266024 464034 266076
rect 464154 266024 464160 266076
rect 464212 266064 464218 266076
rect 591022 266064 591028 266076
rect 464212 266036 591028 266064
rect 464212 266024 464218 266036
rect 591022 266024 591028 266036
rect 591080 266024 591086 266076
rect 198734 265888 198740 265940
rect 198792 265928 198798 265940
rect 199654 265928 199660 265940
rect 198792 265900 199660 265928
rect 198792 265888 198798 265900
rect 199654 265888 199660 265900
rect 199712 265888 199718 265940
rect 218054 265888 218060 265940
rect 218112 265928 218118 265940
rect 218790 265928 218796 265940
rect 218112 265900 218796 265928
rect 218112 265888 218118 265900
rect 218790 265888 218796 265900
rect 218848 265888 218854 265940
rect 389082 265888 389088 265940
rect 389140 265928 389146 265940
rect 470594 265928 470600 265940
rect 389140 265900 470600 265928
rect 389140 265888 389146 265900
rect 470594 265888 470600 265900
rect 470652 265888 470658 265940
rect 470778 265888 470784 265940
rect 470836 265928 470842 265940
rect 601694 265928 601700 265940
rect 470836 265900 601700 265928
rect 470836 265888 470842 265900
rect 601694 265888 601700 265900
rect 601752 265888 601758 265940
rect 362586 265752 362592 265804
rect 362644 265792 362650 265804
rect 428274 265792 428280 265804
rect 362644 265764 428280 265792
rect 362644 265752 362650 265764
rect 428274 265752 428280 265764
rect 428332 265752 428338 265804
rect 437658 265752 437664 265804
rect 437716 265792 437722 265804
rect 523678 265792 523684 265804
rect 437716 265764 523684 265792
rect 437716 265752 437722 265764
rect 523678 265752 523684 265764
rect 523736 265752 523742 265804
rect 384666 265616 384672 265668
rect 384724 265656 384730 265668
rect 461394 265656 461400 265668
rect 384724 265628 461400 265656
rect 384724 265616 384730 265628
rect 461394 265616 461400 265628
rect 461452 265616 461458 265668
rect 461578 265616 461584 265668
rect 461636 265656 461642 265668
rect 495894 265656 495900 265668
rect 461636 265628 495900 265656
rect 461636 265616 461642 265628
rect 495894 265616 495900 265628
rect 495952 265616 495958 265668
rect 499482 265616 499488 265668
rect 499540 265656 499546 265668
rect 648614 265656 648620 265668
rect 499540 265628 648620 265656
rect 499540 265616 499546 265628
rect 648614 265616 648620 265628
rect 648672 265616 648678 265668
rect 669314 265548 669320 265600
rect 669372 265588 669378 265600
rect 675478 265588 675484 265600
rect 669372 265560 675484 265588
rect 669372 265548 669378 265560
rect 675478 265548 675484 265560
rect 675536 265548 675542 265600
rect 404538 265480 404544 265532
rect 404596 265520 404602 265532
rect 442258 265520 442264 265532
rect 404596 265492 442264 265520
rect 404596 265480 404602 265492
rect 442258 265480 442264 265492
rect 442316 265480 442322 265532
rect 444282 265480 444288 265532
rect 444340 265520 444346 265532
rect 559282 265520 559288 265532
rect 444340 265492 559288 265520
rect 444340 265480 444346 265492
rect 559282 265480 559288 265492
rect 559340 265480 559346 265532
rect 665266 265412 665272 265464
rect 665324 265452 665330 265464
rect 675478 265452 675484 265464
rect 665324 265424 675484 265452
rect 665324 265412 665330 265424
rect 675478 265412 675484 265424
rect 675536 265412 675542 265464
rect 442074 265344 442080 265396
rect 442132 265384 442138 265396
rect 552658 265384 552664 265396
rect 442132 265356 552664 265384
rect 442132 265344 442138 265356
rect 552658 265344 552664 265356
rect 552716 265344 552722 265396
rect 417786 265208 417792 265260
rect 417844 265248 417850 265260
rect 516410 265248 516416 265260
rect 417844 265220 516416 265248
rect 417844 265208 417850 265220
rect 516410 265208 516416 265220
rect 516468 265208 516474 265260
rect 665082 265208 665088 265260
rect 665140 265248 665146 265260
rect 675294 265248 675300 265260
rect 665140 265220 675300 265248
rect 665140 265208 665146 265220
rect 675294 265208 675300 265220
rect 675352 265208 675358 265260
rect 439866 265072 439872 265124
rect 439924 265112 439930 265124
rect 537754 265112 537760 265124
rect 439924 265084 537760 265112
rect 439924 265072 439930 265084
rect 537754 265072 537760 265084
rect 537812 265072 537818 265124
rect 664254 265072 664260 265124
rect 664312 265112 664318 265124
rect 664312 265084 669452 265112
rect 664312 265072 664318 265084
rect 669424 265044 669452 265084
rect 675478 265044 675484 265056
rect 669424 265016 675484 265044
rect 675478 265004 675484 265016
rect 675536 265004 675542 265056
rect 386138 264936 386144 264988
rect 386196 264976 386202 264988
rect 467282 264976 467288 264988
rect 386196 264948 467288 264976
rect 386196 264936 386202 264948
rect 467282 264936 467288 264948
rect 467340 264936 467346 264988
rect 477402 264936 477408 264988
rect 477460 264976 477466 264988
rect 612734 264976 612740 264988
rect 477460 264948 612740 264976
rect 477460 264936 477466 264948
rect 612734 264936 612740 264948
rect 612792 264936 612798 264988
rect 664254 264936 664260 264988
rect 664312 264976 664318 264988
rect 664312 264948 669314 264976
rect 664312 264936 664318 264948
rect 669286 264920 669314 264948
rect 669286 264880 669320 264920
rect 669314 264868 669320 264880
rect 669372 264868 669378 264920
rect 435450 264732 435456 264784
rect 435508 264772 435514 264784
rect 545114 264772 545120 264784
rect 435508 264744 545120 264772
rect 435508 264732 435514 264744
rect 545114 264732 545120 264744
rect 545172 264732 545178 264784
rect 453114 264596 453120 264648
rect 453172 264636 453178 264648
rect 574094 264636 574100 264648
rect 453172 264608 574100 264636
rect 453172 264596 453178 264608
rect 574094 264596 574100 264608
rect 574152 264596 574158 264648
rect 471882 264460 471888 264512
rect 471940 264500 471946 264512
rect 603074 264500 603080 264512
rect 471940 264472 603080 264500
rect 471940 264460 471946 264472
rect 603074 264460 603080 264472
rect 603132 264460 603138 264512
rect 491018 264324 491024 264376
rect 491076 264364 491082 264376
rect 491570 264364 491576 264376
rect 491076 264336 491576 264364
rect 491076 264324 491082 264336
rect 491570 264324 491576 264336
rect 491628 264324 491634 264376
rect 497642 264324 497648 264376
rect 497700 264364 497706 264376
rect 643738 264364 643744 264376
rect 497700 264336 643744 264364
rect 497700 264324 497706 264336
rect 643738 264324 643744 264336
rect 643796 264324 643802 264376
rect 51902 264188 51908 264240
rect 51960 264228 51966 264240
rect 655514 264228 655520 264240
rect 51960 264200 655520 264228
rect 51960 264188 51966 264200
rect 655514 264188 655520 264200
rect 655572 264188 655578 264240
rect 507118 264052 507124 264104
rect 507176 264092 507182 264104
rect 600590 264092 600596 264104
rect 507176 264064 600596 264092
rect 507176 264052 507182 264064
rect 600590 264052 600596 264064
rect 600648 264052 600654 264104
rect 666186 263576 666192 263628
rect 666244 263616 666250 263628
rect 675478 263616 675484 263628
rect 666244 263588 675484 263616
rect 666244 263576 666250 263588
rect 675478 263576 675484 263588
rect 675536 263576 675542 263628
rect 666370 262488 666376 262540
rect 666428 262528 666434 262540
rect 675478 262528 675484 262540
rect 666428 262500 675484 262528
rect 666428 262488 666434 262500
rect 675478 262488 675484 262500
rect 675536 262488 675542 262540
rect 669406 262080 669412 262132
rect 669464 262120 669470 262132
rect 675478 262120 675484 262132
rect 669464 262092 675484 262120
rect 669464 262080 669470 262092
rect 675478 262080 675484 262092
rect 675536 262080 675542 262132
rect 511534 261468 511540 261520
rect 511592 261508 511598 261520
rect 568574 261508 568580 261520
rect 511592 261480 568580 261508
rect 511592 261468 511598 261480
rect 568574 261468 568580 261480
rect 568632 261468 568638 261520
rect 675846 260992 675852 261044
rect 675904 261032 675910 261044
rect 676398 261032 676404 261044
rect 675904 261004 676404 261032
rect 675904 260992 675910 261004
rect 676398 260992 676404 261004
rect 676456 260992 676462 261044
rect 673362 260448 673368 260500
rect 673420 260488 673426 260500
rect 675478 260488 675484 260500
rect 673420 260460 675484 260488
rect 673420 260448 673426 260460
rect 675478 260448 675484 260460
rect 675536 260448 675542 260500
rect 669130 259836 669136 259888
rect 669188 259876 669194 259888
rect 675478 259876 675484 259888
rect 669188 259848 675484 259876
rect 669188 259836 669194 259848
rect 675478 259836 675484 259848
rect 675536 259836 675542 259888
rect 671890 259632 671896 259684
rect 671948 259672 671954 259684
rect 675478 259672 675484 259684
rect 671948 259644 675484 259672
rect 671948 259632 671954 259644
rect 675478 259632 675484 259644
rect 675536 259632 675542 259684
rect 510982 259428 510988 259480
rect 511040 259468 511046 259480
rect 514018 259468 514024 259480
rect 511040 259440 514024 259468
rect 511040 259428 511046 259440
rect 514018 259428 514024 259440
rect 514076 259428 514082 259480
rect 673086 258816 673092 258868
rect 673144 258856 673150 258868
rect 675478 258856 675484 258868
rect 673144 258828 675484 258856
rect 673144 258816 673150 258828
rect 675478 258816 675484 258828
rect 675536 258816 675542 258868
rect 672718 258408 672724 258460
rect 672776 258448 672782 258460
rect 675478 258448 675484 258460
rect 672776 258420 675484 258448
rect 672776 258408 672782 258420
rect 675478 258408 675484 258420
rect 675536 258408 675542 258460
rect 35802 258204 35808 258256
rect 35860 258244 35866 258256
rect 40034 258244 40040 258256
rect 35860 258216 40040 258244
rect 35860 258204 35866 258216
rect 40034 258204 40040 258216
rect 40092 258204 40098 258256
rect 35802 257116 35808 257168
rect 35860 257156 35866 257168
rect 39574 257156 39580 257168
rect 35860 257128 39580 257156
rect 35860 257116 35866 257128
rect 39574 257116 39580 257128
rect 39632 257116 39638 257168
rect 40402 256952 40408 256964
rect 36004 256924 40408 256952
rect 35802 256844 35808 256896
rect 35860 256884 35866 256896
rect 36004 256884 36032 256924
rect 40402 256912 40408 256924
rect 40460 256912 40466 256964
rect 35860 256856 36032 256884
rect 35860 256844 35866 256856
rect 42058 256844 42064 256896
rect 42116 256884 42122 256896
rect 49510 256884 49516 256896
rect 42116 256856 49516 256884
rect 42116 256844 42122 256856
rect 49510 256844 49516 256856
rect 49568 256844 49574 256896
rect 41690 256816 41696 256828
rect 40604 256788 41696 256816
rect 35618 256708 35624 256760
rect 35676 256748 35682 256760
rect 40604 256748 40632 256788
rect 41690 256776 41696 256788
rect 41748 256776 41754 256828
rect 35676 256720 40632 256748
rect 35676 256708 35682 256720
rect 510798 256708 510804 256760
rect 510856 256748 510862 256760
rect 567194 256748 567200 256760
rect 510856 256720 567200 256748
rect 510856 256708 510862 256720
rect 567194 256708 567200 256720
rect 567252 256708 567258 256760
rect 675846 256708 675852 256760
rect 675904 256748 675910 256760
rect 683114 256748 683120 256760
rect 675904 256720 683120 256748
rect 675904 256708 675910 256720
rect 683114 256708 683120 256720
rect 683172 256708 683178 256760
rect 35802 255688 35808 255740
rect 35860 255728 35866 255740
rect 41414 255728 41420 255740
rect 35860 255700 41420 255728
rect 35860 255688 35866 255700
rect 41414 255688 41420 255700
rect 41472 255688 41478 255740
rect 41690 255524 41696 255536
rect 41386 255496 41696 255524
rect 35618 255416 35624 255468
rect 35676 255456 35682 255468
rect 41386 255456 41414 255496
rect 41690 255484 41696 255496
rect 41748 255484 41754 255536
rect 42058 255484 42064 255536
rect 42116 255524 42122 255536
rect 42886 255524 42892 255536
rect 42116 255496 42892 255524
rect 42116 255484 42122 255496
rect 42886 255484 42892 255496
rect 42944 255484 42950 255536
rect 35676 255428 41414 255456
rect 35676 255416 35682 255428
rect 35802 255280 35808 255332
rect 35860 255320 35866 255332
rect 41690 255320 41696 255332
rect 35860 255292 41696 255320
rect 35860 255280 35866 255292
rect 41690 255280 41696 255292
rect 41748 255280 41754 255332
rect 42058 255280 42064 255332
rect 42116 255320 42122 255332
rect 45554 255320 45560 255332
rect 42116 255292 45560 255320
rect 42116 255280 42122 255292
rect 45554 255280 45560 255292
rect 45612 255280 45618 255332
rect 35526 254532 35532 254584
rect 35584 254572 35590 254584
rect 39298 254572 39304 254584
rect 35584 254544 39304 254572
rect 35584 254532 35590 254544
rect 39298 254532 39304 254544
rect 39356 254532 39362 254584
rect 39942 254368 39948 254380
rect 36004 254340 39948 254368
rect 35802 254260 35808 254312
rect 35860 254300 35866 254312
rect 36004 254300 36032 254340
rect 39942 254328 39948 254340
rect 40000 254328 40006 254380
rect 35860 254272 36032 254300
rect 35860 254260 35866 254272
rect 40310 254164 40316 254176
rect 36004 254136 40316 254164
rect 35342 254056 35348 254108
rect 35400 254096 35406 254108
rect 36004 254096 36032 254136
rect 40310 254124 40316 254136
rect 40368 254124 40374 254176
rect 35400 254068 36032 254096
rect 35400 254056 35406 254068
rect 35158 253920 35164 253972
rect 35216 253960 35222 253972
rect 41690 253960 41696 253972
rect 35216 253932 41696 253960
rect 35216 253920 35222 253932
rect 41690 253920 41696 253932
rect 41748 253920 41754 253972
rect 42058 253920 42064 253972
rect 42116 253960 42122 253972
rect 43806 253960 43812 253972
rect 42116 253932 43812 253960
rect 42116 253920 42122 253932
rect 43806 253920 43812 253932
rect 43864 253920 43870 253972
rect 669590 253172 669596 253224
rect 669648 253212 669654 253224
rect 675478 253212 675484 253224
rect 669648 253184 675484 253212
rect 669648 253172 669654 253184
rect 675478 253172 675484 253184
rect 675536 253172 675542 253224
rect 35802 252832 35808 252884
rect 35860 252872 35866 252884
rect 41690 252872 41696 252884
rect 35860 252844 41696 252872
rect 35860 252832 35866 252844
rect 41690 252832 41696 252844
rect 41748 252832 41754 252884
rect 42058 252832 42064 252884
rect 42116 252872 42122 252884
rect 42702 252872 42708 252884
rect 42116 252844 42708 252872
rect 42116 252832 42122 252844
rect 42702 252832 42708 252844
rect 42760 252832 42766 252884
rect 35618 252696 35624 252748
rect 35676 252736 35682 252748
rect 41690 252736 41696 252748
rect 35676 252708 41696 252736
rect 35676 252696 35682 252708
rect 41690 252696 41696 252708
rect 41748 252696 41754 252748
rect 35802 252560 35808 252612
rect 35860 252600 35866 252612
rect 41506 252600 41512 252612
rect 35860 252572 41512 252600
rect 35860 252560 35866 252572
rect 41506 252560 41512 252572
rect 41564 252560 41570 252612
rect 511902 252560 511908 252612
rect 511960 252600 511966 252612
rect 559558 252600 559564 252612
rect 511960 252572 559564 252600
rect 511960 252560 511966 252572
rect 559558 252560 559564 252572
rect 559616 252560 559622 252612
rect 35802 251608 35808 251660
rect 35860 251648 35866 251660
rect 40586 251648 40592 251660
rect 35860 251620 40592 251648
rect 35860 251608 35866 251620
rect 40586 251608 40592 251620
rect 40644 251608 40650 251660
rect 35802 251336 35808 251388
rect 35860 251376 35866 251388
rect 41322 251376 41328 251388
rect 35860 251348 41328 251376
rect 35860 251336 35866 251348
rect 41322 251336 41328 251348
rect 41380 251336 41386 251388
rect 35618 251200 35624 251252
rect 35676 251240 35682 251252
rect 41506 251240 41512 251252
rect 35676 251212 41512 251240
rect 35676 251200 35682 251212
rect 41506 251200 41512 251212
rect 41564 251200 41570 251252
rect 511534 250452 511540 250504
rect 511592 250492 511598 250504
rect 571334 250492 571340 250504
rect 511592 250464 571340 250492
rect 511592 250452 511598 250464
rect 571334 250452 571340 250464
rect 571392 250452 571398 250504
rect 669406 250384 669412 250436
rect 669464 250424 669470 250436
rect 672902 250424 672908 250436
rect 669464 250396 672908 250424
rect 669464 250384 669470 250396
rect 672902 250384 672908 250396
rect 672960 250384 672966 250436
rect 35802 250180 35808 250232
rect 35860 250220 35866 250232
rect 39390 250220 39396 250232
rect 35860 250192 39396 250220
rect 35860 250180 35866 250192
rect 39390 250180 39396 250192
rect 39448 250180 39454 250232
rect 40126 250016 40132 250028
rect 36004 249988 40132 250016
rect 35618 249908 35624 249960
rect 35676 249948 35682 249960
rect 36004 249948 36032 249988
rect 40126 249976 40132 249988
rect 40184 249976 40190 250028
rect 35676 249920 36032 249948
rect 35676 249908 35682 249920
rect 35434 249772 35440 249824
rect 35492 249812 35498 249824
rect 39574 249812 39580 249824
rect 35492 249784 39580 249812
rect 35492 249772 35498 249784
rect 39574 249772 39580 249784
rect 39632 249772 39638 249824
rect 35526 248684 35532 248736
rect 35584 248724 35590 248736
rect 39942 248724 39948 248736
rect 35584 248696 39948 248724
rect 35584 248684 35590 248696
rect 39942 248684 39948 248696
rect 40000 248684 40006 248736
rect 35802 248412 35808 248464
rect 35860 248452 35866 248464
rect 40126 248452 40132 248464
rect 35860 248424 40132 248452
rect 35860 248412 35866 248424
rect 40126 248412 40132 248424
rect 40184 248412 40190 248464
rect 674834 247868 674840 247920
rect 674892 247908 674898 247920
rect 675386 247908 675392 247920
rect 674892 247880 675392 247908
rect 674892 247868 674898 247880
rect 675386 247868 675392 247880
rect 675444 247868 675450 247920
rect 35802 247528 35808 247580
rect 35860 247568 35866 247580
rect 41506 247568 41512 247580
rect 35860 247540 41512 247568
rect 35860 247528 35866 247540
rect 41506 247528 41512 247540
rect 41564 247528 41570 247580
rect 42150 247460 42156 247512
rect 42208 247500 42214 247512
rect 129090 247500 129096 247512
rect 42208 247472 129096 247500
rect 42208 247460 42214 247472
rect 129090 247460 129096 247472
rect 129148 247460 129154 247512
rect 35618 247324 35624 247376
rect 35676 247364 35682 247376
rect 40126 247364 40132 247376
rect 35676 247336 40132 247364
rect 35676 247324 35682 247336
rect 40126 247324 40132 247336
rect 40184 247324 40190 247376
rect 35618 247188 35624 247240
rect 35676 247228 35682 247240
rect 41046 247228 41052 247240
rect 35676 247200 41052 247228
rect 35676 247188 35682 247200
rect 41046 247188 41052 247200
rect 41104 247188 41110 247240
rect 510982 247120 510988 247172
rect 511040 247160 511046 247172
rect 512638 247160 512644 247172
rect 511040 247132 512644 247160
rect 511040 247120 511046 247132
rect 512638 247120 512644 247132
rect 512696 247120 512702 247172
rect 35434 247052 35440 247104
rect 35492 247092 35498 247104
rect 41506 247092 41512 247104
rect 35492 247064 41512 247092
rect 35492 247052 35498 247064
rect 41506 247052 41512 247064
rect 41564 247052 41570 247104
rect 42058 247052 42064 247104
rect 42116 247092 42122 247104
rect 128998 247092 129004 247104
rect 42116 247064 129004 247092
rect 42116 247052 42122 247064
rect 128998 247052 129004 247064
rect 129056 247052 129062 247104
rect 674466 246984 674472 247036
rect 674524 247024 674530 247036
rect 675386 247024 675392 247036
rect 674524 246996 675392 247024
rect 674524 246984 674530 246996
rect 675386 246984 675392 246996
rect 675444 246984 675450 247036
rect 510798 246304 510804 246356
rect 510856 246344 510862 246356
rect 570046 246344 570052 246356
rect 510856 246316 570052 246344
rect 510856 246304 510862 246316
rect 570046 246304 570052 246316
rect 570104 246304 570110 246356
rect 663702 244876 663708 244928
rect 663760 244916 663766 244928
rect 669314 244916 669320 244928
rect 663760 244888 669320 244916
rect 663760 244876 663766 244888
rect 669314 244876 669320 244888
rect 669372 244876 669378 244928
rect 511258 242156 511264 242208
rect 511316 242196 511322 242208
rect 632698 242196 632704 242208
rect 511316 242168 632704 242196
rect 511316 242156 511322 242168
rect 632698 242156 632704 242168
rect 632756 242156 632762 242208
rect 673086 241680 673092 241732
rect 673144 241720 673150 241732
rect 675294 241720 675300 241732
rect 673144 241692 675300 241720
rect 673144 241680 673150 241692
rect 675294 241680 675300 241692
rect 675352 241680 675358 241732
rect 673362 241544 673368 241596
rect 673420 241584 673426 241596
rect 673420 241556 675340 241584
rect 673420 241544 673426 241556
rect 666370 241408 666376 241460
rect 666428 241448 666434 241460
rect 674926 241448 674932 241460
rect 666428 241420 674932 241448
rect 666428 241408 666434 241420
rect 674926 241408 674932 241420
rect 674984 241408 674990 241460
rect 675312 241120 675340 241556
rect 675294 241068 675300 241120
rect 675352 241068 675358 241120
rect 511902 240728 511908 240780
rect 511960 240768 511966 240780
rect 629938 240768 629944 240780
rect 511960 240740 629944 240768
rect 511960 240728 511966 240740
rect 629938 240728 629944 240740
rect 629996 240728 630002 240780
rect 42242 240048 42248 240100
rect 42300 240088 42306 240100
rect 45186 240088 45192 240100
rect 42300 240060 45192 240088
rect 42300 240048 42306 240060
rect 45186 240048 45192 240060
rect 45244 240048 45250 240100
rect 514018 238144 514024 238196
rect 514076 238184 514082 238196
rect 568758 238184 568764 238196
rect 514076 238156 568764 238184
rect 514076 238144 514082 238156
rect 568758 238144 568764 238156
rect 568816 238144 568822 238196
rect 674834 238076 674840 238128
rect 674892 238116 674898 238128
rect 675294 238116 675300 238128
rect 674892 238088 675300 238116
rect 674892 238076 674898 238088
rect 675294 238076 675300 238088
rect 675352 238076 675358 238128
rect 512638 238008 512644 238060
rect 512696 238048 512702 238060
rect 633434 238048 633440 238060
rect 512696 238020 633440 238048
rect 512696 238008 512702 238020
rect 633434 238008 633440 238020
rect 633492 238008 633498 238060
rect 42334 235900 42340 235952
rect 42392 235940 42398 235952
rect 44358 235940 44364 235952
rect 42392 235912 44364 235940
rect 42392 235900 42398 235912
rect 44358 235900 44364 235912
rect 44416 235900 44422 235952
rect 42334 234540 42340 234592
rect 42392 234580 42398 234592
rect 44542 234580 44548 234592
rect 42392 234552 44548 234580
rect 42392 234540 42398 234552
rect 44542 234540 44548 234552
rect 44600 234540 44606 234592
rect 510890 233996 510896 234048
rect 510948 234036 510954 234048
rect 577498 234036 577504 234048
rect 510948 234008 577504 234036
rect 510948 233996 510954 234008
rect 577498 233996 577504 234008
rect 577556 233996 577562 234048
rect 511074 233860 511080 233912
rect 511132 233900 511138 233912
rect 631318 233900 631324 233912
rect 511132 233872 631324 233900
rect 511132 233860 511138 233872
rect 631318 233860 631324 233872
rect 631376 233860 631382 233912
rect 42334 232024 42340 232076
rect 42392 232064 42398 232076
rect 45830 232064 45836 232076
rect 42392 232036 45836 232064
rect 42392 232024 42398 232036
rect 45830 232024 45836 232036
rect 45888 232024 45894 232076
rect 157334 231888 157340 231940
rect 157392 231928 157398 231940
rect 164878 231928 164884 231940
rect 157392 231900 164884 231928
rect 157392 231888 157398 231900
rect 164878 231888 164884 231900
rect 164936 231888 164942 231940
rect 190454 231888 190460 231940
rect 190512 231928 190518 231940
rect 191374 231928 191380 231940
rect 190512 231900 191380 231928
rect 190512 231888 190518 231900
rect 191374 231888 191380 231900
rect 191432 231888 191438 231940
rect 42334 231752 42340 231804
rect 42392 231792 42398 231804
rect 43622 231792 43628 231804
rect 42392 231764 43628 231792
rect 42392 231752 42398 231764
rect 43622 231752 43628 231764
rect 43680 231752 43686 231804
rect 54478 231752 54484 231804
rect 54536 231792 54542 231804
rect 641898 231792 641904 231804
rect 54536 231764 641904 231792
rect 54536 231752 54542 231764
rect 641898 231752 641904 231764
rect 641956 231752 641962 231804
rect 53098 231616 53104 231668
rect 53156 231656 53162 231668
rect 641714 231656 641720 231668
rect 53156 231628 641720 231656
rect 53156 231616 53162 231628
rect 641714 231616 641720 231628
rect 641772 231616 641778 231668
rect 46198 231480 46204 231532
rect 46256 231520 46262 231532
rect 643094 231520 643100 231532
rect 46256 231492 643100 231520
rect 46256 231480 46262 231492
rect 643094 231480 643100 231492
rect 643152 231480 643158 231532
rect 47578 231344 47584 231396
rect 47636 231384 47642 231396
rect 645854 231384 645860 231396
rect 47636 231356 645860 231384
rect 47636 231344 47642 231356
rect 645854 231344 645860 231356
rect 645912 231344 645918 231396
rect 51718 231208 51724 231260
rect 51776 231248 51782 231260
rect 650362 231248 650368 231260
rect 51776 231220 650368 231248
rect 51776 231208 51782 231220
rect 650362 231208 650368 231220
rect 650420 231208 650426 231260
rect 44818 231072 44824 231124
rect 44876 231112 44882 231124
rect 644474 231112 644480 231124
rect 44876 231084 644480 231112
rect 44876 231072 44882 231084
rect 644474 231072 644480 231084
rect 644532 231072 644538 231124
rect 129182 230936 129188 230988
rect 129240 230976 129246 230988
rect 661310 230976 661316 230988
rect 129240 230948 661316 230976
rect 129240 230936 129246 230948
rect 661310 230936 661316 230948
rect 661368 230936 661374 230988
rect 120718 230868 120724 230920
rect 120776 230908 120782 230920
rect 123294 230908 123300 230920
rect 120776 230880 123300 230908
rect 120776 230868 120782 230880
rect 123294 230868 123300 230880
rect 123352 230868 123358 230920
rect 176746 230840 176752 230852
rect 176626 230812 176752 230840
rect 99282 230732 99288 230784
rect 99340 230772 99346 230784
rect 176010 230772 176016 230784
rect 99340 230744 176016 230772
rect 99340 230732 99346 230744
rect 176010 230732 176016 230744
rect 176068 230732 176074 230784
rect 176470 230732 176476 230784
rect 176528 230772 176534 230784
rect 176626 230772 176654 230812
rect 176746 230800 176752 230812
rect 176804 230800 176810 230852
rect 178310 230800 178316 230852
rect 178368 230840 178374 230852
rect 185026 230840 185032 230852
rect 178368 230812 185032 230840
rect 178368 230800 178374 230812
rect 185026 230800 185032 230812
rect 185084 230800 185090 230852
rect 176528 230744 176654 230772
rect 176528 230732 176534 230744
rect 475194 230732 475200 230784
rect 475252 230772 475258 230784
rect 479978 230772 479984 230784
rect 475252 230744 479984 230772
rect 475252 230732 475258 230744
rect 479978 230732 479984 230744
rect 480036 230732 480042 230784
rect 481266 230732 481272 230784
rect 481324 230772 481330 230784
rect 489822 230772 489828 230784
rect 481324 230744 489828 230772
rect 481324 230732 481330 230744
rect 489822 230732 489828 230744
rect 489880 230732 489886 230784
rect 113082 230596 113088 230648
rect 113140 230636 113146 230648
rect 186682 230636 186688 230648
rect 113140 230608 186688 230636
rect 113140 230596 113146 230608
rect 186682 230596 186688 230608
rect 186740 230596 186746 230648
rect 194778 230596 194784 230648
rect 194836 230636 194842 230648
rect 195974 230636 195980 230648
rect 194836 230608 195980 230636
rect 194836 230596 194842 230608
rect 195974 230596 195980 230608
rect 196032 230596 196038 230648
rect 450538 230596 450544 230648
rect 450596 230636 450602 230648
rect 510614 230636 510620 230648
rect 450596 230608 510620 230636
rect 450596 230596 450602 230608
rect 510614 230596 510620 230608
rect 510672 230596 510678 230648
rect 123294 230460 123300 230512
rect 123352 230500 123358 230512
rect 147122 230500 147128 230512
rect 123352 230472 147128 230500
rect 123352 230460 123358 230472
rect 147122 230460 147128 230472
rect 147180 230460 147186 230512
rect 206002 230500 206008 230512
rect 154546 230472 206008 230500
rect 42150 230392 42156 230444
rect 42208 230432 42214 230444
rect 43070 230432 43076 230444
rect 42208 230404 43076 230432
rect 42208 230392 42214 230404
rect 43070 230392 43076 230404
rect 43128 230392 43134 230444
rect 107562 230392 107568 230444
rect 107620 230432 107626 230444
rect 107620 230404 115796 230432
rect 107620 230392 107626 230404
rect 42334 230256 42340 230308
rect 42392 230296 42398 230308
rect 43254 230296 43260 230308
rect 42392 230268 43260 230296
rect 42392 230256 42398 230268
rect 43254 230256 43260 230268
rect 43312 230256 43318 230308
rect 90358 230256 90364 230308
rect 90416 230296 90422 230308
rect 115768 230296 115796 230404
rect 117866 230392 117872 230444
rect 117924 230432 117930 230444
rect 123110 230432 123116 230444
rect 117924 230404 123116 230432
rect 117924 230392 117930 230404
rect 123110 230392 123116 230404
rect 123168 230392 123174 230444
rect 154546 230432 154574 230472
rect 206002 230460 206008 230472
rect 206060 230460 206066 230512
rect 441890 230500 441896 230512
rect 441586 230472 441896 230500
rect 147784 230404 154574 230432
rect 147490 230324 147496 230376
rect 147548 230364 147554 230376
rect 147784 230364 147812 230404
rect 213546 230392 213552 230444
rect 213604 230432 213610 230444
rect 253474 230432 253480 230444
rect 213604 230404 253480 230432
rect 213604 230392 213610 230404
rect 253474 230392 253480 230404
rect 253532 230392 253538 230444
rect 339586 230392 339592 230444
rect 339644 230432 339650 230444
rect 341058 230432 341064 230444
rect 339644 230404 341064 230432
rect 339644 230392 339650 230404
rect 341058 230392 341064 230404
rect 341116 230392 341122 230444
rect 407206 230392 407212 230444
rect 407264 230432 407270 230444
rect 412818 230432 412824 230444
rect 407264 230404 412824 230432
rect 407264 230392 407270 230404
rect 412818 230392 412824 230404
rect 412876 230392 412882 230444
rect 421282 230392 421288 230444
rect 421340 230432 421346 230444
rect 422202 230432 422208 230444
rect 421340 230404 422208 230432
rect 421340 230392 421346 230404
rect 422202 230392 422208 230404
rect 422260 230392 422266 230444
rect 427906 230392 427912 230444
rect 427964 230432 427970 230444
rect 429010 230432 429016 230444
rect 427964 230404 429016 230432
rect 427964 230392 427970 230404
rect 429010 230392 429016 230404
rect 429068 230392 429074 230444
rect 429194 230392 429200 230444
rect 429252 230432 429258 230444
rect 441586 230432 441614 230472
rect 441890 230460 441896 230472
rect 441948 230460 441954 230512
rect 442810 230460 442816 230512
rect 442868 230500 442874 230512
rect 442868 230472 444420 230500
rect 442868 230460 442874 230472
rect 429252 230404 441614 230432
rect 444392 230432 444420 230472
rect 451090 230460 451096 230512
rect 451148 230500 451154 230512
rect 512730 230500 512736 230512
rect 451148 230472 512736 230500
rect 451148 230460 451154 230472
rect 512730 230460 512736 230472
rect 512788 230460 512794 230512
rect 450722 230432 450728 230444
rect 444392 230404 450728 230432
rect 429252 230392 429258 230404
rect 450722 230392 450728 230404
rect 450780 230392 450786 230444
rect 147548 230336 147812 230364
rect 147548 230324 147554 230336
rect 159542 230324 159548 230376
rect 159600 230364 159606 230376
rect 167178 230364 167184 230376
rect 159600 230336 167184 230364
rect 159600 230324 159606 230336
rect 167178 230324 167184 230336
rect 167236 230324 167242 230376
rect 167822 230324 167828 230376
rect 167880 230364 167886 230376
rect 171594 230364 171600 230376
rect 167880 230336 171600 230364
rect 167880 230324 167886 230336
rect 171594 230324 171600 230336
rect 171652 230324 171658 230376
rect 200666 230324 200672 230376
rect 200724 230364 200730 230376
rect 200724 230336 203472 230364
rect 200724 230324 200730 230336
rect 147030 230296 147036 230308
rect 90416 230268 103514 230296
rect 115768 230268 147036 230296
rect 90416 230256 90422 230268
rect 103486 230160 103514 230268
rect 147030 230256 147036 230268
rect 147088 230256 147094 230308
rect 149330 230256 149336 230308
rect 149388 230296 149394 230308
rect 156322 230296 156328 230308
rect 149388 230268 156328 230296
rect 149388 230256 149394 230268
rect 156322 230256 156328 230268
rect 156380 230256 156386 230308
rect 171778 230256 171784 230308
rect 171836 230296 171842 230308
rect 200482 230296 200488 230308
rect 171836 230268 200488 230296
rect 171836 230256 171842 230268
rect 200482 230256 200488 230268
rect 200540 230256 200546 230308
rect 203444 230228 203472 230336
rect 204162 230324 204168 230376
rect 204220 230364 204226 230376
rect 205450 230364 205456 230376
rect 204220 230336 205456 230364
rect 204220 230324 204226 230336
rect 205450 230324 205456 230336
rect 205508 230324 205514 230376
rect 205726 230324 205732 230376
rect 205784 230364 205790 230376
rect 207658 230364 207664 230376
rect 205784 230336 207664 230364
rect 205784 230324 205790 230336
rect 207658 230324 207664 230336
rect 207716 230324 207722 230376
rect 298738 230324 298744 230376
rect 298796 230364 298802 230376
rect 299842 230364 299848 230376
rect 298796 230336 299848 230364
rect 298796 230324 298802 230336
rect 299842 230324 299848 230336
rect 299900 230324 299906 230376
rect 313458 230324 313464 230376
rect 313516 230364 313522 230376
rect 313918 230364 313924 230376
rect 313516 230336 313924 230364
rect 313516 230324 313522 230336
rect 313918 230324 313924 230336
rect 313976 230324 313982 230376
rect 319438 230324 319444 230376
rect 319496 230364 319502 230376
rect 321370 230364 321376 230376
rect 319496 230336 321376 230364
rect 319496 230324 319502 230336
rect 321370 230324 321376 230336
rect 321428 230324 321434 230376
rect 328822 230324 328828 230376
rect 328880 230364 328886 230376
rect 329650 230364 329656 230376
rect 328880 230336 329656 230364
rect 328880 230324 328886 230336
rect 329650 230324 329656 230336
rect 329708 230324 329714 230376
rect 331858 230324 331864 230376
rect 331916 230364 331922 230376
rect 333054 230364 333060 230376
rect 331916 230336 333060 230364
rect 331916 230324 331922 230336
rect 333054 230324 333060 230336
rect 333112 230324 333118 230376
rect 333514 230324 333520 230376
rect 333572 230364 333578 230376
rect 334526 230364 334532 230376
rect 333572 230336 334532 230364
rect 333572 230324 333578 230336
rect 334526 230324 334532 230336
rect 334584 230324 334590 230376
rect 335722 230324 335728 230376
rect 335780 230364 335786 230376
rect 337194 230364 337200 230376
rect 335780 230336 337200 230364
rect 335780 230324 335786 230336
rect 337194 230324 337200 230336
rect 337252 230324 337258 230376
rect 337378 230324 337384 230376
rect 337436 230364 337442 230376
rect 338298 230364 338304 230376
rect 337436 230336 338304 230364
rect 337436 230324 337442 230336
rect 338298 230324 338304 230336
rect 338356 230324 338362 230376
rect 342346 230324 342352 230376
rect 342404 230364 342410 230376
rect 343266 230364 343272 230376
rect 342404 230336 343272 230364
rect 342404 230324 342410 230336
rect 343266 230324 343272 230336
rect 343324 230324 343330 230376
rect 344002 230324 344008 230376
rect 344060 230364 344066 230376
rect 344922 230364 344928 230376
rect 344060 230336 344928 230364
rect 344060 230324 344066 230336
rect 344922 230324 344928 230336
rect 344980 230324 344986 230376
rect 348970 230324 348976 230376
rect 349028 230364 349034 230376
rect 352558 230364 352564 230376
rect 349028 230336 352564 230364
rect 349028 230324 349034 230336
rect 352558 230324 352564 230336
rect 352616 230324 352622 230376
rect 356146 230324 356152 230376
rect 356204 230364 356210 230376
rect 357250 230364 357256 230376
rect 356204 230336 357256 230364
rect 356204 230324 356210 230336
rect 357250 230324 357256 230336
rect 357308 230324 357314 230376
rect 360562 230324 360568 230376
rect 360620 230364 360626 230376
rect 362678 230364 362684 230376
rect 360620 230336 362684 230364
rect 360620 230324 360626 230336
rect 362678 230324 362684 230336
rect 362736 230324 362742 230376
rect 364426 230324 364432 230376
rect 364484 230364 364490 230376
rect 365438 230364 365444 230376
rect 364484 230336 365444 230364
rect 364484 230324 364490 230336
rect 365438 230324 365444 230336
rect 365496 230324 365502 230376
rect 367186 230324 367192 230376
rect 367244 230364 367250 230376
rect 368290 230364 368296 230376
rect 367244 230336 368296 230364
rect 367244 230324 367250 230336
rect 368290 230324 368296 230336
rect 368348 230324 368354 230376
rect 368842 230324 368848 230376
rect 368900 230364 368906 230376
rect 369762 230364 369768 230376
rect 368900 230336 369768 230364
rect 368900 230324 368906 230336
rect 369762 230324 369768 230336
rect 369820 230324 369826 230376
rect 371050 230324 371056 230376
rect 371108 230364 371114 230376
rect 372062 230364 372068 230376
rect 371108 230336 372068 230364
rect 371108 230324 371114 230336
rect 372062 230324 372068 230336
rect 372120 230324 372126 230376
rect 378226 230324 378232 230376
rect 378284 230364 378290 230376
rect 379330 230364 379336 230376
rect 378284 230336 379336 230364
rect 378284 230324 378290 230336
rect 379330 230324 379336 230336
rect 379388 230324 379394 230376
rect 385402 230324 385408 230376
rect 385460 230364 385466 230376
rect 386322 230364 386328 230376
rect 385460 230336 386328 230364
rect 385460 230324 385466 230336
rect 386322 230324 386328 230336
rect 386380 230324 386386 230376
rect 387058 230324 387064 230376
rect 387116 230364 387122 230376
rect 388438 230364 388444 230376
rect 387116 230336 388444 230364
rect 387116 230324 387122 230336
rect 388438 230324 388444 230336
rect 388496 230324 388502 230376
rect 403066 230324 403072 230376
rect 403124 230364 403130 230376
rect 404262 230364 404268 230376
rect 403124 230336 404268 230364
rect 403124 230324 403130 230336
rect 404262 230324 404268 230336
rect 404320 230324 404326 230376
rect 405826 230324 405832 230376
rect 405884 230364 405890 230376
rect 407022 230364 407028 230376
rect 405884 230336 407028 230364
rect 405884 230324 405890 230336
rect 407022 230324 407028 230336
rect 407080 230324 407086 230376
rect 413554 230324 413560 230376
rect 413612 230364 413618 230376
rect 418798 230364 418804 230376
rect 413612 230336 418804 230364
rect 413612 230324 413618 230336
rect 418798 230324 418804 230336
rect 418856 230324 418862 230376
rect 441706 230324 441712 230376
rect 441764 230364 441770 230376
rect 442902 230364 442908 230376
rect 441764 230336 442908 230364
rect 441764 230324 441770 230336
rect 442902 230324 442908 230336
rect 442960 230324 442966 230376
rect 443362 230324 443368 230376
rect 443420 230364 443426 230376
rect 444190 230364 444196 230376
rect 443420 230336 444196 230364
rect 443420 230324 443426 230336
rect 444190 230324 444196 230336
rect 444248 230324 444254 230376
rect 208026 230256 208032 230308
rect 208084 230296 208090 230308
rect 240226 230296 240232 230308
rect 208084 230268 240232 230296
rect 208084 230256 208090 230268
rect 240226 230256 240232 230268
rect 240284 230256 240290 230308
rect 244918 230256 244924 230308
rect 244976 230296 244982 230308
rect 246850 230296 246856 230308
rect 244976 230268 246856 230296
rect 244976 230256 244982 230268
rect 246850 230256 246856 230268
rect 246908 230256 246914 230308
rect 255958 230256 255964 230308
rect 256016 230296 256022 230308
rect 279970 230296 279976 230308
rect 256016 230268 279976 230296
rect 256016 230256 256022 230268
rect 279970 230256 279976 230268
rect 280028 230256 280034 230308
rect 285306 230256 285312 230308
rect 285364 230296 285370 230308
rect 291010 230296 291016 230308
rect 285364 230268 291016 230296
rect 285364 230256 285370 230268
rect 291010 230256 291016 230268
rect 291068 230256 291074 230308
rect 339034 230256 339040 230308
rect 339092 230296 339098 230308
rect 339862 230296 339868 230308
rect 339092 230268 339868 230296
rect 339092 230256 339098 230268
rect 339862 230256 339868 230268
rect 339920 230256 339926 230308
rect 390370 230256 390376 230308
rect 390428 230296 390434 230308
rect 399386 230296 399392 230308
rect 390428 230268 399392 230296
rect 390428 230256 390434 230268
rect 399386 230256 399392 230268
rect 399444 230256 399450 230308
rect 413278 230296 413284 230308
rect 411180 230268 413284 230296
rect 204898 230228 204904 230240
rect 157720 230200 166994 230228
rect 203444 230200 204904 230228
rect 122926 230160 122932 230172
rect 103486 230132 122932 230160
rect 122926 230120 122932 230132
rect 122984 230120 122990 230172
rect 123110 230120 123116 230172
rect 123168 230160 123174 230172
rect 157720 230160 157748 230200
rect 123168 230132 157748 230160
rect 166966 230160 166994 230200
rect 204898 230188 204904 230200
rect 204956 230188 204962 230240
rect 297634 230228 297640 230240
rect 296686 230200 297640 230228
rect 186130 230160 186136 230172
rect 166966 230132 186136 230160
rect 123168 230120 123174 230132
rect 186130 230120 186136 230132
rect 186188 230120 186194 230172
rect 186268 230120 186274 230172
rect 186326 230160 186332 230172
rect 187786 230160 187792 230172
rect 186326 230132 187792 230160
rect 186326 230120 186332 230132
rect 187786 230120 187792 230132
rect 187844 230120 187850 230172
rect 189902 230120 189908 230172
rect 189960 230160 189966 230172
rect 189960 230132 191236 230160
rect 189960 230120 189966 230132
rect 83458 229984 83464 230036
rect 83516 230024 83522 230036
rect 157288 230024 157294 230036
rect 83516 229996 157294 230024
rect 83516 229984 83522 229996
rect 157288 229984 157294 229996
rect 157346 229984 157352 230036
rect 162118 229984 162124 230036
rect 162176 230024 162182 230036
rect 171778 230024 171784 230036
rect 162176 229996 171784 230024
rect 162176 229984 162182 229996
rect 171778 229984 171784 229996
rect 171836 229984 171842 230036
rect 171962 229984 171968 230036
rect 172020 230024 172026 230036
rect 174538 230024 174544 230036
rect 172020 229996 174544 230024
rect 172020 229984 172026 229996
rect 174538 229984 174544 229996
rect 174596 229984 174602 230036
rect 174906 229984 174912 230036
rect 174964 230024 174970 230036
rect 176378 230024 176384 230036
rect 174964 229996 176384 230024
rect 174964 229984 174970 229996
rect 176378 229984 176384 229996
rect 176436 229984 176442 230036
rect 176562 229984 176568 230036
rect 176620 230024 176626 230036
rect 190362 230024 190368 230036
rect 176620 229996 190368 230024
rect 176620 229984 176626 229996
rect 190362 229984 190368 229996
rect 190420 229984 190426 230036
rect 191208 230024 191236 230132
rect 191374 230120 191380 230172
rect 191432 230160 191438 230172
rect 194410 230160 194416 230172
rect 191432 230132 194416 230160
rect 191432 230120 191438 230132
rect 194410 230120 194416 230132
rect 194468 230120 194474 230172
rect 194594 230120 194600 230172
rect 194652 230160 194658 230172
rect 198826 230160 198832 230172
rect 194652 230132 198832 230160
rect 194652 230120 194658 230132
rect 198826 230120 198832 230132
rect 198884 230120 198890 230172
rect 199194 230120 199200 230172
rect 199252 230160 199258 230172
rect 203242 230160 203248 230172
rect 199252 230132 203248 230160
rect 199252 230120 199258 230132
rect 203242 230120 203248 230132
rect 203300 230120 203306 230172
rect 205542 230120 205548 230172
rect 205600 230160 205606 230172
rect 244642 230160 244648 230172
rect 205600 230132 244648 230160
rect 205600 230120 205606 230132
rect 244642 230120 244648 230132
rect 244700 230120 244706 230172
rect 247770 230120 247776 230172
rect 247828 230160 247834 230172
rect 275554 230160 275560 230172
rect 247828 230132 275560 230160
rect 247828 230120 247834 230132
rect 275554 230120 275560 230132
rect 275612 230120 275618 230172
rect 279786 230120 279792 230172
rect 279844 230160 279850 230172
rect 296686 230160 296714 230200
rect 297634 230188 297640 230200
rect 297692 230188 297698 230240
rect 313918 230188 313924 230240
rect 313976 230228 313982 230240
rect 315298 230228 315304 230240
rect 313976 230200 315304 230228
rect 313976 230188 313982 230200
rect 315298 230188 315304 230200
rect 315356 230188 315362 230240
rect 341242 230188 341248 230240
rect 341300 230228 341306 230240
rect 343818 230228 343824 230240
rect 341300 230200 343824 230228
rect 341300 230188 341306 230200
rect 343818 230188 343824 230200
rect 343876 230188 343882 230240
rect 355042 230188 355048 230240
rect 355100 230228 355106 230240
rect 360838 230228 360844 230240
rect 355100 230200 360844 230228
rect 355100 230188 355106 230200
rect 360838 230188 360844 230200
rect 360896 230188 360902 230240
rect 378778 230188 378784 230240
rect 378836 230228 378842 230240
rect 380158 230228 380164 230240
rect 378836 230200 380164 230228
rect 378836 230188 378842 230200
rect 380158 230188 380164 230200
rect 380216 230188 380222 230240
rect 380986 230188 380992 230240
rect 381044 230228 381050 230240
rect 389726 230228 389732 230240
rect 381044 230200 389732 230228
rect 381044 230188 381050 230200
rect 389726 230188 389732 230200
rect 389784 230188 389790 230240
rect 404722 230188 404728 230240
rect 404780 230228 404786 230240
rect 411180 230228 411208 230268
rect 413278 230256 413284 230268
rect 413336 230256 413342 230308
rect 420178 230256 420184 230308
rect 420236 230296 420242 230308
rect 434898 230296 434904 230308
rect 420236 230268 434904 230296
rect 420236 230256 420242 230268
rect 434898 230256 434904 230268
rect 434956 230256 434962 230308
rect 435082 230256 435088 230308
rect 435140 230296 435146 230308
rect 436002 230296 436008 230308
rect 435140 230268 436008 230296
rect 435140 230256 435146 230268
rect 436002 230256 436008 230268
rect 436060 230256 436066 230308
rect 446122 230256 446128 230308
rect 446180 230296 446186 230308
rect 505738 230296 505744 230308
rect 446180 230268 505744 230296
rect 446180 230256 446186 230268
rect 505738 230256 505744 230268
rect 505796 230256 505802 230308
rect 404780 230200 411208 230228
rect 404780 230188 404786 230200
rect 279844 230132 296714 230160
rect 279844 230120 279850 230132
rect 344554 230120 344560 230172
rect 344612 230160 344618 230172
rect 349798 230160 349804 230172
rect 344612 230132 349804 230160
rect 344612 230120 344618 230132
rect 349798 230120 349804 230132
rect 349856 230120 349862 230172
rect 369394 230120 369400 230172
rect 369452 230160 369458 230172
rect 371878 230160 371884 230172
rect 369452 230132 371884 230160
rect 369452 230120 369458 230132
rect 371878 230120 371884 230132
rect 371936 230120 371942 230172
rect 372706 230120 372712 230172
rect 372764 230160 372770 230172
rect 392210 230160 392216 230172
rect 372764 230132 373994 230160
rect 372764 230120 372770 230132
rect 297358 230052 297364 230104
rect 297416 230092 297422 230104
rect 299290 230092 299296 230104
rect 297416 230064 299296 230092
rect 297416 230052 297422 230064
rect 299290 230052 299296 230064
rect 299348 230052 299354 230104
rect 320818 230052 320824 230104
rect 320876 230092 320882 230104
rect 321922 230092 321928 230104
rect 320876 230064 321928 230092
rect 320876 230052 320882 230064
rect 321922 230052 321928 230064
rect 321980 230052 321986 230104
rect 340690 230052 340696 230104
rect 340748 230092 340754 230104
rect 344278 230092 344284 230104
rect 340748 230064 344284 230092
rect 340748 230052 340754 230064
rect 344278 230052 344284 230064
rect 344336 230052 344342 230104
rect 357434 230052 357440 230104
rect 357492 230092 357498 230104
rect 363598 230092 363604 230104
rect 357492 230064 363604 230092
rect 357492 230052 357498 230064
rect 363598 230052 363604 230064
rect 363656 230052 363662 230104
rect 196618 230024 196624 230036
rect 191208 229996 196624 230024
rect 196618 229984 196624 229996
rect 196676 229984 196682 230036
rect 196802 229984 196808 230036
rect 196860 230024 196866 230036
rect 235810 230024 235816 230036
rect 196860 229996 235816 230024
rect 196860 229984 196866 229996
rect 235810 229984 235816 229996
rect 235868 229984 235874 230036
rect 241606 229984 241612 230036
rect 241664 230024 241670 230036
rect 271138 230024 271144 230036
rect 241664 229996 271144 230024
rect 241664 229984 241670 229996
rect 271138 229984 271144 229996
rect 271196 229984 271202 230036
rect 275646 229984 275652 230036
rect 275704 230024 275710 230036
rect 293218 230024 293224 230036
rect 275704 229996 293224 230024
rect 275704 229984 275710 229996
rect 293218 229984 293224 229996
rect 293276 229984 293282 230036
rect 367738 229984 367744 230036
rect 367796 230024 367802 230036
rect 370866 230024 370872 230036
rect 367796 229996 370872 230024
rect 367796 229984 367802 229996
rect 370866 229984 370872 229996
rect 370924 229984 370930 230036
rect 190656 229928 191052 229956
rect 77938 229848 77944 229900
rect 77996 229888 78002 229900
rect 133046 229888 133052 229900
rect 77996 229860 133052 229888
rect 77996 229848 78002 229860
rect 133046 229848 133052 229860
rect 133104 229848 133110 229900
rect 133230 229848 133236 229900
rect 133288 229888 133294 229900
rect 182818 229888 182824 229900
rect 133288 229860 182824 229888
rect 133288 229848 133294 229860
rect 182818 229848 182824 229860
rect 182876 229848 182882 229900
rect 183462 229848 183468 229900
rect 183520 229888 183526 229900
rect 190656 229888 190684 229928
rect 183520 229860 190684 229888
rect 191024 229888 191052 229928
rect 231394 229888 231400 229900
rect 191024 229860 231400 229888
rect 183520 229848 183526 229860
rect 231394 229848 231400 229860
rect 231452 229848 231458 229900
rect 233234 229848 233240 229900
rect 233292 229888 233298 229900
rect 266722 229888 266728 229900
rect 233292 229860 266728 229888
rect 233292 229848 233298 229860
rect 266722 229848 266728 229860
rect 266780 229848 266786 229900
rect 266998 229848 267004 229900
rect 267056 229888 267062 229900
rect 288802 229888 288808 229900
rect 267056 229860 288808 229888
rect 267056 229848 267062 229860
rect 288802 229848 288808 229860
rect 288860 229848 288866 229900
rect 338482 229848 338488 229900
rect 338540 229888 338546 229900
rect 339310 229888 339316 229900
rect 338540 229860 339316 229888
rect 338540 229848 338546 229860
rect 339310 229848 339316 229860
rect 339368 229848 339374 229900
rect 359458 229848 359464 229900
rect 359516 229888 359522 229900
rect 369118 229888 369124 229900
rect 359516 229860 369124 229888
rect 359516 229848 359522 229860
rect 369118 229848 369124 229860
rect 369176 229848 369182 229900
rect 373966 229888 373994 230132
rect 389928 230132 392216 230160
rect 374362 229984 374368 230036
rect 374420 230024 374426 230036
rect 377398 230024 377404 230036
rect 374420 229996 377404 230024
rect 374420 229984 374426 229996
rect 377398 229984 377404 229996
rect 377456 229984 377462 230036
rect 379146 229984 379152 230036
rect 379204 230024 379210 230036
rect 389928 230024 389956 230132
rect 392210 230120 392216 230132
rect 392268 230120 392274 230172
rect 392394 230120 392400 230172
rect 392452 230160 392458 230172
rect 394970 230160 394976 230172
rect 392452 230132 394976 230160
rect 392452 230120 392458 230132
rect 394970 230120 394976 230132
rect 395028 230120 395034 230172
rect 411346 230120 411352 230172
rect 411404 230160 411410 230172
rect 414842 230160 414848 230172
rect 411404 230132 414848 230160
rect 411404 230120 411410 230132
rect 414842 230120 414848 230132
rect 414900 230120 414906 230172
rect 415210 230120 415216 230172
rect 415268 230160 415274 230172
rect 441706 230160 441712 230172
rect 415268 230132 441712 230160
rect 415268 230120 415274 230132
rect 441706 230120 441712 230132
rect 441764 230120 441770 230172
rect 441890 230120 441896 230172
rect 441948 230160 441954 230172
rect 447502 230160 447508 230172
rect 441948 230132 447508 230160
rect 441948 230120 441954 230132
rect 447502 230120 447508 230132
rect 447560 230120 447566 230172
rect 455506 230120 455512 230172
rect 455564 230160 455570 230172
rect 456702 230160 456708 230172
rect 455564 230132 456708 230160
rect 455564 230120 455570 230132
rect 456702 230120 456708 230132
rect 456760 230120 456766 230172
rect 457162 230120 457168 230172
rect 457220 230160 457226 230172
rect 458082 230160 458088 230172
rect 457220 230132 458088 230160
rect 457220 230120 457226 230132
rect 458082 230120 458088 230132
rect 458140 230120 458146 230172
rect 458450 230120 458456 230172
rect 458508 230160 458514 230172
rect 475194 230160 475200 230172
rect 458508 230132 475200 230160
rect 458508 230120 458514 230132
rect 475194 230120 475200 230132
rect 475252 230120 475258 230172
rect 476482 230120 476488 230172
rect 476540 230160 476546 230172
rect 479518 230160 479524 230172
rect 476540 230132 479524 230160
rect 476540 230120 476546 230132
rect 479518 230120 479524 230132
rect 479576 230120 479582 230172
rect 479978 230120 479984 230172
rect 480036 230160 480042 230172
rect 481358 230160 481364 230172
rect 480036 230132 481364 230160
rect 480036 230120 480042 230132
rect 481358 230120 481364 230132
rect 481416 230120 481422 230172
rect 482554 230120 482560 230172
rect 482612 230160 482618 230172
rect 541986 230160 541992 230172
rect 482612 230132 541992 230160
rect 482612 230120 482618 230132
rect 541986 230120 541992 230132
rect 542044 230120 542050 230172
rect 379204 229996 389956 230024
rect 379204 229984 379210 229996
rect 392026 229984 392032 230036
rect 392084 230024 392090 230036
rect 396718 230024 396724 230036
rect 392084 229996 396724 230024
rect 392084 229984 392090 229996
rect 396718 229984 396724 229996
rect 396776 229984 396782 230036
rect 398742 229984 398748 230036
rect 398800 230024 398806 230036
rect 398800 229996 413968 230024
rect 398800 229984 398806 229996
rect 382274 229888 382280 229900
rect 373966 229860 382280 229888
rect 382274 229848 382280 229860
rect 382332 229848 382338 229900
rect 391198 229888 391204 229900
rect 382476 229860 391204 229888
rect 300578 229780 300584 229832
rect 300636 229820 300642 229832
rect 301498 229820 301504 229832
rect 300636 229792 301504 229820
rect 300636 229780 300642 229792
rect 301498 229780 301504 229792
rect 301556 229780 301562 229832
rect 67542 229712 67548 229764
rect 67600 229752 67606 229764
rect 149330 229752 149336 229764
rect 67600 229724 149336 229752
rect 67600 229712 67606 229724
rect 149330 229712 149336 229724
rect 149388 229712 149394 229764
rect 150986 229712 150992 229764
rect 151044 229752 151050 229764
rect 154114 229752 154120 229764
rect 151044 229724 154120 229752
rect 151044 229712 151050 229724
rect 154114 229712 154120 229724
rect 154172 229712 154178 229764
rect 154574 229712 154580 229764
rect 154632 229752 154638 229764
rect 157978 229752 157984 229764
rect 154632 229724 157984 229752
rect 154632 229712 154638 229724
rect 157978 229712 157984 229724
rect 158036 229712 158042 229764
rect 158162 229712 158168 229764
rect 158220 229752 158226 229764
rect 160738 229752 160744 229764
rect 158220 229724 160744 229752
rect 158220 229712 158226 229724
rect 160738 229712 160744 229724
rect 160796 229712 160802 229764
rect 161106 229712 161112 229764
rect 161164 229752 161170 229764
rect 163498 229752 163504 229764
rect 161164 229724 163504 229752
rect 161164 229712 161170 229724
rect 163498 229712 163504 229724
rect 163556 229712 163562 229764
rect 163958 229712 163964 229764
rect 164016 229752 164022 229764
rect 171778 229752 171784 229764
rect 164016 229724 171784 229752
rect 164016 229712 164022 229724
rect 171778 229712 171784 229724
rect 171836 229712 171842 229764
rect 171962 229712 171968 229764
rect 172020 229752 172026 229764
rect 218146 229752 218152 229764
rect 172020 229724 218152 229752
rect 172020 229712 172026 229724
rect 218146 229712 218152 229724
rect 218204 229712 218210 229764
rect 220538 229712 220544 229764
rect 220596 229752 220602 229764
rect 257890 229752 257896 229764
rect 220596 229724 257896 229752
rect 220596 229712 220602 229724
rect 257890 229712 257896 229724
rect 257948 229712 257954 229764
rect 261570 229712 261576 229764
rect 261628 229752 261634 229764
rect 284386 229752 284392 229764
rect 261628 229724 284392 229752
rect 261628 229712 261634 229724
rect 284386 229712 284392 229724
rect 284444 229712 284450 229764
rect 289722 229712 289728 229764
rect 289780 229752 289786 229764
rect 289780 229724 296714 229752
rect 289780 229712 289786 229724
rect 296686 229684 296714 229724
rect 305638 229712 305644 229764
rect 305696 229752 305702 229764
rect 313090 229752 313096 229764
rect 305696 229724 313096 229752
rect 305696 229712 305702 229724
rect 313090 229712 313096 229724
rect 313148 229712 313154 229764
rect 342898 229712 342904 229764
rect 342956 229752 342962 229764
rect 348418 229752 348424 229764
rect 342956 229724 348424 229752
rect 342956 229712 342962 229724
rect 348418 229712 348424 229724
rect 348476 229712 348482 229764
rect 361666 229712 361672 229764
rect 361724 229752 361730 229764
rect 373994 229752 374000 229764
rect 361724 229724 374000 229752
rect 361724 229712 361730 229724
rect 373994 229712 374000 229724
rect 374052 229712 374058 229764
rect 377122 229712 377128 229764
rect 377180 229752 377186 229764
rect 382476 229752 382504 229860
rect 391198 229848 391204 229860
rect 391256 229848 391262 229900
rect 391474 229848 391480 229900
rect 391532 229888 391538 229900
rect 392578 229888 392584 229900
rect 391532 229860 392584 229888
rect 391532 229848 391538 229860
rect 392578 229848 392584 229860
rect 392636 229848 392642 229900
rect 400858 229848 400864 229900
rect 400916 229888 400922 229900
rect 413940 229888 413968 229996
rect 414106 229984 414112 230036
rect 414164 230024 414170 230036
rect 415302 230024 415308 230036
rect 414164 229996 415308 230024
rect 414164 229984 414170 229996
rect 415302 229984 415308 229996
rect 415360 229984 415366 230036
rect 416314 229984 416320 230036
rect 416372 230024 416378 230036
rect 416372 229996 422294 230024
rect 416372 229984 416378 229996
rect 416038 229888 416044 229900
rect 400916 229860 412634 229888
rect 413940 229860 416044 229888
rect 400916 229848 400922 229860
rect 391658 229752 391664 229764
rect 377180 229724 382504 229752
rect 383626 229724 391664 229752
rect 377180 229712 377186 229724
rect 304258 229684 304264 229696
rect 296686 229656 304264 229684
rect 304258 229644 304264 229656
rect 304316 229644 304322 229696
rect 122926 229576 122932 229628
rect 122984 229616 122990 229628
rect 132862 229616 132868 229628
rect 122984 229588 132868 229616
rect 122984 229576 122990 229588
rect 132862 229576 132868 229588
rect 132920 229576 132926 229628
rect 194778 229616 194784 229628
rect 133432 229588 194784 229616
rect 130102 229440 130108 229492
rect 130160 229480 130166 229492
rect 133230 229480 133236 229492
rect 130160 229452 133236 229480
rect 130160 229440 130166 229452
rect 133230 229440 133236 229452
rect 133288 229440 133294 229492
rect 126882 229304 126888 229356
rect 126940 229344 126946 229356
rect 133432 229344 133460 229588
rect 194778 229576 194784 229588
rect 194836 229576 194842 229628
rect 195238 229576 195244 229628
rect 195296 229616 195302 229628
rect 200482 229616 200488 229628
rect 195296 229588 200488 229616
rect 195296 229576 195302 229588
rect 200482 229576 200488 229588
rect 200540 229576 200546 229628
rect 201218 229576 201224 229628
rect 201276 229616 201282 229628
rect 226978 229616 226984 229628
rect 201276 229588 226984 229616
rect 201276 229576 201282 229588
rect 226978 229576 226984 229588
rect 227036 229576 227042 229628
rect 230658 229576 230664 229628
rect 230716 229616 230722 229628
rect 262306 229616 262312 229628
rect 230716 229588 262312 229616
rect 230716 229576 230722 229588
rect 262306 229576 262312 229588
rect 262364 229576 262370 229628
rect 313182 229576 313188 229628
rect 313240 229616 313246 229628
rect 319714 229616 319720 229628
rect 313240 229588 319720 229616
rect 313240 229576 313246 229588
rect 319714 229576 319720 229588
rect 319772 229576 319778 229628
rect 374914 229576 374920 229628
rect 374972 229616 374978 229628
rect 383626 229616 383654 229724
rect 391658 229712 391664 229724
rect 391716 229712 391722 229764
rect 392946 229712 392952 229764
rect 393004 229752 393010 229764
rect 399570 229752 399576 229764
rect 393004 229724 399576 229752
rect 393004 229712 393010 229724
rect 399570 229712 399576 229724
rect 399628 229712 399634 229764
rect 412606 229752 412634 229860
rect 416038 229848 416044 229860
rect 416096 229848 416102 229900
rect 419074 229848 419080 229900
rect 419132 229888 419138 229900
rect 422266 229888 422294 229996
rect 424042 229984 424048 230036
rect 424100 230024 424106 230036
rect 429194 230024 429200 230036
rect 424100 229996 429200 230024
rect 424100 229984 424106 229996
rect 429194 229984 429200 229996
rect 429252 229984 429258 230036
rect 429378 229984 429384 230036
rect 429436 230024 429442 230036
rect 446766 230024 446772 230036
rect 429436 229996 446772 230024
rect 429436 229984 429442 229996
rect 446766 229984 446772 229996
rect 446824 229984 446830 230036
rect 448146 229984 448152 230036
rect 448204 230024 448210 230036
rect 507118 230024 507124 230036
rect 448204 229996 507124 230024
rect 448204 229984 448210 229996
rect 507118 229984 507124 229996
rect 507176 229984 507182 230036
rect 427078 229888 427084 229900
rect 419132 229860 420684 229888
rect 422266 229860 427084 229888
rect 419132 229848 419138 229860
rect 420178 229752 420184 229764
rect 412606 229724 420184 229752
rect 420178 229712 420184 229724
rect 420236 229712 420242 229764
rect 420656 229752 420684 229860
rect 427078 229848 427084 229860
rect 427136 229848 427142 229900
rect 428458 229848 428464 229900
rect 428516 229888 428522 229900
rect 473446 229888 473452 229900
rect 428516 229860 473452 229888
rect 428516 229848 428522 229860
rect 473446 229848 473452 229860
rect 473504 229848 473510 229900
rect 475194 229848 475200 229900
rect 475252 229888 475258 229900
rect 484026 229888 484032 229900
rect 475252 229860 484032 229888
rect 475252 229848 475258 229860
rect 484026 229848 484032 229860
rect 484084 229848 484090 229900
rect 484210 229848 484216 229900
rect 484268 229888 484274 229900
rect 487338 229888 487344 229900
rect 484268 229860 487344 229888
rect 484268 229848 484274 229860
rect 487338 229848 487344 229860
rect 487396 229848 487402 229900
rect 487522 229848 487528 229900
rect 487580 229888 487586 229900
rect 487580 229860 499344 229888
rect 487580 229848 487586 229860
rect 428090 229752 428096 229764
rect 420656 229724 428096 229752
rect 428090 229712 428096 229724
rect 428148 229712 428154 229764
rect 438946 229712 438952 229764
rect 439004 229752 439010 229764
rect 484854 229752 484860 229764
rect 439004 229724 484860 229752
rect 439004 229712 439010 229724
rect 484854 229712 484860 229724
rect 484912 229712 484918 229764
rect 485038 229712 485044 229764
rect 485096 229752 485102 229764
rect 495388 229752 495394 229764
rect 485096 229724 495394 229752
rect 485096 229712 485102 229724
rect 495388 229712 495394 229724
rect 495446 229712 495452 229764
rect 499316 229752 499344 229860
rect 499482 229848 499488 229900
rect 499540 229888 499546 229900
rect 551922 229888 551928 229900
rect 499540 229860 551928 229888
rect 499540 229848 499546 229860
rect 551922 229848 551928 229860
rect 551980 229848 551986 229900
rect 558178 229752 558184 229764
rect 499316 229724 558184 229752
rect 558178 229712 558184 229724
rect 558236 229712 558242 229764
rect 499114 229684 499120 229696
rect 495728 229656 499120 229684
rect 374972 229588 383654 229616
rect 374972 229576 374978 229588
rect 389266 229576 389272 229628
rect 389324 229616 389330 229628
rect 390462 229616 390468 229628
rect 389324 229588 390468 229616
rect 389324 229576 389330 229588
rect 390462 229576 390468 229588
rect 390520 229576 390526 229628
rect 394234 229576 394240 229628
rect 394292 229616 394298 229628
rect 400858 229616 400864 229628
rect 394292 229588 400864 229616
rect 394292 229576 394298 229588
rect 400858 229576 400864 229588
rect 400916 229576 400922 229628
rect 407482 229576 407488 229628
rect 407540 229616 407546 229628
rect 424318 229616 424324 229628
rect 407540 229588 424324 229616
rect 407540 229576 407546 229588
rect 424318 229576 424324 229588
rect 424376 229576 424382 229628
rect 425698 229576 425704 229628
rect 425756 229616 425762 229628
rect 425756 229588 428688 229616
rect 425756 229576 425762 229588
rect 126940 229316 133460 229344
rect 133524 229452 152780 229480
rect 126940 229304 126946 229316
rect 133046 229168 133052 229220
rect 133104 229208 133110 229220
rect 133524 229208 133552 229452
rect 133690 229304 133696 229356
rect 133748 229344 133754 229356
rect 152550 229344 152556 229356
rect 133748 229316 152556 229344
rect 133748 229304 133754 229316
rect 152550 229304 152556 229316
rect 152608 229304 152614 229356
rect 152752 229344 152780 229452
rect 153010 229440 153016 229492
rect 153068 229480 153074 229492
rect 162118 229480 162124 229492
rect 153068 229452 162124 229480
rect 153068 229440 153074 229452
rect 162118 229440 162124 229452
rect 162176 229440 162182 229492
rect 163590 229440 163596 229492
rect 163648 229480 163654 229492
rect 165706 229480 165712 229492
rect 163648 229452 165712 229480
rect 163648 229440 163654 229452
rect 165706 229440 165712 229452
rect 165764 229440 165770 229492
rect 166994 229440 167000 229492
rect 167052 229480 167058 229492
rect 171594 229480 171600 229492
rect 167052 229452 171600 229480
rect 167052 229440 167058 229452
rect 171594 229440 171600 229452
rect 171652 229440 171658 229492
rect 171778 229440 171784 229492
rect 171836 229480 171842 229492
rect 200666 229480 200672 229492
rect 171836 229452 200672 229480
rect 171836 229440 171842 229452
rect 200666 229440 200672 229452
rect 200724 229440 200730 229492
rect 200850 229440 200856 229492
rect 200908 229480 200914 229492
rect 208026 229480 208032 229492
rect 200908 229452 208032 229480
rect 200908 229440 200914 229452
rect 208026 229440 208032 229452
rect 208084 229440 208090 229492
rect 208210 229440 208216 229492
rect 208268 229480 208274 229492
rect 209314 229480 209320 229492
rect 208268 229452 209320 229480
rect 208268 229440 208274 229452
rect 209314 229440 209320 229452
rect 209372 229440 209378 229492
rect 211154 229440 211160 229492
rect 211212 229480 211218 229492
rect 220906 229480 220912 229492
rect 211212 229452 220912 229480
rect 211212 229440 211218 229452
rect 220906 229440 220912 229452
rect 220964 229440 220970 229492
rect 225966 229440 225972 229492
rect 226024 229480 226030 229492
rect 229738 229480 229744 229492
rect 226024 229452 229744 229480
rect 226024 229440 226030 229452
rect 229738 229440 229744 229452
rect 229796 229440 229802 229492
rect 249058 229480 249064 229492
rect 238726 229452 249064 229480
rect 156322 229344 156328 229356
rect 152752 229316 156328 229344
rect 156322 229304 156328 229316
rect 156380 229304 156386 229356
rect 156874 229304 156880 229356
rect 156932 229344 156938 229356
rect 200068 229344 200074 229356
rect 156932 229316 200074 229344
rect 156932 229304 156938 229316
rect 200068 229304 200074 229316
rect 200126 229304 200132 229356
rect 200482 229304 200488 229356
rect 200540 229344 200546 229356
rect 213730 229344 213736 229356
rect 200540 229316 213736 229344
rect 200540 229304 200546 229316
rect 213730 229304 213736 229316
rect 213788 229304 213794 229356
rect 220814 229304 220820 229356
rect 220872 229344 220878 229356
rect 225322 229344 225328 229356
rect 220872 229316 225328 229344
rect 220872 229304 220878 229316
rect 225322 229304 225328 229316
rect 225380 229304 225386 229356
rect 226978 229304 226984 229356
rect 227036 229344 227042 229356
rect 236362 229344 236368 229356
rect 227036 229316 236368 229344
rect 227036 229304 227042 229316
rect 236362 229304 236368 229316
rect 236420 229304 236426 229356
rect 133104 229180 133552 229208
rect 133104 229168 133110 229180
rect 133874 229168 133880 229220
rect 133932 229208 133938 229220
rect 147306 229208 147312 229220
rect 133932 229180 147312 229208
rect 133932 229168 133938 229180
rect 147306 229168 147312 229180
rect 147364 229168 147370 229220
rect 147674 229168 147680 229220
rect 147732 229208 147738 229220
rect 157288 229208 157294 229220
rect 147732 229180 157294 229208
rect 147732 229168 147738 229180
rect 157288 229168 157294 229180
rect 157346 229168 157352 229220
rect 157610 229168 157616 229220
rect 157668 229208 157674 229220
rect 195238 229208 195244 229220
rect 157668 229180 195244 229208
rect 157668 229168 157674 229180
rect 195238 229168 195244 229180
rect 195296 229168 195302 229220
rect 196526 229168 196532 229220
rect 196584 229208 196590 229220
rect 201034 229208 201040 229220
rect 196584 229180 201040 229208
rect 196584 229168 196590 229180
rect 201034 229168 201040 229180
rect 201092 229168 201098 229220
rect 201402 229168 201408 229220
rect 201460 229208 201466 229220
rect 208210 229208 208216 229220
rect 201460 229180 208216 229208
rect 201460 229168 201466 229180
rect 208210 229168 208216 229180
rect 208268 229168 208274 229220
rect 208394 229168 208400 229220
rect 208452 229208 208458 229220
rect 216490 229208 216496 229220
rect 208452 229180 216496 229208
rect 208452 229168 208458 229180
rect 216490 229168 216496 229180
rect 216548 229168 216554 229220
rect 222930 229168 222936 229220
rect 222988 229208 222994 229220
rect 238726 229208 238754 229452
rect 249058 229440 249064 229452
rect 249116 229440 249122 229492
rect 385954 229440 385960 229492
rect 386012 229480 386018 229492
rect 392394 229480 392400 229492
rect 386012 229452 392400 229480
rect 386012 229440 386018 229452
rect 392394 229440 392400 229452
rect 392452 229440 392458 229492
rect 396994 229440 397000 229492
rect 397052 229480 397058 229492
rect 397052 229452 402974 229480
rect 397052 229440 397058 229452
rect 290458 229372 290464 229424
rect 290516 229412 290522 229424
rect 295426 229412 295432 229424
rect 290516 229384 295432 229412
rect 290516 229372 290522 229384
rect 295426 229372 295432 229384
rect 295484 229372 295490 229424
rect 372522 229372 372528 229424
rect 372580 229412 372586 229424
rect 374546 229412 374552 229424
rect 372580 229384 374552 229412
rect 372580 229372 372586 229384
rect 374546 229372 374552 229384
rect 374604 229372 374610 229424
rect 402946 229412 402974 229452
rect 405274 229440 405280 229492
rect 405332 229480 405338 229492
rect 428458 229480 428464 229492
rect 405332 229452 428464 229480
rect 405332 229440 405338 229452
rect 428458 229440 428464 229452
rect 428516 229440 428522 229492
rect 428660 229480 428688 229588
rect 428826 229576 428832 229628
rect 428884 229616 428890 229628
rect 441890 229616 441896 229628
rect 428884 229588 441896 229616
rect 428884 229576 428890 229588
rect 441890 229576 441896 229588
rect 441948 229576 441954 229628
rect 444466 229576 444472 229628
rect 444524 229616 444530 229628
rect 495434 229616 495440 229628
rect 444524 229588 495440 229616
rect 444524 229576 444530 229588
rect 495434 229576 495440 229588
rect 495492 229576 495498 229628
rect 429746 229480 429752 229492
rect 428660 229452 429752 229480
rect 429746 229440 429752 229452
rect 429804 229440 429810 229492
rect 434898 229440 434904 229492
rect 434956 229480 434962 229492
rect 439498 229480 439504 229492
rect 434956 229452 439504 229480
rect 434956 229440 434962 229452
rect 439498 229440 439504 229452
rect 439556 229440 439562 229492
rect 441706 229440 441712 229492
rect 441764 229480 441770 229492
rect 450538 229480 450544 229492
rect 441764 229452 450544 229480
rect 441764 229440 441770 229452
rect 450538 229440 450544 229452
rect 450596 229440 450602 229492
rect 450722 229440 450728 229492
rect 450780 229480 450786 229492
rect 495728 229480 495756 229656
rect 499114 229644 499120 229656
rect 499172 229644 499178 229696
rect 499850 229576 499856 229628
rect 499908 229616 499914 229628
rect 499908 229588 502748 229616
rect 499908 229576 499914 229588
rect 450780 229452 495756 229480
rect 450780 229440 450786 229452
rect 495894 229440 495900 229492
rect 495952 229480 495958 229492
rect 499482 229480 499488 229492
rect 495952 229452 499488 229480
rect 495952 229440 495958 229452
rect 499482 229440 499488 229452
rect 499540 229440 499546 229492
rect 499666 229440 499672 229492
rect 499724 229480 499730 229492
rect 502518 229480 502524 229492
rect 499724 229452 502524 229480
rect 499724 229440 499730 229452
rect 502518 229440 502524 229452
rect 502576 229440 502582 229492
rect 502720 229480 502748 229588
rect 502978 229576 502984 229628
rect 503036 229616 503042 229628
rect 511258 229616 511264 229628
rect 503036 229588 511264 229616
rect 503036 229576 503042 229588
rect 511258 229576 511264 229588
rect 511316 229576 511322 229628
rect 504174 229480 504180 229492
rect 502720 229452 504180 229480
rect 504174 229440 504180 229452
rect 504232 229440 504238 229492
rect 504358 229440 504364 229492
rect 504416 229480 504422 229492
rect 507486 229480 507492 229492
rect 504416 229452 507492 229480
rect 504416 229440 504422 229452
rect 507486 229440 507492 229452
rect 507544 229440 507550 229492
rect 404630 229412 404636 229424
rect 402946 229384 404636 229412
rect 404630 229372 404636 229384
rect 404688 229372 404694 229424
rect 396442 229304 396448 229356
rect 396500 229344 396506 229356
rect 397362 229344 397368 229356
rect 396500 229316 397368 229344
rect 396500 229304 396506 229316
rect 397362 229304 397368 229316
rect 397420 229304 397426 229356
rect 412818 229304 412824 229356
rect 412876 229344 412882 229356
rect 421558 229344 421564 229356
rect 412876 229316 421564 229344
rect 412876 229304 412882 229316
rect 421558 229304 421564 229316
rect 421616 229304 421622 229356
rect 421834 229304 421840 229356
rect 421892 229344 421898 229356
rect 451182 229344 451188 229356
rect 421892 229316 451188 229344
rect 421892 229304 421898 229316
rect 451182 229304 451188 229316
rect 451240 229304 451246 229356
rect 453298 229304 453304 229356
rect 453356 229344 453362 229356
rect 455874 229344 455880 229356
rect 453356 229316 455880 229344
rect 453356 229304 453362 229316
rect 455874 229304 455880 229316
rect 455932 229304 455938 229356
rect 456058 229304 456064 229356
rect 456116 229344 456122 229356
rect 458450 229344 458456 229356
rect 456116 229316 458456 229344
rect 456116 229304 456122 229316
rect 458450 229304 458456 229316
rect 458508 229304 458514 229356
rect 458818 229304 458824 229356
rect 458876 229344 458882 229356
rect 480162 229344 480168 229356
rect 458876 229316 480168 229344
rect 458876 229304 458882 229316
rect 480162 229304 480168 229316
rect 480220 229304 480226 229356
rect 480530 229304 480536 229356
rect 480588 229344 480594 229356
rect 481726 229344 481732 229356
rect 480588 229316 481732 229344
rect 480588 229304 480594 229316
rect 481726 229304 481732 229316
rect 481784 229304 481790 229356
rect 484854 229304 484860 229356
rect 484912 229344 484918 229356
rect 489546 229344 489552 229356
rect 484912 229316 489552 229344
rect 484912 229304 484918 229316
rect 489546 229304 489552 229316
rect 489604 229304 489610 229356
rect 490006 229344 490012 229356
rect 489748 229316 490012 229344
rect 334066 229236 334072 229288
rect 334124 229276 334130 229288
rect 335722 229276 335728 229288
rect 334124 229248 335728 229276
rect 334124 229236 334130 229248
rect 335722 229236 335728 229248
rect 335780 229236 335786 229288
rect 350626 229236 350632 229288
rect 350684 229276 350690 229288
rect 355318 229276 355324 229288
rect 350684 229248 355324 229276
rect 350684 229236 350690 229248
rect 355318 229236 355324 229248
rect 355376 229236 355382 229288
rect 390186 229236 390192 229288
rect 390244 229276 390250 229288
rect 393958 229276 393964 229288
rect 390244 229248 393964 229276
rect 390244 229236 390250 229248
rect 393958 229236 393964 229248
rect 394016 229236 394022 229288
rect 399202 229236 399208 229288
rect 399260 229276 399266 229288
rect 404998 229276 405004 229288
rect 399260 229248 405004 229276
rect 399260 229236 399266 229248
rect 404998 229236 405004 229248
rect 405056 229236 405062 229288
rect 222988 229180 238754 229208
rect 222988 229168 222994 229180
rect 422938 229168 422944 229220
rect 422996 229208 423002 229220
rect 429378 229208 429384 229220
rect 422996 229180 429384 229208
rect 422996 229168 423002 229180
rect 429378 229168 429384 229180
rect 429436 229168 429442 229220
rect 429746 229168 429752 229220
rect 429804 229208 429810 229220
rect 446950 229208 446956 229220
rect 429804 229180 446956 229208
rect 429804 229168 429810 229180
rect 446950 229168 446956 229180
rect 447008 229168 447014 229220
rect 448330 229168 448336 229220
rect 448388 229208 448394 229220
rect 463694 229208 463700 229220
rect 448388 229180 463700 229208
rect 448388 229168 448394 229180
rect 463694 229168 463700 229180
rect 463752 229168 463758 229220
rect 464154 229168 464160 229220
rect 464212 229208 464218 229220
rect 466362 229208 466368 229220
rect 464212 229180 466368 229208
rect 464212 229168 464218 229180
rect 466362 229168 466368 229180
rect 466420 229168 466426 229220
rect 466546 229168 466552 229220
rect 466604 229208 466610 229220
rect 470778 229208 470784 229220
rect 466604 229180 470784 229208
rect 466604 229168 466610 229180
rect 470778 229168 470784 229180
rect 470836 229168 470842 229220
rect 473446 229168 473452 229220
rect 473504 229208 473510 229220
rect 476390 229208 476396 229220
rect 473504 229180 476396 229208
rect 473504 229168 473510 229180
rect 476390 229168 476396 229180
rect 476448 229168 476454 229220
rect 479242 229168 479248 229220
rect 479300 229208 479306 229220
rect 485038 229208 485044 229220
rect 479300 229180 485044 229208
rect 479300 229168 479306 229180
rect 485038 229168 485044 229180
rect 485096 229168 485102 229220
rect 485866 229168 485872 229220
rect 485924 229208 485930 229220
rect 489748 229208 489776 229316
rect 490006 229304 490012 229316
rect 490064 229304 490070 229356
rect 490190 229304 490196 229356
rect 490248 229344 490254 229356
rect 536834 229344 536840 229356
rect 490248 229316 536840 229344
rect 490248 229304 490254 229316
rect 536834 229304 536840 229316
rect 536892 229304 536898 229356
rect 485924 229180 489776 229208
rect 485924 229168 485930 229180
rect 489914 229168 489920 229220
rect 489972 229208 489978 229220
rect 533338 229208 533344 229220
rect 489972 229180 533344 229208
rect 489972 229168 489978 229180
rect 533338 229168 533344 229180
rect 533396 229168 533402 229220
rect 304074 229100 304080 229152
rect 304132 229140 304138 229152
rect 308674 229140 308680 229152
rect 304132 229112 308680 229140
rect 304132 229100 304138 229112
rect 308674 229100 308680 229112
rect 308732 229100 308738 229152
rect 322750 229100 322756 229152
rect 322808 229140 322814 229152
rect 326338 229140 326344 229152
rect 322808 229112 326344 229140
rect 322808 229100 322814 229112
rect 326338 229100 326344 229112
rect 326396 229100 326402 229152
rect 335170 229100 335176 229152
rect 335228 229140 335234 229152
rect 335906 229140 335912 229152
rect 335228 229112 335912 229140
rect 335228 229100 335234 229112
rect 335906 229100 335912 229112
rect 335964 229100 335970 229152
rect 87598 229032 87604 229084
rect 87656 229072 87662 229084
rect 147490 229072 147496 229084
rect 87656 229044 147496 229072
rect 87656 229032 87662 229044
rect 147490 229032 147496 229044
rect 147548 229032 147554 229084
rect 147628 229032 147634 229084
rect 147686 229072 147692 229084
rect 152458 229072 152464 229084
rect 147686 229044 152464 229072
rect 147686 229032 147692 229044
rect 152458 229032 152464 229044
rect 152516 229032 152522 229084
rect 152918 229032 152924 229084
rect 152976 229072 152982 229084
rect 185854 229072 185860 229084
rect 152976 229044 185860 229072
rect 152976 229032 152982 229044
rect 185854 229032 185860 229044
rect 185912 229032 185918 229084
rect 188982 229032 188988 229084
rect 189040 229072 189046 229084
rect 195238 229072 195244 229084
rect 189040 229044 195244 229072
rect 189040 229032 189046 229044
rect 195238 229032 195244 229044
rect 195296 229032 195302 229084
rect 195698 229032 195704 229084
rect 195756 229072 195762 229084
rect 195756 229044 197032 229072
rect 195756 229032 195762 229044
rect 119982 228896 119988 228948
rect 120040 228936 120046 228948
rect 189718 228936 189724 228948
rect 120040 228908 189724 228936
rect 120040 228896 120046 228908
rect 189718 228896 189724 228908
rect 189776 228896 189782 228948
rect 194226 228896 194232 228948
rect 194284 228936 194290 228948
rect 196802 228936 196808 228948
rect 194284 228908 196808 228936
rect 194284 228896 194290 228908
rect 196802 228896 196808 228908
rect 196860 228896 196866 228948
rect 197004 228936 197032 229044
rect 198642 229032 198648 229084
rect 198700 229072 198706 229084
rect 201218 229072 201224 229084
rect 198700 229044 201224 229072
rect 198700 229032 198706 229044
rect 201218 229032 201224 229044
rect 201276 229032 201282 229084
rect 212258 229032 212264 229084
rect 212316 229072 212322 229084
rect 251818 229072 251824 229084
rect 212316 229044 251824 229072
rect 212316 229032 212322 229044
rect 251818 229032 251824 229044
rect 251876 229032 251882 229084
rect 262030 229032 262036 229084
rect 262088 229072 262094 229084
rect 284938 229072 284944 229084
rect 262088 229044 284944 229072
rect 262088 229032 262094 229044
rect 284938 229032 284944 229044
rect 284996 229032 285002 229084
rect 361114 229032 361120 229084
rect 361172 229072 361178 229084
rect 373534 229072 373540 229084
rect 361172 229044 373540 229072
rect 361172 229032 361178 229044
rect 373534 229032 373540 229044
rect 373592 229032 373598 229084
rect 382274 229032 382280 229084
rect 382332 229072 382338 229084
rect 382332 229044 388668 229072
rect 382332 229032 382338 229044
rect 202414 228936 202420 228948
rect 197004 228908 202420 228936
rect 202414 228896 202420 228908
rect 202472 228896 202478 228948
rect 202598 228896 202604 228948
rect 202656 228936 202662 228948
rect 245194 228936 245200 228948
rect 202656 228908 245200 228936
rect 202656 228896 202662 228908
rect 245194 228896 245200 228908
rect 245252 228896 245258 228948
rect 245470 228896 245476 228948
rect 245528 228936 245534 228948
rect 273898 228936 273904 228948
rect 245528 228908 273904 228936
rect 245528 228896 245534 228908
rect 273898 228896 273904 228908
rect 273956 228896 273962 228948
rect 286686 228896 286692 228948
rect 286744 228936 286750 228948
rect 300946 228936 300952 228948
rect 286744 228908 300952 228936
rect 286744 228896 286750 228908
rect 300946 228896 300952 228908
rect 301004 228896 301010 228948
rect 373258 228896 373264 228948
rect 373316 228936 373322 228948
rect 388438 228936 388444 228948
rect 373316 228908 388444 228936
rect 373316 228896 373322 228908
rect 388438 228896 388444 228908
rect 388496 228896 388502 228948
rect 388640 228936 388668 229044
rect 391198 229032 391204 229084
rect 391256 229072 391262 229084
rect 397730 229072 397736 229084
rect 391256 229044 397736 229072
rect 391256 229032 391262 229044
rect 397730 229032 397736 229044
rect 397788 229032 397794 229084
rect 407758 229032 407764 229084
rect 407816 229072 407822 229084
rect 429930 229072 429936 229084
rect 407816 229044 429936 229072
rect 407816 229032 407822 229044
rect 429930 229032 429936 229044
rect 429988 229032 429994 229084
rect 430114 229032 430120 229084
rect 430172 229072 430178 229084
rect 457438 229072 457444 229084
rect 430172 229044 457444 229072
rect 430172 229032 430178 229044
rect 457438 229032 457444 229044
rect 457496 229032 457502 229084
rect 459922 229032 459928 229084
rect 459980 229072 459986 229084
rect 525978 229072 525984 229084
rect 459980 229044 525984 229072
rect 459980 229032 459986 229044
rect 525978 229032 525984 229044
rect 526036 229032 526042 229084
rect 391842 228936 391848 228948
rect 388640 228908 391848 228936
rect 391842 228896 391848 228908
rect 391900 228896 391906 228948
rect 400674 228936 400680 228948
rect 393286 228908 400680 228936
rect 110322 228760 110328 228812
rect 110380 228800 110386 228812
rect 183094 228800 183100 228812
rect 110380 228772 183100 228800
rect 110380 228760 110386 228772
rect 183094 228760 183100 228772
rect 183152 228760 183158 228812
rect 183278 228760 183284 228812
rect 183336 228800 183342 228812
rect 225966 228800 225972 228812
rect 183336 228772 225972 228800
rect 183336 228760 183342 228772
rect 225966 228760 225972 228772
rect 226024 228760 226030 228812
rect 238570 228760 238576 228812
rect 238628 228800 238634 228812
rect 269482 228800 269488 228812
rect 238628 228772 269488 228800
rect 238628 228760 238634 228772
rect 269482 228760 269488 228772
rect 269540 228760 269546 228812
rect 275830 228760 275836 228812
rect 275888 228800 275894 228812
rect 293770 228800 293776 228812
rect 275888 228772 293776 228800
rect 275888 228760 275894 228772
rect 293770 228760 293776 228772
rect 293828 228760 293834 228812
rect 295150 228760 295156 228812
rect 295208 228800 295214 228812
rect 307018 228800 307024 228812
rect 295208 228772 307024 228800
rect 295208 228760 295214 228772
rect 307018 228760 307024 228772
rect 307076 228760 307082 228812
rect 352834 228760 352840 228812
rect 352892 228800 352898 228812
rect 361022 228800 361028 228812
rect 352892 228772 361028 228800
rect 352892 228760 352898 228772
rect 361022 228760 361028 228772
rect 361080 228760 361086 228812
rect 362218 228760 362224 228812
rect 362276 228800 362282 228812
rect 376754 228800 376760 228812
rect 362276 228772 376760 228800
rect 362276 228760 362282 228772
rect 376754 228760 376760 228772
rect 376812 228760 376818 228812
rect 377674 228760 377680 228812
rect 377732 228800 377738 228812
rect 393286 228800 393314 228908
rect 400674 228896 400680 228908
rect 400732 228896 400738 228948
rect 401962 228896 401968 228948
rect 402020 228936 402026 228948
rect 437106 228936 437112 228948
rect 402020 228908 437112 228936
rect 402020 228896 402026 228908
rect 437106 228896 437112 228908
rect 437164 228896 437170 228948
rect 439498 228896 439504 228948
rect 439556 228936 439562 228948
rect 465258 228936 465264 228948
rect 439556 228908 465264 228936
rect 439556 228896 439562 228908
rect 465258 228896 465264 228908
rect 465316 228896 465322 228948
rect 477586 228896 477592 228948
rect 477644 228936 477650 228948
rect 495388 228936 495394 228948
rect 477644 228908 495394 228936
rect 477644 228896 477650 228908
rect 495388 228896 495394 228908
rect 495446 228896 495452 228948
rect 495986 228896 495992 228948
rect 496044 228936 496050 228948
rect 507946 228936 507952 228948
rect 496044 228908 507952 228936
rect 496044 228896 496050 228908
rect 507946 228896 507952 228908
rect 508004 228896 508010 228948
rect 508130 228896 508136 228948
rect 508188 228936 508194 228948
rect 552198 228936 552204 228948
rect 508188 228908 552204 228936
rect 508188 228896 508194 228908
rect 552198 228896 552204 228908
rect 552256 228896 552262 228948
rect 495544 228840 495756 228868
rect 377732 228772 393314 228800
rect 377732 228760 377738 228772
rect 397546 228760 397552 228812
rect 397604 228800 397610 228812
rect 407758 228800 407764 228812
rect 397604 228772 407764 228800
rect 397604 228760 397610 228772
rect 407758 228760 407764 228772
rect 407816 228760 407822 228812
rect 423490 228760 423496 228812
rect 423548 228800 423554 228812
rect 468018 228800 468024 228812
rect 423548 228772 468024 228800
rect 423548 228760 423554 228772
rect 468018 228760 468024 228772
rect 468076 228760 468082 228812
rect 468202 228760 468208 228812
rect 468260 228800 468266 228812
rect 495544 228800 495572 228840
rect 468260 228772 495572 228800
rect 495728 228800 495756 228840
rect 538398 228800 538404 228812
rect 495728 228772 538404 228800
rect 468260 228760 468266 228772
rect 538398 228760 538404 228772
rect 538456 228760 538462 228812
rect 85482 228624 85488 228676
rect 85540 228664 85546 228676
rect 85540 228636 167132 228664
rect 85540 228624 85546 228636
rect 100662 228488 100668 228540
rect 100720 228528 100726 228540
rect 166902 228528 166908 228540
rect 100720 228500 166908 228528
rect 100720 228488 100726 228500
rect 166902 228488 166908 228500
rect 166960 228488 166966 228540
rect 167104 228528 167132 228636
rect 167822 228624 167828 228676
rect 167880 228664 167886 228676
rect 171962 228664 171968 228676
rect 167880 228636 171968 228664
rect 167880 228624 167886 228636
rect 171962 228624 171968 228636
rect 172020 228624 172026 228676
rect 172422 228624 172428 228676
rect 172480 228664 172486 228676
rect 213822 228664 213828 228676
rect 172480 228636 213828 228664
rect 172480 228624 172486 228636
rect 213822 228624 213828 228636
rect 213880 228624 213886 228676
rect 226978 228664 226984 228676
rect 214576 228636 226984 228664
rect 169018 228528 169024 228540
rect 167104 228500 169024 228528
rect 169018 228488 169024 228500
rect 169076 228488 169082 228540
rect 171594 228488 171600 228540
rect 171652 228528 171658 228540
rect 193030 228528 193036 228540
rect 171652 228500 193036 228528
rect 171652 228488 171658 228500
rect 193030 228488 193036 228500
rect 193088 228488 193094 228540
rect 195238 228488 195244 228540
rect 195296 228528 195302 228540
rect 214576 228528 214604 228636
rect 226978 228624 226984 228636
rect 227036 228624 227042 228676
rect 231670 228624 231676 228676
rect 231728 228664 231734 228676
rect 266170 228664 266176 228676
rect 231728 228636 266176 228664
rect 231728 228624 231734 228636
rect 266170 228624 266176 228636
rect 266228 228624 266234 228676
rect 266354 228624 266360 228676
rect 266412 228664 266418 228676
rect 287146 228664 287152 228676
rect 266412 228636 287152 228664
rect 266412 228624 266418 228636
rect 287146 228624 287152 228636
rect 287204 228624 287210 228676
rect 292482 228624 292488 228676
rect 292540 228664 292546 228676
rect 304810 228664 304816 228676
rect 292540 228636 304816 228664
rect 292540 228624 292546 228636
rect 304810 228624 304816 228636
rect 304868 228624 304874 228676
rect 315666 228624 315672 228676
rect 315724 228664 315730 228676
rect 320266 228664 320272 228676
rect 315724 228636 320272 228664
rect 315724 228624 315730 228636
rect 320266 228624 320272 228636
rect 320324 228624 320330 228676
rect 349522 228624 349528 228676
rect 349580 228664 349586 228676
rect 359458 228664 359464 228676
rect 349580 228636 359464 228664
rect 349580 228624 349586 228636
rect 359458 228624 359464 228636
rect 359516 228624 359522 228676
rect 370498 228624 370504 228676
rect 370556 228664 370562 228676
rect 387058 228664 387064 228676
rect 370556 228636 387064 228664
rect 370556 228624 370562 228636
rect 387058 228624 387064 228636
rect 387116 228624 387122 228676
rect 393130 228624 393136 228676
rect 393188 228664 393194 228676
rect 424042 228664 424048 228676
rect 393188 228636 424048 228664
rect 393188 228624 393194 228636
rect 424042 228624 424048 228636
rect 424100 228624 424106 228676
rect 426802 228624 426808 228676
rect 426860 228664 426866 228676
rect 475194 228664 475200 228676
rect 426860 228636 475200 228664
rect 426860 228624 426866 228636
rect 475194 228624 475200 228636
rect 475252 228624 475258 228676
rect 475378 228624 475384 228676
rect 475436 228664 475442 228676
rect 495618 228664 495624 228676
rect 475436 228636 495624 228664
rect 475436 228624 475442 228636
rect 495618 228624 495624 228636
rect 495676 228624 495682 228676
rect 495802 228624 495808 228676
rect 495860 228664 495866 228676
rect 495860 228636 507716 228664
rect 495860 228624 495866 228636
rect 195296 228500 214604 228528
rect 195296 228488 195302 228500
rect 214742 228488 214748 228540
rect 214800 228528 214806 228540
rect 248506 228528 248512 228540
rect 214800 228500 248512 228528
rect 214800 228488 214806 228500
rect 248506 228488 248512 228500
rect 248564 228488 248570 228540
rect 253566 228488 253572 228540
rect 253624 228528 253630 228540
rect 278866 228528 278872 228540
rect 253624 228500 278872 228528
rect 253624 228488 253630 228500
rect 278866 228488 278872 228500
rect 278924 228488 278930 228540
rect 285582 228488 285588 228540
rect 285640 228528 285646 228540
rect 300394 228528 300400 228540
rect 285640 228500 300400 228528
rect 285640 228488 285646 228500
rect 300394 228488 300400 228500
rect 300452 228488 300458 228540
rect 300762 228488 300768 228540
rect 300820 228528 300826 228540
rect 309778 228528 309784 228540
rect 300820 228500 309784 228528
rect 300820 228488 300826 228500
rect 309778 228488 309784 228500
rect 309836 228488 309842 228540
rect 325602 228488 325608 228540
rect 325660 228528 325666 228540
rect 328362 228528 328368 228540
rect 325660 228500 328368 228528
rect 325660 228488 325666 228500
rect 328362 228488 328368 228500
rect 328420 228488 328426 228540
rect 353386 228488 353392 228540
rect 353444 228528 353450 228540
rect 364426 228528 364432 228540
rect 353444 228500 364432 228528
rect 353444 228488 353450 228500
rect 364426 228488 364432 228500
rect 364484 228488 364490 228540
rect 364978 228488 364984 228540
rect 365036 228528 365042 228540
rect 376386 228528 376392 228540
rect 365036 228500 376392 228528
rect 365036 228488 365042 228500
rect 376386 228488 376392 228500
rect 376444 228488 376450 228540
rect 376754 228488 376760 228540
rect 376812 228528 376818 228540
rect 377674 228528 377680 228540
rect 376812 228500 377680 228528
rect 376812 228488 376818 228500
rect 377674 228488 377680 228500
rect 377732 228488 377738 228540
rect 386506 228488 386512 228540
rect 386564 228528 386570 228540
rect 414198 228528 414204 228540
rect 386564 228500 414204 228528
rect 386564 228488 386570 228500
rect 414198 228488 414204 228500
rect 414256 228488 414262 228540
rect 414842 228488 414848 228540
rect 414900 228528 414906 228540
rect 451458 228528 451464 228540
rect 414900 228500 451464 228528
rect 414900 228488 414906 228500
rect 451458 228488 451464 228500
rect 451516 228488 451522 228540
rect 451642 228488 451648 228540
rect 451700 228528 451706 228540
rect 505048 228528 505054 228540
rect 451700 228500 505054 228528
rect 451700 228488 451706 228500
rect 505048 228488 505054 228500
rect 505106 228488 505112 228540
rect 505186 228488 505192 228540
rect 505244 228528 505250 228540
rect 507486 228528 507492 228540
rect 505244 228500 507492 228528
rect 505244 228488 505250 228500
rect 507486 228488 507492 228500
rect 507544 228488 507550 228540
rect 507688 228528 507716 228636
rect 507946 228624 507952 228676
rect 508004 228664 508010 228676
rect 548334 228664 548340 228676
rect 508004 228636 548340 228664
rect 508004 228624 508010 228636
rect 548334 228624 548340 228636
rect 548392 228624 548398 228676
rect 548518 228528 548524 228540
rect 507688 228500 548524 228528
rect 548518 228488 548524 228500
rect 548576 228488 548582 228540
rect 49142 228352 49148 228404
rect 49200 228392 49206 228404
rect 653214 228392 653220 228404
rect 49200 228364 653220 228392
rect 49200 228352 49206 228364
rect 653214 228352 653220 228364
rect 653272 228352 653278 228404
rect 96430 228216 96436 228268
rect 96488 228256 96494 228268
rect 96488 228228 151584 228256
rect 96488 228216 96494 228228
rect 69566 228080 69572 228132
rect 69624 228120 69630 228132
rect 147950 228120 147956 228132
rect 69624 228092 147956 228120
rect 69624 228080 69630 228092
rect 147950 228080 147956 228092
rect 148008 228080 148014 228132
rect 149238 228080 149244 228132
rect 149296 228120 149302 228132
rect 151354 228120 151360 228132
rect 149296 228092 151360 228120
rect 149296 228080 149302 228092
rect 151354 228080 151360 228092
rect 151412 228080 151418 228132
rect 151556 228120 151584 228228
rect 152458 228216 152464 228268
rect 152516 228256 152522 228268
rect 171594 228256 171600 228268
rect 152516 228228 171600 228256
rect 152516 228216 152522 228228
rect 171594 228216 171600 228228
rect 171652 228216 171658 228268
rect 208394 228256 208400 228268
rect 171796 228228 208400 228256
rect 159818 228120 159824 228132
rect 151556 228092 159824 228120
rect 159818 228080 159824 228092
rect 159876 228080 159882 228132
rect 160002 228080 160008 228132
rect 160060 228120 160066 228132
rect 171796 228120 171824 228228
rect 208394 228216 208400 228228
rect 208452 228216 208458 228268
rect 213822 228216 213828 228268
rect 213880 228256 213886 228268
rect 220814 228256 220820 228268
rect 213880 228228 220820 228256
rect 213880 228216 213886 228228
rect 220814 228216 220820 228228
rect 220872 228216 220878 228268
rect 222010 228216 222016 228268
rect 222068 228256 222074 228268
rect 258442 228256 258448 228268
rect 222068 228228 258448 228256
rect 222068 228216 222074 228228
rect 258442 228216 258448 228228
rect 258500 228216 258506 228268
rect 376386 228216 376392 228268
rect 376444 228256 376450 228268
rect 382642 228256 382648 228268
rect 376444 228228 382648 228256
rect 376444 228216 376450 228228
rect 382642 228216 382648 228228
rect 382700 228216 382706 228268
rect 388438 228216 388444 228268
rect 388496 228256 388502 228268
rect 394234 228256 394240 228268
rect 388496 228228 394240 228256
rect 388496 228216 388502 228228
rect 394234 228216 394240 228228
rect 394292 228216 394298 228268
rect 400306 228216 400312 228268
rect 400364 228256 400370 228268
rect 432598 228256 432604 228268
rect 400364 228228 432604 228256
rect 400364 228216 400370 228228
rect 432598 228216 432604 228228
rect 432656 228216 432662 228268
rect 434530 228216 434536 228268
rect 434588 228256 434594 228268
rect 442442 228256 442448 228268
rect 434588 228228 442448 228256
rect 434588 228216 434594 228228
rect 442442 228216 442448 228228
rect 442500 228216 442506 228268
rect 446766 228216 446772 228268
rect 446824 228256 446830 228268
rect 466178 228256 466184 228268
rect 446824 228228 466184 228256
rect 446824 228216 446830 228228
rect 466178 228216 466184 228228
rect 466236 228216 466242 228268
rect 466362 228216 466368 228268
rect 466420 228256 466426 228268
rect 531682 228256 531688 228268
rect 466420 228228 531688 228256
rect 466420 228216 466426 228228
rect 531682 228216 531688 228228
rect 531740 228216 531746 228268
rect 160060 228092 171824 228120
rect 160060 228080 160066 228092
rect 171962 228080 171968 228132
rect 172020 228120 172026 228132
rect 211154 228120 211160 228132
rect 172020 228092 211160 228120
rect 172020 228080 172026 228092
rect 211154 228080 211160 228092
rect 211212 228080 211218 228132
rect 456518 228080 456524 228132
rect 456576 228120 456582 228132
rect 520918 228120 520924 228132
rect 456576 228092 520924 228120
rect 456576 228080 456582 228092
rect 520918 228080 520924 228092
rect 520976 228080 520982 228132
rect 133506 227944 133512 227996
rect 133564 227984 133570 227996
rect 147490 227984 147496 227996
rect 133564 227956 147496 227984
rect 133564 227944 133570 227956
rect 147490 227944 147496 227956
rect 147548 227944 147554 227996
rect 147674 227944 147680 227996
rect 147732 227984 147738 227996
rect 204162 227984 204168 227996
rect 147732 227956 204168 227984
rect 147732 227944 147738 227956
rect 204162 227944 204168 227956
rect 204220 227944 204226 227996
rect 205266 227944 205272 227996
rect 205324 227984 205330 227996
rect 214742 227984 214748 227996
rect 205324 227956 214748 227984
rect 205324 227944 205330 227956
rect 214742 227944 214748 227956
rect 214800 227944 214806 227996
rect 454954 227944 454960 227996
rect 455012 227984 455018 227996
rect 517790 227984 517796 227996
rect 455012 227956 517796 227984
rect 455012 227944 455018 227956
rect 517790 227944 517796 227956
rect 517848 227944 517854 227996
rect 310330 227876 310336 227928
rect 310388 227916 310394 227928
rect 316402 227916 316408 227928
rect 310388 227888 316408 227916
rect 310388 227876 310394 227888
rect 316402 227876 316408 227888
rect 316460 227876 316466 227928
rect 136542 227808 136548 227860
rect 136600 227848 136606 227860
rect 196526 227848 196532 227860
rect 136600 227820 196532 227848
rect 136600 227808 136606 227820
rect 196526 227808 196532 227820
rect 196584 227808 196590 227860
rect 201034 227808 201040 227860
rect 201092 227848 201098 227860
rect 222562 227848 222568 227860
rect 201092 227820 222568 227848
rect 201092 227808 201098 227820
rect 222562 227808 222568 227820
rect 222620 227808 222626 227860
rect 226242 227808 226248 227860
rect 226300 227848 226306 227860
rect 230658 227848 230664 227860
rect 226300 227820 230664 227848
rect 226300 227808 226306 227820
rect 230658 227808 230664 227820
rect 230716 227808 230722 227860
rect 236638 227808 236644 227860
rect 236696 227848 236702 227860
rect 238018 227848 238024 227860
rect 236696 227820 238024 227848
rect 236696 227808 236702 227820
rect 238018 227808 238024 227820
rect 238076 227808 238082 227860
rect 240042 227808 240048 227860
rect 240100 227848 240106 227860
rect 241606 227848 241612 227860
rect 240100 227820 241612 227848
rect 240100 227808 240106 227820
rect 241606 227808 241612 227820
rect 241664 227808 241670 227860
rect 259270 227808 259276 227860
rect 259328 227848 259334 227860
rect 261570 227848 261576 227860
rect 259328 227820 261576 227848
rect 259328 227808 259334 227820
rect 261570 227808 261576 227820
rect 261628 227808 261634 227860
rect 436738 227808 436744 227860
rect 436796 227848 436802 227860
rect 436796 227820 481220 227848
rect 436796 227808 436802 227820
rect 249058 227740 249064 227792
rect 249116 227780 249122 227792
rect 251266 227780 251272 227792
rect 249116 227752 251272 227780
rect 249116 227740 249122 227752
rect 251266 227740 251272 227752
rect 251324 227740 251330 227792
rect 251726 227740 251732 227792
rect 251784 227780 251790 227792
rect 255682 227780 255688 227792
rect 251784 227752 255688 227780
rect 251784 227740 251790 227752
rect 255682 227740 255688 227752
rect 255740 227740 255746 227792
rect 308766 227740 308772 227792
rect 308824 227780 308830 227792
rect 315482 227780 315488 227792
rect 308824 227752 315488 227780
rect 308824 227740 308830 227752
rect 315482 227740 315488 227752
rect 315540 227740 315546 227792
rect 317046 227740 317052 227792
rect 317104 227780 317110 227792
rect 320542 227780 320548 227792
rect 317104 227752 320548 227780
rect 317104 227740 317110 227752
rect 320542 227740 320548 227752
rect 320600 227740 320606 227792
rect 321462 227740 321468 227792
rect 321520 227780 321526 227792
rect 324682 227780 324688 227792
rect 321520 227752 324688 227780
rect 321520 227740 321526 227752
rect 324682 227740 324688 227752
rect 324740 227740 324746 227792
rect 345106 227740 345112 227792
rect 345164 227780 345170 227792
rect 352834 227780 352840 227792
rect 345164 227752 352840 227780
rect 345164 227740 345170 227752
rect 352834 227740 352840 227752
rect 352892 227740 352898 227792
rect 394786 227740 394792 227792
rect 394844 227780 394850 227792
rect 402238 227780 402244 227792
rect 394844 227752 402244 227780
rect 394844 227740 394850 227752
rect 402238 227740 402244 227752
rect 402296 227740 402302 227792
rect 111702 227672 111708 227724
rect 111760 227712 111766 227724
rect 183922 227712 183928 227724
rect 111760 227684 183928 227712
rect 111760 227672 111766 227684
rect 183922 227672 183928 227684
rect 183980 227672 183986 227724
rect 196618 227672 196624 227724
rect 196676 227712 196682 227724
rect 207106 227712 207112 227724
rect 196676 227684 207112 227712
rect 196676 227672 196682 227684
rect 207106 227672 207112 227684
rect 207164 227672 207170 227724
rect 209590 227672 209596 227724
rect 209648 227712 209654 227724
rect 276658 227712 276664 227724
rect 209648 227684 248414 227712
rect 209648 227672 209654 227684
rect 248386 227644 248414 227684
rect 255884 227684 276664 227712
rect 249610 227644 249616 227656
rect 248386 227616 249616 227644
rect 249610 227604 249616 227616
rect 249668 227604 249674 227656
rect 251082 227604 251088 227656
rect 251140 227644 251146 227656
rect 255884 227644 255912 227684
rect 276658 227672 276664 227684
rect 276716 227672 276722 227724
rect 429562 227672 429568 227724
rect 429620 227712 429626 227724
rect 476206 227712 476212 227724
rect 429620 227684 476212 227712
rect 429620 227672 429626 227684
rect 476206 227672 476212 227684
rect 476264 227672 476270 227724
rect 481192 227712 481220 227820
rect 481358 227808 481364 227860
rect 481416 227848 481422 227860
rect 489868 227848 489874 227860
rect 481416 227820 489874 227848
rect 481416 227808 481422 227820
rect 489868 227808 489874 227820
rect 489926 227808 489932 227860
rect 630674 227780 630680 227792
rect 490024 227752 504956 227780
rect 487614 227712 487620 227724
rect 481192 227684 487620 227712
rect 487614 227672 487620 227684
rect 487672 227672 487678 227724
rect 489546 227672 489552 227724
rect 489604 227712 489610 227724
rect 490024 227712 490052 227752
rect 489604 227684 490052 227712
rect 504928 227712 504956 227752
rect 505066 227752 630680 227780
rect 505066 227712 505094 227752
rect 630674 227740 630680 227752
rect 630732 227740 630738 227792
rect 504928 227684 505094 227712
rect 489604 227672 489610 227684
rect 251140 227616 255912 227644
rect 251140 227604 251146 227616
rect 93762 227536 93768 227588
rect 93820 227576 93826 227588
rect 173986 227576 173992 227588
rect 93820 227548 173992 227576
rect 93820 227536 93826 227548
rect 173986 227536 173992 227548
rect 174044 227536 174050 227588
rect 184198 227536 184204 227588
rect 184256 227576 184262 227588
rect 198274 227576 198280 227588
rect 184256 227548 198280 227576
rect 184256 227536 184262 227548
rect 198274 227536 198280 227548
rect 198332 227536 198338 227588
rect 199470 227536 199476 227588
rect 199528 227576 199534 227588
rect 205542 227576 205548 227588
rect 199528 227548 205548 227576
rect 199528 227536 199534 227548
rect 205542 227536 205548 227548
rect 205600 227536 205606 227588
rect 205910 227536 205916 227588
rect 205968 227576 205974 227588
rect 247402 227576 247408 227588
rect 205968 227548 247408 227576
rect 205968 227536 205974 227548
rect 247402 227536 247408 227548
rect 247460 227536 247466 227588
rect 256510 227536 256516 227588
rect 256568 227576 256574 227588
rect 276106 227576 276112 227588
rect 256568 227548 276112 227576
rect 256568 227536 256574 227548
rect 276106 227536 276112 227548
rect 276164 227536 276170 227588
rect 395338 227536 395344 227588
rect 395396 227576 395402 227588
rect 427354 227576 427360 227588
rect 395396 227548 427360 227576
rect 395396 227536 395402 227548
rect 427354 227536 427360 227548
rect 427412 227536 427418 227588
rect 461578 227536 461584 227588
rect 461636 227576 461642 227588
rect 527818 227576 527824 227588
rect 461636 227548 527824 227576
rect 461636 227536 461642 227548
rect 527818 227536 527824 227548
rect 527876 227536 527882 227588
rect 68922 227400 68928 227452
rect 68980 227440 68986 227452
rect 154574 227440 154580 227452
rect 68980 227412 154580 227440
rect 68980 227400 68986 227412
rect 154574 227400 154580 227412
rect 154632 227400 154638 227452
rect 155678 227400 155684 227452
rect 155736 227440 155742 227452
rect 155736 227412 162164 227440
rect 155736 227400 155742 227412
rect 73706 227264 73712 227316
rect 73764 227304 73770 227316
rect 160186 227304 160192 227316
rect 73764 227276 160192 227304
rect 73764 227264 73770 227276
rect 160186 227264 160192 227276
rect 160244 227264 160250 227316
rect 162136 227304 162164 227412
rect 166718 227400 166724 227452
rect 166776 227440 166782 227452
rect 167822 227440 167828 227452
rect 166776 227412 167828 227440
rect 166776 227400 166782 227412
rect 167822 227400 167828 227412
rect 167880 227400 167886 227452
rect 176562 227400 176568 227452
rect 176620 227440 176626 227452
rect 176620 227400 176654 227440
rect 182818 227400 182824 227452
rect 182876 227440 182882 227452
rect 233050 227440 233056 227452
rect 182876 227412 233056 227440
rect 182876 227400 182882 227412
rect 233050 227400 233056 227412
rect 233108 227400 233114 227452
rect 234430 227400 234436 227452
rect 234488 227440 234494 227452
rect 268286 227440 268292 227452
rect 234488 227412 268292 227440
rect 234488 227400 234494 227412
rect 268286 227400 268292 227412
rect 268344 227400 268350 227452
rect 374546 227400 374552 227452
rect 374604 227440 374610 227452
rect 390094 227440 390100 227452
rect 374604 227412 390100 227440
rect 374604 227400 374610 227412
rect 390094 227400 390100 227412
rect 390152 227400 390158 227452
rect 392210 227400 392216 227452
rect 392268 227440 392274 227452
rect 401686 227440 401692 227452
rect 392268 227412 401692 227440
rect 392268 227400 392274 227412
rect 401686 227400 401692 227412
rect 401744 227400 401750 227452
rect 404078 227400 404084 227452
rect 404136 227440 404142 227452
rect 440602 227440 440608 227452
rect 404136 227412 440608 227440
rect 404136 227400 404142 227412
rect 440602 227400 440608 227412
rect 440660 227400 440666 227452
rect 446950 227400 446956 227452
rect 447008 227440 447014 227452
rect 471238 227440 471244 227452
rect 447008 227412 471244 227440
rect 447008 227400 447014 227412
rect 471238 227400 471244 227412
rect 471296 227400 471302 227452
rect 473722 227400 473728 227452
rect 473780 227440 473786 227452
rect 546586 227440 546592 227452
rect 473780 227412 546592 227440
rect 473780 227400 473786 227412
rect 546586 227400 546592 227412
rect 546644 227400 546650 227452
rect 176626 227304 176654 227400
rect 227530 227304 227536 227316
rect 162136 227276 166994 227304
rect 176626 227276 227536 227304
rect 66162 227128 66168 227180
rect 66220 227168 66226 227180
rect 149514 227168 149520 227180
rect 66220 227140 149520 227168
rect 66220 227128 66226 227140
rect 149514 227128 149520 227140
rect 149572 227128 149578 227180
rect 151722 227168 151728 227180
rect 149716 227140 151728 227168
rect 63402 226992 63408 227044
rect 63460 227032 63466 227044
rect 149716 227032 149744 227140
rect 151722 227128 151728 227140
rect 151780 227128 151786 227180
rect 156690 227128 156696 227180
rect 156748 227168 156754 227180
rect 163958 227168 163964 227180
rect 156748 227140 163964 227168
rect 156748 227128 156754 227140
rect 163958 227128 163964 227140
rect 164016 227128 164022 227180
rect 166966 227168 166994 227276
rect 227530 227264 227536 227276
rect 227588 227264 227594 227316
rect 228818 227264 228824 227316
rect 228876 227304 228882 227316
rect 262858 227304 262864 227316
rect 228876 227276 262864 227304
rect 228876 227264 228882 227276
rect 262858 227264 262864 227276
rect 262916 227264 262922 227316
rect 272426 227264 272432 227316
rect 272484 227304 272490 227316
rect 282178 227304 282184 227316
rect 272484 227276 282184 227304
rect 272484 227264 272490 227276
rect 282178 227264 282184 227276
rect 282236 227264 282242 227316
rect 293770 227264 293776 227316
rect 293828 227304 293834 227316
rect 305362 227304 305368 227316
rect 293828 227276 305368 227304
rect 293828 227264 293834 227276
rect 305362 227264 305368 227276
rect 305420 227264 305426 227316
rect 376570 227264 376576 227316
rect 376628 227304 376634 227316
rect 396718 227304 396724 227316
rect 376628 227276 396724 227304
rect 376628 227264 376634 227276
rect 396718 227264 396724 227276
rect 396776 227264 396782 227316
rect 417970 227264 417976 227316
rect 418028 227304 418034 227316
rect 462130 227304 462136 227316
rect 418028 227276 462136 227304
rect 418028 227264 418034 227276
rect 462130 227264 462136 227276
rect 462188 227264 462194 227316
rect 471514 227264 471520 227316
rect 471572 227304 471578 227316
rect 543458 227304 543464 227316
rect 471572 227276 543464 227304
rect 471572 227264 471578 227276
rect 543458 227264 543464 227276
rect 543516 227264 543522 227316
rect 214282 227168 214288 227180
rect 166966 227140 214288 227168
rect 214282 227128 214288 227140
rect 214340 227128 214346 227180
rect 215202 227128 215208 227180
rect 215260 227168 215266 227180
rect 255130 227168 255136 227180
rect 215260 227140 255136 227168
rect 215260 227128 215266 227140
rect 255130 227128 255136 227140
rect 255188 227128 255194 227180
rect 277210 227128 277216 227180
rect 277268 227168 277274 227180
rect 294322 227168 294328 227180
rect 277268 227140 294328 227168
rect 277268 227128 277274 227140
rect 294322 227128 294328 227140
rect 294380 227128 294386 227180
rect 363874 227128 363880 227180
rect 363932 227168 363938 227180
rect 374638 227168 374644 227180
rect 363932 227140 374644 227168
rect 363932 227128 363938 227140
rect 374638 227128 374644 227140
rect 374696 227128 374702 227180
rect 384298 227128 384304 227180
rect 384356 227168 384362 227180
rect 410610 227168 410616 227180
rect 384356 227140 410616 227168
rect 384356 227128 384362 227140
rect 410610 227128 410616 227140
rect 410668 227128 410674 227180
rect 424594 227128 424600 227180
rect 424652 227168 424658 227180
rect 472158 227168 472164 227180
rect 424652 227140 472164 227168
rect 424652 227128 424658 227140
rect 472158 227128 472164 227140
rect 472216 227128 472222 227180
rect 474274 227128 474280 227180
rect 474332 227168 474338 227180
rect 547506 227168 547512 227180
rect 474332 227140 547512 227168
rect 474332 227128 474338 227140
rect 547506 227128 547512 227140
rect 547564 227128 547570 227180
rect 63460 227004 149744 227032
rect 63460 226992 63466 227004
rect 149882 226992 149888 227044
rect 149940 227032 149946 227044
rect 149940 227004 200114 227032
rect 149940 226992 149946 227004
rect 117222 226856 117228 226908
rect 117280 226896 117286 226908
rect 184842 226896 184848 226908
rect 117280 226868 184848 226896
rect 117280 226856 117286 226868
rect 184842 226856 184848 226868
rect 184900 226856 184906 226908
rect 200086 226896 200114 227004
rect 205450 226992 205456 227044
rect 205508 227032 205514 227044
rect 205910 227032 205916 227044
rect 205508 227004 205916 227032
rect 205508 226992 205514 227004
rect 205910 226992 205916 227004
rect 205968 226992 205974 227044
rect 210970 226992 210976 227044
rect 211028 227032 211034 227044
rect 250162 227032 250168 227044
rect 211028 227004 250168 227032
rect 211028 226992 211034 227004
rect 250162 226992 250168 227004
rect 250220 226992 250226 227044
rect 256142 226992 256148 227044
rect 256200 227032 256206 227044
rect 281626 227032 281632 227044
rect 256200 227004 281632 227032
rect 256200 226992 256206 227004
rect 281626 226992 281632 227004
rect 281684 226992 281690 227044
rect 282730 226992 282736 227044
rect 282788 227032 282794 227044
rect 298186 227032 298192 227044
rect 282788 227004 298192 227032
rect 282788 226992 282794 227004
rect 298186 226992 298192 227004
rect 298244 226992 298250 227044
rect 304626 226992 304632 227044
rect 304684 227032 304690 227044
rect 314746 227032 314752 227044
rect 304684 227004 314752 227032
rect 304684 226992 304690 227004
rect 314746 226992 314752 227004
rect 314804 226992 314810 227044
rect 351730 226992 351736 227044
rect 351788 227032 351794 227044
rect 361574 227032 361580 227044
rect 351788 227004 361580 227032
rect 351788 226992 351794 227004
rect 361574 226992 361580 227004
rect 361632 226992 361638 227044
rect 366634 226992 366640 227044
rect 366692 227032 366698 227044
rect 384298 227032 384304 227044
rect 366692 227004 384304 227032
rect 366692 226992 366698 227004
rect 384298 226992 384304 227004
rect 384356 226992 384362 227044
rect 388162 226992 388168 227044
rect 388220 227032 388226 227044
rect 414934 227032 414940 227044
rect 388220 227004 414940 227032
rect 388220 226992 388226 227004
rect 414934 226992 414940 227004
rect 414992 226992 414998 227044
rect 426250 226992 426256 227044
rect 426308 227032 426314 227044
rect 473722 227032 473728 227044
rect 426308 227004 473728 227032
rect 426308 226992 426314 227004
rect 473722 226992 473728 227004
rect 473780 226992 473786 227044
rect 479794 226992 479800 227044
rect 479852 227032 479858 227044
rect 555694 227032 555700 227044
rect 479852 227004 555700 227032
rect 479852 226992 479858 227004
rect 555694 226992 555700 227004
rect 555752 226992 555758 227044
rect 210694 226896 210700 226908
rect 200086 226868 210700 226896
rect 210694 226856 210700 226868
rect 210752 226856 210758 226908
rect 249610 226856 249616 226908
rect 249668 226896 249674 226908
rect 256510 226896 256516 226908
rect 249668 226868 256516 226896
rect 249668 226856 249674 226868
rect 256510 226856 256516 226868
rect 256568 226856 256574 226908
rect 470778 226856 470784 226908
rect 470836 226896 470842 226908
rect 535914 226896 535920 226908
rect 470836 226868 535920 226896
rect 470836 226856 470842 226868
rect 535914 226856 535920 226868
rect 535972 226856 535978 226908
rect 146110 226720 146116 226772
rect 146168 226760 146174 226772
rect 205726 226760 205732 226772
rect 146168 226732 205732 226760
rect 146168 226720 146174 226732
rect 205726 226720 205732 226732
rect 205784 226720 205790 226772
rect 458634 226720 458640 226772
rect 458692 226760 458698 226772
rect 523494 226760 523500 226772
rect 458692 226732 523500 226760
rect 458692 226720 458698 226732
rect 523494 226720 523500 226732
rect 523552 226720 523558 226772
rect 129550 226584 129556 226636
rect 129608 226624 129614 226636
rect 189902 226624 189908 226636
rect 129608 226596 189908 226624
rect 129608 226584 129614 226596
rect 189902 226584 189908 226596
rect 189960 226584 189966 226636
rect 441890 226584 441896 226636
rect 441948 226624 441954 226636
rect 477586 226624 477592 226636
rect 441948 226596 477592 226624
rect 441948 226584 441954 226596
rect 477586 226584 477592 226596
rect 477644 226584 477650 226636
rect 481726 226584 481732 226636
rect 481784 226624 481790 226636
rect 515950 226624 515956 226636
rect 481784 226596 515956 226624
rect 481784 226584 481790 226596
rect 515950 226584 515956 226596
rect 516008 226584 516014 226636
rect 139302 226448 139308 226500
rect 139360 226488 139366 226500
rect 199286 226488 199292 226500
rect 139360 226460 199292 226488
rect 139360 226448 139366 226460
rect 199286 226448 199292 226460
rect 199344 226448 199350 226500
rect 391658 226380 391664 226432
rect 391716 226420 391722 226432
rect 395062 226420 395068 226432
rect 391716 226392 395068 226420
rect 391716 226380 391722 226392
rect 395062 226380 395068 226392
rect 395120 226380 395126 226432
rect 484026 226380 484032 226432
rect 484084 226420 484090 226432
rect 484084 226392 490052 226420
rect 484084 226380 484090 226392
rect 206094 226312 206100 226364
rect 206152 226352 206158 226364
rect 211522 226352 211528 226364
rect 206152 226324 211528 226352
rect 206152 226312 206158 226324
rect 211522 226312 211528 226324
rect 211580 226312 211586 226364
rect 64782 226244 64788 226296
rect 64840 226284 64846 226296
rect 125686 226284 125692 226296
rect 64840 226256 125692 226284
rect 64840 226244 64846 226256
rect 125686 226244 125692 226256
rect 125744 226244 125750 226296
rect 125870 226244 125876 226296
rect 125928 226284 125934 226296
rect 125928 226256 127756 226284
rect 125928 226244 125934 226256
rect 118602 226108 118608 226160
rect 118660 226148 118666 226160
rect 127728 226148 127756 226256
rect 129366 226244 129372 226296
rect 129424 226284 129430 226296
rect 129424 226256 137324 226284
rect 129424 226244 129430 226256
rect 137094 226148 137100 226160
rect 118660 226120 127664 226148
rect 127728 226120 137100 226148
rect 118660 226108 118666 226120
rect 122742 225972 122748 226024
rect 122800 226012 122806 226024
rect 125870 226012 125876 226024
rect 122800 225984 125876 226012
rect 122800 225972 122806 225984
rect 125870 225972 125876 225984
rect 125928 225972 125934 226024
rect 127636 226012 127664 226120
rect 137094 226108 137100 226120
rect 137152 226108 137158 226160
rect 137296 226148 137324 226256
rect 137462 226244 137468 226296
rect 137520 226284 137526 226296
rect 147950 226284 147956 226296
rect 137520 226256 147956 226284
rect 137520 226244 137526 226256
rect 147950 226244 147956 226256
rect 148008 226244 148014 226296
rect 148336 226256 157196 226284
rect 148336 226148 148364 226256
rect 137296 226120 148364 226148
rect 148502 226108 148508 226160
rect 148560 226148 148566 226160
rect 156506 226148 156512 226160
rect 148560 226120 156512 226148
rect 148560 226108 148566 226120
rect 156506 226108 156512 226120
rect 156564 226108 156570 226160
rect 157168 226148 157196 226256
rect 157288 226244 157294 226296
rect 157346 226284 157352 226296
rect 202138 226284 202144 226296
rect 157346 226256 202144 226284
rect 157346 226244 157352 226256
rect 202138 226244 202144 226256
rect 202196 226244 202202 226296
rect 214374 226244 214380 226296
rect 214432 226284 214438 226296
rect 245746 226284 245752 226296
rect 214432 226256 245752 226284
rect 214432 226244 214438 226256
rect 245746 226244 245752 226256
rect 245804 226244 245810 226296
rect 393682 226244 393688 226296
rect 393740 226284 393746 226296
rect 425698 226284 425704 226296
rect 393740 226256 425704 226284
rect 393740 226244 393746 226256
rect 425698 226244 425704 226256
rect 425756 226244 425762 226296
rect 428090 226244 428096 226296
rect 428148 226284 428154 226296
rect 461302 226284 461308 226296
rect 428148 226256 461308 226284
rect 428148 226244 428154 226256
rect 461302 226244 461308 226256
rect 461360 226244 461366 226296
rect 462682 226244 462688 226296
rect 462740 226284 462746 226296
rect 489868 226284 489874 226296
rect 462740 226256 489874 226284
rect 462740 226244 462746 226256
rect 489868 226244 489874 226256
rect 489926 226244 489932 226296
rect 490024 226284 490052 226392
rect 509602 226380 509608 226432
rect 509660 226420 509666 226432
rect 509660 226392 510016 226420
rect 509660 226380 509666 226392
rect 509988 226284 510016 226392
rect 510154 226380 510160 226432
rect 510212 226420 510218 226432
rect 510212 226392 514754 226420
rect 510212 226380 510218 226392
rect 514570 226284 514576 226296
rect 490024 226256 509924 226284
rect 509988 226256 514576 226284
rect 197722 226148 197728 226160
rect 157168 226120 197728 226148
rect 197722 226108 197728 226120
rect 197780 226108 197786 226160
rect 197906 226108 197912 226160
rect 197964 226148 197970 226160
rect 197964 226120 199976 226148
rect 197964 226108 197970 226120
rect 127636 225984 181668 226012
rect 181640 225944 181668 225984
rect 181990 225972 181996 226024
rect 182048 226012 182054 226024
rect 193306 226012 193312 226024
rect 182048 225984 193312 226012
rect 182048 225972 182054 225984
rect 193306 225972 193312 225984
rect 193364 225972 193370 226024
rect 193674 225972 193680 226024
rect 193732 226012 193738 226024
rect 195698 226012 195704 226024
rect 193732 225984 195704 226012
rect 193732 225972 193738 225984
rect 195698 225972 195704 225984
rect 195756 225972 195762 226024
rect 195882 225972 195888 226024
rect 195940 226012 195946 226024
rect 199286 226012 199292 226024
rect 195940 225984 199292 226012
rect 195940 225972 195946 225984
rect 199286 225972 199292 225984
rect 199344 225972 199350 226024
rect 199948 226012 199976 226120
rect 200114 226108 200120 226160
rect 200172 226148 200178 226160
rect 242986 226148 242992 226160
rect 200172 226120 242992 226148
rect 200172 226108 200178 226120
rect 242986 226108 242992 226120
rect 243044 226108 243050 226160
rect 270126 226108 270132 226160
rect 270184 226148 270190 226160
rect 289906 226148 289912 226160
rect 270184 226120 289912 226148
rect 270184 226108 270190 226120
rect 289906 226108 289912 226120
rect 289964 226108 289970 226160
rect 382090 226108 382096 226160
rect 382148 226148 382154 226160
rect 407482 226148 407488 226160
rect 382148 226120 407488 226148
rect 382148 226108 382154 226120
rect 407482 226108 407488 226120
rect 407540 226108 407546 226160
rect 415762 226108 415768 226160
rect 415820 226148 415826 226160
rect 449158 226148 449164 226160
rect 415820 226120 449164 226148
rect 415820 226108 415826 226120
rect 449158 226108 449164 226120
rect 449216 226108 449222 226160
rect 453850 226108 453856 226160
rect 453908 226148 453914 226160
rect 509896 226148 509924 226256
rect 514570 226244 514576 226256
rect 514628 226244 514634 226296
rect 514726 226284 514754 226392
rect 530578 226284 530584 226296
rect 514726 226256 530584 226284
rect 530578 226244 530584 226256
rect 530636 226244 530642 226296
rect 533338 226244 533344 226296
rect 533396 226284 533402 226296
rect 556706 226284 556712 226296
rect 533396 226256 556712 226284
rect 533396 226244 533402 226256
rect 556706 226244 556712 226256
rect 556764 226244 556770 226296
rect 518894 226148 518900 226160
rect 453908 226120 509832 226148
rect 509896 226120 518900 226148
rect 453908 226108 453914 226120
rect 238294 226012 238300 226024
rect 199948 225984 238300 226012
rect 238294 225972 238300 225984
rect 238352 225972 238358 226024
rect 246850 225972 246856 226024
rect 246908 226012 246914 226024
rect 274450 226012 274456 226024
rect 246908 225984 274456 226012
rect 246908 225972 246914 225984
rect 274450 225972 274456 225984
rect 274508 225972 274514 226024
rect 399754 225972 399760 226024
rect 399812 226012 399818 226024
rect 433978 226012 433984 226024
rect 399812 225984 433984 226012
rect 399812 225972 399818 225984
rect 433978 225972 433984 225984
rect 434036 225972 434042 226024
rect 436554 225972 436560 226024
rect 436612 226012 436618 226024
rect 467282 226012 467288 226024
rect 436612 225984 467288 226012
rect 436612 225972 436618 225984
rect 467282 225972 467288 225984
rect 467340 225972 467346 226024
rect 469306 225972 469312 226024
rect 469364 226012 469370 226024
rect 489868 226012 489874 226024
rect 469364 225984 489874 226012
rect 469364 225972 469370 225984
rect 489868 225972 489874 225984
rect 489926 225972 489932 226024
rect 490006 225972 490012 226024
rect 490064 226012 490070 226024
rect 505048 226012 505054 226024
rect 490064 225984 505054 226012
rect 490064 225972 490070 225984
rect 505048 225972 505054 225984
rect 505106 225972 505112 226024
rect 505186 225972 505192 226024
rect 505244 226012 505250 226024
rect 509602 226012 509608 226024
rect 505244 225984 509608 226012
rect 505244 225972 505250 225984
rect 509602 225972 509608 225984
rect 509660 225972 509666 226024
rect 509804 226012 509832 226120
rect 518894 226108 518900 226120
rect 518952 226108 518958 226160
rect 536834 226108 536840 226160
rect 536892 226148 536898 226160
rect 561766 226148 561772 226160
rect 536892 226120 561772 226148
rect 536892 226108 536898 226120
rect 561766 226108 561772 226120
rect 561824 226108 561830 226160
rect 514570 226012 514576 226024
rect 509804 225984 514576 226012
rect 514570 225972 514576 225984
rect 514628 225972 514634 226024
rect 514708 225972 514714 226024
rect 514766 226012 514772 226024
rect 540238 226012 540244 226024
rect 514766 225984 540244 226012
rect 514766 225972 514772 225984
rect 540238 225972 540244 225984
rect 540296 225972 540302 226024
rect 181640 225916 181852 225944
rect 57882 225836 57888 225888
rect 57940 225876 57946 225888
rect 107562 225876 107568 225888
rect 57940 225848 107568 225876
rect 57940 225836 57946 225848
rect 107562 225836 107568 225848
rect 107620 225836 107626 225888
rect 115290 225836 115296 225888
rect 115348 225876 115354 225888
rect 181824 225876 181852 225916
rect 190178 225876 190184 225888
rect 115348 225848 181484 225876
rect 181824 225848 190184 225876
rect 115348 225836 115354 225848
rect 181456 225808 181484 225848
rect 190178 225836 190184 225848
rect 190236 225836 190242 225888
rect 190362 225836 190368 225888
rect 190420 225876 190426 225888
rect 204530 225876 204536 225888
rect 190420 225848 204536 225876
rect 190420 225836 190426 225848
rect 204530 225836 204536 225848
rect 204588 225836 204594 225888
rect 204714 225836 204720 225888
rect 204772 225876 204778 225888
rect 214558 225876 214564 225888
rect 204772 225848 214564 225876
rect 204772 225836 204778 225848
rect 214558 225836 214564 225848
rect 214616 225836 214622 225888
rect 244182 225836 244188 225888
rect 244240 225876 244246 225888
rect 272242 225876 272248 225888
rect 244240 225848 272248 225876
rect 244240 225836 244246 225848
rect 272242 225836 272248 225848
rect 272300 225836 272306 225888
rect 390922 225836 390928 225888
rect 390980 225876 390986 225888
rect 419718 225876 419724 225888
rect 390980 225848 419724 225876
rect 390980 225836 390986 225848
rect 419718 225836 419724 225848
rect 419776 225836 419782 225888
rect 422386 225836 422392 225888
rect 422444 225876 422450 225888
rect 458634 225876 458640 225888
rect 422444 225848 458640 225876
rect 422444 225836 422450 225848
rect 458634 225836 458640 225848
rect 458692 225836 458698 225888
rect 467650 225836 467656 225888
rect 467708 225876 467714 225888
rect 536834 225876 536840 225888
rect 467708 225848 536840 225876
rect 467708 225836 467714 225848
rect 536834 225836 536840 225848
rect 536892 225836 536898 225888
rect 181456 225780 181760 225808
rect 93578 225700 93584 225752
rect 93636 225740 93642 225752
rect 166350 225740 166356 225752
rect 93636 225712 166356 225740
rect 93636 225700 93642 225712
rect 166350 225700 166356 225712
rect 166408 225700 166414 225752
rect 181254 225740 181260 225752
rect 167104 225712 181260 225740
rect 167104 225672 167132 225712
rect 181254 225700 181260 225712
rect 181312 225700 181318 225752
rect 181732 225740 181760 225780
rect 188614 225740 188620 225752
rect 181732 225712 188620 225740
rect 188614 225700 188620 225712
rect 188672 225700 188678 225752
rect 190408 225700 190414 225752
rect 190466 225740 190472 225752
rect 234154 225740 234160 225752
rect 190466 225712 234160 225740
rect 190466 225700 190472 225712
rect 234154 225700 234160 225712
rect 234212 225700 234218 225752
rect 235902 225700 235908 225752
rect 235960 225740 235966 225752
rect 267274 225740 267280 225752
rect 235960 225712 267280 225740
rect 235960 225700 235966 225712
rect 267274 225700 267280 225712
rect 267332 225700 267338 225752
rect 267642 225700 267648 225752
rect 267700 225740 267706 225752
rect 290182 225740 290188 225752
rect 267700 225712 290188 225740
rect 267700 225700 267706 225712
rect 290182 225700 290188 225712
rect 290240 225700 290246 225752
rect 291010 225700 291016 225752
rect 291068 225740 291074 225752
rect 303154 225740 303160 225752
rect 291068 225712 303160 225740
rect 291068 225700 291074 225712
rect 303154 225700 303160 225712
rect 303212 225700 303218 225752
rect 363322 225700 363328 225752
rect 363380 225740 363386 225752
rect 376846 225740 376852 225752
rect 363380 225712 376852 225740
rect 363380 225700 363386 225712
rect 376846 225700 376852 225712
rect 376904 225700 376910 225752
rect 402514 225700 402520 225752
rect 402572 225740 402578 225752
rect 439038 225740 439044 225752
rect 402572 225712 439044 225740
rect 402572 225700 402578 225712
rect 439038 225700 439044 225712
rect 439096 225700 439102 225752
rect 447502 225700 447508 225752
rect 447560 225740 447566 225752
rect 469306 225740 469312 225752
rect 447560 225712 469312 225740
rect 447560 225700 447566 225712
rect 469306 225700 469312 225712
rect 469364 225700 469370 225752
rect 472618 225700 472624 225752
rect 472676 225740 472682 225752
rect 543734 225740 543740 225752
rect 472676 225712 543740 225740
rect 472676 225700 472682 225712
rect 543734 225700 543740 225712
rect 543792 225700 543798 225752
rect 166966 225644 167132 225672
rect 75730 225564 75736 225616
rect 75788 225604 75794 225616
rect 147766 225604 147772 225616
rect 75788 225576 147772 225604
rect 75788 225564 75794 225576
rect 147766 225564 147772 225576
rect 147824 225564 147830 225616
rect 147950 225564 147956 225616
rect 148008 225604 148014 225616
rect 156966 225604 156972 225616
rect 148008 225576 156972 225604
rect 148008 225564 148014 225576
rect 156966 225564 156972 225576
rect 157024 225564 157030 225616
rect 157150 225564 157156 225616
rect 157208 225604 157214 225616
rect 157288 225604 157294 225616
rect 157208 225576 157294 225604
rect 157208 225564 157214 225576
rect 157288 225564 157294 225576
rect 157346 225564 157352 225616
rect 157426 225564 157432 225616
rect 157484 225604 157490 225616
rect 166966 225604 166994 225644
rect 157484 225576 166994 225604
rect 157484 225564 157490 225576
rect 169018 225564 169024 225616
rect 169076 225604 169082 225616
rect 214190 225604 214196 225616
rect 169076 225576 214196 225604
rect 169076 225564 169082 225576
rect 214190 225564 214196 225576
rect 214248 225564 214254 225616
rect 214558 225564 214564 225616
rect 214616 225604 214622 225616
rect 240778 225604 240784 225616
rect 214616 225576 240784 225604
rect 214616 225564 214622 225576
rect 240778 225564 240784 225576
rect 240836 225564 240842 225616
rect 241146 225564 241152 225616
rect 241204 225604 241210 225616
rect 272794 225604 272800 225616
rect 241204 225576 272800 225604
rect 241204 225564 241210 225576
rect 272794 225564 272800 225576
rect 272852 225564 272858 225616
rect 274542 225564 274548 225616
rect 274600 225604 274606 225616
rect 292114 225604 292120 225616
rect 274600 225576 292120 225604
rect 274600 225564 274606 225576
rect 292114 225564 292120 225576
rect 292172 225564 292178 225616
rect 294966 225564 294972 225616
rect 295024 225604 295030 225616
rect 308122 225604 308128 225616
rect 295024 225576 308128 225604
rect 295024 225564 295030 225576
rect 308122 225564 308128 225576
rect 308180 225564 308186 225616
rect 308950 225564 308956 225616
rect 309008 225604 309014 225616
rect 317506 225604 317512 225616
rect 309008 225576 317512 225604
rect 309008 225564 309014 225576
rect 317506 225564 317512 225576
rect 317564 225564 317570 225616
rect 359274 225564 359280 225616
rect 359332 225604 359338 225616
rect 370222 225604 370228 225616
rect 359332 225576 370228 225604
rect 359332 225564 359338 225576
rect 370222 225564 370228 225576
rect 370280 225564 370286 225616
rect 371602 225564 371608 225616
rect 371660 225604 371666 225616
rect 392578 225604 392584 225616
rect 371660 225576 392584 225604
rect 371660 225564 371666 225576
rect 392578 225564 392584 225576
rect 392636 225564 392642 225616
rect 438394 225564 438400 225616
rect 438452 225604 438458 225616
rect 472618 225604 472624 225616
rect 438452 225576 472624 225604
rect 438452 225564 438458 225576
rect 472618 225564 472624 225576
rect 472676 225564 472682 225616
rect 475930 225564 475936 225616
rect 475988 225604 475994 225616
rect 504726 225604 504732 225616
rect 475988 225576 504732 225604
rect 475988 225564 475994 225576
rect 504726 225564 504732 225576
rect 504784 225564 504790 225616
rect 505186 225564 505192 225616
rect 505244 225604 505250 225616
rect 549898 225604 549904 225616
rect 505244 225576 549904 225604
rect 505244 225564 505250 225576
rect 549898 225564 549904 225576
rect 549956 225564 549962 225616
rect 125226 225428 125232 225480
rect 125284 225468 125290 225480
rect 195514 225468 195520 225480
rect 125284 225440 195520 225468
rect 125284 225428 125290 225440
rect 195514 225428 195520 225440
rect 195572 225428 195578 225480
rect 195698 225428 195704 225480
rect 195756 225468 195762 225480
rect 197722 225468 197728 225480
rect 195756 225440 197728 225468
rect 195756 225428 195762 225440
rect 197722 225428 197728 225440
rect 197780 225428 197786 225480
rect 197906 225428 197912 225480
rect 197964 225468 197970 225480
rect 204714 225468 204720 225480
rect 197964 225440 204720 225468
rect 197964 225428 197970 225440
rect 204714 225428 204720 225440
rect 204772 225428 204778 225480
rect 204898 225428 204904 225480
rect 204956 225468 204962 225480
rect 241882 225468 241888 225480
rect 204956 225440 241888 225468
rect 204956 225428 204962 225440
rect 241882 225428 241888 225440
rect 241940 225428 241946 225480
rect 432874 225428 432880 225480
rect 432932 225468 432938 225480
rect 464522 225468 464528 225480
rect 432932 225440 464528 225468
rect 432932 225428 432938 225440
rect 464522 225428 464528 225440
rect 464580 225428 464586 225480
rect 464706 225428 464712 225480
rect 464764 225468 464770 225480
rect 531958 225468 531964 225480
rect 464764 225440 531964 225468
rect 464764 225428 464770 225440
rect 531958 225428 531964 225440
rect 532016 225428 532022 225480
rect 125686 225292 125692 225344
rect 125744 225332 125750 225344
rect 133874 225332 133880 225344
rect 125744 225304 133880 225332
rect 125744 225292 125750 225304
rect 133874 225292 133880 225304
rect 133932 225292 133938 225344
rect 137094 225292 137100 225344
rect 137152 225332 137158 225344
rect 141602 225332 141608 225344
rect 137152 225304 141608 225332
rect 137152 225292 137158 225304
rect 141602 225292 141608 225304
rect 141660 225292 141666 225344
rect 141786 225292 141792 225344
rect 141844 225332 141850 225344
rect 206554 225332 206560 225344
rect 141844 225304 206560 225332
rect 141844 225292 141850 225304
rect 206554 225292 206560 225304
rect 206612 225292 206618 225344
rect 208026 225292 208032 225344
rect 208084 225332 208090 225344
rect 250714 225332 250720 225344
rect 208084 225304 250720 225332
rect 208084 225292 208090 225304
rect 250714 225292 250720 225304
rect 250772 225292 250778 225344
rect 418522 225292 418528 225344
rect 418580 225332 418586 225344
rect 446398 225332 446404 225344
rect 418580 225304 446404 225332
rect 418580 225292 418586 225304
rect 446398 225292 446404 225304
rect 446456 225292 446462 225344
rect 459370 225292 459376 225344
rect 459428 225332 459434 225344
rect 525058 225332 525064 225344
rect 459428 225304 525064 225332
rect 459428 225292 459434 225304
rect 525058 225292 525064 225304
rect 525116 225292 525122 225344
rect 107562 225156 107568 225208
rect 107620 225196 107626 225208
rect 130102 225196 130108 225208
rect 107620 225168 130108 225196
rect 107620 225156 107626 225168
rect 130102 225156 130108 225168
rect 130160 225156 130166 225208
rect 132402 225156 132408 225208
rect 132460 225196 132466 225208
rect 199654 225196 199660 225208
rect 132460 225168 199660 225196
rect 132460 225156 132466 225168
rect 199654 225156 199660 225168
rect 199712 225156 199718 225208
rect 199838 225156 199844 225208
rect 199896 225196 199902 225208
rect 204898 225196 204904 225208
rect 199896 225168 204904 225196
rect 199896 225156 199902 225168
rect 204898 225156 204904 225168
rect 204956 225156 204962 225208
rect 205082 225156 205088 225208
rect 205140 225196 205146 225208
rect 214374 225196 214380 225208
rect 205140 225168 214380 225196
rect 205140 225156 205146 225168
rect 214374 225156 214380 225168
rect 214432 225156 214438 225208
rect 217318 225156 217324 225208
rect 217376 225196 217382 225208
rect 229186 225196 229192 225208
rect 217376 225168 229192 225196
rect 217376 225156 217382 225168
rect 229186 225156 229192 225168
rect 229244 225156 229250 225208
rect 406378 225156 406384 225208
rect 406436 225196 406442 225208
rect 443914 225196 443920 225208
rect 406436 225168 443920 225196
rect 406436 225156 406442 225168
rect 443914 225156 443920 225168
rect 443972 225156 443978 225208
rect 461118 225156 461124 225208
rect 461176 225196 461182 225208
rect 528462 225196 528468 225208
rect 461176 225168 528468 225196
rect 461176 225156 461182 225168
rect 528462 225156 528468 225168
rect 528520 225156 528526 225208
rect 116946 225020 116952 225072
rect 117004 225060 117010 225072
rect 117866 225060 117872 225072
rect 117004 225032 117872 225060
rect 117004 225020 117010 225032
rect 117866 225020 117872 225032
rect 117924 225020 117930 225072
rect 135070 225020 135076 225072
rect 135128 225060 135134 225072
rect 137462 225060 137468 225072
rect 135128 225032 137468 225060
rect 135128 225020 135134 225032
rect 137462 225020 137468 225032
rect 137520 225020 137526 225072
rect 139118 225020 139124 225072
rect 139176 225060 139182 225072
rect 204346 225060 204352 225072
rect 139176 225032 204352 225060
rect 139176 225020 139182 225032
rect 204346 225020 204352 225032
rect 204404 225020 204410 225072
rect 204530 225020 204536 225072
rect 204588 225060 204594 225072
rect 212074 225060 212080 225072
rect 204588 225032 212080 225060
rect 204588 225020 204594 225032
rect 212074 225020 212080 225032
rect 212132 225020 212138 225072
rect 214190 225020 214196 225072
rect 214248 225060 214254 225072
rect 218698 225060 218704 225072
rect 214248 225032 218704 225060
rect 214248 225020 214254 225032
rect 218698 225020 218704 225032
rect 218756 225020 218762 225072
rect 465994 225020 466000 225072
rect 466052 225060 466058 225072
rect 534994 225060 535000 225072
rect 466052 225032 535000 225060
rect 466052 225020 466058 225032
rect 534994 225020 535000 225032
rect 535052 225020 535058 225072
rect 553394 225060 553400 225072
rect 552584 225032 553400 225060
rect 273162 224952 273168 225004
rect 273220 224992 273226 225004
rect 275646 224992 275652 225004
rect 273220 224964 275652 224992
rect 273220 224952 273226 224964
rect 275646 224952 275652 224964
rect 275704 224952 275710 225004
rect 42426 224884 42432 224936
rect 42484 224924 42490 224936
rect 47118 224924 47124 224936
rect 42484 224896 47124 224924
rect 42484 224884 42490 224896
rect 47118 224884 47124 224896
rect 47176 224884 47182 224936
rect 96246 224884 96252 224936
rect 96304 224924 96310 224936
rect 171594 224924 171600 224936
rect 96304 224896 171600 224924
rect 96304 224884 96310 224896
rect 171594 224884 171600 224896
rect 171652 224884 171658 224936
rect 182266 224924 182272 224936
rect 171796 224896 182272 224924
rect 106182 224748 106188 224800
rect 106240 224788 106246 224800
rect 171796 224788 171824 224896
rect 182266 224884 182272 224896
rect 182324 224884 182330 224936
rect 185394 224884 185400 224936
rect 185452 224924 185458 224936
rect 185452 224896 190454 224924
rect 185452 224884 185458 224896
rect 106240 224760 171824 224788
rect 106240 224748 106246 224760
rect 171962 224748 171968 224800
rect 172020 224788 172026 224800
rect 173434 224788 173440 224800
rect 172020 224760 173440 224788
rect 172020 224748 172026 224760
rect 173434 224748 173440 224760
rect 173492 224748 173498 224800
rect 175090 224748 175096 224800
rect 175148 224788 175154 224800
rect 185578 224788 185584 224800
rect 175148 224760 185584 224788
rect 175148 224748 175154 224760
rect 185578 224748 185584 224760
rect 185636 224748 185642 224800
rect 190426 224788 190454 224896
rect 191466 224884 191472 224936
rect 191524 224924 191530 224936
rect 239674 224924 239680 224936
rect 191524 224896 239680 224924
rect 191524 224884 191530 224896
rect 239674 224884 239680 224896
rect 239732 224884 239738 224936
rect 419994 224884 420000 224936
rect 420052 224924 420058 224936
rect 454862 224924 454868 224936
rect 420052 224896 454868 224924
rect 420052 224884 420058 224896
rect 454862 224884 454868 224896
rect 454920 224884 454926 224936
rect 470962 224884 470968 224936
rect 471020 224924 471026 224936
rect 542354 224924 542360 224936
rect 471020 224896 542360 224924
rect 471020 224884 471026 224896
rect 542354 224884 542360 224896
rect 542412 224884 542418 224936
rect 543734 224884 543740 224936
rect 543792 224924 543798 224936
rect 545022 224924 545028 224936
rect 543792 224896 545028 224924
rect 543792 224884 543798 224896
rect 545022 224884 545028 224896
rect 545080 224924 545086 224936
rect 552584 224924 552612 225032
rect 553394 225020 553400 225032
rect 553452 225020 553458 225072
rect 545080 224896 552612 224924
rect 545080 224884 545086 224896
rect 552750 224884 552756 224936
rect 552808 224924 552814 224936
rect 559006 224924 559012 224936
rect 552808 224896 559012 224924
rect 552808 224884 552814 224896
rect 559006 224884 559012 224896
rect 559064 224884 559070 224936
rect 194778 224788 194784 224800
rect 190426 224760 194784 224788
rect 194778 224748 194784 224760
rect 194836 224748 194842 224800
rect 195238 224748 195244 224800
rect 195296 224788 195302 224800
rect 237466 224788 237472 224800
rect 195296 224760 237472 224788
rect 195296 224748 195302 224760
rect 237466 224748 237472 224760
rect 237524 224748 237530 224800
rect 255222 224748 255228 224800
rect 255280 224788 255286 224800
rect 280522 224788 280528 224800
rect 255280 224760 280528 224788
rect 255280 224748 255286 224760
rect 280522 224748 280528 224760
rect 280580 224748 280586 224800
rect 408586 224748 408592 224800
rect 408644 224788 408650 224800
rect 447226 224788 447232 224800
rect 408644 224760 447232 224788
rect 408644 224748 408650 224760
rect 447226 224748 447232 224760
rect 447284 224748 447290 224800
rect 480346 224748 480352 224800
rect 480404 224788 480410 224800
rect 483658 224788 483664 224800
rect 480404 224760 483664 224788
rect 480404 224748 480410 224760
rect 483658 224748 483664 224760
rect 483716 224748 483722 224800
rect 485866 224748 485872 224800
rect 485924 224788 485930 224800
rect 485924 224760 486096 224788
rect 485924 224748 485930 224760
rect 85298 224612 85304 224664
rect 85356 224652 85362 224664
rect 165982 224652 165988 224664
rect 85356 224624 165988 224652
rect 85356 224612 85362 224624
rect 165982 224612 165988 224624
rect 166040 224612 166046 224664
rect 166258 224612 166264 224664
rect 166316 224652 166322 224664
rect 221642 224652 221648 224664
rect 166316 224624 221648 224652
rect 166316 224612 166322 224624
rect 221642 224612 221648 224624
rect 221700 224612 221706 224664
rect 257338 224652 257344 224664
rect 229066 224624 257344 224652
rect 89622 224476 89628 224528
rect 89680 224516 89686 224528
rect 171226 224516 171232 224528
rect 89680 224488 171232 224516
rect 89680 224476 89686 224488
rect 171226 224476 171232 224488
rect 171284 224476 171290 224528
rect 171594 224476 171600 224528
rect 171652 224516 171658 224528
rect 175642 224516 175648 224528
rect 171652 224488 175648 224516
rect 171652 224476 171658 224488
rect 175642 224476 175648 224488
rect 175700 224476 175706 224528
rect 185394 224516 185400 224528
rect 175844 224488 185400 224516
rect 82722 224340 82728 224392
rect 82780 224380 82786 224392
rect 166534 224380 166540 224392
rect 82780 224352 166540 224380
rect 82780 224340 82786 224352
rect 166534 224340 166540 224352
rect 166592 224340 166598 224392
rect 168190 224340 168196 224392
rect 168248 224380 168254 224392
rect 171962 224380 171968 224392
rect 168248 224352 171968 224380
rect 168248 224340 168254 224352
rect 171962 224340 171968 224352
rect 172020 224340 172026 224392
rect 173250 224340 173256 224392
rect 173308 224380 173314 224392
rect 175844 224380 175872 224488
rect 185394 224476 185400 224488
rect 185452 224476 185458 224528
rect 185578 224476 185584 224528
rect 185636 224516 185642 224528
rect 221274 224516 221280 224528
rect 185636 224488 221280 224516
rect 185636 224476 185642 224488
rect 221274 224476 221280 224488
rect 221332 224476 221338 224528
rect 221458 224476 221464 224528
rect 221516 224516 221522 224528
rect 229066 224516 229094 224624
rect 257338 224612 257344 224624
rect 257396 224612 257402 224664
rect 379882 224612 379888 224664
rect 379940 224652 379946 224664
rect 402974 224652 402980 224664
rect 379940 224624 402980 224652
rect 379940 224612 379946 224624
rect 402974 224612 402980 224624
rect 403032 224612 403038 224664
rect 413002 224612 413008 224664
rect 413060 224652 413066 224664
rect 453850 224652 453856 224664
rect 413060 224624 453856 224652
rect 413060 224612 413066 224624
rect 453850 224612 453856 224624
rect 453908 224612 453914 224664
rect 457714 224612 457720 224664
rect 457772 224652 457778 224664
rect 486068 224652 486096 224760
rect 486234 224748 486240 224800
rect 486292 224788 486298 224800
rect 556522 224788 556528 224800
rect 486292 224760 556528 224788
rect 486292 224748 486298 224760
rect 556522 224748 556528 224760
rect 556580 224748 556586 224800
rect 556706 224748 556712 224800
rect 556764 224788 556770 224800
rect 557350 224788 557356 224800
rect 556764 224760 557356 224788
rect 556764 224748 556770 224760
rect 557350 224748 557356 224760
rect 557408 224748 557414 224800
rect 557810 224748 557816 224800
rect 557868 224788 557874 224800
rect 561490 224788 561496 224800
rect 557868 224760 561496 224788
rect 557868 224748 557874 224760
rect 561490 224748 561496 224760
rect 561548 224748 561554 224800
rect 552750 224652 552756 224664
rect 457772 224624 485636 224652
rect 486068 224624 552756 224652
rect 457772 224612 457778 224624
rect 221516 224488 229094 224516
rect 221516 224476 221522 224488
rect 250898 224476 250904 224528
rect 250956 224516 250962 224528
rect 279418 224516 279424 224528
rect 250956 224488 279424 224516
rect 250956 224476 250962 224488
rect 279418 224476 279424 224488
rect 279476 224476 279482 224528
rect 279970 224476 279976 224528
rect 280028 224516 280034 224528
rect 296530 224516 296536 224528
rect 280028 224488 296536 224516
rect 280028 224476 280034 224488
rect 296530 224476 296536 224488
rect 296588 224476 296594 224528
rect 370866 224476 370872 224528
rect 370924 224516 370930 224528
rect 383470 224516 383476 224528
rect 370924 224488 383476 224516
rect 370924 224476 370930 224488
rect 383470 224476 383476 224488
rect 383528 224476 383534 224528
rect 387610 224476 387616 224528
rect 387668 224516 387674 224528
rect 413278 224516 413284 224528
rect 387668 224488 413284 224516
rect 387668 224476 387674 224488
rect 413278 224476 413284 224488
rect 413336 224476 413342 224528
rect 414658 224476 414664 224528
rect 414716 224516 414722 224528
rect 425882 224516 425888 224528
rect 414716 224488 425888 224516
rect 414716 224476 414722 224488
rect 425882 224476 425888 224488
rect 425940 224476 425946 224528
rect 434162 224476 434168 224528
rect 434220 224516 434226 224528
rect 481818 224516 481824 224528
rect 434220 224488 481824 224516
rect 434220 224476 434226 224488
rect 481818 224476 481824 224488
rect 481876 224476 481882 224528
rect 482002 224476 482008 224528
rect 482060 224516 482066 224528
rect 484854 224516 484860 224528
rect 482060 224488 484860 224516
rect 482060 224476 482066 224488
rect 484854 224476 484860 224488
rect 484912 224476 484918 224528
rect 485608 224516 485636 224624
rect 552750 224612 552756 224624
rect 552808 224612 552814 224664
rect 552934 224612 552940 224664
rect 552992 224652 552998 224664
rect 552992 224624 572714 224652
rect 552992 224612 552998 224624
rect 487982 224516 487988 224528
rect 485608 224488 487988 224516
rect 487982 224476 487988 224488
rect 488040 224476 488046 224528
rect 491938 224476 491944 224528
rect 491996 224516 492002 224528
rect 557810 224516 557816 224528
rect 491996 224488 557816 224516
rect 491996 224476 492002 224488
rect 557810 224476 557816 224488
rect 557868 224476 557874 224528
rect 557994 224476 558000 224528
rect 558052 224516 558058 224528
rect 566458 224516 566464 224528
rect 558052 224488 566464 224516
rect 558052 224476 558058 224488
rect 566458 224476 566464 224488
rect 566516 224476 566522 224528
rect 173308 224352 175872 224380
rect 173308 224340 173314 224352
rect 176010 224340 176016 224392
rect 176068 224380 176074 224392
rect 224218 224380 224224 224392
rect 176068 224352 224224 224380
rect 176068 224340 176074 224352
rect 224218 224340 224224 224352
rect 224276 224340 224282 224392
rect 226058 224340 226064 224392
rect 226116 224380 226122 224392
rect 260374 224380 260380 224392
rect 226116 224352 260380 224380
rect 226116 224340 226122 224352
rect 260374 224340 260380 224352
rect 260432 224340 260438 224392
rect 283282 224380 283288 224392
rect 267706 224352 283288 224380
rect 57238 224204 57244 224256
rect 57296 224244 57302 224256
rect 142108 224244 142114 224256
rect 57296 224216 142114 224244
rect 57296 224204 57302 224216
rect 142108 224204 142114 224216
rect 142166 224204 142172 224256
rect 142246 224204 142252 224256
rect 142304 224244 142310 224256
rect 156690 224244 156696 224256
rect 142304 224216 156696 224244
rect 142304 224204 142310 224216
rect 156690 224204 156696 224216
rect 156748 224204 156754 224256
rect 156966 224204 156972 224256
rect 157024 224244 157030 224256
rect 158530 224244 158536 224256
rect 157024 224216 158536 224244
rect 157024 224204 157030 224216
rect 158530 224204 158536 224216
rect 158588 224204 158594 224256
rect 158714 224204 158720 224256
rect 158772 224244 158778 224256
rect 217594 224244 217600 224256
rect 158772 224216 217600 224244
rect 158772 224204 158778 224216
rect 217594 224204 217600 224216
rect 217652 224204 217658 224256
rect 224586 224204 224592 224256
rect 224644 224244 224650 224256
rect 261754 224244 261760 224256
rect 224644 224216 261760 224244
rect 224644 224204 224650 224216
rect 261754 224204 261760 224216
rect 261812 224204 261818 224256
rect 262674 224204 262680 224256
rect 262732 224244 262738 224256
rect 264514 224244 264520 224256
rect 262732 224216 264520 224244
rect 262732 224204 262738 224216
rect 264514 224204 264520 224216
rect 264572 224204 264578 224256
rect 101398 224068 101404 224120
rect 101456 224108 101462 224120
rect 168374 224108 168380 224120
rect 101456 224080 168380 224108
rect 101456 224068 101462 224080
rect 168374 224068 168380 224080
rect 168432 224068 168438 224120
rect 168558 224068 168564 224120
rect 168616 224108 168622 224120
rect 172238 224108 172244 224120
rect 168616 224080 172244 224108
rect 168616 224068 168622 224080
rect 172238 224068 172244 224080
rect 172296 224068 172302 224120
rect 172606 224068 172612 224120
rect 172664 224108 172670 224120
rect 172664 224080 173250 224108
rect 172664 224068 172670 224080
rect 92106 223932 92112 223984
rect 92164 223972 92170 223984
rect 173066 223972 173072 223984
rect 92164 223944 173072 223972
rect 92164 223932 92170 223944
rect 173066 223932 173072 223944
rect 173124 223932 173130 223984
rect 173222 223972 173250 224080
rect 173434 224068 173440 224120
rect 173492 224108 173498 224120
rect 176010 224108 176016 224120
rect 173492 224080 176016 224108
rect 173492 224068 173498 224080
rect 176010 224068 176016 224080
rect 176068 224068 176074 224120
rect 176378 224068 176384 224120
rect 176436 224108 176442 224120
rect 193858 224108 193864 224120
rect 176436 224080 193864 224108
rect 176436 224068 176442 224080
rect 193858 224068 193864 224080
rect 193916 224068 193922 224120
rect 194778 224068 194784 224120
rect 194836 224108 194842 224120
rect 198642 224108 198648 224120
rect 194836 224080 198648 224108
rect 194836 224068 194842 224080
rect 198642 224068 198648 224080
rect 198700 224068 198706 224120
rect 216490 224068 216496 224120
rect 216548 224108 216554 224120
rect 254026 224108 254032 224120
rect 216548 224080 254032 224108
rect 216548 224068 216554 224080
rect 254026 224068 254032 224080
rect 254084 224068 254090 224120
rect 260190 224068 260196 224120
rect 260248 224108 260254 224120
rect 267706 224108 267734 224352
rect 283282 224340 283288 224352
rect 283340 224340 283346 224392
rect 296622 224340 296628 224392
rect 296680 224380 296686 224392
rect 304074 224380 304080 224392
rect 296680 224352 304080 224380
rect 296680 224340 296686 224352
rect 304074 224340 304080 224352
rect 304132 224340 304138 224392
rect 358446 224340 358452 224392
rect 358504 224380 358510 224392
rect 372706 224380 372712 224392
rect 358504 224352 372712 224380
rect 358504 224340 358510 224352
rect 372706 224340 372712 224352
rect 372764 224340 372770 224392
rect 383010 224340 383016 224392
rect 383068 224380 383074 224392
rect 403434 224380 403440 224392
rect 383068 224352 403440 224380
rect 383068 224340 383074 224352
rect 403434 224340 403440 224352
rect 403492 224340 403498 224392
rect 403618 224340 403624 224392
rect 403676 224380 403682 224392
rect 405366 224380 405372 224392
rect 403676 224352 405372 224380
rect 403676 224340 403682 224352
rect 405366 224340 405372 224352
rect 405424 224340 405430 224392
rect 410794 224340 410800 224392
rect 410852 224380 410858 224392
rect 434162 224380 434168 224392
rect 410852 224352 434168 224380
rect 410852 224340 410858 224352
rect 434162 224340 434168 224352
rect 434220 224340 434226 224392
rect 485038 224380 485044 224392
rect 435560 224352 485044 224380
rect 275278 224204 275284 224256
rect 275336 224244 275342 224256
rect 294782 224244 294788 224256
rect 275336 224216 294788 224244
rect 275336 224204 275342 224216
rect 294782 224204 294788 224216
rect 294840 224204 294846 224256
rect 296438 224204 296444 224256
rect 296496 224244 296502 224256
rect 307294 224244 307300 224256
rect 296496 224216 307300 224244
rect 296496 224204 296502 224216
rect 307294 224204 307300 224216
rect 307352 224204 307358 224256
rect 307478 224204 307484 224256
rect 307536 224244 307542 224256
rect 316678 224244 316684 224256
rect 307536 224216 316684 224244
rect 307536 224204 307542 224216
rect 316678 224204 316684 224216
rect 316736 224204 316742 224256
rect 331214 224204 331220 224256
rect 331272 224244 331278 224256
rect 332134 224244 332140 224256
rect 331272 224216 332140 224244
rect 331272 224204 331278 224216
rect 332134 224204 332140 224216
rect 332192 224204 332198 224256
rect 335722 224204 335728 224256
rect 335780 224244 335786 224256
rect 336274 224244 336280 224256
rect 335780 224216 336280 224244
rect 335780 224204 335786 224216
rect 336274 224204 336280 224216
rect 336332 224204 336338 224256
rect 352282 224204 352288 224256
rect 352340 224244 352346 224256
rect 358078 224244 358084 224256
rect 352340 224216 358084 224244
rect 352340 224204 352346 224216
rect 358078 224204 358084 224216
rect 358136 224204 358142 224256
rect 370406 224204 370412 224256
rect 370464 224244 370470 224256
rect 386782 224244 386788 224256
rect 370464 224216 386788 224244
rect 370464 224204 370470 224216
rect 386782 224204 386788 224216
rect 386840 224204 386846 224256
rect 388806 224204 388812 224256
rect 388864 224244 388870 224256
rect 417418 224244 417424 224256
rect 388864 224216 417424 224244
rect 388864 224204 388870 224216
rect 417418 224204 417424 224216
rect 417476 224204 417482 224256
rect 432322 224204 432328 224256
rect 432380 224244 432386 224256
rect 435358 224244 435364 224256
rect 432380 224216 435364 224244
rect 432380 224204 432386 224216
rect 435358 224204 435364 224216
rect 435416 224204 435422 224256
rect 260248 224080 267734 224108
rect 260248 224068 260254 224080
rect 403434 224068 403440 224120
rect 403492 224108 403498 224120
rect 409138 224108 409144 224120
rect 403492 224080 409144 224108
rect 403492 224068 403498 224080
rect 409138 224068 409144 224080
rect 409196 224068 409202 224120
rect 409690 224068 409696 224120
rect 409748 224108 409754 224120
rect 421834 224108 421840 224120
rect 409748 224080 421840 224108
rect 409748 224068 409754 224080
rect 421834 224068 421840 224080
rect 421892 224068 421898 224120
rect 433794 224068 433800 224120
rect 433852 224108 433858 224120
rect 435560 224108 435588 224352
rect 485038 224340 485044 224352
rect 485096 224340 485102 224392
rect 490742 224340 490748 224392
rect 490800 224380 490806 224392
rect 563974 224380 563980 224392
rect 490800 224352 563980 224380
rect 490800 224340 490806 224352
rect 563974 224340 563980 224352
rect 564032 224340 564038 224392
rect 486786 224312 486792 224324
rect 486068 224284 486792 224312
rect 438210 224204 438216 224256
rect 438268 224244 438274 224256
rect 484670 224244 484676 224256
rect 438268 224216 484676 224244
rect 438268 224204 438274 224216
rect 484670 224204 484676 224216
rect 484728 224204 484734 224256
rect 433852 224080 435588 224108
rect 433852 224068 433858 224080
rect 442626 224068 442632 224120
rect 442684 224108 442690 224120
rect 486068 224108 486096 224284
rect 486786 224272 486792 224284
rect 486844 224272 486850 224324
rect 572686 224312 572714 224624
rect 590930 224408 590936 224460
rect 590988 224448 590994 224460
rect 597554 224448 597560 224460
rect 590988 224420 597560 224448
rect 590988 224408 590994 224420
rect 597554 224408 597560 224420
rect 597612 224408 597618 224460
rect 572686 224284 591344 224312
rect 486970 224204 486976 224256
rect 487028 224244 487034 224256
rect 557994 224244 558000 224256
rect 487028 224216 558000 224244
rect 487028 224204 487034 224216
rect 557994 224204 558000 224216
rect 558052 224204 558058 224256
rect 591114 224176 591120 224188
rect 558196 224148 591120 224176
rect 442684 224080 486096 224108
rect 442684 224068 442690 224080
rect 487982 224068 487988 224120
rect 488040 224108 488046 224120
rect 522574 224108 522580 224120
rect 488040 224080 522580 224108
rect 488040 224068 488046 224080
rect 522574 224068 522580 224080
rect 522632 224068 522638 224120
rect 536834 224000 536840 224052
rect 536892 224040 536898 224052
rect 537478 224040 537484 224052
rect 536892 224012 537484 224040
rect 536892 224000 536898 224012
rect 537478 224000 537484 224012
rect 537536 224040 537542 224052
rect 537536 224012 544240 224040
rect 537536 224000 537542 224012
rect 210418 223972 210424 223984
rect 173222 223944 210424 223972
rect 210418 223932 210424 223944
rect 210476 223932 210482 223984
rect 219342 223972 219348 223984
rect 215266 223944 219348 223972
rect 113818 223796 113824 223848
rect 113876 223836 113882 223848
rect 161842 223836 161848 223848
rect 113876 223808 161848 223836
rect 113876 223796 113882 223808
rect 161842 223796 161848 223808
rect 161900 223796 161906 223848
rect 162486 223796 162492 223848
rect 162544 223836 162550 223848
rect 215266 223836 215294 223944
rect 219342 223932 219348 223944
rect 219400 223932 219406 223984
rect 221274 223932 221280 223984
rect 221332 223972 221338 223984
rect 228634 223972 228640 223984
rect 221332 223944 228640 223972
rect 221332 223932 221338 223944
rect 228634 223932 228640 223944
rect 228692 223932 228698 223984
rect 417602 223932 417608 223984
rect 417660 223972 417666 223984
rect 431218 223972 431224 223984
rect 417660 223944 431224 223972
rect 417660 223932 417666 223944
rect 431218 223932 431224 223944
rect 431276 223932 431282 223984
rect 431770 223932 431776 223984
rect 431828 223972 431834 223984
rect 438302 223972 438308 223984
rect 431828 223944 438308 223972
rect 431828 223932 431834 223944
rect 438302 223932 438308 223944
rect 438360 223932 438366 223984
rect 454402 223932 454408 223984
rect 454460 223972 454466 223984
rect 485682 223972 485688 223984
rect 454460 223944 485688 223972
rect 454460 223932 454466 223944
rect 485682 223932 485688 223944
rect 485740 223932 485746 223984
rect 485866 223932 485872 223984
rect 485924 223972 485930 223984
rect 517606 223972 517612 223984
rect 485924 223944 517612 223972
rect 485924 223932 485930 223944
rect 517606 223932 517612 223944
rect 517664 223972 517670 223984
rect 517664 223944 518894 223972
rect 517664 223932 517670 223944
rect 518866 223904 518894 223944
rect 544010 223904 544016 223916
rect 518866 223876 544016 223904
rect 544010 223864 544016 223876
rect 544068 223864 544074 223916
rect 544212 223904 544240 224012
rect 544378 224000 544384 224052
rect 544436 224040 544442 224052
rect 558196 224040 558224 224148
rect 591114 224136 591120 224148
rect 591172 224136 591178 224188
rect 591316 224176 591344 224284
rect 610434 224272 610440 224324
rect 610492 224312 610498 224324
rect 610492 224284 615494 224312
rect 610492 224272 610498 224284
rect 610802 224176 610808 224188
rect 591316 224148 610808 224176
rect 610802 224136 610808 224148
rect 610860 224136 610866 224188
rect 615466 224176 615494 224284
rect 617702 224176 617708 224188
rect 615466 224148 617708 224176
rect 617702 224136 617708 224148
rect 617760 224136 617766 224188
rect 544436 224012 558224 224040
rect 544436 224000 544442 224012
rect 558546 224000 558552 224052
rect 558604 224040 558610 224052
rect 626718 224040 626724 224052
rect 558604 224012 626724 224040
rect 558604 224000 558610 224012
rect 626718 224000 626724 224012
rect 626776 224000 626782 224052
rect 552934 223904 552940 223916
rect 544212 223876 552940 223904
rect 552934 223864 552940 223876
rect 552992 223864 552998 223916
rect 553394 223864 553400 223916
rect 553452 223904 553458 223916
rect 623774 223904 623780 223916
rect 553452 223876 623780 223904
rect 553452 223864 553458 223876
rect 623774 223864 623780 223876
rect 623832 223864 623838 223916
rect 162544 223808 215294 223836
rect 162544 223796 162550 223808
rect 219342 223796 219348 223848
rect 219400 223836 219406 223848
rect 256326 223836 256332 223848
rect 219400 223808 256332 223836
rect 219400 223796 219406 223808
rect 256326 223796 256332 223808
rect 256384 223796 256390 223848
rect 452746 223796 452752 223848
rect 452804 223836 452810 223848
rect 485682 223836 485688 223848
rect 452804 223808 485688 223836
rect 452804 223796 452810 223808
rect 485682 223796 485688 223808
rect 485740 223796 485746 223848
rect 485866 223796 485872 223848
rect 485924 223836 485930 223848
rect 515122 223836 515128 223848
rect 485924 223808 515128 223836
rect 485924 223796 485930 223808
rect 515122 223796 515128 223808
rect 515180 223836 515186 223848
rect 515180 223808 517008 223836
rect 515180 223796 515186 223808
rect 317230 223728 317236 223780
rect 317288 223768 317294 223780
rect 323578 223768 323584 223780
rect 317288 223740 323584 223768
rect 317288 223728 317294 223740
rect 323578 223728 323584 223740
rect 323636 223728 323642 223780
rect 516980 223768 517008 223808
rect 516980 223740 610664 223768
rect 129734 223660 129740 223712
rect 129792 223700 129798 223712
rect 187234 223700 187240 223712
rect 129792 223672 187240 223700
rect 129792 223660 129798 223672
rect 187234 223660 187240 223672
rect 187292 223660 187298 223712
rect 188798 223660 188804 223712
rect 188856 223700 188862 223712
rect 195238 223700 195244 223712
rect 188856 223672 195244 223700
rect 188856 223660 188862 223672
rect 195238 223660 195244 223672
rect 195296 223660 195302 223712
rect 210418 223660 210424 223712
rect 210476 223700 210482 223712
rect 221090 223700 221096 223712
rect 210476 223672 221096 223700
rect 210476 223660 210482 223672
rect 221090 223660 221096 223672
rect 221148 223660 221154 223712
rect 440050 223660 440056 223712
rect 440108 223700 440114 223712
rect 496078 223700 496084 223712
rect 440108 223672 485728 223700
rect 440108 223660 440114 223672
rect 485700 223632 485728 223672
rect 486436 223672 496084 223700
rect 486436 223632 486464 223672
rect 496078 223660 496084 223672
rect 496136 223660 496142 223712
rect 505002 223660 505008 223712
rect 505060 223700 505066 223712
rect 505060 223672 511488 223700
rect 505060 223660 505066 223672
rect 485700 223604 486464 223632
rect 511460 223632 511488 223672
rect 590930 223632 590936 223644
rect 511460 223604 590936 223632
rect 590930 223592 590936 223604
rect 590988 223592 590994 223644
rect 591114 223592 591120 223644
rect 591172 223632 591178 223644
rect 610434 223632 610440 223644
rect 591172 223604 610440 223632
rect 591172 223592 591178 223604
rect 610434 223592 610440 223604
rect 610492 223592 610498 223644
rect 610636 223632 610664 223740
rect 610802 223728 610808 223780
rect 610860 223768 610866 223780
rect 622578 223768 622584 223780
rect 610860 223740 622584 223768
rect 610860 223728 610866 223740
rect 622578 223728 622584 223740
rect 622636 223728 622642 223780
rect 617058 223632 617064 223644
rect 610636 223604 617064 223632
rect 617058 223592 617064 223604
rect 617116 223592 617122 223644
rect 42242 223524 42248 223576
rect 42300 223564 42306 223576
rect 46934 223564 46940 223576
rect 42300 223536 46940 223564
rect 42300 223524 42306 223536
rect 46934 223524 46940 223536
rect 46992 223524 46998 223576
rect 121086 223524 121092 223576
rect 121144 223564 121150 223576
rect 190546 223564 190552 223576
rect 121144 223536 190552 223564
rect 121144 223524 121150 223536
rect 190546 223524 190552 223536
rect 190604 223524 190610 223576
rect 194410 223524 194416 223576
rect 194468 223564 194474 223576
rect 239122 223564 239128 223576
rect 194468 223536 239128 223564
rect 194468 223524 194474 223536
rect 239122 223524 239128 223536
rect 239180 223524 239186 223576
rect 246666 223524 246672 223576
rect 246724 223564 246730 223576
rect 271690 223564 271696 223576
rect 246724 223536 271696 223564
rect 246724 223524 246730 223536
rect 271690 223524 271696 223536
rect 271748 223524 271754 223576
rect 305914 223524 305920 223576
rect 305972 223564 305978 223576
rect 306466 223564 306472 223576
rect 305972 223536 306472 223564
rect 305972 223524 305978 223536
rect 306466 223524 306472 223536
rect 306524 223524 306530 223576
rect 347866 223524 347872 223576
rect 347924 223564 347930 223576
rect 353662 223564 353668 223576
rect 347924 223536 353668 223564
rect 347924 223524 347930 223536
rect 353662 223524 353668 223536
rect 353720 223524 353726 223576
rect 399386 223524 399392 223576
rect 399444 223564 399450 223576
rect 418246 223564 418252 223576
rect 399444 223536 418252 223564
rect 399444 223524 399450 223536
rect 418246 223524 418252 223536
rect 418304 223524 418310 223576
rect 435634 223524 435640 223576
rect 435692 223564 435698 223576
rect 474642 223564 474648 223576
rect 435692 223536 474648 223564
rect 435692 223524 435698 223536
rect 474642 223524 474648 223536
rect 474700 223524 474706 223576
rect 477034 223524 477040 223576
rect 477092 223564 477098 223576
rect 484118 223564 484124 223576
rect 477092 223536 484124 223564
rect 477092 223524 477098 223536
rect 484118 223524 484124 223536
rect 484176 223524 484182 223576
rect 487062 223524 487068 223576
rect 487120 223564 487126 223576
rect 511258 223564 511264 223576
rect 487120 223536 511264 223564
rect 487120 223524 487126 223536
rect 511258 223524 511264 223536
rect 511316 223524 511322 223576
rect 243814 223496 243820 223508
rect 239324 223468 243820 223496
rect 108666 223388 108672 223440
rect 108724 223428 108730 223440
rect 133138 223428 133144 223440
rect 108724 223400 133144 223428
rect 108724 223388 108730 223400
rect 133138 223388 133144 223400
rect 133196 223388 133202 223440
rect 133782 223388 133788 223440
rect 133840 223428 133846 223440
rect 197170 223428 197176 223440
rect 133840 223400 197176 223428
rect 133840 223388 133846 223400
rect 197170 223388 197176 223400
rect 197228 223388 197234 223440
rect 198090 223388 198096 223440
rect 198148 223428 198154 223440
rect 239324 223428 239352 223468
rect 243814 223456 243820 223468
rect 243872 223456 243878 223508
rect 245286 223456 245292 223508
rect 245344 223496 245350 223508
rect 245344 223468 246528 223496
rect 245344 223456 245350 223468
rect 198148 223400 239352 223428
rect 246500 223428 246528 223468
rect 529382 223456 529388 223508
rect 529440 223496 529446 223508
rect 536098 223496 536104 223508
rect 529440 223468 536104 223496
rect 529440 223456 529446 223468
rect 536098 223456 536104 223468
rect 536156 223456 536162 223508
rect 246500 223400 248414 223428
rect 198148 223388 198154 223400
rect 242158 223320 242164 223372
rect 242216 223360 242222 223372
rect 246298 223360 246304 223372
rect 242216 223332 246304 223360
rect 242216 223320 242222 223332
rect 246298 223320 246304 223332
rect 246356 223320 246362 223372
rect 97902 223252 97908 223304
rect 97960 223292 97966 223304
rect 171410 223292 171416 223304
rect 97960 223264 171416 223292
rect 97960 223252 97966 223264
rect 171410 223252 171416 223264
rect 171468 223252 171474 223304
rect 171594 223252 171600 223304
rect 171652 223292 171658 223304
rect 180610 223292 180616 223304
rect 171652 223264 180616 223292
rect 171652 223252 171658 223264
rect 180610 223252 180616 223264
rect 180668 223252 180674 223304
rect 187326 223252 187332 223304
rect 187384 223292 187390 223304
rect 234706 223292 234712 223304
rect 187384 223264 234712 223292
rect 187384 223252 187390 223264
rect 234706 223252 234712 223264
rect 234764 223252 234770 223304
rect 248386 223292 248414 223400
rect 267458 223388 267464 223440
rect 267516 223428 267522 223440
rect 287698 223428 287704 223440
rect 267516 223400 287704 223428
rect 267516 223388 267522 223400
rect 287698 223388 287704 223400
rect 287756 223388 287762 223440
rect 410242 223388 410248 223440
rect 410300 223428 410306 223440
rect 448054 223428 448060 223440
rect 410300 223400 448060 223428
rect 410300 223388 410306 223400
rect 448054 223388 448060 223400
rect 448112 223388 448118 223440
rect 451274 223388 451280 223440
rect 451332 223428 451338 223440
rect 467098 223428 467104 223440
rect 451332 223400 467104 223428
rect 451332 223388 451338 223400
rect 467098 223388 467104 223400
rect 467156 223388 467162 223440
rect 468754 223388 468760 223440
rect 468812 223428 468818 223440
rect 529198 223428 529204 223440
rect 468812 223400 529204 223428
rect 468812 223388 468818 223400
rect 529198 223388 529204 223400
rect 529256 223388 529262 223440
rect 551922 223388 551928 223440
rect 551980 223428 551986 223440
rect 564802 223428 564808 223440
rect 551980 223400 564808 223428
rect 551980 223388 551986 223400
rect 564802 223388 564808 223400
rect 564860 223388 564866 223440
rect 275002 223292 275008 223304
rect 248386 223264 275008 223292
rect 275002 223252 275008 223264
rect 275060 223252 275066 223304
rect 375466 223252 375472 223304
rect 375524 223292 375530 223304
rect 397822 223292 397828 223304
rect 375524 223264 397828 223292
rect 375524 223252 375530 223264
rect 397822 223252 397828 223264
rect 397880 223252 397886 223304
rect 399570 223252 399576 223304
rect 399628 223292 399634 223304
rect 421558 223292 421564 223304
rect 399628 223264 421564 223292
rect 399628 223252 399634 223264
rect 421558 223252 421564 223264
rect 421616 223252 421622 223304
rect 431586 223252 431592 223304
rect 431644 223292 431650 223304
rect 469858 223292 469864 223304
rect 431644 223264 469864 223292
rect 431644 223252 431650 223264
rect 469858 223252 469864 223264
rect 469916 223252 469922 223304
rect 470410 223252 470416 223304
rect 470468 223292 470474 223304
rect 541618 223292 541624 223304
rect 470468 223264 541624 223292
rect 470468 223252 470474 223264
rect 541618 223252 541624 223264
rect 541676 223252 541682 223304
rect 541986 223252 541992 223304
rect 542044 223292 542050 223304
rect 557994 223292 558000 223304
rect 542044 223264 558000 223292
rect 542044 223252 542050 223264
rect 557994 223252 558000 223264
rect 558052 223252 558058 223304
rect 558196 223264 576854 223292
rect 81342 223116 81348 223168
rect 81400 223156 81406 223168
rect 160462 223156 160468 223168
rect 81400 223128 160468 223156
rect 81400 223116 81406 223128
rect 160462 223116 160468 223128
rect 160520 223116 160526 223168
rect 184474 223156 184480 223168
rect 161308 223128 184480 223156
rect 161308 223088 161336 223128
rect 184474 223116 184480 223128
rect 184532 223116 184538 223168
rect 184842 223116 184848 223168
rect 184900 223156 184906 223168
rect 232498 223156 232504 223168
rect 184900 223128 232504 223156
rect 184900 223116 184906 223128
rect 232498 223116 232504 223128
rect 232556 223116 232562 223168
rect 237006 223116 237012 223168
rect 237064 223156 237070 223168
rect 268102 223156 268108 223168
rect 237064 223128 268108 223156
rect 237064 223116 237070 223128
rect 268102 223116 268108 223128
rect 268160 223116 268166 223168
rect 284202 223116 284208 223168
rect 284260 223156 284266 223168
rect 300578 223156 300584 223168
rect 284260 223128 300584 223156
rect 284260 223116 284266 223128
rect 300578 223116 300584 223128
rect 300636 223116 300642 223168
rect 365714 223116 365720 223168
rect 365772 223156 365778 223168
rect 380158 223156 380164 223168
rect 365772 223128 380164 223156
rect 365772 223116 365778 223128
rect 380158 223116 380164 223128
rect 380216 223116 380222 223168
rect 384114 223116 384120 223168
rect 384172 223156 384178 223168
rect 408310 223156 408316 223168
rect 384172 223128 408316 223156
rect 384172 223116 384178 223128
rect 408310 223116 408316 223128
rect 408368 223116 408374 223168
rect 417234 223116 417240 223168
rect 417292 223156 417298 223168
rect 456886 223156 456892 223168
rect 417292 223128 456892 223156
rect 417292 223116 417298 223128
rect 456886 223116 456892 223128
rect 456944 223116 456950 223168
rect 460474 223116 460480 223168
rect 460532 223156 460538 223168
rect 523218 223156 523224 223168
rect 460532 223128 523224 223156
rect 460532 223116 460538 223128
rect 523218 223116 523224 223128
rect 523276 223116 523282 223168
rect 523678 223116 523684 223168
rect 523736 223156 523742 223168
rect 529014 223156 529020 223168
rect 523736 223128 529020 223156
rect 523736 223116 523742 223128
rect 529014 223116 529020 223128
rect 529072 223116 529078 223168
rect 529198 223116 529204 223168
rect 529256 223156 529262 223168
rect 539226 223156 539232 223168
rect 529256 223128 539232 223156
rect 529256 223116 529262 223128
rect 539226 223116 539232 223128
rect 539284 223116 539290 223168
rect 548334 223116 548340 223168
rect 548392 223156 548398 223168
rect 549070 223156 549076 223168
rect 548392 223128 549076 223156
rect 548392 223116 548398 223128
rect 549070 223116 549076 223128
rect 549128 223116 549134 223168
rect 550634 223116 550640 223168
rect 550692 223156 550698 223168
rect 558196 223156 558224 223264
rect 576826 223156 576854 223264
rect 550692 223128 558224 223156
rect 558288 223128 572714 223156
rect 576826 223128 605834 223156
rect 550692 223116 550698 223128
rect 160664 223060 161336 223088
rect 42610 222980 42616 223032
rect 42668 223020 42674 223032
rect 62758 223020 62764 223032
rect 42668 222992 62764 223020
rect 42668 222980 42674 222992
rect 62758 222980 62764 222992
rect 62816 222980 62822 223032
rect 75546 222980 75552 223032
rect 75604 223020 75610 223032
rect 152274 223020 152280 223032
rect 75604 222992 152280 223020
rect 75604 222980 75610 222992
rect 152274 222980 152280 222992
rect 152332 222980 152338 223032
rect 152458 222980 152464 223032
rect 152516 223020 152522 223032
rect 156414 223020 156420 223032
rect 152516 222992 156420 223020
rect 152516 222980 152522 222992
rect 156414 222980 156420 222992
rect 156472 222980 156478 223032
rect 160664 223020 160692 223060
rect 156616 222992 160692 223020
rect 62022 222844 62028 222896
rect 62080 222884 62086 222896
rect 146662 222884 146668 222896
rect 62080 222856 146668 222884
rect 62080 222844 62086 222856
rect 146662 222844 146668 222856
rect 146720 222844 146726 222896
rect 146938 222844 146944 222896
rect 146996 222884 147002 222896
rect 156616 222884 156644 222992
rect 161474 222980 161480 223032
rect 161532 223020 161538 223032
rect 171594 223020 171600 223032
rect 161532 222992 171600 223020
rect 161532 222980 161538 222992
rect 171594 222980 171600 222992
rect 171652 222980 171658 223032
rect 171778 222980 171784 223032
rect 171836 223020 171842 223032
rect 176194 223020 176200 223032
rect 171836 222992 176200 223020
rect 171836 222980 171842 222992
rect 176194 222980 176200 222992
rect 176252 222980 176258 223032
rect 177942 222980 177948 223032
rect 178000 223020 178006 223032
rect 228082 223020 228088 223032
rect 178000 222992 228088 223020
rect 178000 222980 178006 222992
rect 228082 222980 228088 222992
rect 228140 222980 228146 223032
rect 233050 222980 233056 223032
rect 233108 223020 233114 223032
rect 265066 223020 265072 223032
rect 233108 222992 265072 223020
rect 233108 222980 233114 222992
rect 265066 222980 265072 222992
rect 265124 222980 265130 223032
rect 271782 222980 271788 223032
rect 271840 223020 271846 223032
rect 292666 223020 292672 223032
rect 271840 222992 292672 223020
rect 271840 222980 271846 222992
rect 292666 222980 292672 222992
rect 292724 222980 292730 223032
rect 300578 222980 300584 223032
rect 300636 223020 300642 223032
rect 312538 223020 312544 223032
rect 300636 222992 312544 223020
rect 300636 222980 300642 222992
rect 312538 222980 312544 222992
rect 312596 222980 312602 223032
rect 353938 222980 353944 223032
rect 353996 223020 354002 223032
rect 366082 223020 366088 223032
rect 353996 222992 366088 223020
rect 353996 222980 354002 222992
rect 366082 222980 366088 222992
rect 366140 222980 366146 223032
rect 376018 222980 376024 223032
rect 376076 223020 376082 223032
rect 399202 223020 399208 223032
rect 376076 222992 399208 223020
rect 376076 222980 376082 222992
rect 399202 222980 399208 222992
rect 399260 222980 399266 223032
rect 404630 222980 404636 223032
rect 404688 223020 404694 223032
rect 428182 223020 428188 223032
rect 404688 222992 428188 223020
rect 404688 222980 404694 222992
rect 428182 222980 428188 222992
rect 428240 222980 428246 223032
rect 430666 222980 430672 223032
rect 430724 223020 430730 223032
rect 471422 223020 471428 223032
rect 430724 222992 471428 223020
rect 430724 222980 430730 222992
rect 471422 222980 471428 222992
rect 471480 222980 471486 223032
rect 478690 222980 478696 223032
rect 478748 223020 478754 223032
rect 483014 223020 483020 223032
rect 478748 222992 483020 223020
rect 478748 222980 478754 222992
rect 483014 222980 483020 222992
rect 483072 222980 483078 223032
rect 484118 222980 484124 223032
rect 484176 223020 484182 223032
rect 551554 223020 551560 223032
rect 484176 222992 551560 223020
rect 484176 222980 484182 222992
rect 551554 222980 551560 222992
rect 551612 222980 551618 223032
rect 551738 222980 551744 223032
rect 551796 223020 551802 223032
rect 558288 223020 558316 223128
rect 551796 222992 558316 223020
rect 551796 222980 551802 222992
rect 558546 222980 558552 223032
rect 558604 223020 558610 223032
rect 567746 223020 567752 223032
rect 558604 222992 567752 223020
rect 558604 222980 558610 222992
rect 567746 222980 567752 222992
rect 567804 222980 567810 223032
rect 571426 223020 571432 223032
rect 567948 222992 571432 223020
rect 146996 222856 156644 222884
rect 146996 222844 147002 222856
rect 156782 222844 156788 222896
rect 156840 222884 156846 222896
rect 213178 222884 213184 222896
rect 156840 222856 213184 222884
rect 156840 222844 156846 222856
rect 213178 222844 213184 222856
rect 213236 222844 213242 222896
rect 215938 222844 215944 222896
rect 215996 222884 216002 222896
rect 220262 222884 220268 222896
rect 215996 222856 220268 222884
rect 215996 222844 216002 222856
rect 220262 222844 220268 222856
rect 220320 222844 220326 222896
rect 221274 222844 221280 222896
rect 221332 222884 221338 222896
rect 259546 222884 259552 222896
rect 221332 222856 259552 222884
rect 221332 222844 221338 222856
rect 259546 222844 259552 222856
rect 259604 222844 259610 222896
rect 261846 222844 261852 222896
rect 261904 222884 261910 222896
rect 286042 222884 286048 222896
rect 261904 222856 286048 222884
rect 261904 222844 261910 222856
rect 286042 222844 286048 222856
rect 286100 222844 286106 222896
rect 293218 222844 293224 222896
rect 293276 222884 293282 222896
rect 306098 222884 306104 222896
rect 293276 222856 306104 222884
rect 293276 222844 293282 222856
rect 306098 222844 306104 222856
rect 306156 222844 306162 222896
rect 362678 222844 362684 222896
rect 362736 222884 362742 222896
rect 376018 222884 376024 222896
rect 362736 222856 376024 222884
rect 362736 222844 362742 222856
rect 376018 222844 376024 222856
rect 376076 222844 376082 222896
rect 380434 222844 380440 222896
rect 380492 222884 380498 222896
rect 405826 222884 405832 222896
rect 380492 222856 405832 222884
rect 380492 222844 380498 222856
rect 405826 222844 405832 222856
rect 405884 222844 405890 222896
rect 412450 222844 412456 222896
rect 412508 222884 412514 222896
rect 451458 222884 451464 222896
rect 412508 222856 451464 222884
rect 412508 222844 412514 222856
rect 451458 222844 451464 222856
rect 451516 222844 451522 222896
rect 471974 222844 471980 222896
rect 472032 222884 472038 222896
rect 544194 222884 544200 222896
rect 472032 222856 544200 222884
rect 472032 222844 472038 222856
rect 544194 222844 544200 222856
rect 544252 222844 544258 222896
rect 554038 222884 554044 222896
rect 548536 222856 554044 222884
rect 128262 222708 128268 222760
rect 128320 222748 128326 222760
rect 194962 222748 194968 222760
rect 128320 222720 194968 222748
rect 128320 222708 128326 222720
rect 194962 222708 194968 222720
rect 195020 222708 195026 222760
rect 197262 222708 197268 222760
rect 197320 222748 197326 222760
rect 197320 222720 238754 222748
rect 197320 222708 197326 222720
rect 133138 222572 133144 222624
rect 133196 222612 133202 222624
rect 146938 222612 146944 222624
rect 133196 222584 146944 222612
rect 133196 222572 133202 222584
rect 146938 222572 146944 222584
rect 146996 222572 147002 222624
rect 147122 222572 147128 222624
rect 147180 222612 147186 222624
rect 151262 222612 151268 222624
rect 147180 222584 151268 222612
rect 147180 222572 147186 222584
rect 151262 222572 151268 222584
rect 151320 222572 151326 222624
rect 151446 222572 151452 222624
rect 151504 222612 151510 222624
rect 156414 222612 156420 222624
rect 151504 222584 156420 222612
rect 151504 222572 151510 222584
rect 156414 222572 156420 222584
rect 156472 222572 156478 222624
rect 156598 222572 156604 222624
rect 156656 222612 156662 222624
rect 208762 222612 208768 222624
rect 156656 222584 208768 222612
rect 156656 222572 156662 222584
rect 208762 222572 208768 222584
rect 208820 222572 208826 222624
rect 210326 222572 210332 222624
rect 210384 222612 210390 222624
rect 231946 222612 231952 222624
rect 210384 222584 231952 222612
rect 210384 222572 210390 222584
rect 231946 222572 231952 222584
rect 232004 222572 232010 222624
rect 238726 222612 238754 222720
rect 239306 222708 239312 222760
rect 239364 222748 239370 222760
rect 242434 222748 242440 222760
rect 239364 222720 242440 222748
rect 239364 222708 239370 222720
rect 242434 222708 242440 222720
rect 242492 222708 242498 222760
rect 242802 222708 242808 222760
rect 242860 222748 242866 222760
rect 246666 222748 246672 222760
rect 242860 222720 246672 222748
rect 242860 222708 242866 222720
rect 246666 222708 246672 222720
rect 246724 222708 246730 222760
rect 408034 222708 408040 222760
rect 408092 222748 408098 222760
rect 444742 222748 444748 222760
rect 408092 222720 444748 222748
rect 408092 222708 408098 222720
rect 444742 222708 444748 222720
rect 444800 222708 444806 222760
rect 465810 222708 465816 222760
rect 465868 222748 465874 222760
rect 533522 222748 533528 222760
rect 465868 222720 533528 222748
rect 465868 222708 465874 222720
rect 533522 222708 533528 222720
rect 533580 222708 533586 222760
rect 533798 222708 533804 222760
rect 533856 222708 533862 222760
rect 534166 222708 534172 222760
rect 534224 222748 534230 222760
rect 548536 222748 548564 222856
rect 554038 222844 554044 222856
rect 554096 222844 554102 222896
rect 554682 222844 554688 222896
rect 554740 222884 554746 222896
rect 554740 222856 558500 222884
rect 554740 222844 554746 222856
rect 555418 222748 555424 222760
rect 534224 222720 548564 222748
rect 548628 222720 555424 222748
rect 534224 222708 534230 222720
rect 240962 222612 240968 222624
rect 238726 222584 240968 222612
rect 240962 222572 240968 222584
rect 241020 222572 241026 222624
rect 395246 222572 395252 222624
rect 395304 222612 395310 222624
rect 411622 222612 411628 222624
rect 395304 222584 411628 222612
rect 395304 222572 395310 222584
rect 411622 222572 411628 222584
rect 411680 222572 411686 222624
rect 425330 222572 425336 222624
rect 425388 222612 425394 222624
rect 459002 222612 459008 222624
rect 425388 222584 459008 222612
rect 425388 222572 425394 222584
rect 459002 222572 459008 222584
rect 459060 222572 459066 222624
rect 467466 222572 467472 222624
rect 467524 222612 467530 222624
rect 467524 222584 528876 222612
rect 467524 222572 467530 222584
rect 131022 222436 131028 222488
rect 131080 222476 131086 222488
rect 133782 222476 133788 222488
rect 131080 222448 133788 222476
rect 131080 222436 131086 222448
rect 133782 222436 133788 222448
rect 133840 222436 133846 222488
rect 137646 222436 137652 222488
rect 137704 222476 137710 222488
rect 201586 222476 201592 222488
rect 137704 222448 201592 222476
rect 137704 222436 137710 222448
rect 201586 222436 201592 222448
rect 201644 222436 201650 222488
rect 205634 222436 205640 222488
rect 205692 222476 205698 222488
rect 215662 222476 215668 222488
rect 205692 222448 215668 222476
rect 205692 222436 205698 222448
rect 215662 222436 215668 222448
rect 215720 222436 215726 222488
rect 427722 222436 427728 222488
rect 427780 222476 427786 222488
rect 460198 222476 460204 222488
rect 427780 222448 460204 222476
rect 427780 222436 427786 222448
rect 460198 222436 460204 222448
rect 460256 222436 460262 222488
rect 461946 222436 461952 222488
rect 462004 222476 462010 222488
rect 524874 222476 524880 222488
rect 462004 222448 524880 222476
rect 462004 222436 462010 222448
rect 524874 222436 524880 222448
rect 524932 222436 524938 222488
rect 528848 222476 528876 222584
rect 529014 222572 529020 222624
rect 529072 222612 529078 222624
rect 533816 222612 533844 222708
rect 548628 222612 548656 222720
rect 555418 222708 555424 222720
rect 555476 222708 555482 222760
rect 558472 222748 558500 222856
rect 559558 222844 559564 222896
rect 559616 222884 559622 222896
rect 567948 222884 567976 222992
rect 571426 222980 571432 222992
rect 571484 222980 571490 223032
rect 572686 223020 572714 223128
rect 605806 223020 605834 223128
rect 620462 223020 620468 223032
rect 572686 222992 601694 223020
rect 605806 222992 620468 223020
rect 559616 222856 567976 222884
rect 559616 222844 559622 222856
rect 568114 222844 568120 222896
rect 568172 222884 568178 222896
rect 596818 222884 596824 222896
rect 568172 222856 596824 222884
rect 568172 222844 568178 222856
rect 596818 222844 596824 222856
rect 596876 222844 596882 222896
rect 601666 222884 601694 222992
rect 620462 222980 620468 222992
rect 620520 222980 620526 223032
rect 619174 222884 619180 222896
rect 601666 222856 619180 222884
rect 619174 222844 619180 222856
rect 619232 222844 619238 222896
rect 620278 222844 620284 222896
rect 620336 222884 620342 222896
rect 625338 222884 625344 222896
rect 620336 222856 625344 222884
rect 620336 222844 620342 222856
rect 625338 222844 625344 222856
rect 625396 222844 625402 222896
rect 664622 222844 664628 222896
rect 664680 222884 664686 222896
rect 675478 222884 675484 222896
rect 664680 222856 675484 222884
rect 664680 222844 664686 222856
rect 675478 222844 675484 222856
rect 675536 222844 675542 222896
rect 630950 222748 630956 222760
rect 558472 222720 630956 222748
rect 630950 222708 630956 222720
rect 631008 222708 631014 222760
rect 664806 222708 664812 222760
rect 664864 222748 664870 222760
rect 675294 222748 675300 222760
rect 664864 222720 675300 222748
rect 664864 222708 664870 222720
rect 675294 222708 675300 222720
rect 675352 222708 675358 222760
rect 596634 222612 596640 222624
rect 529072 222584 533844 222612
rect 543706 222584 548656 222612
rect 548720 222584 596640 222612
rect 529072 222572 529078 222584
rect 536098 222504 536104 222556
rect 536156 222544 536162 222556
rect 543706 222544 543734 222584
rect 536156 222516 543734 222544
rect 536156 222504 536162 222516
rect 533522 222476 533528 222488
rect 528848 222448 533528 222476
rect 533522 222436 533528 222448
rect 533580 222436 533586 222488
rect 526714 222408 526720 222420
rect 525076 222380 526720 222408
rect 88978 222300 88984 222352
rect 89036 222340 89042 222352
rect 148870 222340 148876 222352
rect 89036 222312 148876 222340
rect 89036 222300 89042 222312
rect 148870 222300 148876 222312
rect 148928 222300 148934 222352
rect 151768 222300 151774 222352
rect 151826 222340 151832 222352
rect 156598 222340 156604 222352
rect 151826 222312 156604 222340
rect 151826 222300 151832 222312
rect 156598 222300 156604 222312
rect 156656 222300 156662 222352
rect 158990 222300 158996 222352
rect 159048 222340 159054 222352
rect 161290 222340 161296 222352
rect 159048 222312 161296 222340
rect 159048 222300 159054 222312
rect 161290 222300 161296 222312
rect 161348 222300 161354 222352
rect 161428 222300 161434 222352
rect 161486 222340 161492 222352
rect 209866 222340 209872 222352
rect 161486 222312 209872 222340
rect 161486 222300 161492 222312
rect 209866 222300 209872 222312
rect 209924 222300 209930 222352
rect 459186 222300 459192 222352
rect 459244 222340 459250 222352
rect 523034 222340 523040 222352
rect 459244 222312 523040 222340
rect 459244 222300 459250 222312
rect 523034 222300 523040 222312
rect 523092 222300 523098 222352
rect 523218 222300 523224 222352
rect 523276 222340 523282 222352
rect 525076 222340 525104 222380
rect 526714 222368 526720 222380
rect 526772 222368 526778 222420
rect 527634 222368 527640 222420
rect 527692 222408 527698 222420
rect 528462 222408 528468 222420
rect 527692 222380 528468 222408
rect 527692 222368 527698 222380
rect 528462 222368 528468 222380
rect 528520 222368 528526 222420
rect 533982 222368 533988 222420
rect 534040 222408 534046 222420
rect 548720 222408 548748 222584
rect 596634 222572 596640 222584
rect 596692 222572 596698 222624
rect 596818 222572 596824 222624
rect 596876 222612 596882 222624
rect 618714 222612 618720 222624
rect 596876 222584 618720 222612
rect 596876 222572 596882 222584
rect 618714 222572 618720 222584
rect 618772 222572 618778 222624
rect 619174 222572 619180 222624
rect 619232 222612 619238 222624
rect 629294 222612 629300 222624
rect 619232 222584 629300 222612
rect 619232 222572 619238 222584
rect 629294 222572 629300 222584
rect 629352 222572 629358 222624
rect 661678 222572 661684 222624
rect 661736 222612 661742 222624
rect 661736 222584 663794 222612
rect 661736 222572 661742 222584
rect 620278 222476 620284 222488
rect 563026 222448 620284 222476
rect 534040 222380 548748 222408
rect 534040 222368 534046 222380
rect 549898 222368 549904 222420
rect 549956 222408 549962 222420
rect 563026 222408 563054 222448
rect 620278 222436 620284 222448
rect 620336 222436 620342 222488
rect 620462 222436 620468 222488
rect 620520 222476 620526 222488
rect 631226 222476 631232 222488
rect 620520 222448 631232 222476
rect 620520 222436 620526 222448
rect 631226 222436 631232 222448
rect 631284 222436 631290 222488
rect 663766 222476 663794 222584
rect 668394 222572 668400 222624
rect 668452 222612 668458 222624
rect 675110 222612 675116 222624
rect 668452 222584 675116 222612
rect 668452 222572 668458 222584
rect 675110 222572 675116 222584
rect 675168 222572 675174 222624
rect 663766 222448 668716 222476
rect 549956 222380 563054 222408
rect 549956 222368 549962 222380
rect 523276 222312 525104 222340
rect 523276 222300 523282 222312
rect 597002 222300 597008 222352
rect 597060 222340 597066 222352
rect 619726 222340 619732 222352
rect 597060 222312 619732 222340
rect 597060 222300 597066 222312
rect 619726 222300 619732 222312
rect 619784 222300 619790 222352
rect 416038 222232 416044 222284
rect 416096 222272 416102 222284
rect 416096 222244 416820 222272
rect 416096 222232 416102 222244
rect 91278 222096 91284 222148
rect 91336 222136 91342 222148
rect 161566 222136 161572 222148
rect 91336 222108 161572 222136
rect 91336 222096 91342 222108
rect 161566 222096 161572 222108
rect 161624 222096 161630 222148
rect 161750 222096 161756 222148
rect 161808 222136 161814 222148
rect 167638 222136 167644 222148
rect 161808 222108 167644 222136
rect 161808 222096 161814 222108
rect 167638 222096 167644 222108
rect 167696 222096 167702 222148
rect 171594 222096 171600 222148
rect 171652 222136 171658 222148
rect 179690 222136 179696 222148
rect 171652 222108 179696 222136
rect 171652 222096 171658 222108
rect 179690 222096 179696 222108
rect 179748 222096 179754 222148
rect 184658 222096 184664 222148
rect 184716 222136 184722 222148
rect 234982 222136 234988 222148
rect 184716 222108 234988 222136
rect 184716 222096 184722 222108
rect 234982 222096 234988 222108
rect 235040 222096 235046 222148
rect 258166 222096 258172 222148
rect 258224 222136 258230 222148
rect 261018 222136 261024 222148
rect 258224 222108 261024 222136
rect 258224 222096 258230 222108
rect 261018 222096 261024 222108
rect 261076 222096 261082 222148
rect 265986 222096 265992 222148
rect 266044 222136 266050 222148
rect 266998 222136 267004 222148
rect 266044 222108 267004 222136
rect 266044 222096 266050 222108
rect 266998 222096 267004 222108
rect 267056 222096 267062 222148
rect 377398 222096 377404 222148
rect 377456 222136 377462 222148
rect 393406 222136 393412 222148
rect 377456 222108 393412 222136
rect 377456 222096 377462 222108
rect 393406 222096 393412 222108
rect 393464 222096 393470 222148
rect 393958 222096 393964 222148
rect 394016 222136 394022 222148
rect 416590 222136 416596 222148
rect 394016 222108 416596 222136
rect 394016 222096 394022 222108
rect 416590 222096 416596 222108
rect 416648 222096 416654 222148
rect 416792 222136 416820 222244
rect 525168 222244 596864 222272
rect 509252 222176 509372 222204
rect 429746 222136 429752 222148
rect 416792 222108 429752 222136
rect 429746 222096 429752 222108
rect 429804 222096 429810 222148
rect 452562 222096 452568 222148
rect 452620 222136 452626 222148
rect 509252 222136 509280 222176
rect 452620 222108 509280 222136
rect 452620 222096 452626 222108
rect 79686 222028 79692 222080
rect 79744 222068 79750 222080
rect 509344 222068 509372 222176
rect 511258 222164 511264 222216
rect 511316 222204 511322 222216
rect 523678 222204 523684 222216
rect 511316 222176 523684 222204
rect 511316 222164 511322 222176
rect 523678 222164 523684 222176
rect 523736 222164 523742 222216
rect 523862 222164 523868 222216
rect 523920 222204 523926 222216
rect 525168 222204 525196 222244
rect 523920 222176 525196 222204
rect 596836 222204 596864 222244
rect 618346 222204 618352 222216
rect 596836 222176 618352 222204
rect 523920 222164 523926 222176
rect 618346 222164 618352 222176
rect 618404 222164 618410 222216
rect 618714 222164 618720 222216
rect 618772 222204 618778 222216
rect 619910 222204 619916 222216
rect 618772 222176 619916 222204
rect 618772 222164 618778 222176
rect 619910 222164 619916 222176
rect 619968 222164 619974 222216
rect 663058 222164 663064 222216
rect 663116 222204 663122 222216
rect 668394 222204 668400 222216
rect 663116 222176 668400 222204
rect 663116 222164 663122 222176
rect 668394 222164 668400 222176
rect 668452 222164 668458 222216
rect 668688 222204 668716 222448
rect 675478 222204 675484 222216
rect 668688 222176 675484 222204
rect 675478 222164 675484 222176
rect 675536 222164 675542 222216
rect 529382 222096 529388 222148
rect 529440 222136 529446 222148
rect 553302 222136 553308 222148
rect 529440 222108 553308 222136
rect 529440 222096 529446 222108
rect 553302 222096 553308 222108
rect 553360 222096 553366 222148
rect 555970 222096 555976 222148
rect 556028 222136 556034 222148
rect 565722 222136 565728 222148
rect 556028 222108 565728 222136
rect 556028 222096 556034 222108
rect 565722 222096 565728 222108
rect 565780 222136 565786 222148
rect 567654 222136 567660 222148
rect 565780 222108 567660 222136
rect 565780 222096 565786 222108
rect 567654 222096 567660 222108
rect 567712 222096 567718 222148
rect 567838 222096 567844 222148
rect 567896 222136 567902 222148
rect 591298 222136 591304 222148
rect 567896 222108 591304 222136
rect 567896 222096 567902 222108
rect 591298 222096 591304 222108
rect 591356 222096 591362 222148
rect 591482 222096 591488 222148
rect 591540 222136 591546 222148
rect 591540 222108 592172 222136
rect 591540 222096 591546 222108
rect 514294 222068 514300 222080
rect 79744 222040 84194 222068
rect 509344 222040 514300 222068
rect 79744 222028 79750 222040
rect 80514 221892 80520 221944
rect 80572 221932 80578 221944
rect 83458 221932 83464 221944
rect 80572 221904 83464 221932
rect 80572 221892 80578 221904
rect 83458 221892 83464 221904
rect 83516 221892 83522 221944
rect 84166 221864 84194 222040
rect 514294 222028 514300 222040
rect 514352 222028 514358 222080
rect 517790 222028 517796 222080
rect 517848 222068 517854 222080
rect 518434 222068 518440 222080
rect 517848 222040 518440 222068
rect 517848 222028 517854 222040
rect 518434 222028 518440 222040
rect 518492 222068 518498 222080
rect 592144 222068 592172 222108
rect 597830 222068 597836 222080
rect 518492 222040 529244 222068
rect 592144 222040 597836 222068
rect 518492 222028 518498 222040
rect 88794 221960 88800 222012
rect 88852 222000 88858 222012
rect 156598 222000 156604 222012
rect 88852 221972 156604 222000
rect 88852 221960 88858 221972
rect 156598 221960 156604 221972
rect 156656 221960 156662 222012
rect 156782 221960 156788 222012
rect 156840 222000 156846 222012
rect 178126 222000 178132 222012
rect 156840 221972 178132 222000
rect 156840 221960 156846 221972
rect 178126 221960 178132 221972
rect 178184 221960 178190 222012
rect 180058 221960 180064 222012
rect 180116 222000 180122 222012
rect 230474 222000 230480 222012
rect 180116 221972 230480 222000
rect 180116 221960 180122 221972
rect 230474 221960 230480 221972
rect 230532 221960 230538 222012
rect 251910 221960 251916 222012
rect 251968 222000 251974 222012
rect 278038 222000 278044 222012
rect 251968 221972 278044 222000
rect 251968 221960 251974 221972
rect 278038 221960 278044 221972
rect 278096 221960 278102 222012
rect 280890 221960 280896 222012
rect 280948 222000 280954 222012
rect 297358 222000 297364 222012
rect 280948 221972 297364 222000
rect 280948 221960 280954 221972
rect 297358 221960 297364 221972
rect 297416 221960 297422 222012
rect 369762 221960 369768 222012
rect 369820 222000 369826 222012
rect 387610 222000 387616 222012
rect 369820 221972 387616 222000
rect 369820 221960 369826 221972
rect 387610 221960 387616 221972
rect 387668 221960 387674 222012
rect 396902 221960 396908 222012
rect 396960 222000 396966 222012
rect 419902 222000 419908 222012
rect 396960 221972 419908 222000
rect 396960 221960 396966 221972
rect 419902 221960 419908 221972
rect 419960 221960 419966 222012
rect 424318 221960 424324 222012
rect 424376 222000 424382 222012
rect 443086 222000 443092 222012
rect 424376 221972 443092 222000
rect 424376 221960 424382 221972
rect 443086 221960 443092 221972
rect 443144 221960 443150 222012
rect 449894 221960 449900 222012
rect 449952 222000 449958 222012
rect 509188 222000 509194 222012
rect 449952 221972 509194 222000
rect 449952 221960 449958 221972
rect 509188 221960 509194 221972
rect 509246 221960 509252 222012
rect 529216 222000 529244 222040
rect 597830 222028 597836 222040
rect 597888 222028 597894 222080
rect 591988 222000 591994 222012
rect 529216 221972 591994 222000
rect 591988 221960 591994 221972
rect 592046 221960 592052 222012
rect 524064 221904 524414 221932
rect 84166 221836 89116 221864
rect 73890 221688 73896 221740
rect 73948 221728 73954 221740
rect 77938 221728 77944 221740
rect 73948 221700 77944 221728
rect 73948 221688 73954 221700
rect 77938 221688 77944 221700
rect 77996 221688 78002 221740
rect 79318 221728 79324 221740
rect 78140 221700 79324 221728
rect 60642 221552 60648 221604
rect 60700 221592 60706 221604
rect 78140 221592 78168 221700
rect 79318 221688 79324 221700
rect 79376 221688 79382 221740
rect 82998 221688 83004 221740
rect 83056 221728 83062 221740
rect 88794 221728 88800 221740
rect 83056 221700 88800 221728
rect 83056 221688 83062 221700
rect 88794 221688 88800 221700
rect 88852 221688 88858 221740
rect 89088 221728 89116 221836
rect 89254 221824 89260 221876
rect 89312 221864 89318 221876
rect 161428 221864 161434 221876
rect 89312 221836 161434 221864
rect 89312 221824 89318 221836
rect 161428 221824 161434 221836
rect 161486 221824 161492 221876
rect 161566 221824 161572 221876
rect 161624 221864 161630 221876
rect 164418 221864 164424 221876
rect 161624 221836 164424 221864
rect 161624 221824 161630 221836
rect 164418 221824 164424 221836
rect 164476 221824 164482 221876
rect 164602 221824 164608 221876
rect 164660 221864 164666 221876
rect 170398 221864 170404 221876
rect 164660 221836 170404 221864
rect 164660 221824 164666 221836
rect 170398 221824 170404 221836
rect 170456 221824 170462 221876
rect 170766 221824 170772 221876
rect 170824 221864 170830 221876
rect 173710 221864 173716 221876
rect 170824 221836 173716 221864
rect 170824 221824 170830 221836
rect 173710 221824 173716 221836
rect 173768 221824 173774 221876
rect 173894 221824 173900 221876
rect 173952 221864 173958 221876
rect 174722 221864 174728 221876
rect 173952 221836 174728 221864
rect 173952 221824 173958 221836
rect 174722 221824 174728 221836
rect 174780 221824 174786 221876
rect 174906 221824 174912 221876
rect 174964 221864 174970 221876
rect 223942 221864 223948 221876
rect 174964 221836 223948 221864
rect 174964 221824 174970 221836
rect 223942 221824 223948 221836
rect 224000 221824 224006 221876
rect 227070 221824 227076 221876
rect 227128 221864 227134 221876
rect 258166 221864 258172 221876
rect 227128 221836 258172 221864
rect 227128 221824 227134 221836
rect 258166 221824 258172 221836
rect 258224 221824 258230 221876
rect 258626 221864 258632 221876
rect 258368 221836 258632 221864
rect 151906 221728 151912 221740
rect 89088 221700 151912 221728
rect 151906 221688 151912 221700
rect 151964 221688 151970 221740
rect 152274 221688 152280 221740
rect 152332 221728 152338 221740
rect 156414 221728 156420 221740
rect 152332 221700 156420 221728
rect 152332 221688 152338 221700
rect 156414 221688 156420 221700
rect 156472 221688 156478 221740
rect 156598 221688 156604 221740
rect 156656 221728 156662 221740
rect 163590 221728 163596 221740
rect 156656 221700 163596 221728
rect 156656 221688 156662 221700
rect 163590 221688 163596 221700
rect 163648 221688 163654 221740
rect 164050 221688 164056 221740
rect 164108 221728 164114 221740
rect 218882 221728 218888 221740
rect 164108 221700 218888 221728
rect 164108 221688 164114 221700
rect 218882 221688 218888 221700
rect 218940 221688 218946 221740
rect 223758 221688 223764 221740
rect 223816 221728 223822 221740
rect 258368 221728 258396 221836
rect 258626 221824 258632 221836
rect 258684 221824 258690 221876
rect 263502 221824 263508 221876
rect 263560 221864 263566 221876
rect 285122 221864 285128 221876
rect 263560 221836 285128 221864
rect 263560 221824 263566 221836
rect 285122 221824 285128 221836
rect 285180 221824 285186 221876
rect 351546 221824 351552 221876
rect 351604 221864 351610 221876
rect 361206 221864 361212 221876
rect 351604 221836 361212 221864
rect 351604 221824 351610 221836
rect 361206 221824 361212 221836
rect 361264 221824 361270 221876
rect 372062 221824 372068 221876
rect 372120 221864 372126 221876
rect 390922 221864 390928 221876
rect 372120 221836 390928 221864
rect 372120 221824 372126 221836
rect 390922 221824 390928 221836
rect 390980 221824 390986 221876
rect 397362 221824 397368 221876
rect 397420 221864 397426 221876
rect 426526 221864 426532 221876
rect 397420 221836 426532 221864
rect 397420 221824 397426 221836
rect 426526 221824 426532 221836
rect 426584 221824 426590 221876
rect 427078 221824 427084 221876
rect 427136 221864 427142 221876
rect 456334 221864 456340 221876
rect 427136 221836 456340 221864
rect 427136 221824 427142 221836
rect 456334 221824 456340 221836
rect 456392 221824 456398 221876
rect 456702 221824 456708 221876
rect 456760 221864 456766 221876
rect 519262 221864 519268 221876
rect 456760 221836 519268 221864
rect 456760 221824 456766 221836
rect 519262 221824 519268 221836
rect 519320 221824 519326 221876
rect 520918 221824 520924 221876
rect 520976 221864 520982 221876
rect 520976 221836 522436 221864
rect 520976 221824 520982 221836
rect 223816 221700 258396 221728
rect 223816 221688 223822 221700
rect 258534 221688 258540 221740
rect 258592 221728 258598 221740
rect 282454 221728 282460 221740
rect 258592 221700 282460 221728
rect 258592 221688 258598 221700
rect 282454 221688 282460 221700
rect 282512 221688 282518 221740
rect 298462 221728 298468 221740
rect 296686 221700 298468 221728
rect 60700 221564 78168 221592
rect 60700 221552 60706 221564
rect 78858 221552 78864 221604
rect 78916 221592 78922 221604
rect 161428 221592 161434 221604
rect 78916 221564 161434 221592
rect 78916 221552 78922 221564
rect 161428 221552 161434 221564
rect 161486 221552 161492 221604
rect 161566 221552 161572 221604
rect 161624 221592 161630 221604
rect 171778 221592 171784 221604
rect 161624 221564 171784 221592
rect 161624 221552 161630 221564
rect 171778 221552 171784 221564
rect 171836 221552 171842 221604
rect 171962 221552 171968 221604
rect 172020 221592 172026 221604
rect 226426 221592 226432 221604
rect 172020 221564 226432 221592
rect 172020 221552 172026 221564
rect 226426 221552 226432 221564
rect 226484 221552 226490 221604
rect 227898 221552 227904 221604
rect 227956 221592 227962 221604
rect 263778 221592 263784 221604
rect 227956 221564 263784 221592
rect 227956 221552 227962 221564
rect 263778 221552 263784 221564
rect 263836 221552 263842 221604
rect 278406 221552 278412 221604
rect 278464 221592 278470 221604
rect 295702 221592 295708 221604
rect 278464 221564 295708 221592
rect 278464 221552 278470 221564
rect 295702 221552 295708 221564
rect 295760 221552 295766 221604
rect 59354 221416 59360 221468
rect 59412 221456 59418 221468
rect 147030 221456 147036 221468
rect 59412 221428 147036 221456
rect 59412 221416 59418 221428
rect 147030 221416 147036 221428
rect 147088 221416 147094 221468
rect 147214 221416 147220 221468
rect 147272 221456 147278 221468
rect 150710 221456 150716 221468
rect 147272 221428 150716 221456
rect 147272 221416 147278 221428
rect 150710 221416 150716 221428
rect 150768 221416 150774 221468
rect 150894 221416 150900 221468
rect 150952 221456 150958 221468
rect 150952 221428 196204 221456
rect 150952 221416 150958 221428
rect 196176 221388 196204 221428
rect 197722 221416 197728 221468
rect 197780 221456 197786 221468
rect 214006 221456 214012 221468
rect 197780 221428 214012 221456
rect 197780 221416 197786 221428
rect 214006 221416 214012 221428
rect 214064 221416 214070 221468
rect 220630 221416 220636 221468
rect 220688 221456 220694 221468
rect 256786 221456 256792 221468
rect 220688 221428 256792 221456
rect 220688 221416 220694 221428
rect 256786 221416 256792 221428
rect 256844 221416 256850 221468
rect 257706 221416 257712 221468
rect 257764 221456 257770 221468
rect 283190 221456 283196 221468
rect 257764 221428 283196 221456
rect 257764 221416 257770 221428
rect 283190 221416 283196 221428
rect 283248 221416 283254 221468
rect 283374 221416 283380 221468
rect 283432 221456 283438 221468
rect 296686 221456 296714 221700
rect 298462 221688 298468 221700
rect 298520 221688 298526 221740
rect 303246 221688 303252 221740
rect 303304 221728 303310 221740
rect 311986 221728 311992 221740
rect 303304 221700 311992 221728
rect 303304 221688 303310 221700
rect 311986 221688 311992 221700
rect 312044 221688 312050 221740
rect 357342 221688 357348 221740
rect 357400 221728 357406 221740
rect 369394 221728 369400 221740
rect 357400 221700 369400 221728
rect 357400 221688 357406 221700
rect 369394 221688 369400 221700
rect 369452 221688 369458 221740
rect 379974 221688 379980 221740
rect 380032 221728 380038 221740
rect 400030 221728 400036 221740
rect 380032 221700 400036 221728
rect 380032 221688 380038 221700
rect 400030 221688 400036 221700
rect 400088 221688 400094 221740
rect 404262 221688 404268 221740
rect 404320 221728 404326 221740
rect 436462 221728 436468 221740
rect 404320 221700 436468 221728
rect 404320 221688 404326 221700
rect 436462 221688 436468 221700
rect 436520 221688 436526 221740
rect 441522 221688 441528 221740
rect 441580 221728 441586 221740
rect 449894 221728 449900 221740
rect 441580 221700 449900 221728
rect 441580 221688 441586 221700
rect 449894 221688 449900 221700
rect 449952 221688 449958 221740
rect 458082 221688 458088 221740
rect 458140 221728 458146 221740
rect 521746 221728 521752 221740
rect 458140 221700 521752 221728
rect 458140 221688 458146 221700
rect 521746 221688 521752 221700
rect 521804 221688 521810 221740
rect 522408 221728 522436 221836
rect 522574 221824 522580 221876
rect 522632 221864 522638 221876
rect 523862 221864 523868 221876
rect 522632 221836 523868 221864
rect 522632 221824 522638 221836
rect 523862 221824 523868 221836
rect 523920 221824 523926 221876
rect 524064 221728 524092 221904
rect 524386 221864 524414 221904
rect 600314 221864 600320 221876
rect 524386 221836 600320 221864
rect 600314 221824 600320 221836
rect 600372 221824 600378 221876
rect 522408 221700 524092 221728
rect 529750 221688 529756 221740
rect 529808 221728 529814 221740
rect 602246 221728 602252 221740
rect 529808 221700 602252 221728
rect 529808 221688 529814 221700
rect 602246 221688 602252 221700
rect 602304 221688 602310 221740
rect 317414 221620 317420 221672
rect 317472 221660 317478 221672
rect 318794 221660 318800 221672
rect 317472 221632 318800 221660
rect 317472 221620 317478 221632
rect 318794 221620 318800 221632
rect 318852 221620 318858 221672
rect 296898 221552 296904 221604
rect 296956 221592 296962 221604
rect 301774 221592 301780 221604
rect 296956 221564 301780 221592
rect 296956 221552 296962 221564
rect 301774 221552 301780 221564
rect 301832 221552 301838 221604
rect 310054 221592 310060 221604
rect 301976 221564 310060 221592
rect 283432 221428 296714 221456
rect 283432 221416 283438 221428
rect 297450 221416 297456 221468
rect 297508 221456 297514 221468
rect 301976 221456 302004 221564
rect 310054 221552 310060 221564
rect 310112 221552 310118 221604
rect 344922 221552 344928 221604
rect 344980 221592 344986 221604
rect 348694 221592 348700 221604
rect 344980 221564 348700 221592
rect 344980 221552 344986 221564
rect 348694 221552 348700 221564
rect 348752 221552 348758 221604
rect 360010 221552 360016 221604
rect 360068 221592 360074 221604
rect 374362 221592 374368 221604
rect 360068 221564 374368 221592
rect 360068 221552 360074 221564
rect 374362 221552 374368 221564
rect 374420 221552 374426 221604
rect 383194 221552 383200 221604
rect 383252 221592 383258 221604
rect 406654 221592 406660 221604
rect 383252 221564 406660 221592
rect 383252 221552 383258 221564
rect 406654 221552 406660 221564
rect 406712 221552 406718 221604
rect 412266 221552 412272 221604
rect 412324 221592 412330 221604
rect 446950 221592 446956 221604
rect 412324 221564 446956 221592
rect 412324 221552 412330 221564
rect 446950 221552 446956 221564
rect 447008 221552 447014 221604
rect 486602 221552 486608 221604
rect 486660 221592 486666 221604
rect 555970 221592 555976 221604
rect 486660 221564 555976 221592
rect 486660 221552 486666 221564
rect 555970 221552 555976 221564
rect 556028 221552 556034 221604
rect 563238 221592 563244 221604
rect 556172 221564 563244 221592
rect 297508 221428 302004 221456
rect 297508 221416 297514 221428
rect 304902 221416 304908 221468
rect 304960 221456 304966 221468
rect 313642 221456 313648 221468
rect 304960 221428 313648 221456
rect 304960 221416 304966 221428
rect 313642 221416 313648 221428
rect 313700 221416 313706 221468
rect 315758 221416 315764 221468
rect 315816 221456 315822 221468
rect 320818 221456 320824 221468
rect 315816 221428 320824 221456
rect 315816 221416 315822 221428
rect 320818 221416 320824 221428
rect 320876 221416 320882 221468
rect 347590 221416 347596 221468
rect 347648 221456 347654 221468
rect 356146 221456 356152 221468
rect 347648 221428 356152 221456
rect 347648 221416 347654 221428
rect 356146 221416 356152 221428
rect 356204 221416 356210 221468
rect 368290 221416 368296 221468
rect 368348 221456 368354 221468
rect 385954 221456 385960 221468
rect 368348 221428 385960 221456
rect 368348 221416 368354 221428
rect 385954 221416 385960 221428
rect 386012 221416 386018 221468
rect 386322 221416 386328 221468
rect 386380 221456 386386 221468
rect 409966 221456 409972 221468
rect 386380 221428 409972 221456
rect 386380 221416 386386 221428
rect 409966 221416 409972 221428
rect 410024 221416 410030 221468
rect 422202 221416 422208 221468
rect 422260 221456 422266 221468
rect 464614 221456 464620 221468
rect 422260 221428 464620 221456
rect 422260 221416 422266 221428
rect 464614 221416 464620 221428
rect 464672 221416 464678 221468
rect 484486 221416 484492 221468
rect 484544 221456 484550 221468
rect 556172 221456 556200 221564
rect 563238 221552 563244 221564
rect 563296 221592 563302 221604
rect 563296 221564 568068 221592
rect 563296 221552 563302 221564
rect 484544 221428 556200 221456
rect 484544 221416 484550 221428
rect 556338 221416 556344 221468
rect 556396 221456 556402 221468
rect 567838 221456 567844 221468
rect 556396 221428 567844 221456
rect 556396 221416 556402 221428
rect 567838 221416 567844 221428
rect 567896 221416 567902 221468
rect 568040 221456 568068 221564
rect 568298 221552 568304 221604
rect 568356 221592 568362 221604
rect 611354 221592 611360 221604
rect 568356 221564 611360 221592
rect 568356 221552 568362 221564
rect 611354 221552 611360 221564
rect 611412 221552 611418 221604
rect 609974 221456 609980 221468
rect 568040 221428 609980 221456
rect 609974 221416 609980 221428
rect 610032 221416 610038 221468
rect 196176 221360 196296 221388
rect 87138 221280 87144 221332
rect 87196 221320 87202 221332
rect 90358 221320 90364 221332
rect 87196 221292 90364 221320
rect 87196 221280 87202 221292
rect 90358 221280 90364 221292
rect 90416 221280 90422 221332
rect 102042 221280 102048 221332
rect 102100 221320 102106 221332
rect 171594 221320 171600 221332
rect 102100 221292 171600 221320
rect 102100 221280 102106 221292
rect 171594 221280 171600 221292
rect 171652 221280 171658 221332
rect 171778 221280 171784 221332
rect 171836 221320 171842 221332
rect 195606 221320 195612 221332
rect 171836 221292 195612 221320
rect 171836 221280 171842 221292
rect 195606 221280 195612 221292
rect 195664 221280 195670 221332
rect 196268 221320 196296 221360
rect 210050 221320 210056 221332
rect 196268 221292 210056 221320
rect 210050 221280 210056 221292
rect 210108 221280 210114 221332
rect 211338 221280 211344 221332
rect 211396 221320 211402 221332
rect 252646 221320 252652 221332
rect 211396 221292 252652 221320
rect 211396 221280 211402 221292
rect 252646 221280 252652 221292
rect 252704 221280 252710 221332
rect 400858 221280 400864 221332
rect 400916 221320 400922 221332
rect 423214 221320 423220 221332
rect 400916 221292 423220 221320
rect 400916 221280 400922 221292
rect 423214 221280 423220 221292
rect 423272 221280 423278 221332
rect 428458 221280 428464 221332
rect 428516 221320 428522 221332
rect 439774 221320 439780 221332
rect 428516 221292 439780 221320
rect 428516 221280 428522 221292
rect 439774 221280 439780 221292
rect 439832 221280 439838 221332
rect 444926 221280 444932 221332
rect 444984 221320 444990 221332
rect 503530 221320 503536 221332
rect 444984 221292 503536 221320
rect 444984 221280 444990 221292
rect 503530 221280 503536 221292
rect 503588 221280 503594 221332
rect 504542 221280 504548 221332
rect 504600 221320 504606 221332
rect 529382 221320 529388 221332
rect 504600 221292 529388 221320
rect 504600 221280 504606 221292
rect 529382 221280 529388 221292
rect 529440 221280 529446 221332
rect 529566 221280 529572 221332
rect 529624 221320 529630 221332
rect 593966 221320 593972 221332
rect 529624 221292 593972 221320
rect 529624 221280 529630 221292
rect 593966 221280 593972 221292
rect 594024 221280 594030 221332
rect 195808 221224 196112 221252
rect 86310 221144 86316 221196
rect 86368 221184 86374 221196
rect 89254 221184 89260 221196
rect 86368 221156 89260 221184
rect 86368 221144 86374 221156
rect 89254 221144 89260 221156
rect 89312 221144 89318 221196
rect 97718 221144 97724 221196
rect 97776 221184 97782 221196
rect 173710 221184 173716 221196
rect 97776 221156 173716 221184
rect 97776 221144 97782 221156
rect 173710 221144 173716 221156
rect 173768 221144 173774 221196
rect 173894 221144 173900 221196
rect 173952 221184 173958 221196
rect 195808 221184 195836 221224
rect 173952 221156 195836 221184
rect 196084 221184 196112 221224
rect 594150 221212 594156 221264
rect 594208 221252 594214 221264
rect 601050 221252 601056 221264
rect 594208 221224 601056 221252
rect 594208 221212 594214 221224
rect 601050 221212 601056 221224
rect 601108 221212 601114 221264
rect 664254 221212 664260 221264
rect 664312 221252 664318 221264
rect 675478 221252 675484 221264
rect 664312 221224 675484 221252
rect 664312 221212 664318 221224
rect 675478 221212 675484 221224
rect 675536 221212 675542 221264
rect 222746 221184 222752 221196
rect 196084 221156 222752 221184
rect 173952 221144 173958 221156
rect 222746 221144 222752 221156
rect 222804 221144 222810 221196
rect 389726 221144 389732 221196
rect 389784 221184 389790 221196
rect 403342 221184 403348 221196
rect 389784 221156 403348 221184
rect 389784 221144 389790 221156
rect 403342 221144 403348 221156
rect 403400 221144 403406 221196
rect 409506 221144 409512 221196
rect 409564 221184 409570 221196
rect 422294 221184 422300 221196
rect 409564 221156 422300 221184
rect 409564 221144 409570 221156
rect 422294 221144 422300 221156
rect 422352 221144 422358 221196
rect 444282 221144 444288 221196
rect 444340 221184 444346 221196
rect 501046 221184 501052 221196
rect 444340 221156 501052 221184
rect 444340 221144 444346 221156
rect 501046 221144 501052 221156
rect 501104 221144 501110 221196
rect 509234 221144 509240 221196
rect 509292 221184 509298 221196
rect 511074 221184 511080 221196
rect 509292 221156 511080 221184
rect 509292 221144 509298 221156
rect 511074 221144 511080 221156
rect 511132 221144 511138 221196
rect 515950 221076 515956 221128
rect 516008 221116 516014 221128
rect 600866 221116 600872 221128
rect 516008 221088 600872 221116
rect 516008 221076 516014 221088
rect 600866 221076 600872 221088
rect 600924 221076 600930 221128
rect 104526 221008 104532 221060
rect 104584 221048 104590 221060
rect 179414 221048 179420 221060
rect 104584 221020 179420 221048
rect 104584 221008 104590 221020
rect 179414 221008 179420 221020
rect 179472 221008 179478 221060
rect 179874 221008 179880 221060
rect 179932 221048 179938 221060
rect 183462 221048 183468 221060
rect 179932 221020 183468 221048
rect 179932 221008 179938 221020
rect 183462 221008 183468 221020
rect 183520 221008 183526 221060
rect 186498 221008 186504 221060
rect 186556 221048 186562 221060
rect 194226 221048 194232 221060
rect 186556 221020 194232 221048
rect 186556 221008 186562 221020
rect 194226 221008 194232 221020
rect 194284 221008 194290 221060
rect 195606 221008 195612 221060
rect 195664 221048 195670 221060
rect 197722 221048 197728 221060
rect 195664 221020 197728 221048
rect 195664 221008 195670 221020
rect 197722 221008 197728 221020
rect 197780 221008 197786 221060
rect 213362 221008 213368 221060
rect 213420 221048 213426 221060
rect 252094 221048 252100 221060
rect 213420 221020 252100 221048
rect 213420 221008 213426 221020
rect 252094 221008 252100 221020
rect 252152 221008 252158 221060
rect 420178 221008 420184 221060
rect 420236 221048 420242 221060
rect 433150 221048 433156 221060
rect 420236 221020 433156 221048
rect 420236 221008 420242 221020
rect 433150 221008 433156 221020
rect 433208 221008 433214 221060
rect 439958 221008 439964 221060
rect 440016 221048 440022 221060
rect 491202 221048 491208 221060
rect 440016 221020 491208 221048
rect 440016 221008 440022 221020
rect 491202 221008 491208 221020
rect 491260 221008 491266 221060
rect 669038 221008 669044 221060
rect 669096 221048 669102 221060
rect 675478 221048 675484 221060
rect 669096 221020 675484 221048
rect 669096 221008 669102 221020
rect 675478 221008 675484 221020
rect 675536 221008 675542 221060
rect 513558 220940 513564 220992
rect 513616 220980 513622 220992
rect 598934 220980 598940 220992
rect 513616 220952 598940 220980
rect 513616 220940 513622 220952
rect 598934 220940 598940 220952
rect 598992 220940 598998 220992
rect 117774 220872 117780 220924
rect 117832 220912 117838 220924
rect 187970 220912 187976 220924
rect 117832 220884 187976 220912
rect 117832 220872 117838 220884
rect 187970 220872 187976 220884
rect 188028 220872 188034 220924
rect 253842 220872 253848 220924
rect 253900 220912 253906 220924
rect 259822 220912 259828 220924
rect 253900 220884 259828 220912
rect 253900 220872 253906 220884
rect 259822 220872 259828 220884
rect 259880 220872 259886 220924
rect 343450 220872 343456 220924
rect 343508 220912 343514 220924
rect 347038 220912 347044 220924
rect 343508 220884 347044 220912
rect 343508 220872 343514 220884
rect 347038 220872 347044 220884
rect 347096 220872 347102 220924
rect 463694 220872 463700 220924
rect 463752 220912 463758 220924
rect 508590 220912 508596 220924
rect 463752 220884 508596 220912
rect 463752 220872 463758 220884
rect 508590 220872 508596 220884
rect 508648 220912 508654 220924
rect 508648 220884 509234 220912
rect 508648 220872 508654 220884
rect 312998 220804 313004 220856
rect 313056 220844 313062 220856
rect 318242 220844 318248 220856
rect 313056 220816 318248 220844
rect 313056 220804 313062 220816
rect 318242 220804 318248 220816
rect 318300 220804 318306 220856
rect 320634 220804 320640 220856
rect 320692 220844 320698 220856
rect 325786 220844 325792 220856
rect 320692 220816 325792 220844
rect 320692 220804 320698 220816
rect 325786 220804 325792 220816
rect 325844 220804 325850 220856
rect 509206 220844 509234 220884
rect 591114 220844 591120 220856
rect 509206 220816 591120 220844
rect 591114 220804 591120 220816
rect 591172 220804 591178 220856
rect 591298 220804 591304 220856
rect 591356 220844 591362 220856
rect 607214 220844 607220 220856
rect 591356 220816 607220 220844
rect 591356 220804 591362 220816
rect 607214 220804 607220 220816
rect 607272 220804 607278 220856
rect 667474 220804 667480 220856
rect 667532 220844 667538 220856
rect 675294 220844 675300 220856
rect 667532 220816 675300 220844
rect 667532 220804 667538 220816
rect 675294 220804 675300 220816
rect 675352 220804 675358 220856
rect 83182 220736 83188 220788
rect 83240 220776 83246 220788
rect 152090 220776 152096 220788
rect 83240 220748 152096 220776
rect 83240 220736 83246 220748
rect 152090 220736 152096 220748
rect 152148 220736 152154 220788
rect 155862 220736 155868 220788
rect 155920 220776 155926 220788
rect 215386 220776 215392 220788
rect 155920 220748 215392 220776
rect 155920 220736 155926 220748
rect 215386 220736 215392 220748
rect 215444 220736 215450 220788
rect 240318 220736 240324 220788
rect 240376 220776 240382 220788
rect 269758 220776 269764 220788
rect 240376 220748 269764 220776
rect 240376 220736 240382 220748
rect 269758 220736 269764 220748
rect 269816 220736 269822 220788
rect 310514 220736 310520 220788
rect 310572 220776 310578 220788
rect 311158 220776 311164 220788
rect 310572 220748 311164 220776
rect 310572 220736 310578 220748
rect 311158 220736 311164 220748
rect 311216 220736 311222 220788
rect 337930 220736 337936 220788
rect 337988 220776 337994 220788
rect 341242 220776 341248 220788
rect 337988 220748 341248 220776
rect 337988 220736 337994 220748
rect 341242 220736 341248 220748
rect 341300 220736 341306 220788
rect 345842 220736 345848 220788
rect 345900 220776 345906 220788
rect 346394 220776 346400 220788
rect 345900 220748 346400 220776
rect 345900 220736 345906 220748
rect 346394 220736 346400 220748
rect 346452 220736 346458 220788
rect 348418 220736 348424 220788
rect 348476 220776 348482 220788
rect 349522 220776 349528 220788
rect 348476 220748 349528 220776
rect 348476 220736 348482 220748
rect 349522 220736 349528 220748
rect 349580 220736 349586 220788
rect 349798 220736 349804 220788
rect 349856 220776 349862 220788
rect 351178 220776 351184 220788
rect 349856 220748 351184 220776
rect 349856 220736 349862 220748
rect 351178 220736 351184 220748
rect 351236 220736 351242 220788
rect 369118 220736 369124 220788
rect 369176 220776 369182 220788
rect 371878 220776 371884 220788
rect 369176 220748 371884 220776
rect 369176 220736 369182 220748
rect 371878 220736 371884 220748
rect 371936 220736 371942 220788
rect 379330 220736 379336 220788
rect 379388 220776 379394 220788
rect 402514 220776 402520 220788
rect 379388 220748 402520 220776
rect 379388 220736 379394 220748
rect 402514 220736 402520 220748
rect 402572 220736 402578 220788
rect 413462 220736 413468 220788
rect 413520 220776 413526 220788
rect 442258 220776 442264 220788
rect 413520 220748 442264 220776
rect 413520 220736 413526 220748
rect 442258 220736 442264 220748
rect 442316 220736 442322 220788
rect 446214 220736 446220 220788
rect 446272 220776 446278 220788
rect 505002 220776 505008 220788
rect 446272 220748 505008 220776
rect 446272 220736 446278 220748
rect 505002 220736 505008 220748
rect 505060 220776 505066 220788
rect 506014 220776 506020 220788
rect 505060 220748 506020 220776
rect 505060 220736 505066 220748
rect 506014 220736 506020 220748
rect 506072 220736 506078 220788
rect 318150 220668 318156 220720
rect 318208 220708 318214 220720
rect 322198 220708 322204 220720
rect 318208 220680 322204 220708
rect 318208 220668 318214 220680
rect 322198 220668 322204 220680
rect 322256 220668 322262 220720
rect 543706 220680 544148 220708
rect 107838 220600 107844 220652
rect 107896 220640 107902 220652
rect 181530 220640 181536 220652
rect 107896 220612 181536 220640
rect 107896 220600 107902 220612
rect 181530 220600 181536 220612
rect 181588 220600 181594 220652
rect 190638 220600 190644 220652
rect 190696 220640 190702 220652
rect 236454 220640 236460 220652
rect 190696 220612 236460 220640
rect 190696 220600 190702 220612
rect 236454 220600 236460 220612
rect 236512 220600 236518 220652
rect 247862 220600 247868 220652
rect 247920 220640 247926 220652
rect 276934 220640 276940 220652
rect 247920 220612 276940 220640
rect 247920 220600 247926 220612
rect 276934 220600 276940 220612
rect 276992 220600 276998 220652
rect 288342 220600 288348 220652
rect 288400 220640 288406 220652
rect 302418 220640 302424 220652
rect 288400 220612 302424 220640
rect 288400 220600 288406 220612
rect 302418 220600 302424 220612
rect 302476 220600 302482 220652
rect 340598 220600 340604 220652
rect 340656 220640 340662 220652
rect 344554 220640 344560 220652
rect 340656 220612 344560 220640
rect 340656 220600 340662 220612
rect 344554 220600 344560 220612
rect 344612 220600 344618 220652
rect 347222 220600 347228 220652
rect 347280 220640 347286 220652
rect 354490 220640 354496 220652
rect 347280 220612 354496 220640
rect 347280 220600 347286 220612
rect 354490 220600 354496 220612
rect 354548 220600 354554 220652
rect 392762 220600 392768 220652
rect 392820 220640 392826 220652
rect 422478 220640 422484 220652
rect 392820 220612 422484 220640
rect 392820 220600 392826 220612
rect 422478 220600 422484 220612
rect 422536 220600 422542 220652
rect 437290 220600 437296 220652
rect 437348 220640 437354 220652
rect 478782 220640 478788 220652
rect 437348 220612 478788 220640
rect 437348 220600 437354 220612
rect 478782 220600 478788 220612
rect 478840 220600 478846 220652
rect 479518 220600 479524 220652
rect 479576 220640 479582 220652
rect 543550 220640 543556 220652
rect 479576 220612 543556 220640
rect 479576 220600 479582 220612
rect 543550 220600 543556 220612
rect 543608 220600 543614 220652
rect 103422 220464 103428 220516
rect 103480 220504 103486 220516
rect 177022 220504 177028 220516
rect 103480 220476 177028 220504
rect 103480 220464 103486 220476
rect 177022 220464 177028 220476
rect 177080 220464 177086 220516
rect 180702 220464 180708 220516
rect 180760 220504 180766 220516
rect 229922 220504 229928 220516
rect 180760 220476 229928 220504
rect 180760 220464 180766 220476
rect 229922 220464 229928 220476
rect 229980 220464 229986 220516
rect 233694 220464 233700 220516
rect 233752 220504 233758 220516
rect 265342 220504 265348 220516
rect 233752 220476 265348 220504
rect 233752 220464 233758 220476
rect 265342 220464 265348 220476
rect 265400 220464 265406 220516
rect 268470 220464 268476 220516
rect 268528 220504 268534 220516
rect 288986 220504 288992 220516
rect 268528 220476 288992 220504
rect 268528 220464 268534 220476
rect 288986 220464 288992 220476
rect 289044 220464 289050 220516
rect 352558 220464 352564 220516
rect 352616 220504 352622 220516
rect 357802 220504 357808 220516
rect 352616 220476 357808 220504
rect 352616 220464 352622 220476
rect 357802 220464 357808 220476
rect 357860 220464 357866 220516
rect 362862 220464 362868 220516
rect 362920 220504 362926 220516
rect 379330 220504 379336 220516
rect 362920 220476 379336 220504
rect 362920 220464 362926 220476
rect 379330 220464 379336 220476
rect 379388 220464 379394 220516
rect 384666 220464 384672 220516
rect 384724 220504 384730 220516
rect 412450 220504 412456 220516
rect 384724 220476 412456 220504
rect 384724 220464 384730 220476
rect 412450 220464 412456 220476
rect 412508 220464 412514 220516
rect 415302 220464 415308 220516
rect 415360 220504 415366 220516
rect 453022 220504 453028 220516
rect 415360 220476 453028 220504
rect 415360 220464 415366 220476
rect 453022 220464 453028 220476
rect 453080 220464 453086 220516
rect 473170 220464 473176 220516
rect 473228 220504 473234 220516
rect 539042 220504 539048 220516
rect 473228 220476 539048 220504
rect 473228 220464 473234 220476
rect 539042 220464 539048 220476
rect 539100 220464 539106 220516
rect 540790 220464 540796 220516
rect 540848 220504 540854 220516
rect 543706 220504 543734 220680
rect 540848 220476 543734 220504
rect 540848 220464 540854 220476
rect 94590 220328 94596 220380
rect 94648 220368 94654 220380
rect 172882 220368 172888 220380
rect 94648 220340 172888 220368
rect 94648 220328 94654 220340
rect 172882 220328 172888 220340
rect 172940 220328 172946 220380
rect 174078 220328 174084 220380
rect 174136 220368 174142 220380
rect 225506 220368 225512 220380
rect 174136 220340 225512 220368
rect 174136 220328 174142 220340
rect 225506 220328 225512 220340
rect 225564 220328 225570 220380
rect 230382 220328 230388 220380
rect 230440 220368 230446 220380
rect 263042 220368 263048 220380
rect 230440 220340 263048 220368
rect 230440 220328 230446 220340
rect 263042 220328 263048 220340
rect 263100 220328 263106 220380
rect 264330 220328 264336 220380
rect 264388 220368 264394 220380
rect 287882 220368 287888 220380
rect 264388 220340 287888 220368
rect 264388 220328 264394 220340
rect 287882 220328 287888 220340
rect 287940 220328 287946 220380
rect 288526 220328 288532 220380
rect 288584 220368 288590 220380
rect 303706 220368 303712 220380
rect 288584 220340 303712 220368
rect 288584 220328 288590 220340
rect 303706 220328 303712 220340
rect 303764 220328 303770 220380
rect 354306 220328 354312 220380
rect 354364 220368 354370 220380
rect 361758 220368 361764 220380
rect 354364 220340 361764 220368
rect 354364 220328 354370 220340
rect 361758 220328 361764 220340
rect 361816 220328 361822 220380
rect 365438 220328 365444 220380
rect 365496 220368 365502 220380
rect 380986 220368 380992 220380
rect 365496 220340 380992 220368
rect 365496 220328 365502 220340
rect 380986 220328 380992 220340
rect 381044 220328 381050 220380
rect 390462 220328 390468 220380
rect 390520 220368 390526 220380
rect 419074 220368 419080 220380
rect 390520 220340 419080 220368
rect 390520 220328 390526 220340
rect 419074 220328 419080 220340
rect 419132 220328 419138 220380
rect 420546 220328 420552 220380
rect 420604 220368 420610 220380
rect 459830 220368 459836 220380
rect 420604 220340 459836 220368
rect 420604 220328 420610 220340
rect 459830 220328 459836 220340
rect 459888 220328 459894 220380
rect 477770 220328 477776 220380
rect 477828 220368 477834 220380
rect 543826 220368 543832 220380
rect 477828 220340 543832 220368
rect 477828 220328 477834 220340
rect 543826 220328 543832 220340
rect 543884 220328 543890 220380
rect 544120 220368 544148 220680
rect 553348 220668 553354 220720
rect 553406 220708 553412 220720
rect 553406 220680 558224 220708
rect 553406 220668 553412 220680
rect 544378 220600 544384 220652
rect 544436 220640 544442 220652
rect 553118 220640 553124 220652
rect 544436 220612 553124 220640
rect 544436 220600 544442 220612
rect 553118 220600 553124 220612
rect 553176 220600 553182 220652
rect 557994 220504 558000 220516
rect 544396 220476 558000 220504
rect 544396 220368 544424 220476
rect 557994 220464 558000 220476
rect 558052 220464 558058 220516
rect 558196 220504 558224 220680
rect 558362 220668 558368 220720
rect 558420 220708 558426 220720
rect 562778 220708 562784 220720
rect 558420 220680 562784 220708
rect 558420 220668 558426 220680
rect 562778 220668 562784 220680
rect 562836 220668 562842 220720
rect 562962 220668 562968 220720
rect 563020 220708 563026 220720
rect 572530 220708 572536 220720
rect 563020 220680 572536 220708
rect 563020 220668 563026 220680
rect 572530 220668 572536 220680
rect 572588 220668 572594 220720
rect 572668 220600 572674 220652
rect 572726 220640 572732 220652
rect 574554 220640 574560 220652
rect 572726 220612 574560 220640
rect 572726 220600 572732 220612
rect 574554 220600 574560 220612
rect 574612 220600 574618 220652
rect 574738 220600 574744 220652
rect 574796 220640 574802 220652
rect 597002 220640 597008 220652
rect 574796 220612 597008 220640
rect 574796 220600 574802 220612
rect 597002 220600 597008 220612
rect 597060 220600 597066 220652
rect 607766 220504 607772 220516
rect 558196 220476 607772 220504
rect 607766 220464 607772 220476
rect 607824 220464 607830 220516
rect 544120 220340 544424 220368
rect 545758 220328 545764 220380
rect 545816 220368 545822 220380
rect 545816 220340 553716 220368
rect 545816 220328 545822 220340
rect 76374 220192 76380 220244
rect 76432 220232 76438 220244
rect 153930 220232 153936 220244
rect 76432 220204 153936 220232
rect 76432 220192 76438 220204
rect 153930 220192 153936 220204
rect 153988 220192 153994 220244
rect 156046 220232 156052 220244
rect 154132 220204 156052 220232
rect 69750 220056 69756 220108
rect 69808 220096 69814 220108
rect 154132 220096 154160 220204
rect 156046 220192 156052 220204
rect 156104 220192 156110 220244
rect 156230 220192 156236 220244
rect 156288 220232 156294 220244
rect 160646 220232 160652 220244
rect 156288 220204 160652 220232
rect 156288 220192 156294 220204
rect 160646 220192 160652 220204
rect 160704 220192 160710 220244
rect 160830 220192 160836 220244
rect 160888 220232 160894 220244
rect 216858 220232 216864 220244
rect 160888 220204 216864 220232
rect 160888 220192 160894 220204
rect 216858 220192 216864 220204
rect 216916 220192 216922 220244
rect 226886 220192 226892 220244
rect 226944 220232 226950 220244
rect 233418 220232 233424 220244
rect 226944 220204 233424 220232
rect 226944 220192 226950 220204
rect 233418 220192 233424 220204
rect 233476 220192 233482 220244
rect 237834 220192 237840 220244
rect 237892 220232 237898 220244
rect 270586 220232 270592 220244
rect 237892 220204 270592 220232
rect 237892 220192 237898 220204
rect 270586 220192 270592 220204
rect 270644 220192 270650 220244
rect 271598 220192 271604 220244
rect 271656 220232 271662 220244
rect 291378 220232 291384 220244
rect 271656 220204 291384 220232
rect 271656 220192 271662 220204
rect 291378 220192 291384 220204
rect 291436 220192 291442 220244
rect 303430 220192 303436 220244
rect 303488 220232 303494 220244
rect 310790 220232 310796 220244
rect 303488 220204 310796 220232
rect 303488 220192 303494 220204
rect 310790 220192 310796 220204
rect 310848 220192 310854 220244
rect 343266 220192 343272 220244
rect 343324 220232 343330 220244
rect 347866 220232 347872 220244
rect 343324 220204 347872 220232
rect 343324 220192 343330 220204
rect 347866 220192 347872 220204
rect 347924 220192 347930 220244
rect 358262 220192 358268 220244
rect 358320 220232 358326 220244
rect 371050 220232 371056 220244
rect 358320 220204 371056 220232
rect 358320 220192 358326 220204
rect 371050 220192 371056 220204
rect 371108 220192 371114 220244
rect 372062 220192 372068 220244
rect 372120 220232 372126 220244
rect 389266 220232 389272 220244
rect 372120 220204 389272 220232
rect 372120 220192 372126 220204
rect 389266 220192 389272 220204
rect 389324 220192 389330 220244
rect 395706 220192 395712 220244
rect 395764 220232 395770 220244
rect 429010 220232 429016 220244
rect 395764 220204 429016 220232
rect 395764 220192 395770 220204
rect 429010 220192 429016 220204
rect 429068 220192 429074 220244
rect 436002 220192 436008 220244
rect 436060 220232 436066 220244
rect 480254 220232 480260 220244
rect 436060 220204 480260 220232
rect 436060 220192 436066 220204
rect 480254 220192 480260 220204
rect 480312 220192 480318 220244
rect 481542 220192 481548 220244
rect 481600 220232 481606 220244
rect 552934 220232 552940 220244
rect 481600 220204 552940 220232
rect 481600 220192 481606 220204
rect 552934 220192 552940 220204
rect 552992 220192 552998 220244
rect 553688 220232 553716 220340
rect 553854 220328 553860 220380
rect 553912 220368 553918 220380
rect 608870 220368 608876 220380
rect 553912 220340 608876 220368
rect 553912 220328 553918 220340
rect 608870 220328 608876 220340
rect 608928 220328 608934 220380
rect 557810 220232 557816 220244
rect 553688 220204 557816 220232
rect 557810 220192 557816 220204
rect 557868 220192 557874 220244
rect 557994 220192 558000 220244
rect 558052 220232 558058 220244
rect 564618 220232 564624 220244
rect 558052 220204 564624 220232
rect 558052 220192 558058 220204
rect 564618 220192 564624 220204
rect 564676 220192 564682 220244
rect 596634 220192 596640 220244
rect 596692 220232 596698 220244
rect 605006 220232 605012 220244
rect 596692 220204 605012 220232
rect 596692 220192 596698 220204
rect 605006 220192 605012 220204
rect 605064 220192 605070 220244
rect 596450 220164 596456 220176
rect 565188 220136 596456 220164
rect 69808 220068 154160 220096
rect 69808 220056 69814 220068
rect 154298 220056 154304 220108
rect 154356 220096 154362 220108
rect 212626 220096 212632 220108
rect 154356 220068 212632 220096
rect 154356 220056 154362 220068
rect 212626 220056 212632 220068
rect 212684 220056 212690 220108
rect 217134 220056 217140 220108
rect 217192 220096 217198 220108
rect 254302 220096 254308 220108
rect 217192 220068 254308 220096
rect 217192 220056 217198 220068
rect 254302 220056 254308 220068
rect 254360 220056 254366 220108
rect 256878 220056 256884 220108
rect 256936 220096 256942 220108
rect 280706 220096 280712 220108
rect 256936 220068 280712 220096
rect 256936 220056 256942 220068
rect 280706 220056 280712 220068
rect 280764 220056 280770 220108
rect 281258 220056 281264 220108
rect 281316 220096 281322 220108
rect 297082 220096 297088 220108
rect 281316 220068 297088 220096
rect 281316 220056 281322 220068
rect 297082 220056 297088 220068
rect 297140 220056 297146 220108
rect 298278 220056 298284 220108
rect 298336 220096 298342 220108
rect 309226 220096 309232 220108
rect 298336 220068 309232 220096
rect 298336 220056 298342 220068
rect 309226 220056 309232 220068
rect 309284 220056 309290 220108
rect 355962 220056 355968 220108
rect 356020 220096 356026 220108
rect 367738 220096 367744 220108
rect 356020 220068 367744 220096
rect 356020 220056 356026 220068
rect 367738 220056 367744 220068
rect 367796 220056 367802 220108
rect 373718 220056 373724 220108
rect 373776 220096 373782 220108
rect 395890 220096 395896 220108
rect 373776 220068 395896 220096
rect 373776 220056 373782 220068
rect 395890 220056 395896 220068
rect 395948 220056 395954 220108
rect 398558 220056 398564 220108
rect 398616 220096 398622 220108
rect 432322 220096 432328 220108
rect 398616 220068 432328 220096
rect 398616 220056 398622 220068
rect 432322 220056 432328 220068
rect 432380 220056 432386 220108
rect 442902 220056 442908 220108
rect 442960 220096 442966 220108
rect 485728 220096 485734 220108
rect 442960 220068 485734 220096
rect 442960 220056 442966 220068
rect 485728 220056 485734 220068
rect 485786 220056 485792 220108
rect 485866 220056 485872 220108
rect 485924 220096 485930 220108
rect 553394 220096 553400 220108
rect 485924 220068 553400 220096
rect 485924 220056 485930 220068
rect 553394 220056 553400 220068
rect 553452 220056 553458 220108
rect 565188 220096 565216 220136
rect 596450 220124 596456 220136
rect 596508 220124 596514 220176
rect 560266 220068 565216 220096
rect 560266 220028 560294 220068
rect 555620 220000 560294 220028
rect 124398 219920 124404 219972
rect 124456 219960 124462 219972
rect 192478 219960 192484 219972
rect 124456 219932 192484 219960
rect 124456 219920 124462 219932
rect 192478 219920 192484 219932
rect 192536 219920 192542 219972
rect 200574 219920 200580 219972
rect 200632 219960 200638 219972
rect 243262 219960 243268 219972
rect 200632 219932 243268 219960
rect 200632 219920 200638 219932
rect 243262 219920 243268 219932
rect 243320 219920 243326 219972
rect 388622 219920 388628 219972
rect 388680 219960 388686 219972
rect 415762 219960 415768 219972
rect 388680 219932 415768 219960
rect 388680 219920 388686 219932
rect 415762 219920 415768 219932
rect 415820 219920 415826 219972
rect 418798 219920 418804 219972
rect 418856 219960 418862 219972
rect 455506 219960 455512 219972
rect 418856 219932 455512 219960
rect 418856 219920 418862 219932
rect 455506 219920 455512 219932
rect 455564 219920 455570 219972
rect 469490 219920 469496 219972
rect 469548 219960 469554 219972
rect 526438 219960 526444 219972
rect 469548 219932 526444 219960
rect 469548 219920 469554 219932
rect 526438 219920 526444 219932
rect 526496 219920 526502 219972
rect 533338 219892 533344 219904
rect 529032 219864 533344 219892
rect 126054 219784 126060 219836
rect 126112 219824 126118 219836
rect 191282 219824 191288 219836
rect 126112 219796 191288 219824
rect 126112 219784 126118 219796
rect 191282 219784 191288 219796
rect 191340 219784 191346 219836
rect 193030 219784 193036 219836
rect 193088 219824 193094 219836
rect 200850 219824 200856 219836
rect 193088 219796 200856 219824
rect 193088 219784 193094 219796
rect 200850 219784 200856 219796
rect 200908 219784 200914 219836
rect 207198 219784 207204 219836
rect 207256 219824 207262 219836
rect 247494 219824 247500 219836
rect 207256 219796 247500 219824
rect 207256 219784 207262 219796
rect 247494 219784 247500 219796
rect 247552 219784 247558 219836
rect 428826 219784 428832 219836
rect 428884 219824 428890 219836
rect 462314 219824 462320 219836
rect 428884 219796 462320 219824
rect 428884 219784 428890 219796
rect 462314 219784 462320 219796
rect 462372 219784 462378 219836
rect 464982 219784 464988 219836
rect 465040 219824 465046 219836
rect 529032 219824 529060 219864
rect 533338 219852 533344 219864
rect 533396 219892 533402 219904
rect 533396 219864 534074 219892
rect 533396 219852 533402 219864
rect 465040 219796 529060 219824
rect 465040 219784 465046 219796
rect 530854 219756 530860 219768
rect 529262 219728 530860 219756
rect 48958 219648 48964 219700
rect 49016 219688 49022 219700
rect 54202 219688 54208 219700
rect 49016 219660 54208 219688
rect 49016 219648 49022 219660
rect 54202 219648 54208 219660
rect 54260 219648 54266 219700
rect 138290 219648 138296 219700
rect 138348 219688 138354 219700
rect 143626 219688 143632 219700
rect 138348 219660 143632 219688
rect 138348 219648 138354 219660
rect 143626 219648 143632 219660
rect 143684 219648 143690 219700
rect 203518 219688 203524 219700
rect 144288 219660 203524 219688
rect 128446 219580 128452 219632
rect 128504 219620 128510 219632
rect 129734 219620 129740 219632
rect 128504 219592 129740 219620
rect 128504 219580 128510 219592
rect 129734 219580 129740 219592
rect 129792 219580 129798 219632
rect 140958 219512 140964 219564
rect 141016 219552 141022 219564
rect 144288 219552 144316 219660
rect 203518 219648 203524 219660
rect 203576 219648 203582 219700
rect 205358 219648 205364 219700
rect 205416 219688 205422 219700
rect 205818 219688 205824 219700
rect 205416 219660 205824 219688
rect 205416 219648 205422 219660
rect 205818 219648 205824 219660
rect 205876 219648 205882 219700
rect 213914 219648 213920 219700
rect 213972 219688 213978 219700
rect 224402 219688 224408 219700
rect 213972 219660 224408 219688
rect 213972 219648 213978 219660
rect 224402 219648 224408 219660
rect 224460 219648 224466 219700
rect 421374 219648 421380 219700
rect 421432 219688 421438 219700
rect 445570 219688 445576 219700
rect 421432 219660 445576 219688
rect 421432 219648 421438 219660
rect 445570 219648 445576 219660
rect 445628 219648 445634 219700
rect 463510 219648 463516 219700
rect 463568 219688 463574 219700
rect 529262 219688 529290 219728
rect 530854 219716 530860 219728
rect 530912 219716 530918 219768
rect 534046 219756 534074 219864
rect 538674 219852 538680 219904
rect 538732 219892 538738 219904
rect 540790 219892 540796 219904
rect 538732 219864 540796 219892
rect 538732 219852 538738 219864
rect 540790 219852 540796 219864
rect 540848 219852 540854 219904
rect 540974 219852 540980 219904
rect 541032 219892 541038 219904
rect 555620 219892 555648 220000
rect 565354 219988 565360 220040
rect 565412 220028 565418 220040
rect 574738 220028 574744 220040
rect 565412 220000 574744 220028
rect 565412 219988 565418 220000
rect 574738 219988 574744 220000
rect 574796 219988 574802 220040
rect 574922 219988 574928 220040
rect 574980 220028 574986 220040
rect 610158 220028 610164 220040
rect 574980 220000 610164 220028
rect 574980 219988 574986 220000
rect 610158 219988 610164 220000
rect 610216 219988 610222 220040
rect 541032 219864 555648 219892
rect 541032 219852 541038 219864
rect 557810 219852 557816 219904
rect 557868 219892 557874 219904
rect 557868 219864 596864 219892
rect 557868 219852 557874 219864
rect 534046 219728 538904 219756
rect 463568 219660 529290 219688
rect 463568 219648 463574 219660
rect 350258 219580 350264 219632
rect 350316 219620 350322 219632
rect 350316 219592 355732 219620
rect 350316 219580 350322 219592
rect 141016 219524 144316 219552
rect 141016 219512 141022 219524
rect 145006 219512 145012 219564
rect 145064 219552 145070 219564
rect 147398 219552 147404 219564
rect 145064 219524 147404 219552
rect 145064 219512 145070 219524
rect 147398 219512 147404 219524
rect 147456 219512 147462 219564
rect 147582 219512 147588 219564
rect 147640 219552 147646 219564
rect 207842 219552 207848 219564
rect 147640 219524 207848 219552
rect 147640 219512 147646 219524
rect 207842 219512 207848 219524
rect 207900 219512 207906 219564
rect 83182 219484 83188 219496
rect 82004 219456 83188 219484
rect 63126 219376 63132 219428
rect 63184 219416 63190 219428
rect 82004 219416 82032 219456
rect 83182 219444 83188 219456
rect 83240 219444 83246 219496
rect 127544 219456 128768 219484
rect 63184 219388 82032 219416
rect 63184 219376 63190 219388
rect 97074 219376 97080 219428
rect 97132 219416 97138 219428
rect 97994 219416 98000 219428
rect 97132 219388 98000 219416
rect 97132 219376 97138 219388
rect 97994 219376 98000 219388
rect 98052 219376 98058 219428
rect 108298 219376 108304 219428
rect 108356 219416 108362 219428
rect 113818 219416 113824 219428
rect 108356 219388 113824 219416
rect 108356 219376 108362 219388
rect 113818 219376 113824 219388
rect 113876 219376 113882 219428
rect 114462 219376 114468 219428
rect 114520 219416 114526 219428
rect 127544 219416 127572 219456
rect 114520 219388 127572 219416
rect 128740 219416 128768 219456
rect 144454 219444 144460 219496
rect 144512 219484 144518 219496
rect 226886 219484 226892 219496
rect 144512 219456 144914 219484
rect 144512 219444 144518 219456
rect 131666 219416 131672 219428
rect 128740 219388 131672 219416
rect 114520 219376 114526 219388
rect 131666 219376 131672 219388
rect 131724 219376 131730 219428
rect 131850 219376 131856 219428
rect 131908 219416 131914 219428
rect 132402 219416 132408 219428
rect 131908 219388 132408 219416
rect 131908 219376 131914 219388
rect 132402 219376 132408 219388
rect 132460 219376 132466 219428
rect 132678 219376 132684 219428
rect 132736 219416 132742 219428
rect 133414 219416 133420 219428
rect 132736 219388 133420 219416
rect 132736 219376 132742 219388
rect 133414 219376 133420 219388
rect 133472 219376 133478 219428
rect 135990 219376 135996 219428
rect 136048 219416 136054 219428
rect 136542 219416 136548 219428
rect 136048 219388 136548 219416
rect 136048 219376 136054 219388
rect 136542 219376 136548 219388
rect 136600 219376 136606 219428
rect 136818 219376 136824 219428
rect 136876 219416 136882 219428
rect 138290 219416 138296 219428
rect 136876 219388 138296 219416
rect 136876 219376 136882 219388
rect 138290 219376 138296 219388
rect 138348 219376 138354 219428
rect 138474 219376 138480 219428
rect 138532 219416 138538 219428
rect 141142 219416 141148 219428
rect 138532 219388 141148 219416
rect 138532 219376 138538 219388
rect 141142 219376 141148 219388
rect 141200 219376 141206 219428
rect 144886 219416 144914 219456
rect 225248 219456 226892 219484
rect 169202 219416 169208 219428
rect 144886 219388 169208 219416
rect 169202 219376 169208 219388
rect 169260 219376 169266 219428
rect 169938 219376 169944 219428
rect 169996 219416 170002 219428
rect 178586 219416 178592 219428
rect 169996 219388 178592 219416
rect 169996 219376 170002 219388
rect 178586 219376 178592 219388
rect 178644 219376 178650 219428
rect 184014 219376 184020 219428
rect 184072 219416 184078 219428
rect 184934 219416 184940 219428
rect 184072 219388 184940 219416
rect 184072 219376 184078 219388
rect 184934 219376 184940 219388
rect 184992 219376 184998 219428
rect 185302 219376 185308 219428
rect 185360 219416 185366 219428
rect 189718 219416 189724 219428
rect 185360 219388 189724 219416
rect 185360 219376 185366 219388
rect 189718 219376 189724 219388
rect 189776 219376 189782 219428
rect 189902 219376 189908 219428
rect 189960 219416 189966 219428
rect 225248 219416 225276 219456
rect 226886 219444 226892 219456
rect 226944 219444 226950 219496
rect 266648 219456 267642 219484
rect 189960 219388 225276 219416
rect 189960 219376 189966 219388
rect 236178 219376 236184 219428
rect 236236 219416 236242 219428
rect 266648 219416 266676 219456
rect 236236 219388 266676 219416
rect 267614 219416 267642 219456
rect 311526 219444 311532 219496
rect 311584 219484 311590 219496
rect 317690 219484 317696 219496
rect 311584 219456 317696 219484
rect 311584 219444 311590 219456
rect 317690 219444 317696 219456
rect 317748 219444 317754 219496
rect 323026 219484 323032 219496
rect 321572 219456 323032 219484
rect 267918 219416 267924 219428
rect 267614 219388 267924 219416
rect 236236 219376 236242 219388
rect 267918 219376 267924 219388
rect 267976 219376 267982 219428
rect 269298 219376 269304 219428
rect 269356 219416 269362 219428
rect 284938 219416 284944 219428
rect 269356 219388 284944 219416
rect 269356 219376 269362 219388
rect 284938 219376 284944 219388
rect 284996 219376 285002 219428
rect 299934 219376 299940 219428
rect 299992 219416 299998 219428
rect 300854 219416 300860 219428
rect 299992 219388 300860 219416
rect 299992 219376 299998 219388
rect 300854 219376 300860 219388
rect 300912 219376 300918 219428
rect 319806 219376 319812 219428
rect 319864 219416 319870 219428
rect 321572 219416 321600 219456
rect 323026 219444 323032 219456
rect 323084 219444 323090 219496
rect 324038 219444 324044 219496
rect 324096 219484 324102 219496
rect 327810 219484 327816 219496
rect 324096 219456 327816 219484
rect 324096 219444 324102 219456
rect 327810 219444 327816 219456
rect 327868 219444 327874 219496
rect 344278 219444 344284 219496
rect 344336 219484 344342 219496
rect 346210 219484 346216 219496
rect 344336 219456 346216 219484
rect 344336 219444 344342 219456
rect 346210 219444 346216 219456
rect 346268 219444 346274 219496
rect 319864 219388 321600 219416
rect 319864 219376 319870 219388
rect 355704 219348 355732 219592
rect 529382 219580 529388 219632
rect 529440 219620 529446 219632
rect 538674 219620 538680 219632
rect 529440 219592 538680 219620
rect 529440 219580 529446 219592
rect 538674 219580 538680 219592
rect 538732 219580 538738 219632
rect 538876 219620 538904 219728
rect 539042 219716 539048 219768
rect 539100 219756 539106 219768
rect 543826 219756 543832 219768
rect 539100 219728 543832 219756
rect 539100 219716 539106 219728
rect 543826 219716 543832 219728
rect 543884 219716 543890 219768
rect 545206 219716 545212 219768
rect 545264 219756 545270 219768
rect 596634 219756 596640 219768
rect 545264 219728 596640 219756
rect 545264 219716 545270 219728
rect 596634 219716 596640 219728
rect 596692 219716 596698 219768
rect 596836 219756 596864 219864
rect 597002 219852 597008 219904
rect 597060 219892 597066 219904
rect 605926 219892 605932 219904
rect 597060 219864 605932 219892
rect 597060 219852 597066 219864
rect 605926 219852 605932 219864
rect 605984 219852 605990 219904
rect 675478 219824 675484 219836
rect 669286 219796 675484 219824
rect 606110 219756 606116 219768
rect 596836 219728 606116 219756
rect 606110 219716 606116 219728
rect 606168 219716 606174 219768
rect 666186 219716 666192 219768
rect 666244 219756 666250 219768
rect 669286 219756 669314 219796
rect 675478 219784 675484 219796
rect 675536 219784 675542 219836
rect 666244 219728 669314 219756
rect 666244 219716 666250 219728
rect 603902 219620 603908 219632
rect 538876 219592 603908 219620
rect 603902 219580 603908 219592
rect 603960 219580 603966 219632
rect 665082 219580 665088 219632
rect 665140 219620 665146 219632
rect 675294 219620 675300 219632
rect 665140 219592 675300 219620
rect 665140 219580 665146 219592
rect 675294 219580 675300 219592
rect 675352 219580 675358 219632
rect 447686 219512 447692 219564
rect 447744 219552 447750 219564
rect 506842 219552 506848 219564
rect 447744 219524 506848 219552
rect 447744 219512 447750 219524
rect 506842 219512 506848 219524
rect 506900 219512 506906 219564
rect 511074 219444 511080 219496
rect 511132 219484 511138 219496
rect 511132 219456 596312 219484
rect 511132 219444 511138 219456
rect 422294 219376 422300 219428
rect 422352 219416 422358 219428
rect 448882 219416 448888 219428
rect 422352 219388 448888 219416
rect 422352 219376 422358 219388
rect 448882 219376 448888 219388
rect 448940 219376 448946 219428
rect 449158 219376 449164 219428
rect 449216 219416 449222 219428
rect 449216 219388 457300 219416
rect 449216 219376 449222 219388
rect 356974 219348 356980 219360
rect 128326 219320 128584 219348
rect 355704 219320 356980 219348
rect 88978 219280 88984 219292
rect 64846 219252 88984 219280
rect 64598 219104 64604 219156
rect 64656 219144 64662 219156
rect 64846 219144 64874 219252
rect 88978 219240 88984 219252
rect 89036 219240 89042 219292
rect 100386 219240 100392 219292
rect 100444 219280 100450 219292
rect 128326 219280 128354 219320
rect 100444 219252 128354 219280
rect 128556 219280 128584 219320
rect 356974 219308 356980 219320
rect 357032 219308 357038 219360
rect 147214 219280 147220 219292
rect 128556 219252 147220 219280
rect 100444 219240 100450 219252
rect 147214 219240 147220 219252
rect 147272 219240 147278 219292
rect 147398 219240 147404 219292
rect 147456 219280 147462 219292
rect 192478 219280 192484 219292
rect 147456 219252 192484 219280
rect 147456 219240 147462 219252
rect 192478 219240 192484 219252
rect 192536 219240 192542 219292
rect 195606 219240 195612 219292
rect 195664 219280 195670 219292
rect 197906 219280 197912 219292
rect 195664 219252 197912 219280
rect 195664 219240 195670 219252
rect 197906 219240 197912 219252
rect 197964 219240 197970 219292
rect 198918 219240 198924 219292
rect 198976 219280 198982 219292
rect 200022 219280 200028 219292
rect 198976 219252 200028 219280
rect 198976 219240 198982 219252
rect 200022 219240 200028 219252
rect 200080 219240 200086 219292
rect 200206 219240 200212 219292
rect 200264 219280 200270 219292
rect 201034 219280 201040 219292
rect 200264 219252 201040 219280
rect 200264 219240 200270 219252
rect 201034 219240 201040 219252
rect 201092 219240 201098 219292
rect 208854 219240 208860 219292
rect 208912 219280 208918 219292
rect 209590 219280 209596 219292
rect 208912 219252 209596 219280
rect 208912 219240 208918 219252
rect 209590 219240 209596 219252
rect 209648 219240 209654 219292
rect 209774 219240 209780 219292
rect 209832 219280 209838 219292
rect 210326 219280 210332 219292
rect 209832 219252 210332 219280
rect 209832 219240 209838 219252
rect 210326 219240 210332 219252
rect 210384 219240 210390 219292
rect 210510 219240 210516 219292
rect 210568 219280 210574 219292
rect 210970 219280 210976 219292
rect 210568 219252 210976 219280
rect 210568 219240 210574 219252
rect 210970 219240 210976 219252
rect 211028 219240 211034 219292
rect 212994 219240 213000 219292
rect 213052 219280 213058 219292
rect 213546 219280 213552 219292
rect 213052 219252 213552 219280
rect 213052 219240 213058 219252
rect 213546 219240 213552 219252
rect 213604 219240 213610 219292
rect 213730 219240 213736 219292
rect 213788 219280 213794 219292
rect 239306 219280 239312 219292
rect 213788 219252 239312 219280
rect 213788 219240 213794 219252
rect 239306 219240 239312 219252
rect 239364 219240 239370 219292
rect 249426 219240 249432 219292
rect 249484 219280 249490 219292
rect 249484 219252 273668 219280
rect 249484 219240 249490 219252
rect 87598 219144 87604 219156
rect 64656 219116 64874 219144
rect 74506 219116 87604 219144
rect 64656 219104 64662 219116
rect 59814 218968 59820 219020
rect 59872 219008 59878 219020
rect 74506 219008 74534 219116
rect 87598 219104 87604 219116
rect 87656 219104 87662 219156
rect 87966 219104 87972 219156
rect 88024 219144 88030 219156
rect 101398 219144 101404 219156
rect 88024 219116 101404 219144
rect 88024 219104 88030 219116
rect 101398 219104 101404 219116
rect 101456 219104 101462 219156
rect 113634 219104 113640 219156
rect 113692 219144 113698 219156
rect 120902 219144 120908 219156
rect 113692 219116 120908 219144
rect 113692 219104 113698 219116
rect 120902 219104 120908 219116
rect 120960 219104 120966 219156
rect 121914 219104 121920 219156
rect 121972 219144 121978 219156
rect 122742 219144 122748 219156
rect 121972 219116 122748 219144
rect 121972 219104 121978 219116
rect 122742 219104 122748 219116
rect 122800 219104 122806 219156
rect 123570 219104 123576 219156
rect 123628 219144 123634 219156
rect 126422 219144 126428 219156
rect 123628 219116 126428 219144
rect 123628 219104 123634 219116
rect 126422 219104 126428 219116
rect 126480 219104 126486 219156
rect 126606 219104 126612 219156
rect 126664 219144 126670 219156
rect 128492 219144 128498 219156
rect 126664 219116 128498 219144
rect 126664 219104 126670 219116
rect 128492 219104 128498 219116
rect 128550 219104 128556 219156
rect 128630 219104 128636 219156
rect 128688 219144 128694 219156
rect 164418 219144 164424 219156
rect 128688 219116 164424 219144
rect 128688 219104 128694 219116
rect 164418 219104 164424 219116
rect 164476 219104 164482 219156
rect 164602 219104 164608 219156
rect 164660 219144 164666 219156
rect 171594 219144 171600 219156
rect 164660 219116 171600 219144
rect 164660 219104 164666 219116
rect 171594 219104 171600 219116
rect 171652 219104 171658 219156
rect 178402 219144 178408 219156
rect 176626 219116 178408 219144
rect 59872 218980 74534 219008
rect 59872 218968 59878 218980
rect 83826 218968 83832 219020
rect 83884 219008 83890 219020
rect 83884 218980 161612 219008
rect 83884 218968 83890 218980
rect 70578 218832 70584 218884
rect 70636 218872 70642 218884
rect 156414 218872 156420 218884
rect 70636 218844 156420 218872
rect 70636 218832 70642 218844
rect 156414 218832 156420 218844
rect 156472 218832 156478 218884
rect 157518 218832 157524 218884
rect 157576 218872 157582 218884
rect 161382 218872 161388 218884
rect 157576 218844 161388 218872
rect 157576 218832 157582 218844
rect 161382 218832 161388 218844
rect 161440 218832 161446 218884
rect 161584 218872 161612 218980
rect 161750 218968 161756 219020
rect 161808 219008 161814 219020
rect 176626 219008 176654 219116
rect 178402 219104 178408 219116
rect 178460 219104 178466 219156
rect 178586 219104 178592 219156
rect 178644 219144 178650 219156
rect 213914 219144 213920 219156
rect 178644 219116 213920 219144
rect 178644 219104 178650 219116
rect 213914 219104 213920 219116
rect 213972 219104 213978 219156
rect 214650 219104 214656 219156
rect 214708 219144 214714 219156
rect 215202 219144 215208 219156
rect 214708 219116 215208 219144
rect 214708 219104 214714 219116
rect 215202 219104 215208 219116
rect 215260 219104 215266 219156
rect 224218 219104 224224 219156
rect 224276 219144 224282 219156
rect 251726 219144 251732 219156
rect 224276 219116 251732 219144
rect 224276 219104 224282 219116
rect 251726 219104 251732 219116
rect 251784 219104 251790 219156
rect 252738 219104 252744 219156
rect 252796 219144 252802 219156
rect 255958 219144 255964 219156
rect 252796 219116 255964 219144
rect 252796 219104 252802 219116
rect 255958 219104 255964 219116
rect 256016 219104 256022 219156
rect 262858 219104 262864 219156
rect 262916 219144 262922 219156
rect 272426 219144 272432 219156
rect 262916 219116 272432 219144
rect 262916 219104 262922 219116
rect 272426 219104 272432 219116
rect 272484 219104 272490 219156
rect 161808 218980 176654 219008
rect 161808 218968 161814 218980
rect 178586 218968 178592 219020
rect 178644 219008 178650 219020
rect 180058 219008 180064 219020
rect 178644 218980 180064 219008
rect 178644 218968 178650 218980
rect 180058 218968 180064 218980
rect 180116 218968 180122 219020
rect 180242 218968 180248 219020
rect 180300 219008 180306 219020
rect 185762 219008 185768 219020
rect 180300 218980 185768 219008
rect 180300 218968 180306 218980
rect 185762 218968 185768 218980
rect 185820 218968 185826 219020
rect 185946 218968 185952 219020
rect 186004 219008 186010 219020
rect 209130 219008 209136 219020
rect 186004 218980 209136 219008
rect 186004 218968 186010 218980
rect 209130 218968 209136 218980
rect 209188 218968 209194 219020
rect 215938 219008 215944 219020
rect 209332 218980 215944 219008
rect 167362 218872 167368 218884
rect 161584 218844 167368 218872
rect 167362 218832 167368 218844
rect 167420 218832 167426 218884
rect 167546 218832 167552 218884
rect 167604 218872 167610 218884
rect 170122 218872 170128 218884
rect 167604 218844 170128 218872
rect 167604 218832 167610 218844
rect 170122 218832 170128 218844
rect 170180 218832 170186 218884
rect 171594 218832 171600 218884
rect 171652 218872 171658 218884
rect 209332 218872 209360 218980
rect 215938 218968 215944 218980
rect 215996 218968 216002 219020
rect 217962 218968 217968 219020
rect 218020 219008 218026 219020
rect 221458 219008 221464 219020
rect 218020 218980 221464 219008
rect 218020 218968 218026 218980
rect 221458 218968 221464 218980
rect 221516 218968 221522 219020
rect 242618 218968 242624 219020
rect 242676 219008 242682 219020
rect 273438 219008 273444 219020
rect 242676 218980 273444 219008
rect 242676 218968 242682 218980
rect 273438 218968 273444 218980
rect 273496 218968 273502 219020
rect 171652 218844 209360 218872
rect 171652 218832 171658 218844
rect 209682 218832 209688 218884
rect 209740 218872 209746 218884
rect 209740 218844 213960 218872
rect 209740 218832 209746 218844
rect 56502 218696 56508 218748
rect 56560 218736 56566 218748
rect 144914 218736 144920 218748
rect 56560 218708 144920 218736
rect 56560 218696 56566 218708
rect 144914 218696 144920 218708
rect 144972 218696 144978 218748
rect 147398 218736 147404 218748
rect 145070 218708 147404 218736
rect 78030 218560 78036 218612
rect 78088 218600 78094 218612
rect 108298 218600 108304 218612
rect 78088 218572 108304 218600
rect 78088 218560 78094 218572
rect 108298 218560 108304 218572
rect 108356 218560 108362 218612
rect 111978 218560 111984 218612
rect 112036 218600 112042 218612
rect 113082 218600 113088 218612
rect 112036 218572 113088 218600
rect 112036 218560 112042 218572
rect 113082 218560 113088 218572
rect 113140 218560 113146 218612
rect 115768 218572 120212 218600
rect 110138 218424 110144 218476
rect 110196 218464 110202 218476
rect 115768 218464 115796 218572
rect 110196 218436 115796 218464
rect 110196 218424 110202 218436
rect 116118 218424 116124 218476
rect 116176 218464 116182 218476
rect 117222 218464 117228 218476
rect 116176 218436 117228 218464
rect 116176 218424 116182 218436
rect 117222 218424 117228 218436
rect 117280 218424 117286 218476
rect 119430 218424 119436 218476
rect 119488 218464 119494 218476
rect 119982 218464 119988 218476
rect 119488 218436 119988 218464
rect 119488 218424 119494 218436
rect 119982 218424 119988 218436
rect 120040 218424 120046 218476
rect 120184 218464 120212 218572
rect 120350 218560 120356 218612
rect 120408 218600 120414 218612
rect 125502 218600 125508 218612
rect 120408 218572 125508 218600
rect 120408 218560 120414 218572
rect 125502 218560 125508 218572
rect 125560 218560 125566 218612
rect 125686 218560 125692 218612
rect 125744 218600 125750 218612
rect 125744 218572 140912 218600
rect 125744 218560 125750 218572
rect 120718 218464 120724 218476
rect 120184 218436 120724 218464
rect 120718 218424 120724 218436
rect 120776 218424 120782 218476
rect 120902 218424 120908 218476
rect 120960 218464 120966 218476
rect 126606 218464 126612 218476
rect 120960 218436 126612 218464
rect 120960 218424 120966 218436
rect 126606 218424 126612 218436
rect 126664 218424 126670 218476
rect 127710 218424 127716 218476
rect 127768 218464 127774 218476
rect 128262 218464 128268 218476
rect 127768 218436 128268 218464
rect 127768 218424 127774 218436
rect 128262 218424 128268 218436
rect 128320 218424 128326 218476
rect 128538 218424 128544 218476
rect 128596 218464 128602 218476
rect 129274 218464 129280 218476
rect 128596 218436 129280 218464
rect 128596 218424 128602 218436
rect 129274 218424 129280 218436
rect 129332 218424 129338 218476
rect 131666 218424 131672 218476
rect 131724 218464 131730 218476
rect 137922 218464 137928 218476
rect 131724 218436 137928 218464
rect 131724 218424 131730 218436
rect 137922 218424 137928 218436
rect 137980 218424 137986 218476
rect 138474 218424 138480 218476
rect 138532 218464 138538 218476
rect 139118 218464 139124 218476
rect 138532 218436 139124 218464
rect 138532 218424 138538 218436
rect 139118 218424 139124 218436
rect 139176 218424 139182 218476
rect 140130 218424 140136 218476
rect 140188 218464 140194 218476
rect 140682 218464 140688 218476
rect 140188 218436 140688 218464
rect 140188 218424 140194 218436
rect 140682 218424 140688 218436
rect 140740 218424 140746 218476
rect 140884 218464 140912 218572
rect 141142 218560 141148 218612
rect 141200 218600 141206 218612
rect 142246 218600 142252 218612
rect 141200 218572 142252 218600
rect 141200 218560 141206 218572
rect 142246 218560 142252 218572
rect 142304 218560 142310 218612
rect 144454 218600 144460 218612
rect 142448 218572 144460 218600
rect 142448 218464 142476 218572
rect 144454 218560 144460 218572
rect 144512 218560 144518 218612
rect 145070 218600 145098 218708
rect 147398 218696 147404 218708
rect 147456 218696 147462 218748
rect 149238 218696 149244 218748
rect 149296 218736 149302 218748
rect 149296 218708 151308 218736
rect 149296 218696 149302 218708
rect 144656 218572 145098 218600
rect 140884 218436 142476 218464
rect 142614 218424 142620 218476
rect 142672 218464 142678 218476
rect 143442 218464 143448 218476
rect 142672 218436 143448 218464
rect 142672 218424 142678 218436
rect 143442 218424 143448 218436
rect 143500 218424 143506 218476
rect 143626 218424 143632 218476
rect 143684 218464 143690 218476
rect 144656 218464 144684 218572
rect 146754 218560 146760 218612
rect 146812 218600 146818 218612
rect 151078 218600 151084 218612
rect 146812 218572 151084 218600
rect 146812 218560 146818 218572
rect 151078 218560 151084 218572
rect 151136 218560 151142 218612
rect 143684 218436 144684 218464
rect 143684 218424 143690 218436
rect 145098 218424 145104 218476
rect 145156 218464 145162 218476
rect 145926 218464 145932 218476
rect 145156 218436 145932 218464
rect 145156 218424 145162 218436
rect 145926 218424 145932 218436
rect 145984 218424 145990 218476
rect 148410 218424 148416 218476
rect 148468 218464 148474 218476
rect 149882 218464 149888 218476
rect 148468 218436 149888 218464
rect 148468 218424 148474 218436
rect 149882 218424 149888 218436
rect 149940 218424 149946 218476
rect 151280 218464 151308 218708
rect 151906 218696 151912 218748
rect 151964 218736 151970 218748
rect 151964 218708 200068 218736
rect 151964 218696 151970 218708
rect 151446 218560 151452 218612
rect 151504 218600 151510 218612
rect 191926 218600 191932 218612
rect 151504 218572 191932 218600
rect 151504 218560 151510 218572
rect 191926 218560 191932 218572
rect 191984 218560 191990 218612
rect 192294 218560 192300 218612
rect 192352 218600 192358 218612
rect 193766 218600 193772 218612
rect 192352 218572 193772 218600
rect 192352 218560 192358 218572
rect 193766 218560 193772 218572
rect 193824 218560 193830 218612
rect 193950 218560 193956 218612
rect 194008 218600 194014 218612
rect 194410 218600 194416 218612
rect 194008 218572 194416 218600
rect 194008 218560 194014 218572
rect 194410 218560 194416 218572
rect 194468 218560 194474 218612
rect 194778 218560 194784 218612
rect 194836 218600 194842 218612
rect 195882 218600 195888 218612
rect 194836 218572 195888 218600
rect 194836 218560 194842 218572
rect 195882 218560 195888 218572
rect 195940 218560 195946 218612
rect 196250 218560 196256 218612
rect 196308 218600 196314 218612
rect 199838 218600 199844 218612
rect 196308 218572 199844 218600
rect 196308 218560 196314 218572
rect 199838 218560 199844 218572
rect 199896 218560 199902 218612
rect 200040 218600 200068 218708
rect 200206 218696 200212 218748
rect 200264 218736 200270 218748
rect 202874 218736 202880 218748
rect 200264 218708 202880 218736
rect 200264 218696 200270 218708
rect 202874 218696 202880 218708
rect 202932 218696 202938 218748
rect 205496 218696 205502 218748
rect 205554 218736 205560 218748
rect 213730 218736 213736 218748
rect 205554 218708 213736 218736
rect 205554 218696 205560 218708
rect 213730 218696 213736 218708
rect 213788 218696 213794 218748
rect 213932 218736 213960 218844
rect 214098 218832 214104 218884
rect 214156 218872 214162 218884
rect 222838 218872 222844 218884
rect 214156 218844 222844 218872
rect 214156 218832 214162 218844
rect 222838 218832 222844 218844
rect 222896 218832 222902 218884
rect 229554 218832 229560 218884
rect 229612 218872 229618 218884
rect 262674 218872 262680 218884
rect 229612 218844 262680 218872
rect 229612 218832 229618 218844
rect 262674 218832 262680 218844
rect 262732 218832 262738 218884
rect 273640 218872 273668 219252
rect 295794 219240 295800 219292
rect 295852 219280 295858 219292
rect 296714 219280 296720 219292
rect 295852 219252 296720 219280
rect 295852 219240 295858 219252
rect 296714 219240 296720 219252
rect 296772 219240 296778 219292
rect 342254 219240 342260 219292
rect 342312 219280 342318 219292
rect 345382 219280 345388 219292
rect 342312 219252 345388 219280
rect 342312 219240 342318 219252
rect 345382 219240 345388 219252
rect 345440 219240 345446 219292
rect 402238 219240 402244 219292
rect 402296 219280 402302 219292
rect 424870 219280 424876 219292
rect 402296 219252 424876 219280
rect 402296 219240 402302 219252
rect 424870 219240 424876 219252
rect 424928 219240 424934 219292
rect 430850 219280 430856 219292
rect 425762 219252 430856 219280
rect 285858 219104 285864 219156
rect 285916 219144 285922 219156
rect 296898 219144 296904 219156
rect 285916 219116 296904 219144
rect 285916 219104 285922 219116
rect 296898 219104 296904 219116
rect 296956 219104 296962 219156
rect 302418 219104 302424 219156
rect 302476 219144 302482 219156
rect 305638 219144 305644 219156
rect 302476 219116 305644 219144
rect 302476 219104 302482 219116
rect 305638 219104 305644 219116
rect 305696 219104 305702 219156
rect 404998 219104 405004 219156
rect 405056 219144 405062 219156
rect 425762 219144 425790 219252
rect 430850 219240 430856 219252
rect 430908 219240 430914 219292
rect 431218 219240 431224 219292
rect 431276 219280 431282 219292
rect 431276 219252 436784 219280
rect 431276 219240 431282 219252
rect 405056 219116 425790 219144
rect 405056 219104 405062 219116
rect 425882 219104 425888 219156
rect 425940 219144 425946 219156
rect 436756 219144 436784 219252
rect 436922 219240 436928 219292
rect 436980 219280 436986 219292
rect 454678 219280 454684 219292
rect 436980 219252 454684 219280
rect 436980 219240 436986 219252
rect 454678 219240 454684 219252
rect 454736 219240 454742 219292
rect 457272 219280 457300 219388
rect 457438 219376 457444 219428
rect 457496 219416 457502 219428
rect 457496 219388 461072 219416
rect 457496 219376 457502 219388
rect 458818 219280 458824 219292
rect 457272 219252 458824 219280
rect 458818 219240 458824 219252
rect 458876 219240 458882 219292
rect 461044 219280 461072 219388
rect 462314 219376 462320 219428
rect 462372 219416 462378 219428
rect 474550 219416 474556 219428
rect 462372 219388 474556 219416
rect 462372 219376 462378 219388
rect 474550 219376 474556 219388
rect 474608 219376 474614 219428
rect 474734 219376 474740 219428
rect 474792 219416 474798 219428
rect 489362 219416 489368 219428
rect 474792 219388 489368 219416
rect 474792 219376 474798 219388
rect 489362 219376 489368 219388
rect 489420 219376 489426 219428
rect 490190 219348 490196 219360
rect 489518 219320 490196 219348
rect 471054 219280 471060 219292
rect 461044 219252 471060 219280
rect 471054 219240 471060 219252
rect 471112 219240 471118 219292
rect 471422 219240 471428 219292
rect 471480 219280 471486 219292
rect 475746 219280 475752 219292
rect 471480 219252 475752 219280
rect 471480 219240 471486 219252
rect 475746 219240 475752 219252
rect 475804 219240 475810 219292
rect 480254 219240 480260 219292
rect 480312 219280 480318 219292
rect 483566 219280 483572 219292
rect 480312 219252 483572 219280
rect 480312 219240 480318 219252
rect 483566 219240 483572 219252
rect 483624 219240 483630 219292
rect 483750 219240 483756 219292
rect 483808 219280 483814 219292
rect 484302 219280 484308 219292
rect 483808 219252 484308 219280
rect 483808 219240 483814 219252
rect 484302 219240 484308 219252
rect 484360 219240 484366 219292
rect 489518 219280 489546 219320
rect 490190 219308 490196 219320
rect 490248 219308 490254 219360
rect 490374 219308 490380 219360
rect 490432 219348 490438 219360
rect 490432 219320 543872 219348
rect 490432 219308 490438 219320
rect 484872 219252 489546 219280
rect 425940 219116 436692 219144
rect 436756 219116 460060 219144
rect 425940 219104 425946 219116
rect 275646 218968 275652 219020
rect 275704 219008 275710 219020
rect 290458 219008 290464 219020
rect 275704 218980 290464 219008
rect 275704 218968 275710 218980
rect 290458 218968 290464 218980
rect 290516 218968 290522 219020
rect 301590 218968 301596 219020
rect 301648 219008 301654 219020
rect 310514 219008 310520 219020
rect 301648 218980 310520 219008
rect 301648 218968 301654 218980
rect 310514 218968 310520 218980
rect 310572 218968 310578 219020
rect 314010 218968 314016 219020
rect 314068 219008 314074 219020
rect 319438 219008 319444 219020
rect 314068 218980 319444 219008
rect 314068 218968 314074 218980
rect 319438 218968 319444 218980
rect 319496 218968 319502 219020
rect 363598 218968 363604 219020
rect 363656 219008 363662 219020
rect 368566 219008 368572 219020
rect 363656 218980 368572 219008
rect 363656 218968 363662 218980
rect 368566 218968 368572 218980
rect 368624 218968 368630 219020
rect 407022 218968 407028 219020
rect 407080 219008 407086 219020
rect 436278 219008 436284 219020
rect 407080 218980 436284 219008
rect 407080 218968 407086 218980
rect 436278 218968 436284 218980
rect 436336 218968 436342 219020
rect 436664 219008 436692 219116
rect 436922 219008 436928 219020
rect 436664 218980 436928 219008
rect 436922 218968 436928 218980
rect 436980 218968 436986 219020
rect 446398 218968 446404 219020
rect 446456 219008 446462 219020
rect 459646 219008 459652 219020
rect 446456 218980 459652 219008
rect 446456 218968 446462 218980
rect 459646 218968 459652 218980
rect 459704 218968 459710 219020
rect 460032 219008 460060 219116
rect 460198 219104 460204 219156
rect 460256 219144 460262 219156
rect 472894 219144 472900 219156
rect 460256 219116 472900 219144
rect 460256 219104 460262 219116
rect 472894 219104 472900 219116
rect 472952 219104 472958 219156
rect 475102 219104 475108 219156
rect 475160 219144 475166 219156
rect 482830 219144 482836 219156
rect 475160 219116 482836 219144
rect 475160 219104 475166 219116
rect 482830 219104 482836 219116
rect 482888 219104 482894 219156
rect 484872 219144 484900 219252
rect 489822 219172 489828 219224
rect 489880 219212 489886 219224
rect 543844 219212 543872 219320
rect 547506 219308 547512 219360
rect 547564 219348 547570 219360
rect 549438 219348 549444 219360
rect 547564 219320 549444 219348
rect 547564 219308 547570 219320
rect 549438 219308 549444 219320
rect 549496 219308 549502 219360
rect 559834 219308 559840 219360
rect 559892 219348 559898 219360
rect 568022 219348 568028 219360
rect 559892 219320 568028 219348
rect 559892 219308 559898 219320
rect 568022 219308 568028 219320
rect 568080 219308 568086 219360
rect 568206 219308 568212 219360
rect 568264 219348 568270 219360
rect 596284 219348 596312 219456
rect 596450 219444 596456 219496
rect 596508 219484 596514 219496
rect 604546 219484 604552 219496
rect 596508 219456 604552 219484
rect 596508 219444 596514 219456
rect 604546 219444 604552 219456
rect 604604 219444 604610 219496
rect 671890 219444 671896 219496
rect 671948 219484 671954 219496
rect 675478 219484 675484 219496
rect 671948 219456 675484 219484
rect 671948 219444 671954 219456
rect 675478 219444 675484 219456
rect 675536 219444 675542 219496
rect 599118 219348 599124 219360
rect 568264 219320 572714 219348
rect 596284 219320 599124 219348
rect 568264 219308 568270 219320
rect 572686 219280 572714 219320
rect 599118 219308 599124 219320
rect 599176 219308 599182 219360
rect 574738 219280 574744 219292
rect 572686 219252 574744 219280
rect 574738 219240 574744 219252
rect 574796 219240 574802 219292
rect 551738 219212 551744 219224
rect 489880 219184 543734 219212
rect 543844 219184 551744 219212
rect 489880 219172 489886 219184
rect 482986 219116 484900 219144
rect 460474 219008 460480 219020
rect 460032 218980 460480 219008
rect 460474 218968 460480 218980
rect 460532 218968 460538 219020
rect 467282 218968 467288 219020
rect 467340 219008 467346 219020
rect 482986 219008 483014 219116
rect 485038 219104 485044 219156
rect 485096 219144 485102 219156
rect 486142 219144 486148 219156
rect 485096 219116 486148 219144
rect 485096 219104 485102 219116
rect 486142 219104 486148 219116
rect 486200 219104 486206 219156
rect 491478 219036 491484 219088
rect 491536 219076 491542 219088
rect 495250 219076 495256 219088
rect 491536 219048 495256 219076
rect 491536 219036 491542 219048
rect 495250 219036 495256 219048
rect 495308 219036 495314 219088
rect 526438 219036 526444 219088
rect 526496 219076 526502 219088
rect 529382 219076 529388 219088
rect 526496 219048 529388 219076
rect 526496 219036 526502 219048
rect 529382 219036 529388 219048
rect 529440 219036 529446 219088
rect 530118 219036 530124 219088
rect 530176 219076 530182 219088
rect 530578 219076 530584 219088
rect 530176 219048 530584 219076
rect 530176 219036 530182 219048
rect 530578 219036 530584 219048
rect 530636 219036 530642 219088
rect 531958 219036 531964 219088
rect 532016 219076 532022 219088
rect 532510 219076 532516 219088
rect 532016 219048 532516 219076
rect 532016 219036 532022 219048
rect 532510 219036 532516 219048
rect 532568 219036 532574 219088
rect 535914 219036 535920 219088
rect 535972 219076 535978 219088
rect 540974 219076 540980 219088
rect 535972 219048 540980 219076
rect 535972 219036 535978 219048
rect 540974 219036 540980 219048
rect 541032 219036 541038 219088
rect 543706 219076 543734 219184
rect 551738 219172 551744 219184
rect 551796 219172 551802 219224
rect 554866 219104 554872 219156
rect 554924 219144 554930 219156
rect 554924 219116 558408 219144
rect 554924 219104 554930 219116
rect 550634 219076 550640 219088
rect 543706 219048 550640 219076
rect 550634 219036 550640 219048
rect 550692 219036 550698 219088
rect 467340 218980 483014 219008
rect 467340 218968 467346 218980
rect 485406 218968 485412 219020
rect 485464 219008 485470 219020
rect 485464 218980 485774 219008
rect 485464 218968 485470 218980
rect 277578 218872 277584 218884
rect 273640 218844 277584 218872
rect 277578 218832 277584 218844
rect 277636 218832 277642 218884
rect 282546 218832 282552 218884
rect 282604 218872 282610 218884
rect 298738 218872 298744 218884
rect 282604 218844 298744 218872
rect 282604 218832 282610 218844
rect 298738 218832 298744 218844
rect 298796 218832 298802 218884
rect 305730 218832 305736 218884
rect 305788 218872 305794 218884
rect 313826 218872 313832 218884
rect 305788 218844 313832 218872
rect 305788 218832 305794 218844
rect 313826 218832 313832 218844
rect 313884 218832 313890 218884
rect 366726 218832 366732 218884
rect 366784 218872 366790 218884
rect 381814 218872 381820 218884
rect 366784 218844 381820 218872
rect 366784 218832 366790 218844
rect 381814 218832 381820 218844
rect 381872 218832 381878 218884
rect 382182 218832 382188 218884
rect 382240 218872 382246 218884
rect 404998 218872 405004 218884
rect 382240 218844 405004 218872
rect 382240 218832 382246 218844
rect 404998 218832 405004 218844
rect 405056 218832 405062 218884
rect 405366 218832 405372 218884
rect 405424 218872 405430 218884
rect 438118 218872 438124 218884
rect 405424 218844 438124 218872
rect 405424 218832 405430 218844
rect 438118 218832 438124 218844
rect 438176 218832 438182 218884
rect 454862 218832 454868 218884
rect 454920 218872 454926 218884
rect 463786 218872 463792 218884
rect 454920 218844 463792 218872
rect 454920 218832 454926 218844
rect 463786 218832 463792 218844
rect 463844 218832 463850 218884
rect 469858 218832 469864 218884
rect 469916 218872 469922 218884
rect 474918 218872 474924 218884
rect 469916 218844 474924 218872
rect 469916 218832 469922 218844
rect 474918 218832 474924 218844
rect 474976 218832 474982 218884
rect 485406 218872 485412 218884
rect 475672 218844 485412 218872
rect 243538 218736 243544 218748
rect 213932 218708 243544 218736
rect 243538 218696 243544 218708
rect 243596 218696 243602 218748
rect 262674 218696 262680 218748
rect 262732 218736 262738 218748
rect 286042 218736 286048 218748
rect 262732 218708 286048 218736
rect 262732 218696 262738 218708
rect 286042 218696 286048 218708
rect 286100 218696 286106 218748
rect 292298 218696 292304 218748
rect 292356 218736 292362 218748
rect 305914 218736 305920 218748
rect 292356 218708 305920 218736
rect 292356 218696 292362 218708
rect 305914 218696 305920 218708
rect 305972 218696 305978 218748
rect 310698 218696 310704 218748
rect 310756 218736 310762 218748
rect 317414 218736 317420 218748
rect 310756 218708 317420 218736
rect 310756 218696 310762 218708
rect 317414 218696 317420 218708
rect 317472 218696 317478 218748
rect 323118 218696 323124 218748
rect 323176 218736 323182 218748
rect 324682 218736 324688 218748
rect 323176 218708 324688 218736
rect 323176 218696 323182 218708
rect 324682 218696 324688 218708
rect 324740 218696 324746 218748
rect 355318 218696 355324 218748
rect 355376 218736 355382 218748
rect 358630 218736 358636 218748
rect 355376 218708 358636 218736
rect 355376 218696 355382 218708
rect 358630 218696 358636 218708
rect 358688 218696 358694 218748
rect 360838 218696 360844 218748
rect 360896 218736 360902 218748
rect 365254 218736 365260 218748
rect 360896 218708 365260 218736
rect 360896 218696 360902 218708
rect 365254 218696 365260 218708
rect 365312 218696 365318 218748
rect 368106 218696 368112 218748
rect 368164 218736 368170 218748
rect 385126 218736 385132 218748
rect 368164 218708 385132 218736
rect 368164 218696 368170 218708
rect 385126 218696 385132 218708
rect 385184 218696 385190 218748
rect 401318 218696 401324 218748
rect 401376 218736 401382 218748
rect 434806 218736 434812 218748
rect 401376 218708 434812 218736
rect 401376 218696 401382 218708
rect 434806 218696 434812 218708
rect 434864 218696 434870 218748
rect 438302 218696 438308 218748
rect 438360 218736 438366 218748
rect 475102 218736 475108 218748
rect 438360 218708 475108 218736
rect 438360 218696 438366 218708
rect 475102 218696 475108 218708
rect 475160 218696 475166 218748
rect 475672 218736 475700 218844
rect 485406 218832 485412 218844
rect 485464 218832 485470 218884
rect 485746 218872 485774 218980
rect 485866 218968 485872 219020
rect 485924 219008 485930 219020
rect 491294 219008 491300 219020
rect 485924 218980 491300 219008
rect 485924 218968 485930 218980
rect 491294 218968 491300 218980
rect 491352 218968 491358 219020
rect 498378 218968 498384 219020
rect 498436 219008 498442 219020
rect 524322 219008 524328 219020
rect 498436 218980 524328 219008
rect 498436 218968 498442 218980
rect 524322 218968 524328 218980
rect 524380 218968 524386 219020
rect 552198 218968 552204 219020
rect 552256 219008 552262 219020
rect 552382 219008 552388 219020
rect 552256 218980 552388 219008
rect 552256 218968 552262 218980
rect 552382 218968 552388 218980
rect 552440 219008 552446 219020
rect 558178 219008 558184 219020
rect 552440 218980 558184 219008
rect 552440 218968 552446 218980
rect 558178 218968 558184 218980
rect 558236 218968 558242 219020
rect 558380 219008 558408 219116
rect 561766 219104 561772 219156
rect 561824 219144 561830 219156
rect 562318 219144 562324 219156
rect 561824 219116 562324 219144
rect 561824 219104 561830 219116
rect 562318 219104 562324 219116
rect 562376 219144 562382 219156
rect 567470 219144 567476 219156
rect 562376 219116 567476 219144
rect 562376 219104 562382 219116
rect 567470 219104 567476 219116
rect 567528 219104 567534 219156
rect 567654 219104 567660 219156
rect 567712 219144 567718 219156
rect 574922 219144 574928 219156
rect 567712 219116 574928 219144
rect 567712 219104 567718 219116
rect 574922 219104 574928 219116
rect 574980 219104 574986 219156
rect 567838 219008 567844 219020
rect 558380 218980 567844 219008
rect 567838 218968 567844 218980
rect 567896 218968 567902 219020
rect 568022 218968 568028 219020
rect 568080 219008 568086 219020
rect 575290 219008 575296 219020
rect 568080 218980 575296 219008
rect 568080 218968 568086 218980
rect 575290 218968 575296 218980
rect 575348 218968 575354 219020
rect 529566 218872 529572 218884
rect 485746 218844 529572 218872
rect 529566 218832 529572 218844
rect 529624 218832 529630 218884
rect 530578 218832 530584 218884
rect 530636 218872 530642 218884
rect 596082 218872 596088 218884
rect 530636 218844 596088 218872
rect 530636 218832 530642 218844
rect 596082 218832 596088 218844
rect 596140 218832 596146 218884
rect 481174 218736 481180 218748
rect 475580 218708 475700 218736
rect 480272 218708 481180 218736
rect 254394 218628 254400 218680
rect 254452 218668 254458 218680
rect 256142 218668 256148 218680
rect 254452 218640 256148 218668
rect 254452 218628 254458 218640
rect 256142 218628 256148 218640
rect 256200 218628 256206 218680
rect 475580 218668 475608 218708
rect 475442 218640 475608 218668
rect 200040 218572 205634 218600
rect 205606 218532 205634 218572
rect 207842 218560 207848 218612
rect 207900 218600 207906 218612
rect 244918 218600 244924 218612
rect 207900 218572 244924 218600
rect 207900 218560 207906 218572
rect 244918 218560 244924 218572
rect 244976 218560 244982 218612
rect 324774 218560 324780 218612
rect 324832 218600 324838 218612
rect 326062 218600 326068 218612
rect 324832 218572 326068 218600
rect 324832 218560 324838 218572
rect 326062 218560 326068 218572
rect 326120 218560 326126 218612
rect 349154 218560 349160 218612
rect 349212 218600 349218 218612
rect 355318 218600 355324 218612
rect 349212 218572 355324 218600
rect 349212 218560 349218 218572
rect 355318 218560 355324 218572
rect 355376 218560 355382 218612
rect 357158 218560 357164 218612
rect 357216 218600 357222 218612
rect 366910 218600 366916 218612
rect 357216 218572 366916 218600
rect 357216 218560 357222 218572
rect 366910 218560 366916 218572
rect 366968 218560 366974 218612
rect 421834 218560 421840 218612
rect 421892 218600 421898 218612
rect 446398 218600 446404 218612
rect 421892 218572 446404 218600
rect 421892 218560 421898 218572
rect 446398 218560 446404 218572
rect 446456 218560 446462 218612
rect 450538 218560 450544 218612
rect 450596 218600 450602 218612
rect 457162 218600 457168 218612
rect 450596 218572 457168 218600
rect 450596 218560 450602 218572
rect 457162 218560 457168 218572
rect 457220 218560 457226 218612
rect 459002 218560 459008 218612
rect 459060 218600 459066 218612
rect 469582 218600 469588 218612
rect 459060 218572 469588 218600
rect 459060 218560 459066 218572
rect 469582 218560 469588 218572
rect 469640 218560 469646 218612
rect 475442 218600 475470 218640
rect 470566 218572 475470 218600
rect 206094 218532 206100 218544
rect 205606 218504 206100 218532
rect 206094 218492 206100 218504
rect 206152 218492 206158 218544
rect 256050 218492 256056 218544
rect 256108 218532 256114 218544
rect 262858 218532 262864 218544
rect 256108 218504 262864 218532
rect 256108 218492 256114 218504
rect 262858 218492 262864 218504
rect 262916 218492 262922 218544
rect 152458 218464 152464 218476
rect 151280 218436 152464 218464
rect 152458 218424 152464 218436
rect 152516 218424 152522 218476
rect 153212 218436 156184 218464
rect 89438 218288 89444 218340
rect 89496 218328 89502 218340
rect 89496 218300 93854 218328
rect 89496 218288 89502 218300
rect 55674 218152 55680 218204
rect 55732 218192 55738 218204
rect 57238 218192 57244 218204
rect 55732 218164 57244 218192
rect 55732 218152 55738 218164
rect 57238 218152 57244 218164
rect 57296 218152 57302 218204
rect 66438 218152 66444 218204
rect 66496 218192 66502 218204
rect 69566 218192 69572 218204
rect 66496 218164 69572 218192
rect 66496 218152 66502 218164
rect 69566 218152 69572 218164
rect 69624 218152 69630 218204
rect 90450 218152 90456 218204
rect 90508 218192 90514 218204
rect 93826 218192 93854 218300
rect 95418 218288 95424 218340
rect 95476 218328 95482 218340
rect 96246 218328 96252 218340
rect 95476 218300 96252 218328
rect 95476 218288 95482 218300
rect 96246 218288 96252 218300
rect 96304 218288 96310 218340
rect 103698 218288 103704 218340
rect 103756 218328 103762 218340
rect 153212 218328 153240 218436
rect 103756 218300 153240 218328
rect 103756 218288 103762 218300
rect 153378 218288 153384 218340
rect 153436 218328 153442 218340
rect 154114 218328 154120 218340
rect 153436 218300 154120 218328
rect 153436 218288 153442 218300
rect 154114 218288 154120 218300
rect 154172 218288 154178 218340
rect 155034 218288 155040 218340
rect 155092 218328 155098 218340
rect 155954 218328 155960 218340
rect 155092 218300 155960 218328
rect 155092 218288 155098 218300
rect 155954 218288 155960 218300
rect 156012 218288 156018 218340
rect 156156 218328 156184 218436
rect 156690 218424 156696 218476
rect 156748 218464 156754 218476
rect 161290 218464 161296 218476
rect 156748 218436 161296 218464
rect 156748 218424 156754 218436
rect 161290 218424 161296 218436
rect 161348 218424 161354 218476
rect 161474 218424 161480 218476
rect 161532 218464 161538 218476
rect 183554 218464 183560 218476
rect 161532 218436 183560 218464
rect 161532 218424 161538 218436
rect 183554 218424 183560 218436
rect 183612 218424 183618 218476
rect 205450 218464 205456 218476
rect 183940 218436 205456 218464
rect 158990 218328 158996 218340
rect 156156 218300 158996 218328
rect 158990 218288 158996 218300
rect 159048 218288 159054 218340
rect 159174 218288 159180 218340
rect 159232 218328 159238 218340
rect 160002 218328 160008 218340
rect 159232 218300 160008 218328
rect 159232 218288 159238 218300
rect 160002 218288 160008 218300
rect 160060 218288 160066 218340
rect 160186 218288 160192 218340
rect 160244 218328 160250 218340
rect 164786 218328 164792 218340
rect 160244 218300 164792 218328
rect 160244 218288 160250 218300
rect 164786 218288 164792 218300
rect 164844 218288 164850 218340
rect 166626 218288 166632 218340
rect 166684 218328 166690 218340
rect 166684 218300 178172 218328
rect 166684 218288 166690 218300
rect 164970 218220 164976 218272
rect 165028 218260 165034 218272
rect 166258 218260 166264 218272
rect 165028 218232 166264 218260
rect 165028 218220 165034 218232
rect 166258 218220 166264 218232
rect 166316 218220 166322 218272
rect 161474 218192 161480 218204
rect 90508 218164 93762 218192
rect 93826 218164 161480 218192
rect 90508 218152 90514 218164
rect 57330 218016 57336 218068
rect 57388 218056 57394 218068
rect 57882 218056 57888 218068
rect 57388 218028 57888 218056
rect 57388 218016 57394 218028
rect 57882 218016 57888 218028
rect 57940 218016 57946 218068
rect 58158 218016 58164 218068
rect 58216 218056 58222 218068
rect 59354 218056 59360 218068
rect 58216 218028 59360 218056
rect 58216 218016 58222 218028
rect 59354 218016 59360 218028
rect 59412 218016 59418 218068
rect 61470 218016 61476 218068
rect 61528 218056 61534 218068
rect 62022 218056 62028 218068
rect 61528 218028 62028 218056
rect 61528 218016 61534 218028
rect 62022 218016 62028 218028
rect 62080 218016 62086 218068
rect 62298 218016 62304 218068
rect 62356 218056 62362 218068
rect 63402 218056 63408 218068
rect 62356 218028 63408 218056
rect 62356 218016 62362 218028
rect 63402 218016 63408 218028
rect 63460 218016 63466 218068
rect 63954 218016 63960 218068
rect 64012 218056 64018 218068
rect 64782 218056 64788 218068
rect 64012 218028 64788 218056
rect 64012 218016 64018 218028
rect 64782 218016 64788 218028
rect 64840 218016 64846 218068
rect 65610 218016 65616 218068
rect 65668 218056 65674 218068
rect 66162 218056 66168 218068
rect 65668 218028 66168 218056
rect 65668 218016 65674 218028
rect 66162 218016 66168 218028
rect 66220 218016 66226 218068
rect 68094 218016 68100 218068
rect 68152 218056 68158 218068
rect 68738 218056 68744 218068
rect 68152 218028 68744 218056
rect 68152 218016 68158 218028
rect 68738 218016 68744 218028
rect 68796 218016 68802 218068
rect 72234 218016 72240 218068
rect 72292 218056 72298 218068
rect 73706 218056 73712 218068
rect 72292 218028 73712 218056
rect 72292 218016 72298 218028
rect 73706 218016 73712 218028
rect 73764 218016 73770 218068
rect 74718 218016 74724 218068
rect 74776 218056 74782 218068
rect 75546 218056 75552 218068
rect 74776 218028 75552 218056
rect 74776 218016 74782 218028
rect 75546 218016 75552 218028
rect 75604 218016 75610 218068
rect 82170 218016 82176 218068
rect 82228 218056 82234 218068
rect 82722 218056 82728 218068
rect 82228 218028 82728 218056
rect 82228 218016 82234 218028
rect 82722 218016 82728 218028
rect 82780 218016 82786 218068
rect 84654 218016 84660 218068
rect 84712 218056 84718 218068
rect 85298 218056 85304 218068
rect 84712 218028 85304 218056
rect 84712 218016 84718 218028
rect 85298 218016 85304 218028
rect 85356 218016 85362 218068
rect 88794 218016 88800 218068
rect 88852 218056 88858 218068
rect 89622 218056 89628 218068
rect 88852 218028 89628 218056
rect 88852 218016 88858 218028
rect 89622 218016 89628 218028
rect 89680 218016 89686 218068
rect 92934 218016 92940 218068
rect 92992 218056 92998 218068
rect 93578 218056 93584 218068
rect 92992 218028 93584 218056
rect 92992 218016 92998 218028
rect 93578 218016 93584 218028
rect 93636 218016 93642 218068
rect 93734 218056 93762 218164
rect 161474 218152 161480 218164
rect 161532 218152 161538 218204
rect 163314 218152 163320 218204
rect 163372 218192 163378 218204
rect 164602 218192 164608 218204
rect 163372 218164 164608 218192
rect 163372 218152 163378 218164
rect 164602 218152 164608 218164
rect 164660 218152 164666 218204
rect 169110 218152 169116 218204
rect 169168 218192 169174 218204
rect 173894 218192 173900 218204
rect 169168 218164 173900 218192
rect 169168 218152 169174 218164
rect 173894 218152 173900 218164
rect 173952 218152 173958 218204
rect 175734 218152 175740 218204
rect 175792 218192 175798 218204
rect 176562 218192 176568 218204
rect 175792 218164 176568 218192
rect 175792 218152 175798 218164
rect 176562 218152 176568 218164
rect 176620 218152 176626 218204
rect 178144 218192 178172 218300
rect 178402 218288 178408 218340
rect 178460 218328 178466 218340
rect 183940 218328 183968 218436
rect 205450 218424 205456 218436
rect 205508 218424 205514 218476
rect 206370 218424 206376 218476
rect 206428 218464 206434 218476
rect 214098 218464 214104 218476
rect 206428 218436 214104 218464
rect 206428 218424 206434 218436
rect 214098 218424 214104 218436
rect 214156 218424 214162 218476
rect 216306 218424 216312 218476
rect 216364 218464 216370 218476
rect 224218 218464 224224 218476
rect 216364 218436 224224 218464
rect 216364 218424 216370 218436
rect 224218 218424 224224 218436
rect 224276 218424 224282 218476
rect 224402 218424 224408 218476
rect 224460 218464 224466 218476
rect 253842 218464 253848 218476
rect 224460 218436 253848 218464
rect 224460 218424 224466 218436
rect 253842 218424 253848 218436
rect 253900 218424 253906 218476
rect 434162 218424 434168 218476
rect 434220 218464 434226 218476
rect 450538 218464 450544 218476
rect 434220 218436 450544 218464
rect 434220 218424 434226 218436
rect 450538 218424 450544 218436
rect 450596 218424 450602 218476
rect 458634 218424 458640 218476
rect 458692 218464 458698 218476
rect 468754 218464 468760 218476
rect 458692 218436 468760 218464
rect 458692 218424 458698 218436
rect 468754 218424 468760 218436
rect 468812 218424 468818 218476
rect 196250 218328 196256 218340
rect 178460 218300 183968 218328
rect 185596 218300 196256 218328
rect 178460 218288 178466 218300
rect 185596 218192 185624 218300
rect 196250 218288 196256 218300
rect 196308 218288 196314 218340
rect 196434 218288 196440 218340
rect 196492 218328 196498 218340
rect 200206 218328 200212 218340
rect 196492 218300 200212 218328
rect 196492 218288 196498 218300
rect 200206 218288 200212 218300
rect 200264 218288 200270 218340
rect 201402 218288 201408 218340
rect 201460 218328 201466 218340
rect 205450 218328 205456 218340
rect 201460 218300 205456 218328
rect 201460 218288 201466 218300
rect 205450 218288 205456 218300
rect 205508 218288 205514 218340
rect 205634 218288 205640 218340
rect 205692 218328 205698 218340
rect 242158 218328 242164 218340
rect 205692 218300 242164 218328
rect 205692 218288 205698 218300
rect 242158 218288 242164 218300
rect 242216 218288 242222 218340
rect 243538 218288 243544 218340
rect 243596 218328 243602 218340
rect 249058 218328 249064 218340
rect 243596 218300 249064 218328
rect 243596 218288 243602 218300
rect 249058 218288 249064 218300
rect 249116 218288 249122 218340
rect 436278 218288 436284 218340
rect 436336 218328 436342 218340
rect 441430 218328 441436 218340
rect 436336 218300 441436 218328
rect 436336 218288 436342 218300
rect 441430 218288 441436 218300
rect 441488 218288 441494 218340
rect 459830 218288 459836 218340
rect 459888 218328 459894 218340
rect 462958 218328 462964 218340
rect 459888 218300 462964 218328
rect 459888 218288 459894 218300
rect 462958 218288 462964 218300
rect 463016 218288 463022 218340
rect 464798 218288 464804 218340
rect 464856 218328 464862 218340
rect 470566 218328 470594 218572
rect 475746 218560 475752 218612
rect 475804 218600 475810 218612
rect 480272 218600 480300 218708
rect 481174 218696 481180 218708
rect 481232 218696 481238 218748
rect 482646 218696 482652 218748
rect 482704 218736 482710 218748
rect 486970 218736 486976 218748
rect 482704 218708 486976 218736
rect 482704 218696 482710 218708
rect 486970 218696 486976 218708
rect 487028 218696 487034 218748
rect 487890 218696 487896 218748
rect 487948 218736 487954 218748
rect 490374 218736 490380 218748
rect 487948 218708 490380 218736
rect 487948 218696 487954 218708
rect 490374 218696 490380 218708
rect 490432 218696 490438 218748
rect 491294 218696 491300 218748
rect 491352 218736 491358 218748
rect 498378 218736 498384 218748
rect 491352 218708 498384 218736
rect 491352 218696 491358 218708
rect 498378 218696 498384 218708
rect 498436 218696 498442 218748
rect 498746 218696 498752 218748
rect 498804 218736 498810 218748
rect 554682 218736 554688 218748
rect 498804 218708 554688 218736
rect 498804 218696 498810 218708
rect 554682 218696 554688 218708
rect 554740 218696 554746 218748
rect 558178 218696 558184 218748
rect 558236 218736 558242 218748
rect 567654 218736 567660 218748
rect 558236 218708 567660 218736
rect 558236 218696 558242 218708
rect 567654 218696 567660 218708
rect 567712 218696 567718 218748
rect 567838 218696 567844 218748
rect 567896 218736 567902 218748
rect 625062 218736 625068 218748
rect 567896 218708 625068 218736
rect 567896 218696 567902 218708
rect 625062 218696 625068 218708
rect 625120 218696 625126 218748
rect 475804 218572 480300 218600
rect 475804 218560 475810 218572
rect 480438 218560 480444 218612
rect 480496 218600 480502 218612
rect 502978 218600 502984 218612
rect 480496 218572 502984 218600
rect 480496 218560 480502 218572
rect 502978 218560 502984 218572
rect 503036 218560 503042 218612
rect 542354 218560 542360 218612
rect 542412 218600 542418 218612
rect 623314 218600 623320 218612
rect 542412 218572 623320 218600
rect 542412 218560 542418 218572
rect 623314 218560 623320 218572
rect 623372 218560 623378 218612
rect 472618 218424 472624 218476
rect 472676 218464 472682 218476
rect 490328 218464 490334 218476
rect 472676 218436 490334 218464
rect 472676 218424 472682 218436
rect 490328 218424 490334 218436
rect 490386 218424 490392 218476
rect 491294 218424 491300 218476
rect 491352 218464 491358 218476
rect 497734 218464 497740 218476
rect 491352 218436 497740 218464
rect 491352 218424 491358 218436
rect 497734 218424 497740 218436
rect 497792 218464 497798 218476
rect 498746 218464 498752 218476
rect 497792 218436 498752 218464
rect 497792 218424 497798 218436
rect 498746 218424 498752 218436
rect 498804 218424 498810 218476
rect 540054 218424 540060 218476
rect 540112 218464 540118 218476
rect 601694 218464 601700 218476
rect 540112 218436 601700 218464
rect 540112 218424 540118 218436
rect 601694 218424 601700 218436
rect 601752 218424 601758 218476
rect 490484 218368 490696 218396
rect 464856 218300 470594 218328
rect 464856 218288 464862 218300
rect 474918 218288 474924 218340
rect 474976 218328 474982 218340
rect 482002 218328 482008 218340
rect 474976 218300 482008 218328
rect 474976 218288 474982 218300
rect 482002 218288 482008 218300
rect 482060 218288 482066 218340
rect 482186 218288 482192 218340
rect 482244 218328 482250 218340
rect 490484 218328 490512 218368
rect 482244 218300 490512 218328
rect 490668 218328 490696 218368
rect 491938 218328 491944 218340
rect 490668 218300 491944 218328
rect 482244 218288 482250 218300
rect 491938 218288 491944 218300
rect 491996 218328 492002 218340
rect 503346 218328 503352 218340
rect 491996 218300 503352 218328
rect 491996 218288 492002 218300
rect 503346 218288 503352 218300
rect 503404 218288 503410 218340
rect 534994 218288 535000 218340
rect 535052 218328 535058 218340
rect 608502 218328 608508 218340
rect 535052 218300 608508 218328
rect 535052 218288 535058 218300
rect 608502 218288 608508 218300
rect 608560 218288 608566 218340
rect 178144 218164 185624 218192
rect 185762 218152 185768 218204
rect 185820 218192 185826 218204
rect 215202 218192 215208 218204
rect 185820 218164 215208 218192
rect 185820 218152 185826 218164
rect 215202 218152 215208 218164
rect 215260 218152 215266 218204
rect 215478 218152 215484 218204
rect 215536 218192 215542 218204
rect 216490 218192 216496 218204
rect 215536 218164 216496 218192
rect 215536 218152 215542 218164
rect 216490 218152 216496 218164
rect 216548 218152 216554 218204
rect 218790 218152 218796 218204
rect 218848 218192 218854 218204
rect 219342 218192 219348 218204
rect 218848 218164 219348 218192
rect 218848 218152 218854 218164
rect 219342 218152 219348 218164
rect 219400 218152 219406 218204
rect 219618 218152 219624 218204
rect 219676 218192 219682 218204
rect 220354 218192 220360 218204
rect 219676 218164 220360 218192
rect 219676 218152 219682 218164
rect 220354 218152 220360 218164
rect 220412 218152 220418 218204
rect 222930 218152 222936 218204
rect 222988 218192 222994 218204
rect 224402 218192 224408 218204
rect 222988 218164 224408 218192
rect 222988 218152 222994 218164
rect 224402 218152 224408 218164
rect 224460 218152 224466 218204
rect 225414 218152 225420 218204
rect 225472 218192 225478 218204
rect 226058 218192 226064 218204
rect 225472 218164 226064 218192
rect 225472 218152 225478 218164
rect 226058 218152 226064 218164
rect 226116 218152 226122 218204
rect 236638 218192 236644 218204
rect 229066 218164 236644 218192
rect 161658 218084 161664 218136
rect 161716 218124 161722 218136
rect 162486 218124 162492 218136
rect 161716 218096 162492 218124
rect 161716 218084 161722 218096
rect 162486 218084 162492 218096
rect 162544 218084 162550 218136
rect 165798 218084 165804 218136
rect 165856 218124 165862 218136
rect 166810 218124 166816 218136
rect 165856 218096 166816 218124
rect 165856 218084 165862 218096
rect 166810 218084 166816 218096
rect 166868 218084 166874 218136
rect 177390 218084 177396 218136
rect 177448 218124 177454 218136
rect 177942 218124 177948 218136
rect 177448 218096 177948 218124
rect 177448 218084 177454 218096
rect 177942 218084 177948 218096
rect 178000 218084 178006 218136
rect 93734 218028 96660 218056
rect 96632 217852 96660 218028
rect 98730 218016 98736 218068
rect 98788 218056 98794 218068
rect 99282 218056 99288 218068
rect 98788 218028 99288 218056
rect 98788 218016 98794 218028
rect 99282 218016 99288 218028
rect 99340 218016 99346 218068
rect 99558 218016 99564 218068
rect 99616 218056 99622 218068
rect 100662 218056 100668 218068
rect 99616 218028 100668 218056
rect 99616 218016 99622 218028
rect 100662 218016 100668 218028
rect 100720 218016 100726 218068
rect 101214 218016 101220 218068
rect 101272 218056 101278 218068
rect 103422 218056 103428 218068
rect 101272 218028 103428 218056
rect 101272 218016 101278 218028
rect 103422 218016 103428 218028
rect 103480 218016 103486 218068
rect 105354 218016 105360 218068
rect 105412 218056 105418 218068
rect 106182 218056 106188 218068
rect 105412 218028 106188 218056
rect 105412 218016 105418 218028
rect 106182 218016 106188 218028
rect 106240 218016 106246 218068
rect 107010 218016 107016 218068
rect 107068 218056 107074 218068
rect 107562 218056 107568 218068
rect 107068 218028 107568 218056
rect 107068 218016 107074 218028
rect 107562 218016 107568 218028
rect 107620 218016 107626 218068
rect 109494 218016 109500 218068
rect 109552 218056 109558 218068
rect 110322 218056 110328 218068
rect 109552 218028 110328 218056
rect 109552 218016 109558 218028
rect 110322 218016 110328 218028
rect 110380 218016 110386 218068
rect 111150 218016 111156 218068
rect 111208 218056 111214 218068
rect 111702 218056 111708 218068
rect 111208 218028 111708 218056
rect 111208 218016 111214 218028
rect 111702 218016 111708 218028
rect 111760 218016 111766 218068
rect 112806 218016 112812 218068
rect 112864 218056 112870 218068
rect 112864 218028 113174 218056
rect 112864 218016 112870 218028
rect 113146 217988 113174 218028
rect 181530 218016 181536 218068
rect 181588 218056 181594 218068
rect 182818 218056 182824 218068
rect 181588 218028 182824 218056
rect 181588 218016 181594 218028
rect 182818 218016 182824 218028
rect 182876 218016 182882 218068
rect 183002 218016 183008 218068
rect 183060 218056 183066 218068
rect 183060 218028 185532 218056
rect 183060 218016 183066 218028
rect 113146 217960 180794 217988
rect 180766 217920 180794 217960
rect 185118 217920 185124 217932
rect 180766 217892 185124 217920
rect 185118 217880 185124 217892
rect 185176 217880 185182 217932
rect 185504 217920 185532 218028
rect 185670 218016 185676 218068
rect 185728 218056 185734 218068
rect 186130 218056 186136 218068
rect 185728 218028 186136 218056
rect 185728 218016 185734 218028
rect 186130 218016 186136 218028
rect 186188 218016 186194 218068
rect 188154 218016 188160 218068
rect 188212 218056 188218 218068
rect 188798 218056 188804 218068
rect 188212 218028 188804 218056
rect 188212 218016 188218 218028
rect 188798 218016 188804 218028
rect 188856 218016 188862 218068
rect 189810 218016 189816 218068
rect 189868 218056 189874 218068
rect 229066 218056 229094 218164
rect 236638 218152 236644 218164
rect 236696 218152 236702 218204
rect 274266 218152 274272 218204
rect 274324 218192 274330 218204
rect 275278 218192 275284 218204
rect 274324 218164 275284 218192
rect 274324 218152 274330 218164
rect 275278 218152 275284 218164
rect 275336 218152 275342 218204
rect 277578 218152 277584 218204
rect 277636 218192 277642 218204
rect 281258 218192 281264 218204
rect 277636 218164 281264 218192
rect 277636 218152 277642 218164
rect 281258 218152 281264 218164
rect 281316 218152 281322 218204
rect 290826 218152 290832 218204
rect 290884 218192 290890 218204
rect 293218 218192 293224 218204
rect 290884 218164 293224 218192
rect 290884 218152 290890 218164
rect 293218 218152 293224 218164
rect 293276 218152 293282 218204
rect 306558 218152 306564 218204
rect 306616 218192 306622 218204
rect 313458 218192 313464 218204
rect 306616 218164 313464 218192
rect 306616 218152 306622 218164
rect 313458 218152 313464 218164
rect 313516 218152 313522 218204
rect 318978 218152 318984 218204
rect 319036 218192 319042 218204
rect 323302 218192 323308 218204
rect 319036 218164 323308 218192
rect 319036 218152 319042 218164
rect 323302 218152 323308 218164
rect 323360 218152 323366 218204
rect 327258 218152 327264 218204
rect 327316 218192 327322 218204
rect 329926 218192 329932 218204
rect 327316 218164 329932 218192
rect 327316 218152 327322 218164
rect 329926 218152 329932 218164
rect 329984 218152 329990 218204
rect 339310 218152 339316 218204
rect 339368 218192 339374 218204
rect 342898 218192 342904 218204
rect 339368 218164 342904 218192
rect 339368 218152 339374 218164
rect 342898 218152 342904 218164
rect 342956 218152 342962 218204
rect 346026 218152 346032 218204
rect 346084 218192 346090 218204
rect 352006 218192 352012 218204
rect 346084 218164 352012 218192
rect 346084 218152 346090 218164
rect 352006 218152 352012 218164
rect 352064 218152 352070 218204
rect 361022 218152 361028 218204
rect 361080 218192 361086 218204
rect 361942 218192 361948 218204
rect 361080 218164 361948 218192
rect 361080 218152 361086 218164
rect 361942 218152 361948 218164
rect 362000 218152 362006 218204
rect 449894 218152 449900 218204
rect 449952 218192 449958 218204
rect 490558 218192 490564 218204
rect 449952 218164 490564 218192
rect 449952 218152 449958 218164
rect 490558 218152 490564 218164
rect 490616 218152 490622 218204
rect 490926 218152 490932 218204
rect 490984 218192 490990 218204
rect 493686 218192 493692 218204
rect 490984 218164 493692 218192
rect 490984 218152 490990 218164
rect 493686 218152 493692 218164
rect 493744 218152 493750 218204
rect 493870 218152 493876 218204
rect 493928 218192 493934 218204
rect 496906 218192 496912 218204
rect 493928 218164 496912 218192
rect 493928 218152 493934 218164
rect 496906 218152 496912 218164
rect 496964 218152 496970 218204
rect 532510 218152 532516 218204
rect 532568 218192 532574 218204
rect 597186 218192 597192 218204
rect 532568 218164 597192 218192
rect 532568 218152 532574 218164
rect 597186 218152 597192 218164
rect 597244 218152 597250 218204
rect 189868 218028 229094 218056
rect 189868 218016 189874 218028
rect 231210 218016 231216 218068
rect 231268 218056 231274 218068
rect 231670 218056 231676 218068
rect 231268 218028 231676 218056
rect 231268 218016 231274 218028
rect 231670 218016 231676 218028
rect 231728 218016 231734 218068
rect 232038 218016 232044 218068
rect 232096 218056 232102 218068
rect 233050 218056 233056 218068
rect 232096 218028 233056 218056
rect 232096 218016 232102 218028
rect 233050 218016 233056 218028
rect 233108 218016 233114 218068
rect 235350 218016 235356 218068
rect 235408 218056 235414 218068
rect 235902 218056 235908 218068
rect 235408 218028 235908 218056
rect 235408 218016 235414 218028
rect 235902 218016 235908 218028
rect 235960 218016 235966 218068
rect 239490 218016 239496 218068
rect 239548 218056 239554 218068
rect 240042 218056 240048 218068
rect 239548 218028 240048 218056
rect 239548 218016 239554 218028
rect 240042 218016 240048 218028
rect 240100 218016 240106 218068
rect 241974 218016 241980 218068
rect 242032 218056 242038 218068
rect 242802 218056 242808 218068
rect 242032 218028 242808 218056
rect 242032 218016 242038 218028
rect 242802 218016 242808 218028
rect 242860 218016 242866 218068
rect 243630 218016 243636 218068
rect 243688 218056 243694 218068
rect 244182 218056 244188 218068
rect 243688 218028 244188 218056
rect 243688 218016 243694 218028
rect 244182 218016 244188 218028
rect 244240 218016 244246 218068
rect 244458 218016 244464 218068
rect 244516 218056 244522 218068
rect 245286 218056 245292 218068
rect 244516 218028 245292 218056
rect 244516 218016 244522 218028
rect 245286 218016 245292 218028
rect 245344 218016 245350 218068
rect 246114 218016 246120 218068
rect 246172 218056 246178 218068
rect 247586 218056 247592 218068
rect 246172 218028 247592 218056
rect 246172 218016 246178 218028
rect 247586 218016 247592 218028
rect 247644 218016 247650 218068
rect 248598 218016 248604 218068
rect 248656 218056 248662 218068
rect 249610 218056 249616 218068
rect 248656 218028 249616 218056
rect 248656 218016 248662 218028
rect 249610 218016 249616 218028
rect 249668 218016 249674 218068
rect 250254 218016 250260 218068
rect 250312 218056 250318 218068
rect 251174 218056 251180 218068
rect 250312 218028 251180 218056
rect 250312 218016 250318 218028
rect 251174 218016 251180 218028
rect 251232 218016 251238 218068
rect 261018 218016 261024 218068
rect 261076 218056 261082 218068
rect 261846 218056 261852 218068
rect 261076 218028 261852 218056
rect 261076 218016 261082 218028
rect 261846 218016 261852 218028
rect 261904 218016 261910 218068
rect 265158 218016 265164 218068
rect 265216 218056 265222 218068
rect 266262 218056 266268 218068
rect 265216 218028 266268 218056
rect 265216 218016 265222 218028
rect 266262 218016 266268 218028
rect 266320 218016 266326 218068
rect 266814 218016 266820 218068
rect 266872 218056 266878 218068
rect 267458 218056 267464 218068
rect 266872 218028 267464 218056
rect 266872 218016 266878 218028
rect 267458 218016 267464 218028
rect 267516 218016 267522 218068
rect 270954 218016 270960 218068
rect 271012 218056 271018 218068
rect 271874 218056 271880 218068
rect 271012 218028 271880 218056
rect 271012 218016 271018 218028
rect 271874 218016 271880 218028
rect 271932 218016 271938 218068
rect 272610 218016 272616 218068
rect 272668 218056 272674 218068
rect 273162 218056 273168 218068
rect 272668 218028 273168 218056
rect 272668 218016 272674 218028
rect 273162 218016 273168 218028
rect 273220 218016 273226 218068
rect 273438 218016 273444 218068
rect 273496 218056 273502 218068
rect 274542 218056 274548 218068
rect 273496 218028 274548 218056
rect 273496 218016 273502 218028
rect 274542 218016 274548 218028
rect 274600 218016 274606 218068
rect 275094 218016 275100 218068
rect 275152 218056 275158 218068
rect 275830 218056 275836 218068
rect 275152 218028 275836 218056
rect 275152 218016 275158 218028
rect 275830 218016 275836 218028
rect 275888 218016 275894 218068
rect 276750 218016 276756 218068
rect 276808 218056 276814 218068
rect 277210 218056 277216 218068
rect 276808 218028 277216 218056
rect 276808 218016 276814 218028
rect 277210 218016 277216 218028
rect 277268 218016 277274 218068
rect 279234 218016 279240 218068
rect 279292 218056 279298 218068
rect 279786 218056 279792 218068
rect 279292 218028 279792 218056
rect 279292 218016 279298 218028
rect 279786 218016 279792 218028
rect 279844 218016 279850 218068
rect 281718 218016 281724 218068
rect 281776 218056 281782 218068
rect 282730 218056 282736 218068
rect 281776 218028 282736 218056
rect 281776 218016 281782 218028
rect 282730 218016 282736 218028
rect 282788 218016 282794 218068
rect 285030 218016 285036 218068
rect 285088 218056 285094 218068
rect 285582 218056 285588 218068
rect 285088 218028 285588 218056
rect 285088 218016 285094 218028
rect 285582 218016 285588 218028
rect 285640 218016 285646 218068
rect 287514 218016 287520 218068
rect 287572 218056 287578 218068
rect 288526 218056 288532 218068
rect 287572 218028 288532 218056
rect 287572 218016 287578 218028
rect 288526 218016 288532 218028
rect 288584 218016 288590 218068
rect 289170 218016 289176 218068
rect 289228 218056 289234 218068
rect 289722 218056 289728 218068
rect 289228 218028 289728 218056
rect 289228 218016 289234 218028
rect 289722 218016 289728 218028
rect 289780 218016 289786 218068
rect 289998 218016 290004 218068
rect 290056 218056 290062 218068
rect 291010 218056 291016 218068
rect 290056 218028 291016 218056
rect 290056 218016 290062 218028
rect 291010 218016 291016 218028
rect 291068 218016 291074 218068
rect 291654 218016 291660 218068
rect 291712 218056 291718 218068
rect 292482 218056 292488 218068
rect 291712 218028 292488 218056
rect 291712 218016 291718 218028
rect 292482 218016 292488 218028
rect 292540 218016 292546 218068
rect 293310 218016 293316 218068
rect 293368 218056 293374 218068
rect 293770 218056 293776 218068
rect 293368 218028 293776 218056
rect 293368 218016 293374 218028
rect 293770 218016 293776 218028
rect 293828 218016 293834 218068
rect 294138 218016 294144 218068
rect 294196 218056 294202 218068
rect 294966 218056 294972 218068
rect 294196 218028 294972 218056
rect 294196 218016 294202 218028
rect 294966 218016 294972 218028
rect 295024 218016 295030 218068
rect 299106 218016 299112 218068
rect 299164 218056 299170 218068
rect 303430 218056 303436 218068
rect 299164 218028 303436 218056
rect 299164 218016 299170 218028
rect 303430 218016 303436 218028
rect 303488 218016 303494 218068
rect 304074 218016 304080 218068
rect 304132 218056 304138 218068
rect 304626 218056 304632 218068
rect 304132 218028 304632 218056
rect 304132 218016 304138 218028
rect 304626 218016 304632 218028
rect 304684 218016 304690 218068
rect 308214 218016 308220 218068
rect 308272 218056 308278 218068
rect 308766 218056 308772 218068
rect 308272 218028 308772 218056
rect 308272 218016 308278 218028
rect 308766 218016 308772 218028
rect 308824 218016 308830 218068
rect 309870 218016 309876 218068
rect 309928 218056 309934 218068
rect 310330 218056 310336 218068
rect 309928 218028 310336 218056
rect 309928 218016 309934 218028
rect 310330 218016 310336 218028
rect 310388 218016 310394 218068
rect 312354 218016 312360 218068
rect 312412 218056 312418 218068
rect 313274 218056 313280 218068
rect 312412 218028 313280 218056
rect 312412 218016 312418 218028
rect 313274 218016 313280 218028
rect 313332 218016 313338 218068
rect 314838 218016 314844 218068
rect 314896 218056 314902 218068
rect 315574 218056 315580 218068
rect 314896 218028 315580 218056
rect 314896 218016 314902 218028
rect 315574 218016 315580 218028
rect 315632 218016 315638 218068
rect 316494 218016 316500 218068
rect 316552 218056 316558 218068
rect 317046 218056 317052 218068
rect 316552 218028 317052 218056
rect 316552 218016 316558 218028
rect 317046 218016 317052 218028
rect 317104 218016 317110 218068
rect 322290 218016 322296 218068
rect 322348 218056 322354 218068
rect 322750 218056 322756 218068
rect 322348 218028 322756 218056
rect 322348 218016 322354 218028
rect 322750 218016 322756 218028
rect 322808 218016 322814 218068
rect 326430 218016 326436 218068
rect 326488 218056 326494 218068
rect 327626 218056 327632 218068
rect 326488 218028 327632 218056
rect 326488 218016 326494 218028
rect 327626 218016 327632 218028
rect 327684 218016 327690 218068
rect 328086 218016 328092 218068
rect 328144 218056 328150 218068
rect 328546 218056 328552 218068
rect 328144 218028 328552 218056
rect 328144 218016 328150 218028
rect 328546 218016 328552 218028
rect 328604 218016 328610 218068
rect 328914 218016 328920 218068
rect 328972 218056 328978 218068
rect 330110 218056 330116 218068
rect 328972 218028 330116 218056
rect 328972 218016 328978 218028
rect 330110 218016 330116 218028
rect 330168 218016 330174 218068
rect 330570 218016 330576 218068
rect 330628 218056 330634 218068
rect 331214 218056 331220 218068
rect 330628 218028 331220 218056
rect 330628 218016 330634 218028
rect 331214 218016 331220 218028
rect 331272 218016 331278 218068
rect 332226 218016 332232 218068
rect 332284 218056 332290 218068
rect 332686 218056 332692 218068
rect 332284 218028 332692 218056
rect 332284 218016 332290 218028
rect 332686 218016 332692 218028
rect 332744 218016 332750 218068
rect 336550 218016 336556 218068
rect 336608 218056 336614 218068
rect 339586 218056 339592 218068
rect 336608 218028 339592 218056
rect 336608 218016 336614 218028
rect 339586 218016 339592 218028
rect 339644 218016 339650 218068
rect 346394 218016 346400 218068
rect 346452 218056 346458 218068
rect 350350 218056 350356 218068
rect 346452 218028 350356 218056
rect 346452 218016 346458 218028
rect 350350 218016 350356 218028
rect 350408 218016 350414 218068
rect 358078 218016 358084 218068
rect 358136 218056 358142 218068
rect 360286 218056 360292 218068
rect 358136 218028 360292 218056
rect 358136 218016 358142 218028
rect 360286 218016 360292 218028
rect 360344 218016 360350 218068
rect 361758 218016 361764 218068
rect 361816 218056 361822 218068
rect 363598 218056 363604 218068
rect 361816 218028 363604 218056
rect 361816 218016 361822 218028
rect 363598 218016 363604 218028
rect 363656 218016 363662 218068
rect 374638 218016 374644 218068
rect 374696 218056 374702 218068
rect 378502 218056 378508 218068
rect 374696 218028 378508 218056
rect 374696 218016 374702 218028
rect 378502 218016 378508 218028
rect 378560 218016 378566 218068
rect 387058 218016 387064 218068
rect 387116 218056 387122 218068
rect 388438 218056 388444 218068
rect 387116 218028 388444 218056
rect 387116 218016 387122 218028
rect 388438 218016 388444 218028
rect 388496 218016 388502 218068
rect 429930 218016 429936 218068
rect 429988 218056 429994 218068
rect 430666 218056 430672 218068
rect 429988 218028 430672 218056
rect 429988 218016 429994 218028
rect 430666 218016 430672 218028
rect 430724 218016 430730 218068
rect 430850 218016 430856 218068
rect 430908 218056 430914 218068
rect 431494 218056 431500 218068
rect 430908 218028 431500 218056
rect 430908 218016 430914 218028
rect 431494 218016 431500 218028
rect 431552 218016 431558 218068
rect 432598 218016 432604 218068
rect 432656 218056 432662 218068
rect 435634 218056 435640 218068
rect 432656 218028 435640 218056
rect 432656 218016 432662 218028
rect 435634 218016 435640 218028
rect 435692 218016 435698 218068
rect 446950 218016 446956 218068
rect 447008 218056 447014 218068
rect 449710 218056 449716 218068
rect 447008 218028 449716 218056
rect 447008 218016 447014 218028
rect 449710 218016 449716 218028
rect 449768 218016 449774 218068
rect 471054 218016 471060 218068
rect 471112 218056 471118 218068
rect 477862 218056 477868 218068
rect 471112 218028 477868 218056
rect 471112 218016 471118 218028
rect 477862 218016 477868 218028
rect 477920 218016 477926 218068
rect 479610 218016 479616 218068
rect 479668 218056 479674 218068
rect 504358 218056 504364 218068
rect 479668 218028 504364 218056
rect 479668 218016 479674 218028
rect 504358 218016 504364 218028
rect 504416 218016 504422 218068
rect 549438 218016 549444 218068
rect 549496 218056 549502 218068
rect 567654 218056 567660 218068
rect 549496 218028 567660 218056
rect 549496 218016 549502 218028
rect 567654 218016 567660 218028
rect 567712 218016 567718 218068
rect 574186 218016 574192 218068
rect 574244 218056 574250 218068
rect 614114 218056 614120 218068
rect 574244 218028 614120 218056
rect 574244 218016 574250 218028
rect 614114 218016 614120 218028
rect 614172 218016 614178 218068
rect 527818 217948 527824 218000
rect 527876 217988 527882 218000
rect 528370 217988 528376 218000
rect 527876 217960 528376 217988
rect 527876 217948 527882 217960
rect 528370 217948 528376 217960
rect 528428 217948 528434 218000
rect 543826 217948 543832 218000
rect 543884 217988 543890 218000
rect 545850 217988 545856 218000
rect 543884 217960 545856 217988
rect 543884 217948 543890 217960
rect 545850 217948 545856 217960
rect 545908 217988 545914 218000
rect 545908 217960 548472 217988
rect 545908 217948 545914 217960
rect 185946 217920 185952 217932
rect 185504 217892 185952 217920
rect 185946 217880 185952 217892
rect 186004 217880 186010 217932
rect 205450 217880 205456 217932
rect 205508 217920 205514 217932
rect 205634 217920 205640 217932
rect 205508 217892 205640 217920
rect 205508 217880 205514 217892
rect 205634 217880 205640 217892
rect 205692 217880 205698 217932
rect 486510 217880 486516 217932
rect 486568 217920 486574 217932
rect 492766 217920 492772 217932
rect 486568 217892 492772 217920
rect 486568 217880 486574 217892
rect 492766 217880 492772 217892
rect 492824 217880 492830 217932
rect 548444 217920 548472 217960
rect 567838 217948 567844 218000
rect 567896 217988 567902 218000
rect 570138 217988 570144 218000
rect 567896 217960 570144 217988
rect 567896 217948 567902 217960
rect 570138 217948 570144 217960
rect 570196 217948 570202 218000
rect 548444 217892 553394 217920
rect 167270 217852 167276 217864
rect 96632 217824 167276 217852
rect 167270 217812 167276 217824
rect 167328 217812 167334 217864
rect 167454 217812 167460 217864
rect 167512 217852 167518 217864
rect 172606 217852 172612 217864
rect 167512 217824 172612 217852
rect 167512 217812 167518 217824
rect 172606 217812 172612 217824
rect 172664 217812 172670 217864
rect 176562 217812 176568 217864
rect 176620 217852 176626 217864
rect 180242 217852 180248 217864
rect 176620 217824 180248 217852
rect 176620 217812 176626 217824
rect 180242 217812 180248 217824
rect 180300 217812 180306 217864
rect 397638 217812 397644 217864
rect 397696 217852 397702 217864
rect 398374 217852 398380 217864
rect 397696 217824 398380 217852
rect 397696 217812 397702 217824
rect 398374 217812 398380 217824
rect 398432 217812 398438 217864
rect 530854 217812 530860 217864
rect 530912 217852 530918 217864
rect 548150 217852 548156 217864
rect 530912 217824 548156 217852
rect 530912 217812 530918 217824
rect 548150 217812 548156 217824
rect 548208 217812 548214 217864
rect 553366 217852 553394 217892
rect 601970 217852 601976 217864
rect 553366 217824 601976 217852
rect 601970 217812 601976 217824
rect 602028 217812 602034 217864
rect 134334 217676 134340 217728
rect 134392 217716 134398 217728
rect 199102 217716 199108 217728
rect 134392 217688 199108 217716
rect 134392 217676 134398 217688
rect 199102 217676 199108 217688
rect 199160 217676 199166 217728
rect 445386 217676 445392 217728
rect 445444 217716 445450 217728
rect 456058 217716 456064 217728
rect 445444 217688 456064 217716
rect 445444 217676 445450 217688
rect 456058 217676 456064 217688
rect 456116 217676 456122 217728
rect 528370 217676 528376 217728
rect 528428 217716 528434 217728
rect 596634 217716 596640 217728
rect 528428 217688 596640 217716
rect 528428 217676 528434 217688
rect 596634 217676 596640 217688
rect 596692 217676 596698 217728
rect 596818 217676 596824 217728
rect 596876 217716 596882 217728
rect 608318 217716 608324 217728
rect 596876 217688 608324 217716
rect 596876 217676 596882 217688
rect 608318 217676 608324 217688
rect 608376 217676 608382 217728
rect 608502 217676 608508 217728
rect 608560 217716 608566 217728
rect 621658 217716 621664 217728
rect 608560 217688 621664 217716
rect 608560 217676 608566 217688
rect 621658 217676 621664 217688
rect 621716 217676 621722 217728
rect 122742 217540 122748 217592
rect 122800 217580 122806 217592
rect 192110 217580 192116 217592
rect 122800 217552 192116 217580
rect 122800 217540 122806 217552
rect 192110 217540 192116 217552
rect 192168 217540 192174 217592
rect 444098 217540 444104 217592
rect 444156 217580 444162 217592
rect 501874 217580 501880 217592
rect 444156 217552 501880 217580
rect 444156 217540 444162 217552
rect 501874 217540 501880 217552
rect 501932 217540 501938 217592
rect 548150 217540 548156 217592
rect 548208 217580 548214 217592
rect 601510 217580 601516 217592
rect 548208 217552 601516 217580
rect 548208 217540 548214 217552
rect 601510 217540 601516 217552
rect 601568 217540 601574 217592
rect 601694 217540 601700 217592
rect 601752 217580 601758 217592
rect 622762 217580 622768 217592
rect 601752 217552 622768 217580
rect 601752 217540 601758 217552
rect 622762 217540 622768 217552
rect 622820 217540 622826 217592
rect 106182 217404 106188 217456
rect 106240 217444 106246 217456
rect 181162 217444 181168 217456
rect 106240 217416 181168 217444
rect 106240 217404 106246 217416
rect 181162 217404 181168 217416
rect 181220 217404 181226 217456
rect 456058 217404 456064 217456
rect 456116 217444 456122 217456
rect 504358 217444 504364 217456
rect 456116 217416 504364 217444
rect 456116 217404 456122 217416
rect 504358 217404 504364 217416
rect 504416 217404 504422 217456
rect 555694 217404 555700 217456
rect 555752 217444 555758 217456
rect 555752 217416 570000 217444
rect 555752 217404 555758 217416
rect 449526 217336 449532 217388
rect 449584 217376 449590 217388
rect 449584 217348 451274 217376
rect 449584 217336 449590 217348
rect 178034 217308 178040 217320
rect 103486 217280 178040 217308
rect 102824 217200 102830 217252
rect 102882 217240 102888 217252
rect 103486 217240 103514 217280
rect 178034 217268 178040 217280
rect 178092 217268 178098 217320
rect 451246 217308 451274 217348
rect 451246 217280 509234 217308
rect 102882 217212 103514 217240
rect 102882 217200 102888 217212
rect 203012 217200 203018 217252
rect 203070 217240 203076 217252
rect 207842 217240 207848 217252
rect 203070 217212 207848 217240
rect 203070 217200 203076 217212
rect 207842 217200 207848 217212
rect 207900 217200 207906 217252
rect 361574 217200 361580 217252
rect 361632 217240 361638 217252
rect 362816 217240 362822 217252
rect 361632 217212 362822 217240
rect 361632 217200 361638 217212
rect 362816 217200 362822 217212
rect 362874 217200 362880 217252
rect 373994 217200 374000 217252
rect 374052 217240 374058 217252
rect 375236 217240 375242 217252
rect 374052 217212 375242 217240
rect 374052 217200 374058 217212
rect 375236 217200 375242 217212
rect 375294 217200 375300 217252
rect 402974 217200 402980 217252
rect 403032 217240 403038 217252
rect 404216 217240 404222 217252
rect 403032 217212 404222 217240
rect 403032 217200 403038 217212
rect 404216 217200 404222 217212
rect 404274 217200 404280 217252
rect 419718 217200 419724 217252
rect 419776 217240 419782 217252
rect 420776 217240 420782 217252
rect 419776 217212 420782 217240
rect 419776 217200 419782 217212
rect 420776 217200 420782 217212
rect 420834 217200 420840 217252
rect 509206 217240 509234 217280
rect 509372 217240 509378 217252
rect 509206 217212 509378 217240
rect 509372 217200 509378 217212
rect 509430 217200 509436 217252
rect 510614 217200 510620 217252
rect 510672 217240 510678 217252
rect 511856 217240 511862 217252
rect 510672 217212 511862 217240
rect 510672 217200 510678 217212
rect 511856 217200 511862 217212
rect 511914 217200 511920 217252
rect 518894 217200 518900 217252
rect 518952 217240 518958 217252
rect 520136 217240 520142 217252
rect 518952 217212 520142 217240
rect 518952 217200 518958 217212
rect 520136 217200 520142 217212
rect 520194 217200 520200 217252
rect 523034 217200 523040 217252
rect 523092 217240 523098 217252
rect 524276 217240 524282 217252
rect 523092 217212 524282 217240
rect 523092 217200 523098 217212
rect 524276 217200 524282 217212
rect 524334 217200 524340 217252
rect 524874 217200 524880 217252
rect 524932 217240 524938 217252
rect 529244 217240 529250 217252
rect 524932 217212 529250 217240
rect 524932 217200 524938 217212
rect 529244 217200 529250 217212
rect 529302 217200 529308 217252
rect 544148 217200 544154 217252
rect 544206 217240 544212 217252
rect 544562 217240 544568 217252
rect 544206 217212 544568 217240
rect 544206 217200 544212 217212
rect 544562 217200 544568 217212
rect 544620 217200 544626 217252
rect 552934 217200 552940 217252
rect 552992 217240 552998 217252
rect 558224 217240 558230 217252
rect 552992 217212 558230 217240
rect 552992 217200 552998 217212
rect 558224 217200 558230 217212
rect 558282 217240 558288 217252
rect 567838 217240 567844 217252
rect 558282 217212 567844 217240
rect 558282 217200 558288 217212
rect 567838 217200 567844 217212
rect 567896 217200 567902 217252
rect 568574 217200 568580 217252
rect 568632 217240 568638 217252
rect 569816 217240 569822 217252
rect 568632 217212 569822 217240
rect 568632 217200 568638 217212
rect 569816 217200 569822 217212
rect 569874 217200 569880 217252
rect 569972 217240 570000 217416
rect 570138 217404 570144 217456
rect 570196 217444 570202 217456
rect 596818 217444 596824 217456
rect 570196 217416 596824 217444
rect 570196 217404 570202 217416
rect 596818 217404 596824 217416
rect 596876 217404 596882 217456
rect 597002 217404 597008 217456
rect 597060 217444 597066 217456
rect 601326 217444 601332 217456
rect 597060 217416 601332 217444
rect 597060 217404 597066 217416
rect 601326 217404 601332 217416
rect 601384 217404 601390 217456
rect 601648 217404 601654 217456
rect 601706 217444 601712 217456
rect 620554 217444 620560 217456
rect 601706 217416 620560 217444
rect 601706 217404 601712 217416
rect 620554 217404 620560 217416
rect 620612 217404 620618 217456
rect 672350 217336 672356 217388
rect 672408 217376 672414 217388
rect 672902 217376 672908 217388
rect 672408 217348 672908 217376
rect 672408 217336 672414 217348
rect 672902 217336 672908 217348
rect 672960 217336 672966 217388
rect 609054 217308 609060 217320
rect 576826 217280 609060 217308
rect 576826 217240 576854 217280
rect 609054 217268 609060 217280
rect 609112 217268 609118 217320
rect 628834 217308 628840 217320
rect 615466 217280 628840 217308
rect 569972 217212 576854 217240
rect 167270 217132 167276 217184
rect 167328 217172 167334 217184
rect 171226 217172 171232 217184
rect 167328 217144 171232 217172
rect 167328 217132 167334 217144
rect 171226 217132 171232 217144
rect 171284 217132 171290 217184
rect 451274 217132 451280 217184
rect 451332 217172 451338 217184
rect 452240 217172 452246 217184
rect 451332 217144 452246 217172
rect 451332 217132 451338 217144
rect 452240 217132 452246 217144
rect 452298 217132 452304 217184
rect 456886 217132 456892 217184
rect 456944 217172 456950 217184
rect 458036 217172 458042 217184
rect 456944 217144 458042 217172
rect 456944 217132 456950 217144
rect 458036 217132 458042 217144
rect 458094 217132 458100 217184
rect 469306 217132 469312 217184
rect 469364 217172 469370 217184
rect 470456 217172 470462 217184
rect 469364 217144 470462 217172
rect 469364 217132 469370 217144
rect 470456 217132 470462 217144
rect 470514 217132 470520 217184
rect 477586 217132 477592 217184
rect 477644 217172 477650 217184
rect 478736 217172 478742 217184
rect 477644 217144 478742 217172
rect 477644 217132 477650 217144
rect 478736 217132 478742 217144
rect 478794 217132 478800 217184
rect 498194 217132 498200 217184
rect 498252 217172 498258 217184
rect 499436 217172 499442 217184
rect 498252 217144 499442 217172
rect 498252 217132 498258 217144
rect 499436 217132 499442 217144
rect 499494 217132 499500 217184
rect 597002 217132 597008 217184
rect 597060 217172 597066 217184
rect 615466 217172 615494 217280
rect 628834 217268 628840 217280
rect 628892 217268 628898 217320
rect 597060 217144 615494 217172
rect 597060 217132 597066 217144
rect 483566 217064 483572 217116
rect 483624 217104 483630 217116
rect 488672 217104 488678 217116
rect 483624 217076 488678 217104
rect 483624 217064 483630 217076
rect 488672 217064 488678 217076
rect 488730 217104 488736 217116
rect 491386 217104 491392 217116
rect 488730 217076 491392 217104
rect 488730 217064 488736 217076
rect 491386 217064 491392 217076
rect 491444 217064 491450 217116
rect 523448 217064 523454 217116
rect 523506 217104 523512 217116
rect 523678 217104 523684 217116
rect 523506 217076 523684 217104
rect 523506 217064 523512 217076
rect 523678 217064 523684 217076
rect 523736 217104 523742 217116
rect 523736 217076 596864 217104
rect 523736 217064 523742 217076
rect 596836 217036 596864 217076
rect 601786 217036 601792 217048
rect 596836 217008 601792 217036
rect 601786 216996 601792 217008
rect 601844 216996 601850 217048
rect 574278 216928 574284 216980
rect 574336 216968 574342 216980
rect 621106 216968 621112 216980
rect 574336 216940 592034 216968
rect 574336 216928 574342 216940
rect 592006 216900 592034 216940
rect 605806 216940 621112 216968
rect 597002 216900 597008 216912
rect 592006 216872 597008 216900
rect 597002 216860 597008 216872
rect 597060 216860 597066 216912
rect 597186 216792 597192 216844
rect 597244 216832 597250 216844
rect 605806 216832 605834 216940
rect 621106 216928 621112 216940
rect 621164 216928 621170 216980
rect 670602 216928 670608 216980
rect 670660 216968 670666 216980
rect 675386 216968 675392 216980
rect 670660 216940 675392 216968
rect 670660 216928 670666 216940
rect 675386 216928 675392 216940
rect 675444 216928 675450 216980
rect 597244 216804 605834 216832
rect 597244 216792 597250 216804
rect 609606 216792 609612 216844
rect 609664 216832 609670 216844
rect 615678 216832 615684 216844
rect 609664 216804 615684 216832
rect 609664 216792 609670 216804
rect 615678 216792 615684 216804
rect 615736 216792 615742 216844
rect 596082 216656 596088 216708
rect 596140 216696 596146 216708
rect 601602 216696 601608 216708
rect 596140 216668 601608 216696
rect 596140 216656 596146 216668
rect 601602 216656 601608 216668
rect 601660 216656 601666 216708
rect 601970 216656 601976 216708
rect 602028 216696 602034 216708
rect 606754 216696 606760 216708
rect 602028 216668 606760 216696
rect 602028 216656 602034 216668
rect 606754 216656 606760 216668
rect 606812 216656 606818 216708
rect 574922 216316 574928 216368
rect 574980 216356 574986 216368
rect 625522 216356 625528 216368
rect 574980 216328 625528 216356
rect 574980 216316 574986 216328
rect 625522 216316 625528 216328
rect 625580 216316 625586 216368
rect 575290 216180 575296 216232
rect 575348 216220 575354 216232
rect 627178 216220 627184 216232
rect 575348 216192 627184 216220
rect 575348 216180 575354 216192
rect 627178 216180 627184 216192
rect 627236 216180 627242 216232
rect 673362 216112 673368 216164
rect 673420 216152 673426 216164
rect 675386 216152 675392 216164
rect 673420 216124 675392 216152
rect 673420 216112 673426 216124
rect 675386 216112 675392 216124
rect 675444 216112 675450 216164
rect 574922 216044 574928 216096
rect 574980 216084 574986 216096
rect 628282 216084 628288 216096
rect 574980 216056 628288 216084
rect 574980 216044 574986 216056
rect 628282 216044 628288 216056
rect 628340 216044 628346 216096
rect 671982 215976 671988 216028
rect 672040 215976 672046 216028
rect 574554 215908 574560 215960
rect 574612 215948 574618 215960
rect 627914 215948 627920 215960
rect 574612 215920 627920 215948
rect 574612 215908 574618 215920
rect 627914 215908 627920 215920
rect 627972 215908 627978 215960
rect 672000 215472 672028 215976
rect 672258 215568 672264 215620
rect 672316 215608 672322 215620
rect 672316 215580 672488 215608
rect 672316 215568 672322 215580
rect 672166 215472 672172 215484
rect 672000 215444 672172 215472
rect 672166 215432 672172 215444
rect 672224 215432 672230 215484
rect 672258 215228 672264 215280
rect 672316 215268 672322 215280
rect 672460 215268 672488 215580
rect 672316 215240 672488 215268
rect 672316 215228 672322 215240
rect 672350 215092 672356 215144
rect 672408 215132 672414 215144
rect 672902 215132 672908 215144
rect 672408 215104 672908 215132
rect 672408 215092 672414 215104
rect 672902 215092 672908 215104
rect 672960 215092 672966 215144
rect 35526 214684 35532 214736
rect 35584 214724 35590 214736
rect 39758 214724 39764 214736
rect 35584 214696 39764 214724
rect 35584 214684 35590 214696
rect 39758 214684 39764 214696
rect 39816 214684 39822 214736
rect 575106 214684 575112 214736
rect 575164 214724 575170 214736
rect 612274 214724 612280 214736
rect 575164 214696 612280 214724
rect 575164 214684 575170 214696
rect 612274 214684 612280 214696
rect 612332 214684 612338 214736
rect 574738 214548 574744 214600
rect 574796 214588 574802 214600
rect 574796 214560 605834 214588
rect 574796 214548 574802 214560
rect 597830 214412 597836 214464
rect 597888 214452 597894 214464
rect 598474 214452 598480 214464
rect 597888 214424 598480 214452
rect 597888 214412 597894 214424
rect 598474 214412 598480 214424
rect 598532 214412 598538 214464
rect 598934 214412 598940 214464
rect 598992 214452 598998 214464
rect 599578 214452 599584 214464
rect 598992 214424 599584 214452
rect 598992 214412 598998 214424
rect 599578 214412 599584 214424
rect 599636 214412 599642 214464
rect 600314 214412 600320 214464
rect 600372 214452 600378 214464
rect 601234 214452 601240 214464
rect 600372 214424 601240 214452
rect 600372 214412 600378 214424
rect 601234 214412 601240 214424
rect 601292 214412 601298 214464
rect 605806 214452 605834 214560
rect 609974 214548 609980 214600
rect 610032 214588 610038 214600
rect 610618 214588 610624 214600
rect 610032 214560 610624 214588
rect 610032 214548 610038 214560
rect 610618 214548 610624 214560
rect 610676 214548 610682 214600
rect 618346 214548 618352 214600
rect 618404 214588 618410 214600
rect 618898 214588 618904 214600
rect 618404 214560 618904 214588
rect 618404 214548 618410 214560
rect 618898 214548 618904 214560
rect 618956 214548 618962 214600
rect 624418 214452 624424 214464
rect 605806 214424 624424 214452
rect 624418 214412 624424 214424
rect 624476 214412 624482 214464
rect 35802 214276 35808 214328
rect 35860 214316 35866 214328
rect 40678 214316 40684 214328
rect 35860 214288 40684 214316
rect 35860 214276 35866 214288
rect 40678 214276 40684 214288
rect 40736 214276 40742 214328
rect 35342 213936 35348 213988
rect 35400 213976 35406 213988
rect 40218 213976 40224 213988
rect 35400 213948 40224 213976
rect 35400 213936 35406 213948
rect 40218 213936 40224 213948
rect 40276 213936 40282 213988
rect 625154 213936 625160 213988
rect 625212 213976 625218 213988
rect 626074 213976 626080 213988
rect 625212 213948 626080 213976
rect 625212 213936 625218 213948
rect 626074 213936 626080 213948
rect 626132 213936 626138 213988
rect 632698 213868 632704 213920
rect 632756 213908 632762 213920
rect 633434 213908 633440 213920
rect 632756 213880 633440 213908
rect 632756 213868 632762 213880
rect 633434 213868 633440 213880
rect 633492 213868 633498 213920
rect 637206 213868 637212 213920
rect 637264 213908 637270 213920
rect 650914 213908 650920 213920
rect 637264 213880 650920 213908
rect 637264 213868 637270 213880
rect 650914 213868 650920 213880
rect 650972 213868 650978 213920
rect 608318 213732 608324 213784
rect 608376 213772 608382 213784
rect 609514 213772 609520 213784
rect 608376 213744 609520 213772
rect 608376 213732 608382 213744
rect 609514 213732 609520 213744
rect 609572 213732 609578 213784
rect 638862 213732 638868 213784
rect 638920 213772 638926 213784
rect 652478 213772 652484 213784
rect 638920 213744 652484 213772
rect 638920 213732 638926 213744
rect 652478 213732 652484 213744
rect 652536 213732 652542 213784
rect 673086 213664 673092 213716
rect 673144 213704 673150 213716
rect 675478 213704 675484 213716
rect 673144 213676 675484 213704
rect 673144 213664 673150 213676
rect 675478 213664 675484 213676
rect 675536 213664 675542 213716
rect 639966 213596 639972 213648
rect 640024 213636 640030 213648
rect 652754 213636 652760 213648
rect 640024 213608 652760 213636
rect 640024 213596 640030 213608
rect 652754 213596 652760 213608
rect 652812 213596 652818 213648
rect 638310 213460 638316 213512
rect 638368 213500 638374 213512
rect 651466 213500 651472 213512
rect 638368 213472 651472 213500
rect 638368 213460 638374 213472
rect 651466 213460 651472 213472
rect 651524 213460 651530 213512
rect 629938 213392 629944 213444
rect 629996 213432 630002 213444
rect 633802 213432 633808 213444
rect 629996 213404 633808 213432
rect 629996 213392 630002 213404
rect 633802 213392 633808 213404
rect 633860 213392 633866 213444
rect 575474 213324 575480 213376
rect 575532 213364 575538 213376
rect 594794 213364 594800 213376
rect 575532 213336 594800 213364
rect 575532 213324 575538 213336
rect 594794 213324 594800 213336
rect 594852 213324 594858 213376
rect 636654 213324 636660 213376
rect 636712 213364 636718 213376
rect 650822 213364 650828 213376
rect 636712 213336 650828 213364
rect 636712 213324 636718 213336
rect 650822 213324 650828 213336
rect 650880 213324 650886 213376
rect 672902 213256 672908 213308
rect 672960 213296 672966 213308
rect 675478 213296 675484 213308
rect 672960 213268 675484 213296
rect 672960 213256 672966 213268
rect 675478 213256 675484 213268
rect 675536 213256 675542 213308
rect 574370 213188 574376 213240
rect 574428 213228 574434 213240
rect 629938 213228 629944 213240
rect 574428 213200 629944 213228
rect 574428 213188 574434 213200
rect 629938 213188 629944 213200
rect 629996 213188 630002 213240
rect 635550 213188 635556 213240
rect 635608 213228 635614 213240
rect 650086 213228 650092 213240
rect 635608 213200 650092 213228
rect 635608 213188 635614 213200
rect 650086 213188 650092 213200
rect 650144 213188 650150 213240
rect 641530 213052 641536 213104
rect 641588 213092 641594 213104
rect 651834 213092 651840 213104
rect 641588 213064 651840 213092
rect 641588 213052 641594 213064
rect 651834 213052 651840 213064
rect 651892 213052 651898 213104
rect 39298 213024 39304 213036
rect 38626 212996 39304 213024
rect 35802 212916 35808 212968
rect 35860 212956 35866 212968
rect 38626 212956 38654 212996
rect 39298 212984 39304 212996
rect 39356 212984 39362 213036
rect 35860 212928 38654 212956
rect 35860 212916 35866 212928
rect 640242 212916 640248 212968
rect 640300 212956 640306 212968
rect 651098 212956 651104 212968
rect 640300 212928 651104 212956
rect 640300 212916 640306 212928
rect 651098 212916 651104 212928
rect 651156 212916 651162 212968
rect 631410 212712 631416 212764
rect 631468 212752 631474 212764
rect 632698 212752 632704 212764
rect 631468 212724 632704 212752
rect 631468 212712 631474 212724
rect 632698 212712 632704 212724
rect 632756 212712 632762 212764
rect 35802 212644 35808 212696
rect 35860 212684 35866 212696
rect 39758 212684 39764 212696
rect 35860 212656 39764 212684
rect 35860 212644 35866 212656
rect 39758 212644 39764 212656
rect 39816 212644 39822 212696
rect 42150 212644 42156 212696
rect 42208 212684 42214 212696
rect 50982 212684 50988 212696
rect 42208 212656 50988 212684
rect 42208 212644 42214 212656
rect 50982 212644 50988 212656
rect 51040 212644 51046 212696
rect 41230 212616 41236 212628
rect 40052 212588 41236 212616
rect 35618 212508 35624 212560
rect 35676 212548 35682 212560
rect 40052 212548 40080 212588
rect 41230 212576 41236 212588
rect 41288 212576 41294 212628
rect 35676 212520 40080 212548
rect 35676 212508 35682 212520
rect 647234 212372 647240 212424
rect 647292 212412 647298 212424
rect 648154 212412 648160 212424
rect 647292 212384 648160 212412
rect 647292 212372 647298 212384
rect 648154 212372 648160 212384
rect 648212 212372 648218 212424
rect 659654 212372 659660 212424
rect 659712 212412 659718 212424
rect 660298 212412 660304 212424
rect 659712 212384 660304 212412
rect 659712 212372 659718 212384
rect 660298 212372 660304 212384
rect 660356 212372 660362 212424
rect 661310 212372 661316 212424
rect 661368 212412 661374 212424
rect 661954 212412 661960 212424
rect 661368 212384 661960 212412
rect 661368 212372 661374 212384
rect 661954 212372 661960 212384
rect 662012 212372 662018 212424
rect 662414 212372 662420 212424
rect 662472 212412 662478 212424
rect 663058 212412 663064 212424
rect 662472 212384 663064 212412
rect 662472 212372 662478 212384
rect 663058 212372 663064 212384
rect 663116 212372 663122 212424
rect 670970 212032 670976 212084
rect 671028 212072 671034 212084
rect 675478 212072 675484 212084
rect 671028 212044 675484 212072
rect 671028 212032 671034 212044
rect 675478 212032 675484 212044
rect 675536 212032 675542 212084
rect 35802 211556 35808 211608
rect 35860 211596 35866 211608
rect 41230 211596 41236 211608
rect 35860 211568 41236 211596
rect 35860 211556 35866 211568
rect 41230 211556 41236 211568
rect 41288 211556 41294 211608
rect 39666 211392 39672 211404
rect 36004 211364 39672 211392
rect 35802 211284 35808 211336
rect 35860 211324 35866 211336
rect 36004 211324 36032 211364
rect 39666 211352 39672 211364
rect 39724 211352 39730 211404
rect 35860 211296 36032 211324
rect 35860 211284 35866 211296
rect 578326 211284 578332 211336
rect 578384 211324 578390 211336
rect 580626 211324 580632 211336
rect 578384 211296 580632 211324
rect 578384 211284 578390 211296
rect 580626 211284 580632 211296
rect 580684 211284 580690 211336
rect 41046 211256 41052 211268
rect 36096 211228 41052 211256
rect 35618 211148 35624 211200
rect 35676 211188 35682 211200
rect 35676 211160 36032 211188
rect 35676 211148 35682 211160
rect 36004 211120 36032 211160
rect 36096 211120 36124 211228
rect 41046 211216 41052 211228
rect 41104 211216 41110 211268
rect 36004 211092 36124 211120
rect 644474 211012 644480 211064
rect 644532 211052 644538 211064
rect 644842 211052 644848 211064
rect 644532 211024 644848 211052
rect 644532 211012 644538 211024
rect 644842 211012 644848 211024
rect 644900 211012 644906 211064
rect 663794 211012 663800 211064
rect 663852 211052 663858 211064
rect 664162 211052 664168 211064
rect 663852 211024 664168 211052
rect 663852 211012 663858 211024
rect 664162 211012 664168 211024
rect 664220 211012 664226 211064
rect 661770 210672 661776 210724
rect 661828 210712 661834 210724
rect 672534 210712 672540 210724
rect 661828 210684 672540 210712
rect 661828 210672 661834 210684
rect 672534 210672 672540 210684
rect 672592 210672 672598 210724
rect 652202 210536 652208 210588
rect 652260 210576 652266 210588
rect 667290 210576 667296 210588
rect 652260 210548 667296 210576
rect 652260 210536 652266 210548
rect 667290 210536 667296 210548
rect 667348 210536 667354 210588
rect 652018 210400 652024 210452
rect 652076 210440 652082 210452
rect 673914 210440 673920 210452
rect 652076 210412 673920 210440
rect 652076 210400 652082 210412
rect 673914 210400 673920 210412
rect 673972 210400 673978 210452
rect 662138 210264 662144 210316
rect 662196 210304 662202 210316
rect 667474 210304 667480 210316
rect 662196 210276 667480 210304
rect 662196 210264 662202 210276
rect 667474 210264 667480 210276
rect 667532 210264 667538 210316
rect 579522 210060 579528 210112
rect 579580 210100 579586 210112
rect 582282 210100 582288 210112
rect 579580 210072 582288 210100
rect 579580 210060 579586 210072
rect 582282 210060 582288 210072
rect 582340 210060 582346 210112
rect 597554 210060 597560 210112
rect 597612 210100 597618 210112
rect 597922 210100 597928 210112
rect 597612 210072 597928 210100
rect 597612 210060 597618 210072
rect 597922 210060 597928 210072
rect 597980 210060 597986 210112
rect 35618 209924 35624 209976
rect 35676 209964 35682 209976
rect 41690 209964 41696 209976
rect 35676 209936 41696 209964
rect 35676 209924 35682 209936
rect 41690 209924 41696 209936
rect 41748 209924 41754 209976
rect 35802 209788 35808 209840
rect 35860 209828 35866 209840
rect 40034 209828 40040 209840
rect 35860 209800 40040 209828
rect 35860 209788 35866 209800
rect 40034 209788 40040 209800
rect 40092 209788 40098 209840
rect 591298 209788 591304 209840
rect 591356 209828 591362 209840
rect 632146 209828 632152 209840
rect 591356 209800 632152 209828
rect 591356 209788 591362 209800
rect 632146 209788 632152 209800
rect 632204 209788 632210 209840
rect 672258 209380 672264 209432
rect 672316 209380 672322 209432
rect 672276 208956 672304 209380
rect 672258 208904 672264 208956
rect 672316 208904 672322 208956
rect 35802 208632 35808 208684
rect 35860 208672 35866 208684
rect 35860 208644 38654 208672
rect 35860 208632 35866 208644
rect 38626 208604 38654 208644
rect 39666 208604 39672 208616
rect 38626 208576 39672 208604
rect 39666 208564 39672 208576
rect 39724 208564 39730 208616
rect 35618 208360 35624 208412
rect 35676 208400 35682 208412
rect 39574 208400 39580 208412
rect 35676 208372 39580 208400
rect 35676 208360 35682 208372
rect 39574 208360 39580 208372
rect 39632 208360 39638 208412
rect 578878 208224 578884 208276
rect 578936 208264 578942 208276
rect 589458 208264 589464 208276
rect 578936 208236 589464 208264
rect 578936 208224 578942 208236
rect 589458 208224 589464 208236
rect 589516 208224 589522 208276
rect 35802 207272 35808 207324
rect 35860 207312 35866 207324
rect 39758 207312 39764 207324
rect 35860 207284 39764 207312
rect 35860 207272 35866 207284
rect 39758 207272 39764 207284
rect 39816 207272 39822 207324
rect 35526 207000 35532 207052
rect 35584 207040 35590 207052
rect 40310 207040 40316 207052
rect 35584 207012 40316 207040
rect 35584 207000 35590 207012
rect 40310 207000 40316 207012
rect 40368 207000 40374 207052
rect 580626 206932 580632 206984
rect 580684 206972 580690 206984
rect 589550 206972 589556 206984
rect 580684 206944 589556 206972
rect 580684 206932 580690 206944
rect 589550 206932 589556 206944
rect 589608 206932 589614 206984
rect 671706 206728 671712 206780
rect 671764 206728 671770 206780
rect 671724 206644 671752 206728
rect 671706 206592 671712 206644
rect 671764 206592 671770 206644
rect 35802 205912 35808 205964
rect 35860 205952 35866 205964
rect 39390 205952 39396 205964
rect 35860 205924 39396 205952
rect 35860 205912 35866 205924
rect 39390 205912 39396 205924
rect 39448 205912 39454 205964
rect 579522 205776 579528 205828
rect 579580 205816 579586 205828
rect 580994 205816 581000 205828
rect 579580 205788 581000 205816
rect 579580 205776 579586 205788
rect 580994 205776 581000 205788
rect 581052 205776 581058 205828
rect 35618 205640 35624 205692
rect 35676 205680 35682 205692
rect 41138 205680 41144 205692
rect 35676 205652 41144 205680
rect 35676 205640 35682 205652
rect 41138 205640 41144 205652
rect 41196 205640 41202 205692
rect 582282 205504 582288 205556
rect 582340 205544 582346 205556
rect 589458 205544 589464 205556
rect 582340 205516 589464 205544
rect 582340 205504 582346 205516
rect 589458 205504 589464 205516
rect 589516 205504 589522 205556
rect 35802 204824 35808 204876
rect 35860 204864 35866 204876
rect 39942 204864 39948 204876
rect 35860 204836 39948 204864
rect 35860 204824 35866 204836
rect 39942 204824 39948 204836
rect 40000 204824 40006 204876
rect 35618 204620 35624 204672
rect 35676 204660 35682 204672
rect 35676 204632 35894 204660
rect 35676 204620 35682 204632
rect 35866 204592 35894 204632
rect 41690 204592 41696 204604
rect 35866 204564 41696 204592
rect 41690 204552 41696 204564
rect 41748 204552 41754 204604
rect 42058 204552 42064 204604
rect 42116 204592 42122 204604
rect 44358 204592 44364 204604
rect 42116 204564 44364 204592
rect 42116 204552 42122 204564
rect 44358 204552 44364 204564
rect 44416 204552 44422 204604
rect 35526 204416 35532 204468
rect 35584 204456 35590 204468
rect 41690 204456 41696 204468
rect 35584 204428 41696 204456
rect 35584 204416 35590 204428
rect 41690 204416 41696 204428
rect 41748 204416 41754 204468
rect 42058 204416 42064 204468
rect 42116 204456 42122 204468
rect 47578 204456 47584 204468
rect 42116 204428 47584 204456
rect 42116 204416 42122 204428
rect 47578 204416 47584 204428
rect 47636 204416 47642 204468
rect 35802 204280 35808 204332
rect 35860 204320 35866 204332
rect 41690 204320 41696 204332
rect 35860 204292 41696 204320
rect 35860 204280 35866 204292
rect 41690 204280 41696 204292
rect 41748 204280 41754 204332
rect 42058 204280 42064 204332
rect 42116 204320 42122 204332
rect 48958 204320 48964 204332
rect 42116 204292 48964 204320
rect 42116 204280 42122 204292
rect 48958 204280 48964 204292
rect 49016 204280 49022 204332
rect 579706 204212 579712 204264
rect 579764 204252 579770 204264
rect 589458 204252 589464 204264
rect 579764 204224 589464 204252
rect 579764 204212 579770 204224
rect 589458 204212 589464 204224
rect 589516 204212 589522 204264
rect 41230 203232 41236 203244
rect 38626 203204 41236 203232
rect 35618 203124 35624 203176
rect 35676 203164 35682 203176
rect 38626 203164 38654 203204
rect 41230 203192 41236 203204
rect 41288 203192 41294 203244
rect 35676 203136 38654 203164
rect 35676 203124 35682 203136
rect 42058 202988 42064 203040
rect 42116 203028 42122 203040
rect 50338 203028 50344 203040
rect 42116 203000 50344 203028
rect 42116 202988 42122 203000
rect 50338 202988 50344 203000
rect 50396 202988 50402 203040
rect 35802 202852 35808 202904
rect 35860 202892 35866 202904
rect 41690 202892 41696 202904
rect 35860 202864 41696 202892
rect 35860 202852 35866 202864
rect 41690 202852 41696 202864
rect 41748 202852 41754 202904
rect 578326 202852 578332 202904
rect 578384 202892 578390 202904
rect 580258 202892 580264 202904
rect 578384 202864 580264 202892
rect 578384 202852 578390 202864
rect 580258 202852 580264 202864
rect 580316 202852 580322 202904
rect 580994 202784 581000 202836
rect 581052 202824 581058 202836
rect 589458 202824 589464 202836
rect 581052 202796 589464 202824
rect 581052 202784 581058 202796
rect 589458 202784 589464 202796
rect 589516 202784 589522 202836
rect 673362 201832 673368 201884
rect 673420 201872 673426 201884
rect 675386 201872 675392 201884
rect 673420 201844 675392 201872
rect 673420 201832 673426 201844
rect 675386 201832 675392 201844
rect 675444 201832 675450 201884
rect 671982 201288 671988 201340
rect 672040 201328 672046 201340
rect 675202 201328 675208 201340
rect 672040 201300 675208 201328
rect 672040 201288 672046 201300
rect 675202 201288 675208 201300
rect 675260 201288 675266 201340
rect 674834 200880 674840 200932
rect 674892 200920 674898 200932
rect 675294 200920 675300 200932
rect 674892 200892 675300 200920
rect 674892 200880 674898 200892
rect 675294 200880 675300 200892
rect 675352 200880 675358 200932
rect 673086 200472 673092 200524
rect 673144 200512 673150 200524
rect 675018 200512 675024 200524
rect 673144 200484 675024 200512
rect 673144 200472 673150 200484
rect 675018 200472 675024 200484
rect 675076 200472 675082 200524
rect 579154 200132 579160 200184
rect 579212 200172 579218 200184
rect 590562 200172 590568 200184
rect 579212 200144 590568 200172
rect 579212 200132 579218 200144
rect 590562 200132 590568 200144
rect 590620 200132 590626 200184
rect 580258 199996 580264 200048
rect 580316 200036 580322 200048
rect 589458 200036 589464 200048
rect 580316 200008 589464 200036
rect 580316 199996 580322 200008
rect 589458 199996 589464 200008
rect 589516 199996 589522 200048
rect 578878 197344 578884 197396
rect 578936 197384 578942 197396
rect 589458 197384 589464 197396
rect 578936 197356 589464 197384
rect 578936 197344 578942 197356
rect 589458 197344 589464 197356
rect 589516 197344 589522 197396
rect 666922 196664 666928 196716
rect 666980 196704 666986 196716
rect 667842 196704 667848 196716
rect 666980 196676 667848 196704
rect 666980 196664 666986 196676
rect 667842 196664 667848 196676
rect 667900 196664 667906 196716
rect 667658 196528 667664 196580
rect 667716 196568 667722 196580
rect 667716 196540 667888 196568
rect 667716 196528 667722 196540
rect 667860 196376 667888 196540
rect 667842 196324 667848 196376
rect 667900 196324 667906 196376
rect 579522 195984 579528 196036
rect 579580 196024 579586 196036
rect 589550 196024 589556 196036
rect 579580 195996 589556 196024
rect 579580 195984 579586 195996
rect 589550 195984 589556 195996
rect 589608 195984 589614 196036
rect 42426 195644 42432 195696
rect 42484 195684 42490 195696
rect 43806 195684 43812 195696
rect 42484 195656 43812 195684
rect 42484 195644 42490 195656
rect 43806 195644 43812 195656
rect 43864 195644 43870 195696
rect 674466 194488 674472 194540
rect 674524 194528 674530 194540
rect 675110 194528 675116 194540
rect 674524 194500 675116 194528
rect 674524 194488 674530 194500
rect 675110 194488 675116 194500
rect 675168 194488 675174 194540
rect 579522 193808 579528 193860
rect 579580 193848 579586 193860
rect 589550 193848 589556 193860
rect 579580 193820 589556 193848
rect 579580 193808 579586 193820
rect 589550 193808 589556 193820
rect 589608 193808 589614 193860
rect 42426 193128 42432 193180
rect 42484 193168 42490 193180
rect 43622 193168 43628 193180
rect 42484 193140 43628 193168
rect 42484 193128 42490 193140
rect 43622 193128 43628 193140
rect 43680 193128 43686 193180
rect 666922 192244 666928 192296
rect 666980 192284 666986 192296
rect 669314 192284 669320 192296
rect 666980 192256 669320 192284
rect 666980 192244 666986 192256
rect 669314 192244 669320 192256
rect 669372 192244 669378 192296
rect 42426 191768 42432 191820
rect 42484 191808 42490 191820
rect 44542 191808 44548 191820
rect 42484 191780 44548 191808
rect 42484 191768 42490 191780
rect 44542 191768 44548 191780
rect 44600 191768 44606 191820
rect 42426 191632 42432 191684
rect 42484 191672 42490 191684
rect 44358 191672 44364 191684
rect 42484 191644 44364 191672
rect 42484 191632 42490 191644
rect 44358 191632 44364 191644
rect 44416 191632 44422 191684
rect 579522 191088 579528 191140
rect 579580 191128 579586 191140
rect 589458 191128 589464 191140
rect 579580 191100 589464 191128
rect 579580 191088 579586 191100
rect 589458 191088 589464 191100
rect 589516 191088 589522 191140
rect 42426 190340 42432 190392
rect 42484 190380 42490 190392
rect 42978 190380 42984 190392
rect 42484 190352 42984 190380
rect 42484 190340 42490 190352
rect 42978 190340 42984 190352
rect 43036 190340 43042 190392
rect 675846 189728 675852 189780
rect 675904 189768 675910 189780
rect 683114 189768 683120 189780
rect 675904 189740 683120 189768
rect 675904 189728 675910 189740
rect 683114 189728 683120 189740
rect 683172 189728 683178 189780
rect 579522 188980 579528 189032
rect 579580 189020 579586 189032
rect 589458 189020 589464 189032
rect 579580 188992 589464 189020
rect 579580 188980 579586 188992
rect 589458 188980 589464 188992
rect 589516 188980 589522 189032
rect 42426 187620 42432 187672
rect 42484 187660 42490 187672
rect 43438 187660 43444 187672
rect 42484 187632 43444 187660
rect 42484 187620 42490 187632
rect 43438 187620 43444 187632
rect 43496 187620 43502 187672
rect 579522 186940 579528 186992
rect 579580 186980 579586 186992
rect 589458 186980 589464 186992
rect 579580 186952 589464 186980
rect 579580 186940 579586 186952
rect 589458 186940 589464 186952
rect 589516 186940 589522 186992
rect 579430 184900 579436 184952
rect 579488 184940 579494 184952
rect 589458 184940 589464 184952
rect 579488 184912 589464 184940
rect 579488 184900 579494 184912
rect 589458 184900 589464 184912
rect 589516 184900 589522 184952
rect 578510 184764 578516 184816
rect 578568 184804 578574 184816
rect 589642 184804 589648 184816
rect 578568 184776 589648 184804
rect 578568 184764 578574 184776
rect 589642 184764 589648 184776
rect 589700 184764 589706 184816
rect 42426 183472 42432 183524
rect 42484 183512 42490 183524
rect 44174 183512 44180 183524
rect 42484 183484 44180 183512
rect 42484 183472 42490 183484
rect 44174 183472 44180 183484
rect 44232 183472 44238 183524
rect 668210 183472 668216 183524
rect 668268 183512 668274 183524
rect 670970 183512 670976 183524
rect 668268 183484 670976 183512
rect 668268 183472 668274 183484
rect 670970 183472 670976 183484
rect 671028 183472 671034 183524
rect 669222 182860 669228 182912
rect 669280 182900 669286 182912
rect 672350 182900 672356 182912
rect 669280 182872 672356 182900
rect 669280 182860 669286 182872
rect 672350 182860 672356 182872
rect 672408 182860 672414 182912
rect 580902 182180 580908 182232
rect 580960 182220 580966 182232
rect 589458 182220 589464 182232
rect 580960 182192 589464 182220
rect 580960 182180 580966 182192
rect 589458 182180 589464 182192
rect 589516 182180 589522 182232
rect 583110 180820 583116 180872
rect 583168 180860 583174 180872
rect 589458 180860 589464 180872
rect 583168 180832 589464 180860
rect 583168 180820 583174 180832
rect 589458 180820 589464 180832
rect 589516 180820 589522 180872
rect 581730 179392 581736 179444
rect 581788 179432 581794 179444
rect 589458 179432 589464 179444
rect 581788 179404 589464 179432
rect 581788 179392 581794 179404
rect 589458 179392 589464 179404
rect 589516 179392 589522 179444
rect 578326 179324 578332 179376
rect 578384 179364 578390 179376
rect 580902 179364 580908 179376
rect 578384 179336 580908 179364
rect 578384 179324 578390 179336
rect 580902 179324 580908 179336
rect 580960 179324 580966 179376
rect 672534 178236 672540 178288
rect 672592 178276 672598 178288
rect 675478 178276 675484 178288
rect 672592 178248 675484 178276
rect 672592 178236 672598 178248
rect 675478 178236 675484 178248
rect 675536 178236 675542 178288
rect 579706 178032 579712 178084
rect 579764 178072 579770 178084
rect 589458 178072 589464 178084
rect 579764 178044 589464 178072
rect 579764 178032 579770 178044
rect 589458 178032 589464 178044
rect 589516 178032 589522 178084
rect 667106 178032 667112 178084
rect 667164 178072 667170 178084
rect 675294 178072 675300 178084
rect 667164 178044 675300 178072
rect 667164 178032 667170 178044
rect 675294 178032 675300 178044
rect 675352 178032 675358 178084
rect 667934 177896 667940 177948
rect 667992 177936 667998 177948
rect 673178 177936 673184 177948
rect 667992 177908 673184 177936
rect 667992 177896 667998 177908
rect 673178 177896 673184 177908
rect 673236 177896 673242 177948
rect 667750 176808 667756 176860
rect 667808 176848 667814 176860
rect 675294 176848 675300 176860
rect 667808 176820 675300 176848
rect 667808 176808 667814 176820
rect 675294 176808 675300 176820
rect 675352 176808 675358 176860
rect 673270 176672 673276 176724
rect 673328 176712 673334 176724
rect 675478 176712 675484 176724
rect 673328 176684 675484 176712
rect 673328 176672 673334 176684
rect 675478 176672 675484 176684
rect 675536 176672 675542 176724
rect 579522 176604 579528 176656
rect 579580 176644 579586 176656
rect 583110 176644 583116 176656
rect 579580 176616 583116 176644
rect 579580 176604 579586 176616
rect 583110 176604 583116 176616
rect 583168 176604 583174 176656
rect 587158 175312 587164 175364
rect 587216 175352 587222 175364
rect 589274 175352 589280 175364
rect 587216 175324 589280 175352
rect 587216 175312 587222 175324
rect 589274 175312 589280 175324
rect 589332 175312 589338 175364
rect 673086 175176 673092 175228
rect 673144 175216 673150 175228
rect 675478 175216 675484 175228
rect 673144 175188 675484 175216
rect 673144 175176 673150 175188
rect 675478 175176 675484 175188
rect 675536 175176 675542 175228
rect 578694 174836 578700 174888
rect 578752 174876 578758 174888
rect 581730 174876 581736 174888
rect 578752 174848 581736 174876
rect 578752 174836 578758 174848
rect 581730 174836 581736 174848
rect 581788 174836 581794 174888
rect 667934 174700 667940 174752
rect 667992 174740 667998 174752
rect 669958 174740 669964 174752
rect 667992 174712 669964 174740
rect 667992 174700 667998 174712
rect 669958 174700 669964 174712
rect 670016 174700 670022 174752
rect 581730 173136 581736 173188
rect 581788 173176 581794 173188
rect 589458 173176 589464 173188
rect 581788 173148 589464 173176
rect 581788 173136 581794 173148
rect 589458 173136 589464 173148
rect 589516 173136 589522 173188
rect 669406 171912 669412 171964
rect 669464 171952 669470 171964
rect 675478 171952 675484 171964
rect 669464 171924 675484 171952
rect 669464 171912 669470 171924
rect 675478 171912 675484 171924
rect 675536 171912 675542 171964
rect 673362 171164 673368 171216
rect 673420 171204 673426 171216
rect 675478 171204 675484 171216
rect 673420 171176 675484 171204
rect 673420 171164 673426 171176
rect 675478 171164 675484 171176
rect 675536 171164 675542 171216
rect 579798 171096 579804 171148
rect 579856 171136 579862 171148
rect 589458 171136 589464 171148
rect 579856 171108 589464 171136
rect 579856 171096 579862 171108
rect 589458 171096 589464 171108
rect 589516 171096 589522 171148
rect 578878 170348 578884 170400
rect 578936 170388 578942 170400
rect 587158 170388 587164 170400
rect 578936 170360 587164 170388
rect 578936 170348 578942 170360
rect 587158 170348 587164 170360
rect 587216 170348 587222 170400
rect 670602 170280 670608 170332
rect 670660 170320 670666 170332
rect 675478 170320 675484 170332
rect 670660 170292 675484 170320
rect 670660 170280 670666 170292
rect 675478 170280 675484 170292
rect 675536 170280 675542 170332
rect 667934 169668 667940 169720
rect 667992 169708 667998 169720
rect 670142 169708 670148 169720
rect 667992 169680 670148 169708
rect 667992 169668 667998 169680
rect 670142 169668 670148 169680
rect 670200 169668 670206 169720
rect 579246 169532 579252 169584
rect 579304 169572 579310 169584
rect 581730 169572 581736 169584
rect 579304 169544 581736 169572
rect 579304 169532 579310 169544
rect 581730 169532 581736 169544
rect 581788 169532 581794 169584
rect 672350 169056 672356 169108
rect 672408 169096 672414 169108
rect 675478 169096 675484 169108
rect 672408 169068 675484 169096
rect 672408 169056 672414 169068
rect 675478 169056 675484 169068
rect 675536 169056 675542 169108
rect 671982 168648 671988 168700
rect 672040 168688 672046 168700
rect 675478 168688 675484 168700
rect 672040 168660 675484 168688
rect 672040 168648 672046 168660
rect 675478 168648 675484 168660
rect 675536 168648 675542 168700
rect 583018 168376 583024 168428
rect 583076 168416 583082 168428
rect 589458 168416 589464 168428
rect 583076 168388 589464 168416
rect 583076 168376 583082 168388
rect 589458 168376 589464 168388
rect 589516 168376 589522 168428
rect 672534 168240 672540 168292
rect 672592 168280 672598 168292
rect 675478 168280 675484 168292
rect 672592 168252 675484 168280
rect 672592 168240 672598 168252
rect 675478 168240 675484 168252
rect 675536 168240 675542 168292
rect 669958 167832 669964 167884
rect 670016 167872 670022 167884
rect 675478 167872 675484 167884
rect 670016 167844 675484 167872
rect 670016 167832 670022 167844
rect 675478 167832 675484 167844
rect 675536 167832 675542 167884
rect 581638 167016 581644 167068
rect 581696 167056 581702 167068
rect 589458 167056 589464 167068
rect 581696 167028 589464 167056
rect 581696 167016 581702 167028
rect 589458 167016 589464 167028
rect 589516 167016 589522 167068
rect 670970 166880 670976 166932
rect 671028 166920 671034 166932
rect 675386 166920 675392 166932
rect 671028 166892 675392 166920
rect 671028 166880 671034 166892
rect 675386 166880 675392 166892
rect 675444 166880 675450 166932
rect 579522 166268 579528 166320
rect 579580 166308 579586 166320
rect 589734 166308 589740 166320
rect 579580 166280 589740 166308
rect 579580 166268 579586 166280
rect 589734 166268 589740 166280
rect 589792 166268 589798 166320
rect 668026 164908 668032 164960
rect 668084 164948 668090 164960
rect 670326 164948 670332 164960
rect 668084 164920 670332 164948
rect 668084 164908 668090 164920
rect 670326 164908 670332 164920
rect 670384 164908 670390 164960
rect 580258 164228 580264 164280
rect 580316 164268 580322 164280
rect 589458 164268 589464 164280
rect 580316 164240 589464 164268
rect 580316 164228 580322 164240
rect 589458 164228 589464 164240
rect 589516 164228 589522 164280
rect 587342 162868 587348 162920
rect 587400 162908 587406 162920
rect 589734 162908 589740 162920
rect 587400 162880 589740 162908
rect 587400 162868 587406 162880
rect 589734 162868 589740 162880
rect 589792 162868 589798 162920
rect 675846 162664 675852 162716
rect 675904 162704 675910 162716
rect 678238 162704 678244 162716
rect 675904 162676 678244 162704
rect 675904 162664 675910 162676
rect 678238 162664 678244 162676
rect 678296 162664 678302 162716
rect 585962 160080 585968 160132
rect 586020 160120 586026 160132
rect 589458 160120 589464 160132
rect 586020 160092 589464 160120
rect 586020 160080 586026 160092
rect 589458 160080 589464 160092
rect 589516 160080 589522 160132
rect 579522 159944 579528 159996
rect 579580 159984 579586 159996
rect 588538 159984 588544 159996
rect 579580 159956 588544 159984
rect 579580 159944 579586 159956
rect 588538 159944 588544 159956
rect 588596 159944 588602 159996
rect 668578 158312 668584 158364
rect 668636 158352 668642 158364
rect 674098 158352 674104 158364
rect 668636 158324 674104 158352
rect 668636 158312 668642 158324
rect 674098 158312 674104 158324
rect 674156 158312 674162 158364
rect 584398 157360 584404 157412
rect 584456 157400 584462 157412
rect 589458 157400 589464 157412
rect 584456 157372 589464 157400
rect 584456 157360 584462 157372
rect 589458 157360 589464 157372
rect 589516 157360 589522 157412
rect 579246 157292 579252 157344
rect 579304 157332 579310 157344
rect 583018 157332 583024 157344
rect 579304 157304 583024 157332
rect 579304 157292 579310 157304
rect 583018 157292 583024 157304
rect 583076 157292 583082 157344
rect 673362 156952 673368 157004
rect 673420 156992 673426 157004
rect 675110 156992 675116 157004
rect 673420 156964 675116 156992
rect 673420 156952 673426 156964
rect 675110 156952 675116 156964
rect 675168 156952 675174 157004
rect 578694 155456 578700 155508
rect 578752 155496 578758 155508
rect 581638 155496 581644 155508
rect 578752 155468 581644 155496
rect 578752 155456 578758 155468
rect 581638 155456 581644 155468
rect 581696 155456 581702 155508
rect 583202 154572 583208 154624
rect 583260 154612 583266 154624
rect 589366 154612 589372 154624
rect 583260 154584 589372 154612
rect 583260 154572 583266 154584
rect 589366 154572 589372 154584
rect 589424 154572 589430 154624
rect 578326 153416 578332 153468
rect 578384 153456 578390 153468
rect 580258 153456 580264 153468
rect 578384 153428 580264 153456
rect 578384 153416 578390 153428
rect 580258 153416 580264 153428
rect 580316 153416 580322 153468
rect 581822 153212 581828 153264
rect 581880 153252 581886 153264
rect 589458 153252 589464 153264
rect 581880 153224 589464 153252
rect 581880 153212 581886 153224
rect 589458 153212 589464 153224
rect 589516 153212 589522 153264
rect 672350 153144 672356 153196
rect 672408 153184 672414 153196
rect 675110 153184 675116 153196
rect 672408 153156 675116 153184
rect 672408 153144 672414 153156
rect 675110 153144 675116 153156
rect 675168 153144 675174 153196
rect 578418 152464 578424 152516
rect 578476 152504 578482 152516
rect 590102 152504 590108 152516
rect 578476 152476 590108 152504
rect 578476 152464 578482 152476
rect 590102 152464 590108 152476
rect 590160 152464 590166 152516
rect 671982 151716 671988 151768
rect 672040 151756 672046 151768
rect 675110 151756 675116 151768
rect 672040 151728 675116 151756
rect 672040 151716 672046 151728
rect 675110 151716 675116 151728
rect 675168 151716 675174 151768
rect 580626 151036 580632 151088
rect 580684 151076 580690 151088
rect 589734 151076 589740 151088
rect 580684 151048 589740 151076
rect 580684 151036 580690 151048
rect 589734 151036 589740 151048
rect 589792 151036 589798 151088
rect 579522 150356 579528 150408
rect 579580 150396 579586 150408
rect 587342 150396 587348 150408
rect 579580 150368 587348 150396
rect 579580 150356 579586 150368
rect 587342 150356 587348 150368
rect 587400 150356 587406 150408
rect 668762 150220 668768 150272
rect 668820 150260 668826 150272
rect 671246 150260 671252 150272
rect 668820 150232 671252 150260
rect 668820 150220 668826 150232
rect 671246 150220 671252 150232
rect 671304 150220 671310 150272
rect 587158 149064 587164 149116
rect 587216 149104 587222 149116
rect 589274 149104 589280 149116
rect 587216 149076 589280 149104
rect 587216 149064 587222 149076
rect 589274 149064 589280 149076
rect 589332 149064 589338 149116
rect 669406 148996 669412 149048
rect 669464 149036 669470 149048
rect 675294 149036 675300 149048
rect 669464 149008 675300 149036
rect 669464 148996 669470 149008
rect 675294 148996 675300 149008
rect 675352 148996 675358 149048
rect 670602 147568 670608 147620
rect 670660 147608 670666 147620
rect 675110 147608 675116 147620
rect 670660 147580 675116 147608
rect 670660 147568 670666 147580
rect 675110 147568 675116 147580
rect 675168 147568 675174 147620
rect 586882 146276 586888 146328
rect 586940 146316 586946 146328
rect 589458 146316 589464 146328
rect 586940 146288 589464 146316
rect 586940 146276 586946 146288
rect 589458 146276 589464 146288
rect 589516 146276 589522 146328
rect 668762 145528 668768 145580
rect 668820 145568 668826 145580
rect 671430 145568 671436 145580
rect 668820 145540 671436 145568
rect 668820 145528 668826 145540
rect 671430 145528 671436 145540
rect 671488 145528 671494 145580
rect 578786 145392 578792 145444
rect 578844 145432 578850 145444
rect 585962 145432 585968 145444
rect 578844 145404 585968 145432
rect 578844 145392 578850 145404
rect 585962 145392 585968 145404
rect 586020 145392 586026 145444
rect 585778 144916 585784 144968
rect 585836 144956 585842 144968
rect 589458 144956 589464 144968
rect 585836 144928 589464 144956
rect 585836 144916 585842 144928
rect 589458 144916 589464 144928
rect 589516 144916 589522 144968
rect 578878 144168 578884 144220
rect 578936 144208 578942 144220
rect 586882 144208 586888 144220
rect 578936 144180 586888 144208
rect 578936 144168 578942 144180
rect 586882 144168 586888 144180
rect 586940 144168 586946 144220
rect 579246 143420 579252 143472
rect 579304 143460 579310 143472
rect 588722 143460 588728 143472
rect 579304 143432 588728 143460
rect 579304 143420 579310 143432
rect 588722 143420 588728 143432
rect 588780 143420 588786 143472
rect 583754 140768 583760 140820
rect 583812 140808 583818 140820
rect 589458 140808 589464 140820
rect 583812 140780 589464 140808
rect 583812 140768 583818 140780
rect 589458 140768 589464 140780
rect 589516 140768 589522 140820
rect 579522 140564 579528 140616
rect 579580 140604 579586 140616
rect 584398 140604 584404 140616
rect 579580 140576 584404 140604
rect 579580 140564 579586 140576
rect 584398 140564 584404 140576
rect 584456 140564 584462 140616
rect 668670 140428 668676 140480
rect 668728 140468 668734 140480
rect 671614 140468 671620 140480
rect 668728 140440 671620 140468
rect 668728 140428 668734 140440
rect 671614 140428 671620 140440
rect 671672 140428 671678 140480
rect 580258 140020 580264 140072
rect 580316 140060 580322 140072
rect 590286 140060 590292 140072
rect 580316 140032 590292 140060
rect 580316 140020 580322 140032
rect 590286 140020 590292 140032
rect 590344 140020 590350 140072
rect 579062 138660 579068 138712
rect 579120 138700 579126 138712
rect 589918 138700 589924 138712
rect 579120 138672 589924 138700
rect 579120 138660 579126 138672
rect 589918 138660 589924 138672
rect 589976 138660 589982 138712
rect 668762 138388 668768 138440
rect 668820 138428 668826 138440
rect 674282 138428 674288 138440
rect 668820 138400 674288 138428
rect 668820 138388 668826 138400
rect 674282 138388 674288 138400
rect 674340 138388 674346 138440
rect 578326 137844 578332 137896
rect 578384 137884 578390 137896
rect 583202 137884 583208 137896
rect 578384 137856 583208 137884
rect 578384 137844 578390 137856
rect 583202 137844 583208 137856
rect 583260 137844 583266 137896
rect 583018 137232 583024 137284
rect 583076 137272 583082 137284
rect 589458 137272 589464 137284
rect 583076 137244 589464 137272
rect 583076 137232 583082 137244
rect 589458 137232 589464 137244
rect 589516 137232 589522 137284
rect 668762 136484 668768 136536
rect 668820 136524 668826 136536
rect 671798 136524 671804 136536
rect 668820 136496 671804 136524
rect 668820 136484 668826 136496
rect 671798 136484 671804 136496
rect 671856 136484 671862 136536
rect 581638 135260 581644 135312
rect 581696 135300 581702 135312
rect 589458 135300 589464 135312
rect 581696 135272 589464 135300
rect 581696 135260 581702 135272
rect 589458 135260 589464 135272
rect 589516 135260 589522 135312
rect 579338 135124 579344 135176
rect 579396 135164 579402 135176
rect 581822 135164 581828 135176
rect 579396 135136 581828 135164
rect 579396 135124 579402 135136
rect 581822 135124 581828 135136
rect 581880 135124 581886 135176
rect 580442 133900 580448 133952
rect 580500 133940 580506 133952
rect 589458 133940 589464 133952
rect 580500 133912 589464 133940
rect 580500 133900 580506 133912
rect 589458 133900 589464 133912
rect 589516 133900 589522 133952
rect 578326 133764 578332 133816
rect 578384 133804 578390 133816
rect 580626 133804 580632 133816
rect 578384 133776 580632 133804
rect 578384 133764 578390 133776
rect 580626 133764 580632 133776
rect 580684 133764 580690 133816
rect 579246 133424 579252 133476
rect 579304 133464 579310 133476
rect 583754 133464 583760 133476
rect 579304 133436 583760 133464
rect 579304 133424 579310 133436
rect 583754 133424 583760 133436
rect 583812 133424 583818 133476
rect 673914 132948 673920 133000
rect 673972 132988 673978 133000
rect 675478 132988 675484 133000
rect 673972 132960 675484 132988
rect 673972 132948 673978 132960
rect 675478 132948 675484 132960
rect 675536 132948 675542 133000
rect 667474 132744 667480 132796
rect 667532 132784 667538 132796
rect 675478 132784 675484 132796
rect 667532 132756 675484 132784
rect 667532 132744 667538 132756
rect 675478 132744 675484 132756
rect 675536 132744 675542 132796
rect 584766 132472 584772 132524
rect 584824 132512 584830 132524
rect 589458 132512 589464 132524
rect 584824 132484 589464 132512
rect 584824 132472 584830 132484
rect 589458 132472 589464 132484
rect 589516 132472 589522 132524
rect 667290 132472 667296 132524
rect 667348 132512 667354 132524
rect 675294 132512 675300 132524
rect 667348 132484 675300 132512
rect 667348 132472 667354 132484
rect 675294 132472 675300 132484
rect 675352 132472 675358 132524
rect 673362 131248 673368 131300
rect 673420 131288 673426 131300
rect 675294 131288 675300 131300
rect 673420 131260 675300 131288
rect 673420 131248 673426 131260
rect 675294 131248 675300 131260
rect 675352 131248 675358 131300
rect 668762 131112 668768 131164
rect 668820 131152 668826 131164
rect 675478 131152 675484 131164
rect 668820 131124 675484 131152
rect 668820 131112 668826 131124
rect 675478 131112 675484 131124
rect 675536 131112 675542 131164
rect 667934 130908 667940 130960
rect 667992 130948 667998 130960
rect 669774 130948 669780 130960
rect 667992 130920 669780 130948
rect 667992 130908 667998 130920
rect 669774 130908 669780 130920
rect 669832 130908 669838 130960
rect 674098 130840 674104 130892
rect 674156 130880 674162 130892
rect 675478 130880 675484 130892
rect 674156 130852 675484 130880
rect 674156 130840 674162 130852
rect 675478 130840 675484 130852
rect 675536 130840 675542 130892
rect 673086 130228 673092 130280
rect 673144 130268 673150 130280
rect 675478 130268 675484 130280
rect 673144 130240 675484 130268
rect 673144 130228 673150 130240
rect 675478 130228 675484 130240
rect 675536 130228 675542 130280
rect 669130 129888 669136 129940
rect 669188 129928 669194 129940
rect 675478 129928 675484 129940
rect 669188 129900 675484 129928
rect 669188 129888 669194 129900
rect 675478 129888 675484 129900
rect 675536 129888 675542 129940
rect 668578 129752 668584 129804
rect 668636 129792 668642 129804
rect 669130 129792 669136 129804
rect 668636 129764 669136 129792
rect 668636 129752 668642 129764
rect 669130 129752 669136 129764
rect 669188 129752 669194 129804
rect 669222 129004 669228 129056
rect 669280 129044 669286 129056
rect 672718 129044 672724 129056
rect 669280 129016 672724 129044
rect 669280 129004 669286 129016
rect 672718 129004 672724 129016
rect 672776 129004 672782 129056
rect 585962 128324 585968 128376
rect 586020 128364 586026 128376
rect 589458 128364 589464 128376
rect 586020 128336 589464 128364
rect 586020 128324 586026 128336
rect 589458 128324 589464 128336
rect 589516 128324 589522 128376
rect 668946 128324 668952 128376
rect 669004 128364 669010 128376
rect 675478 128364 675484 128376
rect 669004 128336 675484 128364
rect 669004 128324 669010 128336
rect 675478 128324 675484 128336
rect 675536 128324 675542 128376
rect 579522 128188 579528 128240
rect 579580 128228 579586 128240
rect 587158 128228 587164 128240
rect 579580 128200 587164 128228
rect 579580 128188 579586 128200
rect 587158 128188 587164 128200
rect 587216 128188 587222 128240
rect 667934 126148 667940 126200
rect 667992 126188 667998 126200
rect 669590 126188 669596 126200
rect 667992 126160 669596 126188
rect 667992 126148 667998 126160
rect 669590 126148 669596 126160
rect 669648 126148 669654 126200
rect 673178 125944 673184 125996
rect 673236 125984 673242 125996
rect 675478 125984 675484 125996
rect 673236 125956 675484 125984
rect 673236 125944 673242 125956
rect 675478 125944 675484 125956
rect 675536 125944 675542 125996
rect 587342 125604 587348 125656
rect 587400 125644 587406 125656
rect 589274 125644 589280 125656
rect 587400 125616 589280 125644
rect 587400 125604 587406 125616
rect 589274 125604 589280 125616
rect 589332 125604 589338 125656
rect 672718 125604 672724 125656
rect 672776 125644 672782 125656
rect 675478 125644 675484 125656
rect 672776 125616 675484 125644
rect 672776 125604 672782 125616
rect 675478 125604 675484 125616
rect 675536 125604 675542 125656
rect 578418 124856 578424 124908
rect 578476 124896 578482 124908
rect 588538 124896 588544 124908
rect 578476 124868 588544 124896
rect 578476 124856 578482 124868
rect 588538 124856 588544 124868
rect 588596 124856 588602 124908
rect 673914 124720 673920 124772
rect 673972 124760 673978 124772
rect 675478 124760 675484 124772
rect 673972 124732 675484 124760
rect 673972 124720 673978 124732
rect 675478 124720 675484 124732
rect 675536 124720 675542 124772
rect 669222 124108 669228 124160
rect 669280 124148 669286 124160
rect 672902 124148 672908 124160
rect 669280 124120 672908 124148
rect 669280 124108 669286 124120
rect 672902 124108 672908 124120
rect 672960 124108 672966 124160
rect 673362 122952 673368 123004
rect 673420 122992 673426 123004
rect 675294 122992 675300 123004
rect 673420 122964 675300 122992
rect 673420 122952 673426 122964
rect 675294 122952 675300 122964
rect 675352 122952 675358 123004
rect 671338 122816 671344 122868
rect 671396 122856 671402 122868
rect 675478 122856 675484 122868
rect 671396 122828 675484 122856
rect 671396 122816 671402 122828
rect 675478 122816 675484 122828
rect 675536 122816 675542 122868
rect 578878 122612 578884 122664
rect 578936 122652 578942 122664
rect 585778 122652 585784 122664
rect 578936 122624 585784 122652
rect 578936 122612 578942 122624
rect 585778 122612 585784 122624
rect 585836 122612 585842 122664
rect 581822 121456 581828 121508
rect 581880 121496 581886 121508
rect 589458 121496 589464 121508
rect 581880 121468 589464 121496
rect 581880 121456 581886 121468
rect 589458 121456 589464 121468
rect 589516 121456 589522 121508
rect 670142 121456 670148 121508
rect 670200 121496 670206 121508
rect 675294 121496 675300 121508
rect 670200 121468 675300 121496
rect 670200 121456 670206 121468
rect 675294 121456 675300 121468
rect 675352 121456 675358 121508
rect 586146 120708 586152 120760
rect 586204 120748 586210 120760
rect 589918 120748 589924 120760
rect 586204 120720 589924 120748
rect 586204 120708 586210 120720
rect 589918 120708 589924 120720
rect 589976 120708 589982 120760
rect 671522 120708 671528 120760
rect 671580 120748 671586 120760
rect 675478 120748 675484 120760
rect 671580 120720 675484 120748
rect 671580 120708 671586 120720
rect 675478 120708 675484 120720
rect 675536 120708 675542 120760
rect 669130 119212 669136 119264
rect 669188 119252 669194 119264
rect 672534 119252 672540 119264
rect 669188 119224 672540 119252
rect 669188 119212 669194 119224
rect 672534 119212 672540 119224
rect 672592 119212 672598 119264
rect 584582 118668 584588 118720
rect 584640 118708 584646 118720
rect 589458 118708 589464 118720
rect 584640 118680 589464 118708
rect 584640 118668 584646 118680
rect 589458 118668 589464 118680
rect 589516 118668 589522 118720
rect 578510 118260 578516 118312
rect 578568 118300 578574 118312
rect 580258 118300 580264 118312
rect 578568 118272 580264 118300
rect 578568 118260 578574 118272
rect 580258 118260 580264 118272
rect 580316 118260 580322 118312
rect 667934 117784 667940 117836
rect 667992 117824 667998 117836
rect 669958 117824 669964 117836
rect 667992 117796 669964 117824
rect 667992 117784 667998 117796
rect 669958 117784 669964 117796
rect 670016 117784 670022 117836
rect 579062 117308 579068 117360
rect 579120 117348 579126 117360
rect 589458 117348 589464 117360
rect 579120 117320 589464 117348
rect 579120 117308 579126 117320
rect 589458 117308 589464 117320
rect 589516 117308 589522 117360
rect 675846 117240 675852 117292
rect 675904 117280 675910 117292
rect 679618 117280 679624 117292
rect 675904 117252 679624 117280
rect 675904 117240 675910 117252
rect 679618 117240 679624 117252
rect 679676 117240 679682 117292
rect 578878 115948 578884 116000
rect 578936 115988 578942 116000
rect 589458 115988 589464 116000
rect 578936 115960 589464 115988
rect 578936 115948 578942 115960
rect 589458 115948 589464 115960
rect 589516 115948 589522 116000
rect 668394 115812 668400 115864
rect 668452 115852 668458 115864
rect 670970 115852 670976 115864
rect 668452 115824 670976 115852
rect 668452 115812 668458 115824
rect 670970 115812 670976 115824
rect 671028 115812 671034 115864
rect 580626 115200 580632 115252
rect 580684 115240 580690 115252
rect 590286 115240 590292 115252
rect 580684 115212 590292 115240
rect 580684 115200 580690 115212
rect 590286 115200 590292 115212
rect 590344 115200 590350 115252
rect 668394 114316 668400 114368
rect 668452 114356 668458 114368
rect 671338 114356 671344 114368
rect 668452 114328 671344 114356
rect 668452 114316 668458 114328
rect 671338 114316 671344 114328
rect 671396 114316 671402 114368
rect 585778 113160 585784 113212
rect 585836 113200 585842 113212
rect 589458 113200 589464 113212
rect 585836 113172 589464 113200
rect 585836 113160 585842 113172
rect 589458 113160 589464 113172
rect 589516 113160 589522 113212
rect 579522 113092 579528 113144
rect 579580 113132 579586 113144
rect 583018 113132 583024 113144
rect 579580 113104 583024 113132
rect 579580 113092 579586 113104
rect 583018 113092 583024 113104
rect 583076 113092 583082 113144
rect 668026 112888 668032 112940
rect 668084 112928 668090 112940
rect 670142 112928 670148 112940
rect 668084 112900 670148 112928
rect 668084 112888 668090 112900
rect 670142 112888 670148 112900
rect 670200 112888 670206 112940
rect 673178 111732 673184 111784
rect 673236 111772 673242 111784
rect 675110 111772 675116 111784
rect 673236 111744 675116 111772
rect 673236 111732 673242 111744
rect 675110 111732 675116 111744
rect 675168 111732 675174 111784
rect 668762 111596 668768 111648
rect 668820 111636 668826 111648
rect 671522 111636 671528 111648
rect 668820 111608 671528 111636
rect 668820 111596 668826 111608
rect 671522 111596 671528 111608
rect 671580 111596 671586 111648
rect 579522 111188 579528 111240
rect 579580 111228 579586 111240
rect 586146 111228 586152 111240
rect 579580 111200 586152 111228
rect 579580 111188 579586 111200
rect 586146 111188 586152 111200
rect 586204 111188 586210 111240
rect 672718 111120 672724 111172
rect 672776 111160 672782 111172
rect 675386 111160 675392 111172
rect 672776 111132 675392 111160
rect 672776 111120 672782 111132
rect 675386 111120 675392 111132
rect 675444 111120 675450 111172
rect 587158 110440 587164 110492
rect 587216 110480 587222 110492
rect 589642 110480 589648 110492
rect 587216 110452 589648 110480
rect 587216 110440 587222 110452
rect 589642 110440 589648 110452
rect 589700 110440 589706 110492
rect 584398 109012 584404 109064
rect 584456 109052 584462 109064
rect 589458 109052 589464 109064
rect 584456 109024 589464 109052
rect 584456 109012 584462 109024
rect 589458 109012 589464 109024
rect 589516 109012 589522 109064
rect 579246 108740 579252 108792
rect 579304 108780 579310 108792
rect 581638 108780 581644 108792
rect 579304 108752 581644 108780
rect 579304 108740 579310 108752
rect 581638 108740 581644 108752
rect 581696 108740 581702 108792
rect 583202 107652 583208 107704
rect 583260 107692 583266 107704
rect 589458 107692 589464 107704
rect 583260 107664 589464 107692
rect 583260 107652 583266 107664
rect 589458 107652 589464 107664
rect 589516 107652 589522 107704
rect 669222 107652 669228 107704
rect 669280 107692 669286 107704
rect 674098 107692 674104 107704
rect 669280 107664 674104 107692
rect 669280 107652 669286 107664
rect 674098 107652 674104 107664
rect 674156 107652 674162 107704
rect 579246 107176 579252 107228
rect 579304 107216 579310 107228
rect 584766 107216 584772 107228
rect 579304 107188 584772 107216
rect 579304 107176 579310 107188
rect 584766 107176 584772 107188
rect 584824 107176 584830 107228
rect 673914 106972 673920 107024
rect 673972 107012 673978 107024
rect 675294 107012 675300 107024
rect 673972 106984 675300 107012
rect 673972 106972 673978 106984
rect 675294 106972 675300 106984
rect 675352 106972 675358 107024
rect 578326 106768 578332 106820
rect 578384 106808 578390 106820
rect 580442 106808 580448 106820
rect 578384 106780 580448 106808
rect 578384 106768 578390 106780
rect 580442 106768 580448 106780
rect 580500 106768 580506 106820
rect 580258 106292 580264 106344
rect 580316 106332 580322 106344
rect 589458 106332 589464 106344
rect 580316 106304 589464 106332
rect 580316 106292 580322 106304
rect 589458 106292 589464 106304
rect 589516 106292 589522 106344
rect 583018 104864 583024 104916
rect 583076 104904 583082 104916
rect 589458 104904 589464 104916
rect 583076 104876 589464 104904
rect 583076 104864 583082 104876
rect 589458 104864 589464 104876
rect 589516 104864 589522 104916
rect 581638 103504 581644 103556
rect 581696 103544 581702 103556
rect 589458 103544 589464 103556
rect 581696 103516 589464 103544
rect 581696 103504 581702 103516
rect 589458 103504 589464 103516
rect 589516 103504 589522 103556
rect 579522 103368 579528 103420
rect 579580 103408 579586 103420
rect 591298 103408 591304 103420
rect 579580 103380 591304 103408
rect 579580 103368 579586 103380
rect 591298 103368 591304 103380
rect 591356 103368 591362 103420
rect 579522 99288 579528 99340
rect 579580 99328 579586 99340
rect 588906 99328 588912 99340
rect 579580 99300 588912 99328
rect 579580 99288 579586 99300
rect 588906 99288 588912 99300
rect 588964 99288 588970 99340
rect 625062 99152 625068 99204
rect 625120 99192 625126 99204
rect 634446 99192 634452 99204
rect 625120 99164 634452 99192
rect 625120 99152 625126 99164
rect 634446 99152 634452 99164
rect 634504 99152 634510 99204
rect 623682 99016 623688 99068
rect 623740 99056 623746 99068
rect 632146 99056 632152 99068
rect 623740 99028 632152 99056
rect 623740 99016 623746 99028
rect 632146 99016 632152 99028
rect 632204 99016 632210 99068
rect 629754 98880 629760 98932
rect 629812 98920 629818 98932
rect 640978 98920 640984 98932
rect 629812 98892 640984 98920
rect 629812 98880 629818 98892
rect 640978 98880 640984 98892
rect 641036 98880 641042 98932
rect 621658 98744 621664 98796
rect 621716 98784 621722 98796
rect 628374 98784 628380 98796
rect 621716 98756 628380 98784
rect 621716 98744 621722 98756
rect 628374 98744 628380 98756
rect 628432 98744 628438 98796
rect 629018 98744 629024 98796
rect 629076 98784 629082 98796
rect 640242 98784 640248 98796
rect 629076 98756 640248 98784
rect 629076 98744 629082 98756
rect 640242 98744 640248 98756
rect 640300 98744 640306 98796
rect 622302 98608 622308 98660
rect 622360 98648 622366 98660
rect 629478 98648 629484 98660
rect 622360 98620 629484 98648
rect 622360 98608 622366 98620
rect 629478 98608 629484 98620
rect 629536 98608 629542 98660
rect 630490 98608 630496 98660
rect 630548 98648 630554 98660
rect 642082 98648 642088 98660
rect 630548 98620 642088 98648
rect 630548 98608 630554 98620
rect 642082 98608 642088 98620
rect 642140 98608 642146 98660
rect 588538 97996 588544 98048
rect 588596 98036 588602 98048
rect 589366 98036 589372 98048
rect 588596 98008 589372 98036
rect 588596 97996 588602 98008
rect 589366 97996 589372 98008
rect 589424 97996 589430 98048
rect 577498 97928 577504 97980
rect 577556 97968 577562 97980
rect 577556 97940 586514 97968
rect 577556 97928 577562 97940
rect 586486 97696 586514 97940
rect 594058 97928 594064 97980
rect 594116 97968 594122 97980
rect 596174 97968 596180 97980
rect 594116 97940 596180 97968
rect 594116 97928 594122 97940
rect 596174 97928 596180 97940
rect 596232 97928 596238 97980
rect 620186 97928 620192 97980
rect 620244 97968 620250 97980
rect 626074 97968 626080 97980
rect 620244 97940 626080 97968
rect 620244 97928 620250 97940
rect 626074 97928 626080 97940
rect 626132 97928 626138 97980
rect 626810 97928 626816 97980
rect 626868 97968 626874 97980
rect 636378 97968 636384 97980
rect 626868 97940 636384 97968
rect 626868 97928 626874 97940
rect 636378 97928 636384 97940
rect 636436 97928 636442 97980
rect 659746 97968 659752 97980
rect 644446 97940 659752 97968
rect 592678 97792 592684 97844
rect 592736 97832 592742 97844
rect 597554 97832 597560 97844
rect 592736 97804 597560 97832
rect 592736 97792 592742 97804
rect 597554 97792 597560 97804
rect 597612 97792 597618 97844
rect 625890 97792 625896 97844
rect 625948 97832 625954 97844
rect 635274 97832 635280 97844
rect 625948 97804 635280 97832
rect 625948 97792 625954 97804
rect 635274 97792 635280 97804
rect 635332 97792 635338 97844
rect 643002 97792 643008 97844
rect 643060 97832 643066 97844
rect 644446 97832 644474 97940
rect 659746 97928 659752 97940
rect 659804 97928 659810 97980
rect 659930 97928 659936 97980
rect 659988 97968 659994 97980
rect 665726 97968 665732 97980
rect 659988 97940 665732 97968
rect 659988 97928 659994 97940
rect 665726 97928 665732 97940
rect 665784 97928 665790 97980
rect 643060 97804 644474 97832
rect 643060 97792 643066 97804
rect 647142 97792 647148 97844
rect 647200 97832 647206 97844
rect 661954 97832 661960 97844
rect 647200 97804 661960 97832
rect 647200 97792 647206 97804
rect 661954 97792 661960 97804
rect 662012 97792 662018 97844
rect 595254 97696 595260 97708
rect 586486 97668 595260 97696
rect 595254 97656 595260 97668
rect 595312 97696 595318 97708
rect 595622 97696 595628 97708
rect 595312 97668 595628 97696
rect 595312 97656 595318 97668
rect 595622 97656 595628 97668
rect 595680 97656 595686 97708
rect 623130 97656 623136 97708
rect 623188 97696 623194 97708
rect 630674 97696 630680 97708
rect 623188 97668 630680 97696
rect 623188 97656 623194 97668
rect 630674 97656 630680 97668
rect 630732 97656 630738 97708
rect 632698 97656 632704 97708
rect 632756 97696 632762 97708
rect 632756 97668 633204 97696
rect 632756 97656 632762 97668
rect 595438 97520 595444 97572
rect 595496 97560 595502 97572
rect 598934 97560 598940 97572
rect 595496 97532 598940 97560
rect 595496 97520 595502 97532
rect 598934 97520 598940 97532
rect 598992 97520 598998 97572
rect 624602 97520 624608 97572
rect 624660 97560 624666 97572
rect 632974 97560 632980 97572
rect 624660 97532 632980 97560
rect 624660 97520 624666 97532
rect 632974 97520 632980 97532
rect 633032 97520 633038 97572
rect 633176 97560 633204 97668
rect 633342 97656 633348 97708
rect 633400 97696 633406 97708
rect 643922 97696 643928 97708
rect 633400 97668 643928 97696
rect 633400 97656 633406 97668
rect 643922 97656 643928 97668
rect 643980 97656 643986 97708
rect 655422 97656 655428 97708
rect 655480 97696 655486 97708
rect 662506 97696 662512 97708
rect 655480 97668 662512 97696
rect 655480 97656 655486 97668
rect 662506 97656 662512 97668
rect 662564 97656 662570 97708
rect 644750 97560 644756 97572
rect 633176 97532 644756 97560
rect 644750 97520 644756 97532
rect 644808 97520 644814 97572
rect 658826 97560 658832 97572
rect 649966 97532 658832 97560
rect 627546 97384 627552 97436
rect 627604 97424 627610 97436
rect 637574 97424 637580 97436
rect 627604 97396 637580 97424
rect 627604 97384 627610 97396
rect 637574 97384 637580 97396
rect 637632 97384 637638 97436
rect 639322 97384 639328 97436
rect 639380 97424 639386 97436
rect 646498 97424 646504 97436
rect 639380 97396 646504 97424
rect 639380 97384 639386 97396
rect 646498 97384 646504 97396
rect 646556 97384 646562 97436
rect 649966 97424 649994 97532
rect 658826 97520 658832 97532
rect 658884 97520 658890 97572
rect 649276 97396 649994 97424
rect 591298 97248 591304 97300
rect 591356 97288 591362 97300
rect 600406 97288 600412 97300
rect 591356 97260 600412 97288
rect 591356 97248 591362 97260
rect 600406 97248 600412 97260
rect 600464 97248 600470 97300
rect 605466 97248 605472 97300
rect 605524 97288 605530 97300
rect 611906 97288 611912 97300
rect 605524 97260 611912 97288
rect 605524 97248 605530 97260
rect 611906 97248 611912 97260
rect 611964 97248 611970 97300
rect 628190 97248 628196 97300
rect 628248 97288 628254 97300
rect 639046 97288 639052 97300
rect 628248 97260 639052 97288
rect 628248 97248 628254 97260
rect 639046 97248 639052 97260
rect 639104 97248 639110 97300
rect 641530 97248 641536 97300
rect 641588 97288 641594 97300
rect 643002 97288 643008 97300
rect 641588 97260 643008 97288
rect 641588 97248 641594 97260
rect 643002 97248 643008 97260
rect 643060 97248 643066 97300
rect 644290 97248 644296 97300
rect 644348 97288 644354 97300
rect 649276 97288 649304 97396
rect 658182 97384 658188 97436
rect 658240 97424 658246 97436
rect 663058 97424 663064 97436
rect 658240 97396 663064 97424
rect 658240 97384 658246 97396
rect 663058 97384 663064 97396
rect 663116 97384 663122 97436
rect 644348 97260 649304 97288
rect 644348 97248 644354 97260
rect 656802 97248 656808 97300
rect 656860 97288 656866 97300
rect 661402 97288 661408 97300
rect 656860 97260 661408 97288
rect 656860 97248 656866 97260
rect 661402 97248 661408 97260
rect 661460 97248 661466 97300
rect 654778 97180 654784 97232
rect 654836 97220 654842 97232
rect 655238 97220 655244 97232
rect 654836 97192 655244 97220
rect 654836 97180 654842 97192
rect 655238 97180 655244 97192
rect 655296 97180 655302 97232
rect 634170 97112 634176 97164
rect 634228 97152 634234 97164
rect 643462 97152 643468 97164
rect 634228 97124 643468 97152
rect 634228 97112 634234 97124
rect 643462 97112 643468 97124
rect 643520 97112 643526 97164
rect 656710 97044 656716 97096
rect 656768 97084 656774 97096
rect 656768 97056 659654 97084
rect 656768 97044 656774 97056
rect 612642 96976 612648 97028
rect 612700 97016 612706 97028
rect 613378 97016 613384 97028
rect 612700 96988 613384 97016
rect 612700 96976 612706 96988
rect 613378 96976 613384 96988
rect 613436 96976 613442 97028
rect 601694 96908 601700 96960
rect 601752 96948 601758 96960
rect 602614 96948 602620 96960
rect 601752 96920 602620 96948
rect 601752 96908 601758 96920
rect 602614 96908 602620 96920
rect 602672 96908 602678 96960
rect 606202 96908 606208 96960
rect 606260 96948 606266 96960
rect 606938 96948 606944 96960
rect 606260 96920 606944 96948
rect 606260 96908 606266 96920
rect 606938 96908 606944 96920
rect 606996 96908 607002 96960
rect 614022 96908 614028 96960
rect 614080 96948 614086 96960
rect 614758 96948 614764 96960
rect 614080 96920 614764 96948
rect 614080 96908 614086 96920
rect 614758 96908 614764 96920
rect 614816 96908 614822 96960
rect 615770 96908 615776 96960
rect 615828 96948 615834 96960
rect 616782 96948 616788 96960
rect 615828 96920 616788 96948
rect 615828 96908 615834 96920
rect 616782 96908 616788 96920
rect 616840 96908 616846 96960
rect 617242 96908 617248 96960
rect 617300 96948 617306 96960
rect 617886 96948 617892 96960
rect 617300 96920 617892 96948
rect 617300 96908 617306 96920
rect 617886 96908 617892 96920
rect 617944 96908 617950 96960
rect 646682 96908 646688 96960
rect 646740 96948 646746 96960
rect 647142 96948 647148 96960
rect 646740 96920 647148 96948
rect 646740 96908 646746 96920
rect 647142 96908 647148 96920
rect 647200 96908 647206 96960
rect 650362 96908 650368 96960
rect 650420 96948 650426 96960
rect 658274 96948 658280 96960
rect 650420 96920 658280 96948
rect 650420 96908 650426 96920
rect 658274 96908 658280 96920
rect 658332 96908 658338 96960
rect 659626 96948 659654 97056
rect 660114 96948 660120 96960
rect 659626 96920 660120 96948
rect 660114 96908 660120 96920
rect 660172 96908 660178 96960
rect 609146 96840 609152 96892
rect 609204 96880 609210 96892
rect 609698 96880 609704 96892
rect 609204 96852 609704 96880
rect 609204 96840 609210 96852
rect 609698 96840 609704 96852
rect 609756 96840 609762 96892
rect 612090 96840 612096 96892
rect 612148 96880 612154 96892
rect 612642 96880 612648 96892
rect 612148 96852 612648 96880
rect 612148 96840 612154 96852
rect 612642 96840 612648 96852
rect 612700 96840 612706 96892
rect 618714 96840 618720 96892
rect 618772 96880 618778 96892
rect 626258 96880 626264 96892
rect 618772 96852 626264 96880
rect 618772 96840 618778 96852
rect 626258 96840 626264 96852
rect 626316 96840 626322 96892
rect 613562 96772 613568 96824
rect 613620 96812 613626 96824
rect 614022 96812 614028 96824
rect 613620 96784 614028 96812
rect 613620 96772 613626 96784
rect 614022 96772 614028 96784
rect 614080 96772 614086 96824
rect 651834 96772 651840 96824
rect 651892 96812 651898 96824
rect 659562 96812 659568 96824
rect 651892 96784 659568 96812
rect 651892 96772 651898 96784
rect 659562 96772 659568 96784
rect 659620 96772 659626 96824
rect 642818 96744 642824 96756
rect 642100 96716 642824 96744
rect 578602 96568 578608 96620
rect 578660 96608 578666 96620
rect 587342 96608 587348 96620
rect 578660 96580 587348 96608
rect 578660 96568 578666 96580
rect 587342 96568 587348 96580
rect 587400 96568 587406 96620
rect 635642 96568 635648 96620
rect 635700 96608 635706 96620
rect 642100 96608 642128 96716
rect 642818 96704 642824 96716
rect 642876 96704 642882 96756
rect 645210 96704 645216 96756
rect 645268 96744 645274 96756
rect 645762 96744 645768 96756
rect 645268 96716 645768 96744
rect 645268 96704 645274 96716
rect 645762 96704 645768 96716
rect 645820 96704 645826 96756
rect 651098 96636 651104 96688
rect 651156 96676 651162 96688
rect 654318 96676 654324 96688
rect 651156 96648 654324 96676
rect 651156 96636 651162 96648
rect 654318 96636 654324 96648
rect 654376 96636 654382 96688
rect 635700 96580 642128 96608
rect 635700 96568 635706 96580
rect 642266 96568 642272 96620
rect 642324 96608 642330 96620
rect 643278 96608 643284 96620
rect 642324 96580 643284 96608
rect 642324 96568 642330 96580
rect 643278 96568 643284 96580
rect 643336 96568 643342 96620
rect 650914 96608 650920 96620
rect 643434 96580 650920 96608
rect 638586 96432 638592 96484
rect 638644 96472 638650 96484
rect 643434 96472 643462 96580
rect 650914 96568 650920 96580
rect 650972 96568 650978 96620
rect 638644 96444 643462 96472
rect 638644 96432 638650 96444
rect 653306 96432 653312 96484
rect 653364 96472 653370 96484
rect 663978 96472 663984 96484
rect 653364 96444 663984 96472
rect 653364 96432 653370 96444
rect 663978 96432 663984 96444
rect 664036 96432 664042 96484
rect 631226 96296 631232 96348
rect 631284 96336 631290 96348
rect 642634 96336 642640 96348
rect 631284 96308 642640 96336
rect 631284 96296 631290 96308
rect 642634 96296 642640 96308
rect 642692 96296 642698 96348
rect 642818 96296 642824 96348
rect 642876 96336 642882 96348
rect 648798 96336 648804 96348
rect 642876 96308 648804 96336
rect 642876 96296 642882 96308
rect 648798 96296 648804 96308
rect 648856 96296 648862 96348
rect 652570 96296 652576 96348
rect 652628 96336 652634 96348
rect 665358 96336 665364 96348
rect 652628 96308 665364 96336
rect 652628 96296 652634 96308
rect 665358 96296 665364 96308
rect 665416 96296 665422 96348
rect 620922 96228 620928 96280
rect 620980 96268 620986 96280
rect 626442 96268 626448 96280
rect 620980 96240 626448 96268
rect 620980 96228 620986 96240
rect 626442 96228 626448 96240
rect 626500 96228 626506 96280
rect 631870 96160 631876 96212
rect 631928 96200 631934 96212
rect 644474 96200 644480 96212
rect 631928 96172 644480 96200
rect 631928 96160 631934 96172
rect 644474 96160 644480 96172
rect 644532 96160 644538 96212
rect 648614 96160 648620 96212
rect 648672 96200 648678 96212
rect 663794 96200 663800 96212
rect 648672 96172 663800 96200
rect 648672 96160 648678 96172
rect 663794 96160 663800 96172
rect 663852 96160 663858 96212
rect 586514 96024 586520 96076
rect 586572 96064 586578 96076
rect 590102 96064 590108 96076
rect 586572 96036 590108 96064
rect 586572 96024 586578 96036
rect 590102 96024 590108 96036
rect 590160 96024 590166 96076
rect 610618 96024 610624 96076
rect 610676 96064 610682 96076
rect 621658 96064 621664 96076
rect 610676 96036 621664 96064
rect 610676 96024 610682 96036
rect 621658 96024 621664 96036
rect 621716 96024 621722 96076
rect 637850 96024 637856 96076
rect 637908 96064 637914 96076
rect 660666 96064 660672 96076
rect 637908 96036 660672 96064
rect 637908 96024 637914 96036
rect 660666 96024 660672 96036
rect 660724 96024 660730 96076
rect 608410 95888 608416 95940
rect 608468 95928 608474 95940
rect 620278 95928 620284 95940
rect 608468 95900 620284 95928
rect 608468 95888 608474 95900
rect 620278 95888 620284 95900
rect 620336 95888 620342 95940
rect 640794 95888 640800 95940
rect 640852 95928 640858 95940
rect 665174 95928 665180 95940
rect 640852 95900 665180 95928
rect 640852 95888 640858 95900
rect 665174 95888 665180 95900
rect 665232 95888 665238 95940
rect 640058 95752 640064 95804
rect 640116 95792 640122 95804
rect 652018 95792 652024 95804
rect 640116 95764 652024 95792
rect 640116 95752 640122 95764
rect 652018 95752 652024 95764
rect 652076 95752 652082 95804
rect 634722 95616 634728 95668
rect 634780 95656 634786 95668
rect 643094 95656 643100 95668
rect 634780 95628 643100 95656
rect 634780 95616 634786 95628
rect 643094 95616 643100 95628
rect 643152 95616 643158 95668
rect 645578 95616 645584 95668
rect 645636 95656 645642 95668
rect 656158 95656 656164 95668
rect 645636 95628 656164 95656
rect 645636 95616 645642 95628
rect 656158 95616 656164 95628
rect 656216 95616 656222 95668
rect 659194 95616 659200 95668
rect 659252 95656 659258 95668
rect 664162 95656 664168 95668
rect 659252 95628 664168 95656
rect 659252 95616 659258 95628
rect 664162 95616 664168 95628
rect 664220 95616 664226 95668
rect 616506 95140 616512 95192
rect 616564 95180 616570 95192
rect 622670 95180 622676 95192
rect 616564 95152 622676 95180
rect 616564 95140 616570 95152
rect 622670 95140 622676 95152
rect 622728 95140 622734 95192
rect 643738 94596 643744 94648
rect 643796 94636 643802 94648
rect 653398 94636 653404 94648
rect 643796 94608 653404 94636
rect 643796 94596 643802 94608
rect 653398 94596 653404 94608
rect 653456 94596 653462 94648
rect 607674 94460 607680 94512
rect 607732 94500 607738 94512
rect 624970 94500 624976 94512
rect 607732 94472 624976 94500
rect 607732 94460 607738 94472
rect 624970 94460 624976 94472
rect 625028 94460 625034 94512
rect 642910 94460 642916 94512
rect 642968 94500 642974 94512
rect 663242 94500 663248 94512
rect 642968 94472 663248 94500
rect 642968 94460 642974 94472
rect 663242 94460 663248 94472
rect 663300 94460 663306 94512
rect 649626 93984 649632 94036
rect 649684 94024 649690 94036
rect 650638 94024 650644 94036
rect 649684 93996 650644 94024
rect 649684 93984 649690 93996
rect 650638 93984 650644 93996
rect 650696 93984 650702 94036
rect 579522 93780 579528 93832
rect 579580 93820 579586 93832
rect 586514 93820 586520 93832
rect 579580 93792 586520 93820
rect 579580 93780 579586 93792
rect 586514 93780 586520 93792
rect 586572 93780 586578 93832
rect 619542 93780 619548 93832
rect 619600 93820 619606 93832
rect 626442 93820 626448 93832
rect 619600 93792 626448 93820
rect 619600 93780 619606 93792
rect 626442 93780 626448 93792
rect 626500 93780 626506 93832
rect 643278 93780 643284 93832
rect 643336 93820 643342 93832
rect 643336 93792 644474 93820
rect 643336 93780 643342 93792
rect 644446 93752 644474 93792
rect 654134 93752 654140 93764
rect 644446 93724 654140 93752
rect 654134 93712 654140 93724
rect 654192 93712 654198 93764
rect 609698 93100 609704 93152
rect 609756 93140 609762 93152
rect 618898 93140 618904 93152
rect 609756 93112 618904 93140
rect 609756 93100 609762 93112
rect 618898 93100 618904 93112
rect 618956 93100 618962 93152
rect 618070 92420 618076 92472
rect 618128 92460 618134 92472
rect 625430 92460 625436 92472
rect 618128 92432 625436 92460
rect 618128 92420 618134 92432
rect 625430 92420 625436 92432
rect 625488 92420 625494 92472
rect 650914 92420 650920 92472
rect 650972 92460 650978 92472
rect 654318 92460 654324 92472
rect 650972 92432 654324 92460
rect 650972 92420 650978 92432
rect 654318 92420 654324 92432
rect 654376 92420 654382 92472
rect 579522 90992 579528 91044
rect 579580 91032 579586 91044
rect 585962 91032 585968 91044
rect 579580 91004 585968 91032
rect 579580 90992 579586 91004
rect 585962 90992 585968 91004
rect 586020 90992 586026 91044
rect 611262 90992 611268 91044
rect 611320 91032 611326 91044
rect 617334 91032 617340 91044
rect 611320 91004 617340 91032
rect 611320 90992 611326 91004
rect 617334 90992 617340 91004
rect 617392 90992 617398 91044
rect 617886 90992 617892 91044
rect 617944 91032 617950 91044
rect 626442 91032 626448 91044
rect 617944 91004 626448 91032
rect 617944 90992 617950 91004
rect 626442 90992 626448 91004
rect 626500 90992 626506 91044
rect 646498 90992 646504 91044
rect 646556 91032 646562 91044
rect 654134 91032 654140 91044
rect 646556 91004 654140 91032
rect 646556 90992 646562 91004
rect 654134 90992 654140 91004
rect 654192 90992 654198 91044
rect 622670 89632 622676 89684
rect 622728 89672 622734 89684
rect 626442 89672 626448 89684
rect 622728 89644 626448 89672
rect 622728 89632 622734 89644
rect 626442 89632 626448 89644
rect 626500 89632 626506 89684
rect 578510 89564 578516 89616
rect 578568 89604 578574 89616
rect 580626 89604 580632 89616
rect 578568 89576 580632 89604
rect 578568 89564 578574 89576
rect 580626 89564 580632 89576
rect 580684 89564 580690 89616
rect 647142 88952 647148 89004
rect 647200 88992 647206 89004
rect 656894 88992 656900 89004
rect 647200 88964 656900 88992
rect 647200 88952 647206 88964
rect 656894 88952 656900 88964
rect 656952 88952 656958 89004
rect 656158 88748 656164 88800
rect 656216 88788 656222 88800
rect 657446 88788 657452 88800
rect 656216 88760 657452 88788
rect 656216 88748 656222 88760
rect 657446 88748 657452 88760
rect 657504 88748 657510 88800
rect 662322 88748 662328 88800
rect 662380 88788 662386 88800
rect 664162 88788 664168 88800
rect 662380 88760 664168 88788
rect 662380 88748 662386 88760
rect 664162 88748 664168 88760
rect 664220 88748 664226 88800
rect 607306 88272 607312 88324
rect 607364 88312 607370 88324
rect 626442 88312 626448 88324
rect 607364 88284 626448 88312
rect 607364 88272 607370 88284
rect 626442 88272 626448 88284
rect 626500 88272 626506 88324
rect 655238 88272 655244 88324
rect 655296 88312 655302 88324
rect 658458 88312 658464 88324
rect 655296 88284 658464 88312
rect 655296 88272 655302 88284
rect 658458 88272 658464 88284
rect 658516 88272 658522 88324
rect 617334 88136 617340 88188
rect 617392 88176 617398 88188
rect 625614 88176 625620 88188
rect 617392 88148 625620 88176
rect 617392 88136 617398 88148
rect 625614 88136 625620 88148
rect 625672 88136 625678 88188
rect 656526 87252 656532 87304
rect 656584 87292 656590 87304
rect 662506 87292 662512 87304
rect 656584 87264 662512 87292
rect 656584 87252 656590 87264
rect 662506 87252 662512 87264
rect 662564 87252 662570 87304
rect 645762 87116 645768 87168
rect 645820 87156 645826 87168
rect 660666 87156 660672 87168
rect 645820 87128 660672 87156
rect 645820 87116 645826 87128
rect 660666 87116 660672 87128
rect 660724 87116 660730 87168
rect 648338 86980 648344 87032
rect 648396 87020 648402 87032
rect 656526 87020 656532 87032
rect 648396 86992 656532 87020
rect 648396 86980 648402 86992
rect 656526 86980 656532 86992
rect 656584 86980 656590 87032
rect 579522 86912 579528 86964
rect 579580 86952 579586 86964
rect 588722 86952 588728 86964
rect 579580 86924 588728 86952
rect 579580 86912 579586 86924
rect 588722 86912 588728 86924
rect 588780 86912 588786 86964
rect 656710 86912 656716 86964
rect 656768 86952 656774 86964
rect 659562 86952 659568 86964
rect 656768 86924 659568 86952
rect 656768 86912 656774 86924
rect 659562 86912 659568 86924
rect 659620 86912 659626 86964
rect 653398 86708 653404 86760
rect 653456 86748 653462 86760
rect 661402 86748 661408 86760
rect 653456 86720 661408 86748
rect 653456 86708 653462 86720
rect 661402 86708 661408 86720
rect 661460 86708 661466 86760
rect 652018 86572 652024 86624
rect 652076 86612 652082 86624
rect 660114 86612 660120 86624
rect 652076 86584 660120 86612
rect 652076 86572 652082 86584
rect 660114 86572 660120 86584
rect 660172 86572 660178 86624
rect 650638 86436 650644 86488
rect 650696 86476 650702 86488
rect 658826 86476 658832 86488
rect 650696 86448 658832 86476
rect 650696 86436 650702 86448
rect 658826 86436 658832 86448
rect 658884 86436 658890 86488
rect 621658 86232 621664 86284
rect 621716 86272 621722 86284
rect 626442 86272 626448 86284
rect 621716 86244 626448 86272
rect 621716 86232 621722 86244
rect 626442 86232 626448 86244
rect 626500 86232 626506 86284
rect 609882 85484 609888 85536
rect 609940 85524 609946 85536
rect 626442 85524 626448 85536
rect 609940 85496 626448 85524
rect 609940 85484 609946 85496
rect 626442 85484 626448 85496
rect 626500 85484 626506 85536
rect 620278 84124 620284 84176
rect 620336 84164 620342 84176
rect 626258 84164 626264 84176
rect 620336 84136 626264 84164
rect 620336 84124 620342 84136
rect 626258 84124 626264 84136
rect 626316 84124 626322 84176
rect 579338 83988 579344 84040
rect 579396 84028 579402 84040
rect 581822 84028 581828 84040
rect 579396 84000 581828 84028
rect 579396 83988 579402 84000
rect 581822 83988 581828 84000
rect 581880 83988 581886 84040
rect 618898 83988 618904 84040
rect 618956 84028 618962 84040
rect 618956 84000 625154 84028
rect 618956 83988 618962 84000
rect 625126 83960 625154 84000
rect 626442 83960 626448 83972
rect 625126 83932 626448 83960
rect 626442 83920 626448 83932
rect 626500 83920 626506 83972
rect 579522 81336 579528 81388
rect 579580 81376 579586 81388
rect 584582 81376 584588 81388
rect 579580 81348 584588 81376
rect 579580 81336 579586 81348
rect 584582 81336 584588 81348
rect 584640 81336 584646 81388
rect 628558 80928 628564 80980
rect 628616 80968 628622 80980
rect 642450 80968 642456 80980
rect 628616 80940 642456 80968
rect 628616 80928 628622 80940
rect 642450 80928 642456 80940
rect 642508 80928 642514 80980
rect 612642 80792 612648 80844
rect 612700 80832 612706 80844
rect 645854 80832 645860 80844
rect 612700 80804 645860 80832
rect 612700 80792 612706 80804
rect 645854 80792 645860 80804
rect 645912 80792 645918 80844
rect 595622 80656 595628 80708
rect 595680 80696 595686 80708
rect 636102 80696 636108 80708
rect 595680 80668 636108 80696
rect 595680 80656 595686 80668
rect 636102 80656 636108 80668
rect 636160 80656 636166 80708
rect 579246 80044 579252 80096
rect 579304 80084 579310 80096
rect 583202 80084 583208 80096
rect 579304 80056 583208 80084
rect 579304 80044 579310 80056
rect 583202 80044 583208 80056
rect 583260 80044 583266 80096
rect 629202 79432 629208 79484
rect 629260 79472 629266 79484
rect 637482 79472 637488 79484
rect 629260 79444 637488 79472
rect 629260 79432 629266 79444
rect 637482 79432 637488 79444
rect 637540 79432 637546 79484
rect 616782 79296 616788 79348
rect 616840 79336 616846 79348
rect 647418 79336 647424 79348
rect 616840 79308 647424 79336
rect 616840 79296 616846 79308
rect 647418 79296 647424 79308
rect 647476 79296 647482 79348
rect 637482 78208 637488 78260
rect 637540 78248 637546 78260
rect 645302 78248 645308 78260
rect 637540 78220 645308 78248
rect 637540 78208 637546 78220
rect 645302 78208 645308 78220
rect 645360 78208 645366 78260
rect 631042 78072 631048 78124
rect 631100 78112 631106 78124
rect 638954 78112 638960 78124
rect 631100 78084 638960 78112
rect 631100 78072 631106 78084
rect 638954 78072 638960 78084
rect 639012 78072 639018 78124
rect 614022 77936 614028 77988
rect 614080 77976 614086 77988
rect 647602 77976 647608 77988
rect 614080 77948 647608 77976
rect 614080 77936 614086 77948
rect 647602 77936 647608 77948
rect 647660 77936 647666 77988
rect 631042 77704 631048 77716
rect 625126 77676 631048 77704
rect 624418 77392 624424 77444
rect 624476 77432 624482 77444
rect 625126 77432 625154 77676
rect 631042 77664 631048 77676
rect 631100 77664 631106 77716
rect 628282 77528 628288 77580
rect 628340 77568 628346 77580
rect 631502 77568 631508 77580
rect 628340 77540 631508 77568
rect 628340 77528 628346 77540
rect 631502 77528 631508 77540
rect 631560 77528 631566 77580
rect 624476 77404 625154 77432
rect 624476 77392 624482 77404
rect 625798 77392 625804 77444
rect 625856 77432 625862 77444
rect 633894 77432 633900 77444
rect 625856 77404 633900 77432
rect 625856 77392 625862 77404
rect 633894 77392 633900 77404
rect 633952 77392 633958 77444
rect 577498 77256 577504 77308
rect 577556 77296 577562 77308
rect 637114 77296 637120 77308
rect 577556 77268 637120 77296
rect 577556 77256 577562 77268
rect 637114 77256 637120 77268
rect 637172 77296 637178 77308
rect 639598 77296 639604 77308
rect 637172 77268 639604 77296
rect 637172 77256 637178 77268
rect 639598 77256 639604 77268
rect 639656 77256 639662 77308
rect 614758 76644 614764 76696
rect 614816 76684 614822 76696
rect 646314 76684 646320 76696
rect 614816 76656 646320 76684
rect 614816 76644 614822 76656
rect 646314 76644 646320 76656
rect 646372 76644 646378 76696
rect 613378 76508 613384 76560
rect 613436 76548 613442 76560
rect 648982 76548 648988 76560
rect 613436 76520 648988 76548
rect 613436 76508 613442 76520
rect 648982 76508 648988 76520
rect 649040 76508 649046 76560
rect 584582 75896 584588 75948
rect 584640 75936 584646 75948
rect 628282 75936 628288 75948
rect 584640 75908 628288 75936
rect 584640 75896 584646 75908
rect 628282 75896 628288 75908
rect 628340 75896 628346 75948
rect 615402 75284 615408 75336
rect 615460 75324 615466 75336
rect 646130 75324 646136 75336
rect 615460 75296 646136 75324
rect 615460 75284 615466 75296
rect 646130 75284 646136 75296
rect 646188 75284 646194 75336
rect 607122 75148 607128 75200
rect 607180 75188 607186 75200
rect 646866 75188 646872 75200
rect 607180 75160 646872 75188
rect 607180 75148 607186 75160
rect 646866 75148 646872 75160
rect 646924 75148 646930 75200
rect 579522 74468 579528 74520
rect 579580 74508 579586 74520
rect 589918 74508 589924 74520
rect 579580 74480 589924 74508
rect 579580 74468 579586 74480
rect 589918 74468 589924 74480
rect 589976 74468 589982 74520
rect 579522 71476 579528 71528
rect 579580 71516 579586 71528
rect 584398 71516 584404 71528
rect 579580 71488 584404 71516
rect 579580 71476 579586 71488
rect 584398 71476 584404 71488
rect 584456 71476 584462 71528
rect 578510 68960 578516 69012
rect 578568 69000 578574 69012
rect 587158 69000 587164 69012
rect 578568 68972 587164 69000
rect 578568 68960 578574 68972
rect 587158 68960 587164 68972
rect 587216 68960 587222 69012
rect 579522 67464 579528 67516
rect 579580 67504 579586 67516
rect 585778 67504 585784 67516
rect 579580 67476 585784 67504
rect 579580 67464 579586 67476
rect 585778 67464 585784 67476
rect 585836 67464 585842 67516
rect 578510 61956 578516 62008
rect 578568 61996 578574 62008
rect 580258 61996 580264 62008
rect 578568 61968 580264 61996
rect 578568 61956 578574 61968
rect 580258 61956 580264 61968
rect 580316 61956 580322 62008
rect 579522 58964 579528 59016
rect 579580 59004 579586 59016
rect 583018 59004 583024 59016
rect 579580 58976 583024 59004
rect 579580 58964 579586 58976
rect 583018 58964 583024 58976
rect 583076 58964 583082 59016
rect 579062 57876 579068 57928
rect 579120 57916 579126 57928
rect 581638 57916 581644 57928
rect 579120 57888 581644 57916
rect 579120 57876 579126 57888
rect 581638 57876 581644 57888
rect 581696 57876 581702 57928
rect 611998 57196 612004 57248
rect 612056 57236 612062 57248
rect 662414 57236 662420 57248
rect 612056 57208 662420 57236
rect 612056 57196 612062 57208
rect 662414 57196 662420 57208
rect 662472 57196 662478 57248
rect 578510 55156 578516 55208
rect 578568 55196 578574 55208
rect 588538 55196 588544 55208
rect 578568 55168 588544 55196
rect 578568 55156 578574 55168
rect 588538 55156 588544 55168
rect 588596 55156 588602 55208
rect 145374 53048 145380 53100
rect 145432 53088 145438 53100
rect 584582 53088 584588 53100
rect 145432 53060 584588 53088
rect 145432 53048 145438 53060
rect 584582 53048 584588 53060
rect 584640 53048 584646 53100
rect 391934 52436 391940 52488
rect 391992 52476 391998 52488
rect 392578 52476 392584 52488
rect 391992 52448 392584 52476
rect 391992 52436 391998 52448
rect 392578 52436 392584 52448
rect 392636 52476 392642 52488
rect 577498 52476 577504 52488
rect 392636 52448 577504 52476
rect 392636 52436 392642 52448
rect 577498 52436 577504 52448
rect 577556 52436 577562 52488
rect 288158 52300 288164 52352
rect 288216 52340 288222 52352
rect 625798 52340 625804 52352
rect 288216 52312 625804 52340
rect 288216 52300 288222 52312
rect 625798 52300 625804 52312
rect 625856 52300 625862 52352
rect 405090 51688 405096 51740
rect 405148 51728 405154 51740
rect 595438 51728 595444 51740
rect 405148 51700 595444 51728
rect 405148 51688 405154 51700
rect 595438 51688 595444 51700
rect 595496 51688 595502 51740
rect 235810 51008 235816 51060
rect 235868 51048 235874 51060
rect 288158 51048 288164 51060
rect 235868 51020 288164 51048
rect 235868 51008 235874 51020
rect 288158 51008 288164 51020
rect 288216 51008 288222 51060
rect 340506 51008 340512 51060
rect 340564 51048 340570 51060
rect 391934 51048 391940 51060
rect 340564 51020 391940 51048
rect 340564 51008 340570 51020
rect 391934 51008 391940 51020
rect 391992 51008 391998 51060
rect 445202 50464 445208 50516
rect 445260 50504 445266 50516
rect 498102 50504 498108 50516
rect 445260 50476 498108 50504
rect 445260 50464 445266 50476
rect 498102 50464 498108 50476
rect 498160 50464 498166 50516
rect 183462 50328 183468 50380
rect 183520 50368 183526 50380
rect 445018 50368 445024 50380
rect 183520 50340 445024 50368
rect 183520 50328 183526 50340
rect 445018 50328 445024 50340
rect 445076 50328 445082 50380
rect 498102 47268 498108 47320
rect 498160 47308 498166 47320
rect 499574 47308 499580 47320
rect 498160 47280 499580 47308
rect 498160 47268 498166 47280
rect 499574 47268 499580 47280
rect 499632 47268 499638 47320
rect 194042 44820 194048 44872
rect 194100 44860 194106 44872
rect 662598 44860 662604 44872
rect 194100 44832 662604 44860
rect 194100 44820 194106 44832
rect 662598 44820 662604 44832
rect 662656 44820 662662 44872
rect 315942 43392 315948 43444
rect 316000 43432 316006 43444
rect 663794 43432 663800 43444
rect 316000 43404 663800 43432
rect 316000 43392 316006 43404
rect 663794 43392 663800 43404
rect 663852 43392 663858 43444
rect 409598 42340 409604 42392
rect 409656 42340 409662 42392
rect 464890 42328 464896 42380
rect 464948 42328 464954 42380
rect 315942 42173 315948 42225
rect 316000 42173 316006 42225
<< via1 >>
rect 366180 1027828 366232 1027880
rect 366548 1027828 366600 1027880
rect 366180 1024360 366232 1024412
rect 366548 1024360 366600 1024412
rect 504548 1007020 504600 1007072
rect 514208 1007020 514260 1007072
rect 554136 1006952 554188 1007004
rect 559656 1006952 559708 1007004
rect 506204 1006884 506256 1006936
rect 514024 1006884 514076 1006936
rect 145748 1006816 145800 1006868
rect 151728 1006816 151780 1006868
rect 428004 1006816 428056 1006868
rect 439504 1006816 439556 1006868
rect 555148 1006816 555200 1006868
rect 562324 1006816 562376 1006868
rect 300124 1006680 300176 1006732
rect 307760 1006680 307812 1006732
rect 357716 1006680 357768 1006732
rect 374000 1006680 374052 1006732
rect 400864 1006680 400916 1006732
rect 430856 1006680 430908 1006732
rect 557172 1006680 557224 1006732
rect 566648 1006680 566700 1006732
rect 144552 1006544 144604 1006596
rect 151452 1006544 151504 1006596
rect 298744 1006544 298796 1006596
rect 306104 1006544 306156 1006596
rect 427176 1006544 427228 1006596
rect 445024 1006544 445076 1006596
rect 94688 1006408 94740 1006460
rect 101128 1006408 101180 1006460
rect 148324 1006408 148376 1006460
rect 249064 1006408 249116 1006460
rect 255320 1006408 255372 1006460
rect 304080 1006408 304132 1006460
rect 152096 1006340 152148 1006392
rect 210424 1006340 210476 1006392
rect 228364 1006340 228416 1006392
rect 94504 1006272 94556 1006324
rect 100300 1006272 100352 1006324
rect 144184 1006272 144236 1006324
rect 150900 1006272 150952 1006324
rect 158260 1006272 158312 1006324
rect 93124 1006136 93176 1006188
rect 99472 1006136 99524 1006188
rect 102784 1006136 102836 1006188
rect 103980 1006136 104032 1006188
rect 106832 1006136 106884 1006188
rect 124864 1006136 124916 1006188
rect 145564 1006136 145616 1006188
rect 151268 1006136 151320 1006188
rect 151452 1006136 151504 1006188
rect 159456 1006136 159508 1006188
rect 160284 1006136 160336 1006188
rect 164884 1006136 164936 1006188
rect 250260 1006272 250312 1006324
rect 254124 1006272 254176 1006324
rect 298928 1006272 298980 1006324
rect 305276 1006272 305328 1006324
rect 208400 1006204 208452 1006256
rect 175924 1006136 175976 1006188
rect 247868 1006136 247920 1006188
rect 253664 1006136 253716 1006188
rect 262680 1006136 262732 1006188
rect 278044 1006136 278096 1006188
rect 300308 1006136 300360 1006188
rect 306932 1006272 306984 1006324
rect 314660 1006408 314712 1006460
rect 319444 1006408 319496 1006460
rect 361396 1006408 361448 1006460
rect 371884 1006408 371936 1006460
rect 423496 1006408 423548 1006460
rect 447140 1006408 447192 1006460
rect 501696 1006408 501748 1006460
rect 518164 1006408 518216 1006460
rect 331864 1006272 331916 1006324
rect 424324 1006272 424376 1006324
rect 438860 1006272 438912 1006324
rect 502156 1006272 502208 1006324
rect 520924 1006408 520976 1006460
rect 552296 1006408 552348 1006460
rect 554780 1006408 554832 1006460
rect 556804 1006408 556856 1006460
rect 569224 1006408 569276 1006460
rect 554320 1006272 554372 1006324
rect 306104 1006136 306156 1006188
rect 311808 1006136 311860 1006188
rect 314660 1006136 314712 1006188
rect 324964 1006136 325016 1006188
rect 365076 1006136 365128 1006188
rect 367744 1006136 367796 1006188
rect 500500 1006136 500552 1006188
rect 505744 1006136 505796 1006188
rect 93308 1006000 93360 1006052
rect 98276 1006000 98328 1006052
rect 101404 1006000 101456 1006052
rect 104808 1006000 104860 1006052
rect 107660 1006000 107712 1006052
rect 126244 1006000 126296 1006052
rect 148876 1006000 148928 1006052
rect 150072 1006000 150124 1006052
rect 158628 1006000 158680 1006052
rect 177304 1006000 177356 1006052
rect 198004 1006000 198056 1006052
rect 201040 1006000 201092 1006052
rect 229744 1006000 229796 1006052
rect 247684 1006000 247736 1006052
rect 250260 1006000 250312 1006052
rect 250444 1006000 250496 1006052
rect 252468 1006000 252520 1006052
rect 261852 1006000 261904 1006052
rect 280804 1006000 280856 1006052
rect 303252 1006000 303304 1006052
rect 304080 1006000 304132 1006052
rect 305276 1006000 305328 1006052
rect 332048 1006000 332100 1006052
rect 354864 1006000 354916 1006052
rect 356704 1006000 356756 1006052
rect 357348 1006000 357400 1006052
rect 376024 1006000 376076 1006052
rect 423496 1006000 423548 1006052
rect 427820 1006000 427872 1006052
rect 429200 1006000 429252 1006052
rect 471244 1006000 471296 1006052
rect 499672 1006000 499724 1006052
rect 502984 1006000 503036 1006052
rect 505376 1006000 505428 1006052
rect 516784 1006136 516836 1006188
rect 551468 1006136 551520 1006188
rect 555424 1006136 555476 1006188
rect 514024 1006000 514076 1006052
rect 522304 1006000 522356 1006052
rect 553124 1006000 553176 1006052
rect 556804 1006000 556856 1006052
rect 562324 1006272 562376 1006324
rect 571984 1006272 572036 1006324
rect 560852 1006136 560904 1006188
rect 563980 1006136 564032 1006188
rect 574744 1006000 574796 1006052
rect 428372 1005796 428424 1005848
rect 440884 1005796 440936 1005848
rect 509056 1005796 509108 1005848
rect 514024 1005796 514076 1005848
rect 360568 1005660 360620 1005712
rect 377404 1005660 377456 1005712
rect 427544 1005660 427596 1005712
rect 359740 1005524 359792 1005576
rect 373264 1005524 373316 1005576
rect 430856 1005524 430908 1005576
rect 433984 1005524 434036 1005576
rect 438860 1005660 438912 1005712
rect 451924 1005660 451976 1005712
rect 555976 1005660 556028 1005712
rect 563060 1005660 563112 1005712
rect 449164 1005524 449216 1005576
rect 505008 1005524 505060 1005576
rect 356520 1005388 356572 1005440
rect 378784 1005388 378836 1005440
rect 431960 1005388 432012 1005440
rect 443644 1005388 443696 1005440
rect 447140 1005388 447192 1005440
rect 457444 1005388 457496 1005440
rect 508228 1005388 508280 1005440
rect 510988 1005388 511040 1005440
rect 554780 1005524 554832 1005576
rect 567844 1005796 567896 1005848
rect 563980 1005660 564032 1005712
rect 570604 1005660 570656 1005712
rect 522488 1005388 522540 1005440
rect 555148 1005388 555200 1005440
rect 573548 1005388 573600 1005440
rect 425520 1005320 425572 1005372
rect 431776 1005320 431828 1005372
rect 263048 1005252 263100 1005304
rect 279424 1005252 279476 1005304
rect 356888 1005252 356940 1005304
rect 381544 1005252 381596 1005304
rect 149704 1005184 149756 1005236
rect 152924 1005184 152976 1005236
rect 304264 1005184 304316 1005236
rect 307300 1005184 307352 1005236
rect 430028 1005184 430080 1005236
rect 432420 1005252 432472 1005304
rect 465724 1005252 465776 1005304
rect 500500 1005252 500552 1005304
rect 519544 1005252 519596 1005304
rect 551100 1005252 551152 1005304
rect 573364 1005252 573416 1005304
rect 432604 1005116 432656 1005168
rect 507032 1005116 507084 1005168
rect 509700 1005116 509752 1005168
rect 151084 1005048 151136 1005100
rect 153752 1005048 153804 1005100
rect 363420 1005048 363472 1005100
rect 364524 1005048 364576 1005100
rect 365076 1005048 365128 1005100
rect 370504 1005048 370556 1005100
rect 424692 1005048 424744 1005100
rect 431500 1005048 431552 1005100
rect 431684 1005048 431736 1005100
rect 434168 1004980 434220 1005032
rect 508228 1004980 508280 1005032
rect 511264 1004980 511316 1005032
rect 149888 1004912 149940 1004964
rect 152924 1004912 152976 1004964
rect 154396 1004912 154448 1004964
rect 160652 1004912 160704 1004964
rect 209228 1004912 209280 1004964
rect 211804 1004912 211856 1004964
rect 305828 1004912 305880 1004964
rect 308956 1004912 309008 1004964
rect 353208 1004912 353260 1004964
rect 355692 1004912 355744 1004964
rect 361396 1004912 361448 1004964
rect 365168 1004912 365220 1004964
rect 429200 1004912 429252 1004964
rect 431914 1004912 431966 1004964
rect 432420 1004844 432472 1004896
rect 438124 1004844 438176 1004896
rect 507860 1004844 507912 1004896
rect 510068 1004844 510120 1004896
rect 151268 1004776 151320 1004828
rect 154120 1004776 154172 1004828
rect 159456 1004776 159508 1004828
rect 162124 1004776 162176 1004828
rect 207204 1004776 207256 1004828
rect 209872 1004776 209924 1004828
rect 304448 1004776 304500 1004828
rect 306932 1004776 306984 1004828
rect 313832 1004776 313884 1004828
rect 316040 1004776 316092 1004828
rect 364248 1004776 364300 1004828
rect 366364 1004776 366416 1004828
rect 430028 1004776 430080 1004828
rect 432236 1004776 432288 1004828
rect 498108 1004776 498160 1004828
rect 499672 1004776 499724 1004828
rect 555976 1004776 556028 1004828
rect 558184 1004776 558236 1004828
rect 94872 1004640 94924 1004692
rect 103152 1004640 103204 1004692
rect 106188 1004640 106240 1004692
rect 108488 1004640 108540 1004692
rect 160652 1004640 160704 1004692
rect 162860 1004640 162912 1004692
rect 209228 1004640 209280 1004692
rect 211160 1004640 211212 1004692
rect 212540 1004640 212592 1004692
rect 217324 1004640 217376 1004692
rect 305644 1004640 305696 1004692
rect 308128 1004640 308180 1004692
rect 315488 1004640 315540 1004692
rect 318064 1004640 318116 1004692
rect 354588 1004640 354640 1004692
rect 355692 1004640 355744 1004692
rect 362592 1004640 362644 1004692
rect 364984 1004640 365036 1004692
rect 431684 1004640 431736 1004692
rect 433524 1004640 433576 1004692
rect 499488 1004640 499540 1004692
rect 501328 1004640 501380 1004692
rect 509056 1004640 509108 1004692
rect 364524 1004504 364576 1004556
rect 366548 1004504 366600 1004556
rect 510344 1004640 510396 1004692
rect 515404 1004640 515456 1004692
rect 557632 1004640 557684 1004692
rect 559564 1004640 559616 1004692
rect 561680 1004640 561732 1004692
rect 566464 1004640 566516 1004692
rect 510804 1004504 510856 1004556
rect 432880 1004028 432932 1004080
rect 462320 1004028 462372 1004080
rect 425520 1003892 425572 1003944
rect 467840 1003892 467892 1003944
rect 505376 1003892 505428 1003944
rect 516600 1003892 516652 1003944
rect 445024 1002804 445076 1002856
rect 454684 1002804 454736 1002856
rect 558828 1002736 558880 1002788
rect 562324 1002736 562376 1002788
rect 424692 1002668 424744 1002720
rect 446220 1002668 446272 1002720
rect 97264 1002600 97316 1002652
rect 102324 1002600 102376 1002652
rect 558000 1002600 558052 1002652
rect 560300 1002600 560352 1002652
rect 106004 1002532 106056 1002584
rect 109500 1002532 109552 1002584
rect 427820 1002532 427872 1002584
rect 468760 1002532 468812 1002584
rect 502524 1002532 502576 1002584
rect 516048 1002532 516100 1002584
rect 563060 1002532 563112 1002584
rect 571248 1002532 571300 1002584
rect 98644 1002464 98696 1002516
rect 101956 1002464 102008 1002516
rect 157432 1002464 157484 1002516
rect 159364 1002464 159416 1002516
rect 203340 1002464 203392 1002516
rect 206376 1002464 206428 1002516
rect 251824 1002464 251876 1002516
rect 255320 1002464 255372 1002516
rect 261024 1002464 261076 1002516
rect 264244 1002464 264296 1002516
rect 108028 1002396 108080 1002448
rect 110420 1002396 110472 1002448
rect 558000 1002396 558052 1002448
rect 561036 1002396 561088 1002448
rect 97448 1002328 97500 1002380
rect 100300 1002328 100352 1002380
rect 158628 1002328 158680 1002380
rect 160376 1002328 160428 1002380
rect 211252 1002328 211304 1002380
rect 215944 1002328 215996 1002380
rect 253112 1002328 253164 1002380
rect 256148 1002328 256200 1002380
rect 310152 1002328 310204 1002380
rect 311900 1002328 311952 1002380
rect 358544 1002328 358596 1002380
rect 360844 1002328 360896 1002380
rect 105636 1002260 105688 1002312
rect 107844 1002260 107896 1002312
rect 108488 1002260 108540 1002312
rect 111064 1002260 111116 1002312
rect 153936 1002260 153988 1002312
rect 155776 1002260 155828 1002312
rect 551928 1002260 551980 1002312
rect 554320 1002260 554372 1002312
rect 560484 1002260 560536 1002312
rect 563060 1002260 563112 1002312
rect 98828 1002192 98880 1002244
rect 101128 1002192 101180 1002244
rect 156604 1002192 156656 1002244
rect 158720 1002192 158772 1002244
rect 204904 1002192 204956 1002244
rect 206376 1002192 206428 1002244
rect 252008 1002192 252060 1002244
rect 254492 1002192 254544 1002244
rect 303068 1002192 303120 1002244
rect 306104 1002192 306156 1002244
rect 359372 1002192 359424 1002244
rect 500684 1002192 500736 1002244
rect 503352 1002192 503404 1002244
rect 104808 1002124 104860 1002176
rect 106372 1002124 106424 1002176
rect 106832 1002124 106884 1002176
rect 109040 1002124 109092 1002176
rect 152648 1002124 152700 1002176
rect 154580 1002124 154632 1002176
rect 96528 1002056 96580 1002108
rect 99104 1002056 99156 1002108
rect 100208 1002056 100260 1002108
rect 103152 1002056 103204 1002108
rect 109684 1002056 109736 1002108
rect 111892 1002056 111944 1002108
rect 148968 1002056 149020 1002108
rect 150900 1002056 150952 1002108
rect 154948 1002056 155000 1002108
rect 157340 1002056 157392 1002108
rect 211252 1002056 211304 1002108
rect 213184 1002056 213236 1002108
rect 250996 1002056 251048 1002108
rect 253296 1002056 253348 1002108
rect 253480 1002056 253532 1002108
rect 256148 1002056 256200 1002108
rect 263508 1002056 263560 1002108
rect 265624 1002056 265676 1002108
rect 307024 1002056 307076 1002108
rect 308956 1002056 309008 1002108
rect 310980 1002056 311032 1002108
rect 313280 1002056 313332 1002108
rect 106004 1001988 106056 1002040
rect 107752 1001988 107804 1002040
rect 152464 1001988 152516 1002040
rect 153752 1001988 153804 1002040
rect 358728 1001988 358780 1002040
rect 560024 1002124 560076 1002176
rect 562508 1002124 562560 1002176
rect 360568 1002056 360620 1002108
rect 363604 1002056 363656 1002108
rect 433340 1002056 433392 1002108
rect 436744 1002056 436796 1002108
rect 502248 1002056 502300 1002108
rect 504180 1002056 504232 1002108
rect 509884 1002056 509936 1002108
rect 512644 1002056 512696 1002108
rect 553308 1001988 553360 1002040
rect 553952 1001988 554004 1002040
rect 560852 1001988 560904 1002040
rect 565084 1001988 565136 1002040
rect 96344 1001920 96396 1001972
rect 98276 1001920 98328 1001972
rect 100024 1001920 100076 1001972
rect 101956 1001920 102008 1001972
rect 108856 1001920 108908 1001972
rect 112076 1001920 112128 1001972
rect 147588 1001920 147640 1001972
rect 149244 1001920 149296 1001972
rect 154580 1001920 154632 1001972
rect 155776 1001920 155828 1001972
rect 157800 1001920 157852 1001972
rect 160192 1001920 160244 1001972
rect 195336 1001920 195388 1001972
rect 203892 1001920 203944 1001972
rect 204168 1001920 204220 1001972
rect 205548 1001920 205600 1001972
rect 212080 1001920 212132 1001972
rect 213920 1001920 213972 1001972
rect 249708 1001920 249760 1001972
rect 252468 1001920 252520 1001972
rect 261024 1001920 261076 1001972
rect 263600 1001920 263652 1001972
rect 263876 1001920 263928 1001972
rect 267004 1001920 267056 1001972
rect 302884 1001920 302936 1001972
rect 306104 1001920 306156 1001972
rect 308404 1001920 308456 1001972
rect 309784 1001920 309836 1001972
rect 312636 1001920 312688 1001972
rect 314660 1001920 314712 1001972
rect 351828 1001920 351880 1001972
rect 354036 1001920 354088 1001972
rect 355968 1001920 356020 1001972
rect 357348 1001920 357400 1001972
rect 360200 1001920 360252 1001972
rect 362224 1001920 362276 1001972
rect 365904 1001920 365956 1001972
rect 369124 1001920 369176 1001972
rect 419448 1001920 419500 1001972
rect 421472 1001920 421524 1001972
rect 425060 1001920 425112 1001972
rect 426348 1001920 426400 1001972
rect 426532 1001920 426584 1001972
rect 427820 1001920 427872 1001972
rect 428372 1001920 428424 1001972
rect 431224 1001920 431276 1001972
rect 467840 1001920 467892 1001972
rect 472624 1001920 472676 1001972
rect 496728 1001920 496780 1001972
rect 498476 1001920 498528 1001972
rect 500868 1001920 500920 1001972
rect 502524 1001920 502576 1001972
rect 503352 1001920 503404 1001972
rect 504364 1001920 504416 1001972
rect 506204 1001920 506256 1001972
rect 507860 1001920 507912 1001972
rect 558828 1001920 558880 1001972
rect 560392 1001920 560444 1001972
rect 439504 1001172 439556 1001224
rect 446404 1001172 446456 1001224
rect 500684 1001172 500736 1001224
rect 520004 1001172 520056 1001224
rect 298468 1000424 298520 1000476
rect 309140 1000424 309192 1000476
rect 92664 999744 92716 999796
rect 98828 999744 98880 999796
rect 427820 999744 427872 999796
rect 437480 999744 437532 999796
rect 446220 999744 446272 999796
rect 459560 999744 459612 999796
rect 195980 999132 196032 999184
rect 203524 999132 203576 999184
rect 249340 999132 249392 999184
rect 250444 999132 250496 999184
rect 301044 999132 301096 999184
rect 303068 999132 303120 999184
rect 374000 999132 374052 999184
rect 381728 999132 381780 999184
rect 438124 999064 438176 999116
rect 443460 999064 443512 999116
rect 449164 999064 449216 999116
rect 451740 999064 451792 999116
rect 516600 999064 516652 999116
rect 520188 999064 520240 999116
rect 300860 998996 300912 999048
rect 304448 998996 304500 999048
rect 451924 998996 451976 999048
rect 456800 998996 456852 999048
rect 199844 998792 199896 998844
rect 199384 998656 199436 998708
rect 204352 998656 204404 998708
rect 196624 998520 196676 998572
rect 202696 998520 202748 998572
rect 371884 998792 371936 998844
rect 383108 998792 383160 998844
rect 443644 998724 443696 998776
rect 445760 998724 445812 998776
rect 353208 998656 353260 998708
rect 372896 998656 372948 998708
rect 553308 998588 553360 998640
rect 555148 998588 555200 998640
rect 206284 998520 206336 998572
rect 355968 998520 356020 998572
rect 376300 998520 376352 998572
rect 516784 998520 516836 998572
rect 522948 998520 523000 998572
rect 555424 998520 555476 998572
rect 568488 998520 568540 998572
rect 195520 998384 195572 998436
rect 204168 998384 204220 998436
rect 360844 998384 360896 998436
rect 383292 998384 383344 998436
rect 446404 998384 446456 998436
rect 472440 998384 472492 998436
rect 502248 998384 502300 998436
rect 517060 998384 517112 998436
rect 553124 998384 553176 998436
rect 569868 998384 569920 998436
rect 92296 998248 92348 998300
rect 94872 998248 94924 998300
rect 202144 998180 202196 998232
rect 205548 998180 205600 998232
rect 258172 998112 258224 998164
rect 259460 998112 259512 998164
rect 378784 998112 378836 998164
rect 381268 998112 381320 998164
rect 195152 997772 195204 997824
rect 202696 998044 202748 998096
rect 260196 998044 260248 998096
rect 262864 998044 262916 998096
rect 376024 998044 376076 998096
rect 378416 998044 378468 998096
rect 591120 998044 591172 998096
rect 625804 998044 625856 998096
rect 254584 997976 254636 998028
rect 257344 997976 257396 998028
rect 198648 997908 198700 997960
rect 200672 997908 200724 997960
rect 200856 997908 200908 997960
rect 203524 997908 203576 997960
rect 259828 997908 259880 997960
rect 262220 997908 262272 997960
rect 520004 997908 520056 997960
rect 523868 997908 523920 997960
rect 549168 997908 549220 997960
rect 551100 997908 551152 997960
rect 621020 997908 621072 997960
rect 625620 997908 625672 997960
rect 246856 997840 246908 997892
rect 249064 997840 249116 997892
rect 254768 997840 254820 997892
rect 256976 997840 257028 997892
rect 200028 997772 200080 997824
rect 201868 997772 201920 997824
rect 202328 997772 202380 997824
rect 204720 997772 204772 997824
rect 260196 997772 260248 997824
rect 260932 997772 260984 997824
rect 298100 997772 298152 997824
rect 302884 997772 302936 997824
rect 303252 997772 303304 997824
rect 305828 997772 305880 997824
rect 522488 997772 522540 997824
rect 524052 997772 524104 997824
rect 547788 997772 547840 997824
rect 550272 997772 550324 997824
rect 551284 997772 551336 997824
rect 552296 997772 552348 997824
rect 591304 997772 591356 997824
rect 625252 997772 625304 997824
rect 92480 997704 92532 997756
rect 106372 997704 106424 997756
rect 144828 997704 144880 997756
rect 153936 997704 153988 997756
rect 246672 997704 246724 997756
rect 254768 997704 254820 997756
rect 362224 997704 362276 997756
rect 372528 997704 372580 997756
rect 431224 997704 431276 997756
rect 439872 997704 439924 997756
rect 500868 997704 500920 997756
rect 516692 997704 516744 997756
rect 164884 997636 164936 997688
rect 170312 997636 170364 997688
rect 551928 997636 551980 997688
rect 621020 997636 621072 997688
rect 359464 997568 359516 997620
rect 372344 997568 372396 997620
rect 425060 997568 425112 997620
rect 439688 997568 439740 997620
rect 514208 997568 514260 997620
rect 516876 997568 516928 997620
rect 558184 997500 558236 997552
rect 590568 997500 590620 997552
rect 574744 997364 574796 997416
rect 591304 997364 591356 997416
rect 144368 997296 144420 997348
rect 149888 997296 149940 997348
rect 551284 997296 551336 997348
rect 572720 997296 572772 997348
rect 200212 997228 200264 997280
rect 203340 997228 203392 997280
rect 319444 997160 319496 997212
rect 332600 997160 332652 997212
rect 556804 997160 556856 997212
rect 570236 997160 570288 997212
rect 573548 997160 573600 997212
rect 622400 997160 622452 997212
rect 318064 997024 318116 997076
rect 349160 997024 349212 997076
rect 363604 997024 363656 997076
rect 372712 997024 372764 997076
rect 437480 997024 437532 997076
rect 448520 997024 448572 997076
rect 457444 997024 457496 997076
rect 471796 997024 471848 997076
rect 567844 997024 567896 997076
rect 618168 997024 618220 997076
rect 106924 996888 106976 996940
rect 111892 996888 111944 996940
rect 566648 996888 566700 996940
rect 590568 996888 590620 996940
rect 571248 996752 571300 996804
rect 591120 996752 591172 996804
rect 421012 996412 421064 996464
rect 425060 996412 425112 996464
rect 366548 996208 366600 996260
rect 375472 996208 375524 996260
rect 504364 996208 504416 996260
rect 510988 996208 511040 996260
rect 516048 996208 516100 996260
rect 523684 996208 523736 996260
rect 109500 996072 109552 996124
rect 158720 996072 158772 996124
rect 159364 996072 159416 996124
rect 208400 996072 208452 996124
rect 229744 996072 229796 996124
rect 262220 996072 262272 996124
rect 262864 996072 262916 996124
rect 313280 996072 313332 996124
rect 364984 996072 365036 996124
rect 432236 996072 432288 996124
rect 471244 996072 471296 996124
rect 507860 996072 507912 996124
rect 509700 996072 509752 996124
rect 560392 996072 560444 996124
rect 572720 996072 572772 996124
rect 625436 996072 625488 996124
rect 126244 995936 126296 995988
rect 160376 995936 160428 995988
rect 162124 995936 162176 995988
rect 210056 995936 210108 995988
rect 213184 995936 213236 995988
rect 261116 995936 261168 995988
rect 264244 995936 264296 995988
rect 281908 995936 281960 995988
rect 298652 995936 298704 995988
rect 314660 995936 314712 995988
rect 365168 995936 365220 995988
rect 432052 995936 432104 995988
rect 434168 995936 434220 995988
rect 510804 995936 510856 995988
rect 511264 995936 511316 995988
rect 563060 995936 563112 995988
rect 124864 995800 124916 995852
rect 160192 995800 160244 995852
rect 175924 995800 175976 995852
rect 211160 995800 211212 995852
rect 228364 995800 228416 995852
rect 263600 995800 263652 995852
rect 278044 995800 278096 995852
rect 316040 995800 316092 995852
rect 366364 995800 366416 995852
rect 433524 995800 433576 995852
rect 433984 995800 434036 995852
rect 504364 995800 504416 995852
rect 510068 995800 510120 995852
rect 554136 995800 554188 995852
rect 618168 995800 618220 995852
rect 625252 995800 625304 995852
rect 143448 995528 143500 995580
rect 146944 995528 146996 995580
rect 195244 995528 195296 995580
rect 204904 995528 204956 995580
rect 298100 995528 298152 995580
rect 310612 995528 310664 995580
rect 324964 995528 325016 995580
rect 364984 995528 365036 995580
rect 375472 995528 375524 995580
rect 111064 995392 111116 995444
rect 144552 995392 144604 995444
rect 89628 995324 89680 995376
rect 92480 995324 92532 995376
rect 142068 995256 142120 995308
rect 152648 995392 152700 995444
rect 211804 995392 211856 995444
rect 260932 995392 260984 995444
rect 281908 995392 281960 995444
rect 194324 995324 194376 995376
rect 195520 995324 195572 995376
rect 294696 995324 294748 995376
rect 146944 995256 146996 995308
rect 152464 995256 152516 995308
rect 242072 995256 242124 995308
rect 246856 995256 246908 995308
rect 280804 995188 280856 995240
rect 298652 995392 298704 995444
rect 295248 995256 295300 995308
rect 298468 995256 298520 995308
rect 383292 995528 383344 995580
rect 385040 995528 385092 995580
rect 440884 995528 440936 995580
rect 472256 995528 472308 995580
rect 472440 995528 472492 995580
rect 473360 995528 473412 995580
rect 524052 995528 524104 995580
rect 524788 995528 524840 995580
rect 625252 995528 625304 995580
rect 625620 995528 625672 995580
rect 625804 995528 625856 995580
rect 626540 995528 626592 995580
rect 381728 995392 381780 995444
rect 388628 995392 388680 995444
rect 432604 995392 432656 995444
rect 506480 995392 506532 995444
rect 523868 995392 523920 995444
rect 525340 995392 525392 995444
rect 400864 995324 400916 995376
rect 523684 995256 523736 995308
rect 529020 995392 529072 995444
rect 77668 995120 77720 995172
rect 97264 995120 97316 995172
rect 137928 995120 137980 995172
rect 144184 995120 144236 995172
rect 242716 995120 242768 995172
rect 253480 995120 253532 995172
rect 296628 995120 296680 995172
rect 305644 995188 305696 995240
rect 489736 995188 489788 995240
rect 377404 995120 377456 995172
rect 384672 995120 384724 995172
rect 294696 995052 294748 995104
rect 296444 995052 296496 995104
rect 77024 994984 77076 995036
rect 102784 994984 102836 995036
rect 181444 994984 181496 995036
rect 207020 994984 207072 995036
rect 232872 994984 232924 995036
rect 258080 994984 258132 995036
rect 358728 994984 358780 995036
rect 398840 994984 398892 995036
rect 129740 994916 129792 994968
rect 155960 994916 156012 994968
rect 282828 994916 282880 994968
rect 311900 994916 311952 994968
rect 422944 994916 422996 994968
rect 522304 995120 522356 995172
rect 560576 995392 560628 995444
rect 622400 995392 622452 995444
rect 640708 995324 640760 995376
rect 571984 995256 572036 995308
rect 625252 995256 625304 995308
rect 625436 995256 625488 995308
rect 631508 995256 631560 995308
rect 569868 995120 569920 995172
rect 630128 995120 630180 995172
rect 633992 995120 634044 995172
rect 499488 994984 499540 995036
rect 530032 994984 530084 995036
rect 555148 994984 555200 995036
rect 625114 994984 625166 995036
rect 625252 994984 625304 995036
rect 629576 994984 629628 995036
rect 635188 994984 635240 995036
rect 78312 994848 78364 994900
rect 101404 994848 101456 994900
rect 180156 994848 180208 994900
rect 209872 994848 209924 994900
rect 232228 994848 232280 994900
rect 242900 994848 242952 994900
rect 244556 994848 244608 994900
rect 259460 994848 259512 994900
rect 372712 994848 372764 994900
rect 397000 994848 397052 994900
rect 502984 994848 503036 994900
rect 538036 994848 538088 994900
rect 573364 994848 573416 994900
rect 639512 994848 639564 994900
rect 128452 994780 128504 994832
rect 154580 994780 154632 994832
rect 284116 994780 284168 994832
rect 298100 994780 298152 994832
rect 448520 994780 448572 994832
rect 81348 994712 81400 994764
rect 98644 994712 98696 994764
rect 180616 994712 180668 994764
rect 202144 994712 202196 994764
rect 235908 994712 235960 994764
rect 242716 994712 242768 994764
rect 243084 994712 243136 994764
rect 255964 994712 256016 994764
rect 356704 994712 356756 994764
rect 378600 994712 378652 994764
rect 129096 994644 129148 994696
rect 151084 994644 151136 994696
rect 285956 994644 286008 994696
rect 308404 994644 308456 994696
rect 90272 994576 90324 994628
rect 93308 994576 93360 994628
rect 135904 994508 135956 994560
rect 142068 994508 142120 994560
rect 180616 994440 180668 994492
rect 195980 994576 196032 994628
rect 231584 994576 231636 994628
rect 183284 994440 183336 994492
rect 195244 994440 195296 994492
rect 234528 994440 234580 994492
rect 243360 994440 243412 994492
rect 243728 994576 243780 994628
rect 253112 994576 253164 994628
rect 372896 994576 372948 994628
rect 393964 994712 394016 994764
rect 459560 994644 459612 994696
rect 484124 994644 484176 994696
rect 486608 994780 486660 994832
rect 489736 994780 489788 994832
rect 505744 994712 505796 994764
rect 533988 994712 534040 994764
rect 487804 994644 487856 994696
rect 283472 994508 283524 994560
rect 296628 994508 296680 994560
rect 257344 994440 257396 994492
rect 378600 994440 378652 994492
rect 397644 994576 397696 994628
rect 504548 994576 504600 994628
rect 539232 994712 539284 994764
rect 569224 994712 569276 994764
rect 639052 994712 639104 994764
rect 625160 994576 625212 994628
rect 630864 994576 630916 994628
rect 468760 994508 468812 994560
rect 482928 994508 482980 994560
rect 565084 994508 565136 994560
rect 592040 994508 592092 994560
rect 132132 994372 132184 994424
rect 143448 994372 143500 994424
rect 472256 994372 472308 994424
rect 485964 994372 486016 994424
rect 549168 994372 549220 994424
rect 667940 994372 667992 994424
rect 235264 994304 235316 994356
rect 243728 994304 243780 994356
rect 88708 994236 88760 994288
rect 121736 994236 121788 994288
rect 140136 994236 140188 994288
rect 186504 994236 186556 994288
rect 207756 994236 207808 994288
rect 213920 994236 213972 994288
rect 294880 994236 294932 994288
rect 381176 994236 381228 994288
rect 425060 994236 425112 994288
rect 446128 994236 446180 994288
rect 547788 994236 547840 994288
rect 666560 994236 666612 994288
rect 243360 994168 243412 994220
rect 244556 994168 244608 994220
rect 265624 994100 265676 994152
rect 267740 994100 267792 994152
rect 568488 994100 568540 994152
rect 635832 994100 635884 994152
rect 496728 993284 496780 993336
rect 666744 993284 666796 993336
rect 351828 993148 351880 993200
rect 667388 993148 667440 993200
rect 51724 993012 51776 993064
rect 107936 993012 107988 993064
rect 148968 993012 149020 993064
rect 652760 993012 652812 993064
rect 46204 992876 46256 992928
rect 107752 992876 107804 992928
rect 147588 992876 147640 992928
rect 652484 992876 652536 992928
rect 512644 991856 512696 991908
rect 527640 991856 527692 991908
rect 563704 991856 563756 991908
rect 576308 991856 576360 991908
rect 267004 991720 267056 991772
rect 284300 991720 284352 991772
rect 367744 991720 367796 991772
rect 415032 991720 415084 991772
rect 419448 991720 419500 991772
rect 666928 991720 666980 991772
rect 73436 991584 73488 991636
rect 112076 991584 112128 991636
rect 198648 991584 198700 991636
rect 650920 991584 650972 991636
rect 50344 991448 50396 991500
rect 110420 991448 110472 991500
rect 138296 991448 138348 991500
rect 162860 991448 162912 991500
rect 200028 991448 200080 991500
rect 651472 991448 651524 991500
rect 562508 990224 562560 990276
rect 672724 990224 672776 990276
rect 48964 990088 49016 990140
rect 109040 990088 109092 990140
rect 249708 990088 249760 990140
rect 650092 990088 650144 990140
rect 422208 988864 422260 988916
rect 668308 988864 668360 988916
rect 250996 988728 251048 988780
rect 650736 988728 650788 988780
rect 562324 987640 562376 987692
rect 658924 987640 658976 987692
rect 354588 987504 354640 987556
rect 668124 987504 668176 987556
rect 96344 987368 96396 987420
rect 651104 987368 651156 987420
rect 203156 986620 203208 986672
rect 207756 986620 207808 986672
rect 217324 986620 217376 986672
rect 219440 986620 219492 986672
rect 566464 986212 566516 986264
rect 608784 986212 608836 986264
rect 370504 986076 370556 986128
rect 397828 986076 397880 986128
rect 465724 986076 465776 986128
rect 495164 986076 495216 986128
rect 515404 986076 515456 986128
rect 543832 986076 543884 986128
rect 559564 986076 559616 986128
rect 89628 985940 89680 985992
rect 106924 985940 106976 985992
rect 215944 985940 215996 985992
rect 235632 985940 235684 985992
rect 279424 985940 279476 985992
rect 300492 985940 300544 985992
rect 369124 985940 369176 985992
rect 414112 985940 414164 985992
rect 415032 985940 415084 985992
rect 430304 985940 430356 985992
rect 436744 985940 436796 985992
rect 478972 985940 479024 985992
rect 514024 985940 514076 985992
rect 560116 985940 560168 985992
rect 570604 986076 570656 986128
rect 624976 986076 625028 986128
rect 669964 985940 670016 985992
rect 560944 985124 560996 985176
rect 671344 985124 671396 985176
rect 498108 984988 498160 985040
rect 667664 984988 667716 985040
rect 331864 984852 331916 984904
rect 664444 984852 664496 984904
rect 332048 984716 332100 984768
rect 665824 984716 665876 984768
rect 96528 984580 96580 984632
rect 651840 984580 651892 984632
rect 55864 975672 55916 975724
rect 62120 975672 62172 975724
rect 651656 975672 651708 975724
rect 661684 975672 661736 975724
rect 42524 969416 42576 969468
rect 55864 969416 55916 969468
rect 42248 966832 42300 966884
rect 42708 966832 42760 966884
rect 673276 966288 673328 966340
rect 675116 966288 675168 966340
rect 42432 964656 42484 964708
rect 42892 964656 42944 964708
rect 42432 963840 42484 963892
rect 44180 963840 44232 963892
rect 42432 963432 42484 963484
rect 43076 963432 43128 963484
rect 42432 961868 42484 961920
rect 44456 961868 44508 961920
rect 47584 961868 47636 961920
rect 62120 961868 62172 961920
rect 651656 961868 651708 961920
rect 663064 961868 663116 961920
rect 674288 961868 674340 961920
rect 675116 961868 675168 961920
rect 42432 959080 42484 959132
rect 43260 959080 43312 959132
rect 42432 958264 42484 958316
rect 44640 958264 44692 958316
rect 674104 957856 674156 957908
rect 675116 957856 675168 957908
rect 660304 957720 660356 957772
rect 675300 957312 675352 957364
rect 673092 956360 673144 956412
rect 675116 956360 675168 956412
rect 37924 952212 37976 952264
rect 41696 952212 41748 952264
rect 675852 949424 675904 949476
rect 678244 949424 678296 949476
rect 675944 948744 675996 948796
rect 682384 948744 682436 948796
rect 651656 948064 651708 948116
rect 671528 948064 671580 948116
rect 43536 945956 43588 946008
rect 62120 945956 62172 946008
rect 663064 941808 663116 941860
rect 675484 941808 675536 941860
rect 41236 941468 41288 941520
rect 41696 941468 41748 941520
rect 43444 941332 43496 941384
rect 48964 941332 49016 941384
rect 43628 941196 43680 941248
rect 50344 941196 50396 941248
rect 41236 940380 41288 940432
rect 41604 940380 41656 940432
rect 41236 939972 41288 940024
rect 41696 939972 41748 940024
rect 43444 939768 43496 939820
rect 51724 939768 51776 939820
rect 671528 938680 671580 938732
rect 675300 938680 675352 938732
rect 41236 938544 41288 938596
rect 41420 938544 41472 938596
rect 672724 938544 672776 938596
rect 675484 938544 675536 938596
rect 41052 938408 41104 938460
rect 41420 938408 41472 938460
rect 661684 938408 661736 938460
rect 675484 938408 675536 938460
rect 672724 937524 672776 937576
rect 675484 937524 675536 937576
rect 671344 937320 671396 937372
rect 675484 937320 675536 937372
rect 658924 937184 658976 937236
rect 675300 937184 675352 937236
rect 672540 937048 672592 937100
rect 674932 937048 674984 937100
rect 44640 936980 44692 937032
rect 62120 936980 62172 937032
rect 651656 936980 651708 937032
rect 660304 936980 660356 937032
rect 669964 935892 670016 935944
rect 675484 935892 675536 935944
rect 670976 935756 671028 935808
rect 675484 935756 675536 935808
rect 671804 935620 671856 935672
rect 675300 935620 675352 935672
rect 673276 933036 673328 933088
rect 675484 933036 675536 933088
rect 42984 932900 43036 932952
rect 54484 932900 54536 932952
rect 672908 932900 672960 932952
rect 675300 932900 675352 932952
rect 42800 931540 42852 931592
rect 53104 931540 53156 931592
rect 674104 931404 674156 931456
rect 675484 931404 675536 931456
rect 673092 930112 673144 930164
rect 675484 930112 675536 930164
rect 678244 930044 678296 930096
rect 683120 930044 683172 930096
rect 673276 928752 673328 928804
rect 675484 928752 675536 928804
rect 670608 927392 670660 927444
rect 675484 927392 675536 927444
rect 47584 923244 47636 923296
rect 62120 923244 62172 923296
rect 651656 921816 651708 921868
rect 663064 921816 663116 921868
rect 50344 909440 50396 909492
rect 62120 909440 62172 909492
rect 651656 909440 651708 909492
rect 671344 909440 671396 909492
rect 46204 896996 46256 897048
rect 62120 896996 62172 897048
rect 651656 895636 651708 895688
rect 664628 895636 664680 895688
rect 42432 884688 42484 884740
rect 62120 884688 62172 884740
rect 651656 881832 651708 881884
rect 671528 881832 671580 881884
rect 670424 879044 670476 879096
rect 675300 879044 675352 879096
rect 43444 870816 43496 870868
rect 62120 870816 62172 870868
rect 651656 869388 651708 869440
rect 658924 869388 658976 869440
rect 671528 868980 671580 869032
rect 675024 868980 675076 869032
rect 673828 868028 673880 868080
rect 675116 868028 675168 868080
rect 671160 866668 671212 866720
rect 675116 866668 675168 866720
rect 674840 865376 674892 865428
rect 670056 865240 670108 865292
rect 674840 865240 674892 865292
rect 675300 865036 675352 865088
rect 51908 858372 51960 858424
rect 62120 858372 62172 858424
rect 651656 855584 651708 855636
rect 659108 855584 659160 855636
rect 44824 844568 44876 844620
rect 62120 844568 62172 844620
rect 651656 841780 651708 841832
rect 661868 841780 661920 841832
rect 55864 832124 55916 832176
rect 62120 832124 62172 832176
rect 651656 829404 651708 829456
rect 660304 829404 660356 829456
rect 51724 818320 51776 818372
rect 62120 818320 62172 818372
rect 35808 817096 35860 817148
rect 40684 817096 40736 817148
rect 35624 816960 35676 817012
rect 40224 816960 40276 817012
rect 35808 816212 35860 816264
rect 39580 816212 39632 816264
rect 35624 815940 35676 815992
rect 41696 815940 41748 815992
rect 35808 815804 35860 815856
rect 41604 815804 41656 815856
rect 35440 815600 35492 815652
rect 41696 815600 41748 815652
rect 42064 815600 42116 815652
rect 50344 815600 50396 815652
rect 651656 815600 651708 815652
rect 661684 815600 661736 815652
rect 35808 814580 35860 814632
rect 39764 814512 39816 814564
rect 35808 814376 35860 814428
rect 41696 814376 41748 814428
rect 42064 814376 42116 814428
rect 42892 814376 42944 814428
rect 35624 814240 35676 814292
rect 41696 814240 41748 814292
rect 42064 814240 42116 814292
rect 44180 814240 44232 814292
rect 41052 812948 41104 813000
rect 41420 812948 41472 813000
rect 41328 811724 41380 811776
rect 41696 811724 41748 811776
rect 40776 810704 40828 810756
rect 41696 810704 41748 810756
rect 42064 810568 42116 810620
rect 42616 810568 42668 810620
rect 41328 807304 41380 807356
rect 41696 807304 41748 807356
rect 42064 807304 42116 807356
rect 48964 807304 49016 807356
rect 50344 805944 50396 805996
rect 62120 805944 62172 805996
rect 651656 803224 651708 803276
rect 663248 803224 663300 803276
rect 32404 802544 32456 802596
rect 41696 802544 41748 802596
rect 31668 802272 31720 802324
rect 39764 802272 39816 802324
rect 36544 801592 36596 801644
rect 40316 801592 40368 801644
rect 33784 801048 33836 801100
rect 40592 801048 40644 801100
rect 43628 799008 43680 799060
rect 47584 799008 47636 799060
rect 42524 798328 42576 798380
rect 42248 798124 42300 798176
rect 44640 796288 44692 796340
rect 42248 795608 42300 795660
rect 47768 793568 47820 793620
rect 62120 793568 62172 793620
rect 651656 789352 651708 789404
rect 660488 789352 660540 789404
rect 669780 789352 669832 789404
rect 674932 789352 674984 789404
rect 674932 788672 674984 788724
rect 675300 788196 675352 788248
rect 670792 787992 670844 788044
rect 675116 787992 675168 788044
rect 672172 786632 672224 786684
rect 675116 786632 675168 786684
rect 674472 783844 674524 783896
rect 675208 783844 675260 783896
rect 670240 783708 670292 783760
rect 675392 783708 675444 783760
rect 674012 782620 674064 782672
rect 675208 782620 675260 782672
rect 669044 782484 669096 782536
rect 675300 782484 675352 782536
rect 56232 780036 56284 780088
rect 62120 780036 62172 780088
rect 674288 779152 674340 779204
rect 675300 779152 675352 779204
rect 660304 778948 660356 779000
rect 675116 778948 675168 779000
rect 674104 778336 674156 778388
rect 675300 778336 675352 778388
rect 671528 776976 671580 777028
rect 675300 776976 675352 777028
rect 651656 775548 651708 775600
rect 663432 775548 663484 775600
rect 674932 775412 674984 775464
rect 675300 775412 675352 775464
rect 35808 774324 35860 774376
rect 40040 774324 40092 774376
rect 35532 773372 35584 773424
rect 40868 773372 40920 773424
rect 35808 773236 35860 773288
rect 35808 773100 35860 773152
rect 41696 773100 41748 773152
rect 42064 773100 42116 773152
rect 44456 773100 44508 773152
rect 41696 772964 41748 773016
rect 42064 772964 42116 773016
rect 55864 772964 55916 773016
rect 35348 772828 35400 772880
rect 51908 772828 51960 772880
rect 41696 772692 41748 772744
rect 42064 772692 42116 772744
rect 675852 772080 675904 772132
rect 683212 772080 683264 772132
rect 35900 772012 35952 772064
rect 39764 772012 39816 772064
rect 35532 771876 35584 771928
rect 39856 771876 39908 771928
rect 35716 771604 35768 771656
rect 35900 771536 35952 771588
rect 35348 771400 35400 771452
rect 39120 771400 39172 771452
rect 675852 771264 675904 771316
rect 681004 771264 681056 771316
rect 35808 770448 35860 770500
rect 41420 770448 41472 770500
rect 35624 770176 35676 770228
rect 41696 770244 41748 770296
rect 42064 770244 42116 770296
rect 43260 770244 43312 770296
rect 35440 770040 35492 770092
rect 41696 770040 41748 770092
rect 42064 770040 42116 770092
rect 44548 770040 44600 770092
rect 35808 768952 35860 769004
rect 39856 768952 39908 769004
rect 35532 768816 35584 768868
rect 39304 768816 39356 768868
rect 35348 768680 35400 768732
rect 40040 768680 40092 768732
rect 35808 767320 35860 767372
rect 36544 767320 36596 767372
rect 43628 767320 43680 767372
rect 62120 767320 62172 767372
rect 35808 766300 35860 766352
rect 40408 766164 40460 766216
rect 35808 765892 35860 765944
rect 41696 765960 41748 766012
rect 42064 765892 42116 765944
rect 45008 765892 45060 765944
rect 40040 765348 40092 765400
rect 41696 765348 41748 765400
rect 673644 765280 673696 765332
rect 674104 765280 674156 765332
rect 35808 764668 35860 764720
rect 40408 764668 40460 764720
rect 35808 763648 35860 763700
rect 37924 763648 37976 763700
rect 35624 763240 35676 763292
rect 41512 763240 41564 763292
rect 651656 763240 651708 763292
rect 660304 763172 660356 763224
rect 35808 761880 35860 761932
rect 40500 761880 40552 761932
rect 673828 761880 673880 761932
rect 673828 761744 673880 761796
rect 671344 761540 671396 761592
rect 675484 761540 675536 761592
rect 673644 761404 673696 761456
rect 674012 761404 674064 761456
rect 664628 760520 664680 760572
rect 675484 760520 675536 760572
rect 663064 760384 663116 760436
rect 675300 760384 675352 760436
rect 672540 760248 672592 760300
rect 675484 760248 675536 760300
rect 671988 759840 672040 759892
rect 675484 759840 675536 759892
rect 672724 759500 672776 759552
rect 675484 759500 675536 759552
rect 36544 759024 36596 759076
rect 41420 759024 41472 759076
rect 672632 759024 672684 759076
rect 675484 759024 675536 759076
rect 670976 758684 671028 758736
rect 675484 758684 675536 758736
rect 671804 758344 671856 758396
rect 675300 758344 675352 758396
rect 35164 758276 35216 758328
rect 40408 758276 40460 758328
rect 671804 758208 671856 758260
rect 675484 758208 675536 758260
rect 37924 757732 37976 757784
rect 41696 757732 41748 757784
rect 671344 757392 671396 757444
rect 675484 757392 675536 757444
rect 670056 755012 670108 755064
rect 675484 755012 675536 755064
rect 43812 754876 43864 754928
rect 45008 754876 45060 754928
rect 670424 754604 670476 754656
rect 675484 754604 675536 754656
rect 42432 754468 42484 754520
rect 45192 754468 45244 754520
rect 50528 753516 50580 753568
rect 62120 753516 62172 753568
rect 671160 753380 671212 753432
rect 675484 753380 675536 753432
rect 673828 752972 673880 753024
rect 675484 752972 675536 753024
rect 673000 752088 673052 752140
rect 673368 752088 673420 752140
rect 672356 751748 672408 751800
rect 675484 751748 675536 751800
rect 672356 751272 672408 751324
rect 675484 751272 675536 751324
rect 675852 751068 675904 751120
rect 683120 751068 683172 751120
rect 669964 750048 670016 750100
rect 675484 750048 675536 750100
rect 652024 749368 652076 749420
rect 659292 749368 659344 749420
rect 673736 748824 673788 748876
rect 674104 748824 674156 748876
rect 673920 748688 673972 748740
rect 42248 748552 42300 748604
rect 43260 748552 43312 748604
rect 674104 748348 674156 748400
rect 42248 747124 42300 747176
rect 42248 746852 42300 746904
rect 42248 745288 42300 745340
rect 669596 745220 669648 745272
rect 675300 745220 675352 745272
rect 42248 745084 42300 745136
rect 669228 743792 669280 743844
rect 669596 743792 669648 743844
rect 666100 742432 666152 742484
rect 675300 742432 675352 742484
rect 674840 741616 674892 741668
rect 675484 741616 675536 741668
rect 56048 741072 56100 741124
rect 62120 741072 62172 741124
rect 673000 738420 673052 738472
rect 675116 738420 675168 738472
rect 651656 735564 651708 735616
rect 664628 735564 664680 735616
rect 663432 734816 663484 734868
rect 675300 734748 675352 734800
rect 675024 734680 675076 734732
rect 675300 734544 675352 734596
rect 42432 731144 42484 731196
rect 56232 731144 56284 731196
rect 41144 730056 41196 730108
rect 41696 730056 41748 730108
rect 42064 730056 42116 730108
rect 50344 730056 50396 730108
rect 675208 728968 675260 729020
rect 675024 728764 675076 728816
rect 674380 728356 674432 728408
rect 675484 728356 675536 728408
rect 41052 727540 41104 727592
rect 41696 727608 41748 727660
rect 42064 727608 42116 727660
rect 42892 727608 42944 727660
rect 41328 727404 41380 727456
rect 41696 727472 41748 727524
rect 42064 727472 42116 727524
rect 44272 727472 44324 727524
rect 40868 727268 40920 727320
rect 41696 727268 41748 727320
rect 42064 727268 42116 727320
rect 44548 727268 44600 727320
rect 51908 727268 51960 727320
rect 62120 727268 62172 727320
rect 676036 726792 676088 726844
rect 683120 726792 683172 726844
rect 675852 726520 675904 726572
rect 683488 726520 683540 726572
rect 41328 726180 41380 726232
rect 41696 726180 41748 726232
rect 42064 726180 42116 726232
rect 42524 726180 42576 726232
rect 41144 726044 41196 726096
rect 41604 726044 41656 726096
rect 651656 723120 651708 723172
rect 659476 723120 659528 723172
rect 31760 720264 31812 720316
rect 40040 720264 40092 720316
rect 675852 719652 675904 719704
rect 683304 719652 683356 719704
rect 43444 719108 43496 719160
rect 55864 719108 55916 719160
rect 659108 716252 659160 716304
rect 675484 716252 675536 716304
rect 35164 715640 35216 715692
rect 39212 715640 39264 715692
rect 672632 715776 672684 715828
rect 672356 715572 672408 715624
rect 37924 715368 37976 715420
rect 41512 715368 41564 715420
rect 671988 715300 672040 715352
rect 674840 715300 674892 715352
rect 33784 715232 33836 715284
rect 41696 715232 41748 715284
rect 661868 715096 661920 715148
rect 675484 715096 675536 715148
rect 670976 714960 671028 715012
rect 50712 714824 50764 714876
rect 62120 714824 62172 714876
rect 658924 714824 658976 714876
rect 675300 714824 675352 714876
rect 675484 714824 675536 714876
rect 672356 714484 672408 714536
rect 675484 714484 675536 714536
rect 40684 714212 40736 714264
rect 41696 714212 41748 714264
rect 42064 714212 42116 714264
rect 42708 714212 42760 714264
rect 671160 714008 671212 714060
rect 675484 714008 675536 714060
rect 671804 713668 671856 713720
rect 675484 713668 675536 713720
rect 676036 713396 676088 713448
rect 677692 713396 677744 713448
rect 671896 713192 671948 713244
rect 675484 713192 675536 713244
rect 671528 712852 671580 712904
rect 675484 712852 675536 712904
rect 671712 712376 671764 712428
rect 675484 712376 675536 712428
rect 51724 712240 51776 712292
rect 672172 712036 672224 712088
rect 675484 712036 675536 712088
rect 670792 711220 670844 711272
rect 675484 711220 675536 711272
rect 42248 711084 42300 711136
rect 673092 709996 673144 710048
rect 675300 709996 675352 710048
rect 669044 709724 669096 709776
rect 675484 709724 675536 709776
rect 669780 709588 669832 709640
rect 675484 709588 675536 709640
rect 651656 709316 651708 709368
rect 663064 709316 663116 709368
rect 670240 708772 670292 708824
rect 675484 708772 675536 708824
rect 671528 708364 671580 708416
rect 675484 708364 675536 708416
rect 674104 707548 674156 707600
rect 675484 707548 675536 707600
rect 42248 706528 42300 706580
rect 43260 706528 43312 706580
rect 672264 706256 672316 706308
rect 675484 706256 675536 706308
rect 675852 705304 675904 705356
rect 683120 705304 683172 705356
rect 670148 705032 670200 705084
rect 675484 705032 675536 705084
rect 42248 704216 42300 704268
rect 42248 704012 42300 704064
rect 42156 702856 42208 702908
rect 42708 702856 42760 702908
rect 51724 701020 51776 701072
rect 62120 701020 62172 701072
rect 42064 700544 42116 700596
rect 42616 700544 42668 700596
rect 672080 698436 672132 698488
rect 675208 698436 675260 698488
rect 673092 697076 673144 697128
rect 675116 697076 675168 697128
rect 651656 696940 651708 696992
rect 661868 696940 661920 696992
rect 674288 694764 674340 694816
rect 675116 694764 675168 694816
rect 674472 694152 674524 694204
rect 675392 694152 675444 694204
rect 666284 692792 666336 692844
rect 675116 692792 675168 692844
rect 659476 689256 659528 689308
rect 674932 689256 674984 689308
rect 674104 689120 674156 689172
rect 675116 689120 675168 689172
rect 43812 688644 43864 688696
rect 62120 688644 62172 688696
rect 42524 687692 42576 687744
rect 50528 687692 50580 687744
rect 43444 687352 43496 687404
rect 51908 687352 51960 687404
rect 40960 687216 41012 687268
rect 41696 687216 41748 687268
rect 42064 687216 42116 687268
rect 56048 687216 56100 687268
rect 672632 687216 672684 687268
rect 675116 687216 675168 687268
rect 41696 686060 41748 686112
rect 42064 686060 42116 686112
rect 45192 686060 45244 686112
rect 41328 685992 41380 686044
rect 41144 685856 41196 685908
rect 41696 685856 41748 685908
rect 42064 685856 42116 685908
rect 45008 685856 45060 685908
rect 669780 685856 669832 685908
rect 674840 685856 674892 685908
rect 40868 684768 40920 684820
rect 41144 684632 41196 684684
rect 41696 684700 41748 684752
rect 42064 684700 42116 684752
rect 43076 684700 43128 684752
rect 41696 684496 41748 684548
rect 42064 684496 42116 684548
rect 44456 684496 44508 684548
rect 41328 683544 41380 683596
rect 41696 683544 41748 683596
rect 42064 683476 42116 683528
rect 42524 683476 42576 683528
rect 42064 683340 42116 683392
rect 42800 683340 42852 683392
rect 40776 683272 40828 683324
rect 41696 683272 41748 683324
rect 41144 683136 41196 683188
rect 41696 683136 41748 683188
rect 42064 683136 42116 683188
rect 42892 683136 42944 683188
rect 651656 683136 651708 683188
rect 658924 683136 658976 683188
rect 41328 682456 41380 682508
rect 675852 682388 675904 682440
rect 683212 682388 683264 682440
rect 41328 682252 41380 682304
rect 676036 682252 676088 682304
rect 683396 682252 683448 682304
rect 42064 676336 42116 676388
rect 50344 676336 50396 676388
rect 42064 675588 42116 675640
rect 42708 675588 42760 675640
rect 34428 675452 34480 675504
rect 39764 675452 39816 675504
rect 47768 674840 47820 674892
rect 62120 674840 62172 674892
rect 31024 672664 31076 672716
rect 40408 672664 40460 672716
rect 36544 672052 36596 672104
rect 41696 672052 41748 672104
rect 663248 670828 663300 670880
rect 675484 671100 675536 671152
rect 661684 670692 661736 670744
rect 675484 670692 675536 670744
rect 674012 670352 674064 670404
rect 675484 670352 675536 670404
rect 670976 669740 671028 669792
rect 675484 669740 675536 669792
rect 671160 669604 671212 669656
rect 675484 669604 675536 669656
rect 660488 669468 660540 669520
rect 674012 669468 674064 669520
rect 651656 669332 651708 669384
rect 662052 669332 662104 669384
rect 671160 669332 671212 669384
rect 674840 669332 674892 669384
rect 671804 668516 671856 668568
rect 675484 668516 675536 668568
rect 671528 667700 671580 667752
rect 675484 667700 675536 667752
rect 671620 667564 671672 667616
rect 674012 667564 674064 667616
rect 670976 667224 671028 667276
rect 675484 667224 675536 667276
rect 42248 667088 42300 667140
rect 43444 667088 43496 667140
rect 43444 666544 43496 666596
rect 45192 666544 45244 666596
rect 669596 666068 669648 666120
rect 675484 666068 675536 666120
rect 666100 665184 666152 665236
rect 675484 665184 675536 665236
rect 42248 664844 42300 664896
rect 43444 664844 43496 664896
rect 672908 664028 672960 664080
rect 674840 664028 674892 664080
rect 669228 663892 669280 663944
rect 675484 663892 675536 663944
rect 668584 663756 668636 663808
rect 675484 663756 675536 663808
rect 42248 663484 42300 663536
rect 42708 663484 42760 663536
rect 673828 663212 673880 663264
rect 675484 663212 675536 663264
rect 42248 662804 42300 662856
rect 43260 662804 43312 662856
rect 670424 662804 670476 662856
rect 675484 662804 675536 662856
rect 43444 662396 43496 662448
rect 62120 662396 62172 662448
rect 671344 661580 671396 661632
rect 675484 661580 675536 661632
rect 671344 661104 671396 661156
rect 675484 661104 675536 661156
rect 670332 659880 670384 659932
rect 675484 659880 675536 659932
rect 675852 659812 675904 659864
rect 683120 659812 683172 659864
rect 42156 657364 42208 657416
rect 42616 657364 42668 657416
rect 651656 656888 651708 656940
rect 661684 656888 661736 656940
rect 665456 654236 665508 654288
rect 675392 654236 675444 654288
rect 672908 651380 672960 651432
rect 675392 651380 675444 651432
rect 669228 650020 669280 650072
rect 674840 650020 674892 650072
rect 671712 649068 671764 649120
rect 675392 649068 675444 649120
rect 674840 648592 674892 648644
rect 675392 648592 675444 648644
rect 51908 647844 51960 647896
rect 62120 647844 62172 647896
rect 665272 647708 665324 647760
rect 670792 647708 670844 647760
rect 35808 644716 35860 644768
rect 38844 644716 38896 644768
rect 35532 644444 35584 644496
rect 41236 644444 41288 644496
rect 662052 643696 662104 643748
rect 670792 643628 670844 643680
rect 35808 643492 35860 643544
rect 40316 643492 40368 643544
rect 35532 643220 35584 643272
rect 41696 643288 41748 643340
rect 42064 643288 42116 643340
rect 44272 643288 44324 643340
rect 35348 643084 35400 643136
rect 41696 643084 41748 643136
rect 42064 643084 42116 643136
rect 51724 643084 51776 643136
rect 651656 643084 651708 643136
rect 664812 643084 664864 643136
rect 35808 642132 35860 642184
rect 39028 642200 39080 642252
rect 35440 641860 35492 641912
rect 39672 641928 39724 641980
rect 670792 641860 670844 641912
rect 675300 641860 675352 641912
rect 35624 641724 35676 641776
rect 39764 641724 39816 641776
rect 666100 641724 666152 641776
rect 670792 641724 670844 641776
rect 42064 640908 42116 640960
rect 42892 640908 42944 640960
rect 35808 640704 35860 640756
rect 39856 640704 39908 640756
rect 35532 640432 35584 640484
rect 41696 640432 41748 640484
rect 35348 640296 35400 640348
rect 41696 640296 41748 640348
rect 42064 640296 42116 640348
rect 43168 640296 43220 640348
rect 670792 640024 670844 640076
rect 675300 640024 675352 640076
rect 35808 639072 35860 639124
rect 40224 639072 40276 639124
rect 673460 639004 673512 639056
rect 675300 639004 675352 639056
rect 35532 638936 35584 638988
rect 40040 638936 40092 638988
rect 34428 638188 34480 638240
rect 41696 638188 41748 638240
rect 42064 638120 42116 638172
rect 42708 638120 42760 638172
rect 35532 637916 35584 637968
rect 41696 637916 41748 637968
rect 42064 637848 42116 637900
rect 43628 637848 43680 637900
rect 35808 637712 35860 637764
rect 41512 637712 41564 637764
rect 675852 637440 675904 637492
rect 679624 637440 679676 637492
rect 674380 636896 674432 636948
rect 675484 636828 675536 636880
rect 35808 636352 35860 636404
rect 41328 636352 41380 636404
rect 49148 636216 49200 636268
rect 62120 636216 62172 636268
rect 675852 636148 675904 636200
rect 682384 636148 682436 636200
rect 35808 635060 35860 635112
rect 39764 635060 39816 635112
rect 35624 634788 35676 634840
rect 39304 634788 39356 634840
rect 35808 633632 35860 633684
rect 41696 633632 41748 633684
rect 42064 633632 42116 633684
rect 51724 633632 51776 633684
rect 35624 633428 35676 633480
rect 41696 633428 41748 633480
rect 42064 633428 42116 633480
rect 50528 633428 50580 633480
rect 33784 630028 33836 630080
rect 41696 630028 41748 630080
rect 42064 629960 42116 630012
rect 42708 629960 42760 630012
rect 32404 629892 32456 629944
rect 41696 629892 41748 629944
rect 652024 629280 652076 629332
rect 659108 629280 659160 629332
rect 50712 626628 50764 626680
rect 42616 626492 42668 626544
rect 659292 625404 659344 625456
rect 675300 625404 675352 625456
rect 664628 625268 664680 625320
rect 675484 625268 675536 625320
rect 660304 625132 660356 625184
rect 675116 625132 675168 625184
rect 671528 624248 671580 624300
rect 675484 624248 675536 624300
rect 671160 624044 671212 624096
rect 675300 624044 675352 624096
rect 671160 623908 671212 623960
rect 675484 623908 675536 623960
rect 43812 623772 43864 623824
rect 47768 623772 47820 623824
rect 62120 623772 62172 623824
rect 670792 623772 670844 623824
rect 675116 623772 675168 623824
rect 42340 623364 42392 623416
rect 671620 622820 671672 622872
rect 675484 622820 675536 622872
rect 671712 622548 671764 622600
rect 675300 622548 675352 622600
rect 45192 622412 45244 622464
rect 670976 622412 671028 622464
rect 675484 622412 675536 622464
rect 42432 622004 42484 622056
rect 671896 621188 671948 621240
rect 675484 621188 675536 621240
rect 671896 620984 671948 621036
rect 675300 620984 675352 621036
rect 669780 619828 669832 619880
rect 675300 619828 675352 619880
rect 666284 619624 666336 619676
rect 675484 619624 675536 619676
rect 673092 619420 673144 619472
rect 675484 619420 675536 619472
rect 42616 618876 42668 618928
rect 43628 618876 43680 618928
rect 672632 618196 672684 618248
rect 675484 618196 675536 618248
rect 651656 616836 651708 616888
rect 660488 616836 660540 616888
rect 671528 616632 671580 616684
rect 671896 616632 671948 616684
rect 671712 616496 671764 616548
rect 671712 616360 671764 616412
rect 670976 616088 671028 616140
rect 675300 616088 675352 616140
rect 668768 615748 668820 615800
rect 675484 615748 675536 615800
rect 42248 615680 42300 615732
rect 675852 615612 675904 615664
rect 683120 615612 683172 615664
rect 42248 615476 42300 615528
rect 663708 614116 663760 614168
rect 675484 614116 675536 614168
rect 42156 613572 42208 613624
rect 44456 613572 44508 613624
rect 668584 610104 668636 610156
rect 671344 610104 671396 610156
rect 666376 609968 666428 610020
rect 675116 609968 675168 610020
rect 43628 609220 43680 609272
rect 62120 609220 62172 609272
rect 673092 607588 673144 607640
rect 675300 607588 675352 607640
rect 672540 605820 672592 605872
rect 675116 605820 675168 605872
rect 674656 603304 674708 603356
rect 675392 603304 675444 603356
rect 652024 603100 652076 603152
rect 660304 603100 660356 603152
rect 665640 603100 665692 603152
rect 675300 603032 675352 603084
rect 35808 601672 35860 601724
rect 41696 601672 41748 601724
rect 42064 601672 42116 601724
rect 49148 601672 49200 601724
rect 674012 601332 674064 601384
rect 674656 601332 674708 601384
rect 42616 600380 42668 600432
rect 51908 600312 51960 600364
rect 660488 599564 660540 599616
rect 674288 599496 674340 599548
rect 675116 599496 675168 599548
rect 675116 599360 675168 599412
rect 41328 598952 41380 599004
rect 41696 598952 41748 599004
rect 42064 598952 42116 599004
rect 44456 598952 44508 599004
rect 668860 598748 668912 598800
rect 675300 598680 675352 598732
rect 41328 597796 41380 597848
rect 41696 597796 41748 597848
rect 42064 597796 42116 597848
rect 42800 597796 42852 597848
rect 41052 597660 41104 597712
rect 41696 597660 41748 597712
rect 42064 597660 42116 597712
rect 42984 597660 43036 597712
rect 40868 597524 40920 597576
rect 41696 597524 41748 597576
rect 42064 597524 42116 597576
rect 43076 597524 43128 597576
rect 49148 597524 49200 597576
rect 62120 597524 62172 597576
rect 674564 597456 674616 597508
rect 675300 597456 675352 597508
rect 41328 596436 41380 596488
rect 41696 596436 41748 596488
rect 41144 596028 41196 596080
rect 41604 596028 41656 596080
rect 41328 594736 41380 594788
rect 41696 594736 41748 594788
rect 40592 593036 40644 593088
rect 41604 593036 41656 593088
rect 40776 592696 40828 592748
rect 41604 592696 41656 592748
rect 673920 591540 673972 591592
rect 675484 591540 675536 591592
rect 675852 591404 675904 591456
rect 683212 591404 683264 591456
rect 675852 591268 675904 591320
rect 683396 591268 683448 591320
rect 43812 590656 43864 590708
rect 56048 590656 56100 590708
rect 651656 590656 651708 590708
rect 663248 590656 663300 590708
rect 33048 586984 33100 587036
rect 40132 586984 40184 587036
rect 35164 585896 35216 585948
rect 41604 585896 41656 585948
rect 31024 585692 31076 585744
rect 41604 585692 41656 585744
rect 39948 585352 40000 585404
rect 41420 585352 41472 585404
rect 36544 585148 36596 585200
rect 39396 585148 39448 585200
rect 42064 584400 42116 584452
rect 42708 584400 42760 584452
rect 51908 583720 51960 583772
rect 62120 583720 62172 583772
rect 661868 581000 661920 581052
rect 675484 581000 675536 581052
rect 42432 580592 42484 580644
rect 44640 580592 44692 580644
rect 670792 579980 670844 580032
rect 674748 579980 674800 580032
rect 663064 579776 663116 579828
rect 675300 579776 675352 579828
rect 658924 579640 658976 579692
rect 675484 579640 675536 579692
rect 671160 579368 671212 579420
rect 675484 579368 675536 579420
rect 671344 579028 671396 579080
rect 675484 579028 675536 579080
rect 42248 578688 42300 578740
rect 672724 578552 672776 578604
rect 675484 578552 675536 578604
rect 42248 578416 42300 578468
rect 672908 578212 672960 578264
rect 675484 578212 675536 578264
rect 671620 578008 671672 578060
rect 675300 578008 675352 578060
rect 671528 577736 671580 577788
rect 675300 577736 675352 577788
rect 673736 577532 673788 577584
rect 674104 577532 674156 577584
rect 671344 577396 671396 577448
rect 675300 577396 675352 577448
rect 671344 576920 671396 576972
rect 675300 576920 675352 576972
rect 651656 576852 651708 576904
rect 664628 576852 664680 576904
rect 665456 574200 665508 574252
rect 675484 574268 675536 574320
rect 665272 574064 665324 574116
rect 675300 574064 675352 574116
rect 671804 573724 671856 573776
rect 675484 573724 675536 573776
rect 669596 572908 669648 572960
rect 675484 572908 675536 572960
rect 674104 572500 674156 572552
rect 675484 572500 675536 572552
rect 43444 571344 43496 571396
rect 62120 571344 62172 571396
rect 669228 571344 669280 571396
rect 675484 571344 675536 571396
rect 42064 570936 42116 570988
rect 42616 570936 42668 570988
rect 671712 570800 671764 570852
rect 675484 570800 675536 570852
rect 666100 570120 666152 570172
rect 675484 570120 675536 570172
rect 675852 570052 675904 570104
rect 683120 570052 683172 570104
rect 670792 569576 670844 569628
rect 675484 569576 675536 569628
rect 671344 565224 671396 565276
rect 671160 565020 671212 565072
rect 671160 564884 671212 564936
rect 671344 564748 671396 564800
rect 665088 564408 665140 564460
rect 675300 564408 675352 564460
rect 651656 563048 651708 563100
rect 658924 563048 658976 563100
rect 673736 561688 673788 561740
rect 675116 561688 675168 561740
rect 666192 560328 666244 560380
rect 675300 560328 675352 560380
rect 41696 557744 41748 557796
rect 42064 557744 42116 557796
rect 49148 557744 49200 557796
rect 41328 557676 41380 557728
rect 674104 557676 674156 557728
rect 675116 557676 675168 557728
rect 43812 557540 43864 557592
rect 51908 557540 51960 557592
rect 54852 557540 54904 557592
rect 62120 557540 62172 557592
rect 666100 557540 666152 557592
rect 675300 557540 675352 557592
rect 42064 555364 42116 555416
rect 43168 555364 43220 555416
rect 41144 555296 41196 555348
rect 41696 555092 41748 555144
rect 41052 554888 41104 554940
rect 41696 554888 41748 554940
rect 42064 554888 42116 554940
rect 42984 554888 43036 554940
rect 40592 554752 40644 554804
rect 41696 554752 41748 554804
rect 42064 554752 42116 554804
rect 44272 554752 44324 554804
rect 669780 554752 669832 554804
rect 675300 554752 675352 554804
rect 674472 554276 674524 554328
rect 675116 554276 675168 554328
rect 658924 554004 658976 554056
rect 675116 554004 675168 554056
rect 671896 553460 671948 553512
rect 675300 553460 675352 553512
rect 651656 550604 651708 550656
rect 659292 550604 659344 550656
rect 664260 550604 664312 550656
rect 675024 550604 675076 550656
rect 40040 550400 40092 550452
rect 41696 550400 41748 550452
rect 42064 550400 42116 550452
rect 42524 550400 42576 550452
rect 45560 548632 45612 548684
rect 45560 548496 45612 548548
rect 42340 547884 42392 547936
rect 53288 547884 53340 547936
rect 31760 547408 31812 547460
rect 38568 547408 38620 547460
rect 675944 547272 675996 547324
rect 678244 547272 678296 547324
rect 676128 547136 676180 547188
rect 683396 547136 683448 547188
rect 43444 546592 43496 546644
rect 49148 546592 49200 546644
rect 675944 545708 675996 545760
rect 683212 545708 683264 545760
rect 43444 545096 43496 545148
rect 62120 545096 62172 545148
rect 29644 544348 29696 544400
rect 41512 544348 41564 544400
rect 38568 542308 38620 542360
rect 41696 542308 41748 542360
rect 652024 536800 652076 536852
rect 660488 536800 660540 536852
rect 42248 536256 42300 536308
rect 45376 536256 45428 536308
rect 664812 535644 664864 535696
rect 675484 535644 675536 535696
rect 661684 535440 661736 535492
rect 675484 535440 675536 535492
rect 672632 534556 672684 534608
rect 674748 534556 674800 534608
rect 675484 534556 675536 534608
rect 671344 534352 671396 534404
rect 659108 534216 659160 534268
rect 674564 534216 674616 534268
rect 42432 534148 42484 534200
rect 45744 534148 45796 534200
rect 672632 534080 672684 534132
rect 675484 534080 675536 534132
rect 42616 533944 42668 533996
rect 43996 533944 44048 533996
rect 671528 532856 671580 532908
rect 675484 532856 675536 532908
rect 673552 531768 673604 531820
rect 675484 531768 675536 531820
rect 672448 531564 672500 531616
rect 675484 531564 675536 531616
rect 671160 531428 671212 531480
rect 673552 531428 673604 531480
rect 42248 530884 42300 530936
rect 42616 530884 42668 530936
rect 42616 530748 42668 530800
rect 45192 531292 45244 531344
rect 672540 531292 672592 531344
rect 674748 531292 674800 531344
rect 42248 530272 42300 530324
rect 42616 530272 42668 530324
rect 673092 530068 673144 530120
rect 675484 530068 675536 530120
rect 665640 529932 665692 529984
rect 675484 529932 675536 529984
rect 669044 529320 669096 529372
rect 675484 529320 675536 529372
rect 42432 529048 42484 529100
rect 43812 529048 43864 529100
rect 666468 528572 666520 528624
rect 675484 528572 675536 528624
rect 673920 528300 673972 528352
rect 675484 528300 675536 528352
rect 674104 528096 674156 528148
rect 674104 527892 674156 527944
rect 673920 527620 673972 527672
rect 675484 527620 675536 527672
rect 668860 525784 668912 525836
rect 675484 525784 675536 525836
rect 678244 525716 678296 525768
rect 683120 525716 683172 525768
rect 671252 524424 671304 524476
rect 675484 524424 675536 524476
rect 42524 523676 42576 523728
rect 62764 523676 62816 523728
rect 651656 522996 651708 523048
rect 661684 522996 661736 523048
rect 42064 518916 42116 518968
rect 62120 518916 62172 518968
rect 651656 510620 651708 510672
rect 659108 510620 659160 510672
rect 52276 506472 52328 506524
rect 62120 506472 62172 506524
rect 676128 503480 676180 503532
rect 679624 503480 679676 503532
rect 651656 496816 651708 496868
rect 661868 496816 661920 496868
rect 43628 491920 43680 491972
rect 62120 491920 62172 491972
rect 664628 491580 664680 491632
rect 675484 491580 675536 491632
rect 663248 491444 663300 491496
rect 674748 491444 674800 491496
rect 660304 491308 660356 491360
rect 675116 491308 675168 491360
rect 672724 490016 672776 490068
rect 675484 490016 675536 490068
rect 672540 487296 672592 487348
rect 675484 487296 675536 487348
rect 666100 485936 666152 485988
rect 675484 485936 675536 485988
rect 665088 485800 665140 485852
rect 675300 485800 675352 485852
rect 673736 485460 673788 485512
rect 674748 485460 674800 485512
rect 664260 484508 664312 484560
rect 675484 484508 675536 484560
rect 651656 484440 651708 484492
rect 664996 484372 665048 484424
rect 669780 483964 669832 484016
rect 675300 483964 675352 484016
rect 672908 483556 672960 483608
rect 675300 483556 675352 483608
rect 666284 483080 666336 483132
rect 675484 483080 675536 483132
rect 671896 482332 671948 482384
rect 675484 482332 675536 482384
rect 673736 481856 673788 481908
rect 675484 481856 675536 481908
rect 671436 480632 671488 480684
rect 675484 480632 675536 480684
rect 47952 480224 48004 480276
rect 62120 480224 62172 480276
rect 668768 474036 668820 474088
rect 671712 474036 671764 474088
rect 651656 470568 651708 470620
rect 663248 470568 663300 470620
rect 49332 466420 49384 466472
rect 62120 466420 62172 466472
rect 651656 456764 651708 456816
rect 663432 456764 663484 456816
rect 46572 446360 46624 446412
rect 62764 446360 62816 446412
rect 651656 444456 651708 444508
rect 660672 444388 660724 444440
rect 43812 433984 43864 434036
rect 62120 433984 62172 434036
rect 652024 430584 652076 430636
rect 658924 430584 658976 430636
rect 41328 429564 41380 429616
rect 41696 429564 41748 429616
rect 41144 429428 41196 429480
rect 41696 429428 41748 429480
rect 42064 429428 42116 429480
rect 43444 429428 43496 429480
rect 41328 429292 41380 429344
rect 41696 429292 41748 429344
rect 42064 429292 42116 429344
rect 43996 429292 44048 429344
rect 40960 429156 41012 429208
rect 41696 429156 41748 429208
rect 42064 429156 42116 429208
rect 44548 429156 44600 429208
rect 56232 427796 56284 427848
rect 62120 427796 62172 427848
rect 41144 426436 41196 426488
rect 41696 426436 41748 426488
rect 42064 426436 42116 426488
rect 44548 426436 44600 426488
rect 45192 419500 45244 419552
rect 51908 419500 51960 419552
rect 42616 418140 42668 418192
rect 54668 418140 54720 418192
rect 651656 416780 651708 416832
rect 660304 416780 660356 416832
rect 45192 415420 45244 415472
rect 62120 415420 62172 415472
rect 42248 409776 42300 409828
rect 43168 409776 43220 409828
rect 42432 408416 42484 408468
rect 54852 408416 54904 408468
rect 42432 408280 42484 408332
rect 44364 408280 44416 408332
rect 42432 407056 42484 407108
rect 45376 407056 45428 407108
rect 651656 404336 651708 404388
rect 664812 404336 664864 404388
rect 42432 404132 42484 404184
rect 45560 404132 45612 404184
rect 667204 403384 667256 403436
rect 675300 403384 675352 403436
rect 659292 403248 659344 403300
rect 660488 403112 660540 403164
rect 667204 403112 667256 403164
rect 675484 403180 675536 403232
rect 661684 402976 661736 403028
rect 675484 402976 675536 403028
rect 42432 402500 42484 402552
rect 43352 402500 43404 402552
rect 50712 401616 50764 401668
rect 62120 401616 62172 401668
rect 673920 401344 673972 401396
rect 675484 401344 675536 401396
rect 672724 400528 672776 400580
rect 675484 400528 675536 400580
rect 673092 399712 673144 399764
rect 675484 399712 675536 399764
rect 42432 397400 42484 397452
rect 46940 397400 46992 397452
rect 671804 396312 671856 396364
rect 675484 396312 675536 396364
rect 672540 396040 672592 396092
rect 675300 396040 675352 396092
rect 673460 394272 673512 394324
rect 675484 394272 675536 394324
rect 672908 393320 672960 393372
rect 675484 393320 675536 393372
rect 671620 391960 671672 392012
rect 675484 391960 675536 392012
rect 651656 390532 651708 390584
rect 663064 390532 663116 390584
rect 48136 389240 48188 389292
rect 62120 389240 62172 389292
rect 35808 387472 35860 387524
rect 39948 387472 40000 387524
rect 35808 386792 35860 386844
rect 40132 386792 40184 386844
rect 35348 386520 35400 386572
rect 40316 386520 40368 386572
rect 42064 386452 42116 386504
rect 49332 386452 49384 386504
rect 35532 386384 35584 386436
rect 41696 386384 41748 386436
rect 35808 385432 35860 385484
rect 39580 385432 39632 385484
rect 35532 385160 35584 385212
rect 41696 385228 41748 385280
rect 42064 385228 42116 385280
rect 42892 385228 42944 385280
rect 35348 385024 35400 385076
rect 41696 385024 41748 385076
rect 42064 385024 42116 385076
rect 43260 385024 43312 385076
rect 35808 384072 35860 384124
rect 39672 384072 39724 384124
rect 42064 383868 42116 383920
rect 44548 383868 44600 383920
rect 35624 383800 35676 383852
rect 41696 383800 41748 383852
rect 35808 383664 35860 383716
rect 41696 383664 41748 383716
rect 42064 383664 42116 383716
rect 44180 383664 44232 383716
rect 35532 382644 35584 382696
rect 40040 382644 40092 382696
rect 35808 382508 35860 382560
rect 41696 382508 41748 382560
rect 35808 382372 35860 382424
rect 40224 382372 40276 382424
rect 671804 382304 671856 382356
rect 675392 382304 675444 382356
rect 35348 382236 35400 382288
rect 41420 382236 41472 382288
rect 674288 382168 674340 382220
rect 675116 382168 675168 382220
rect 35624 381012 35676 381064
rect 40040 381012 40092 381064
rect 35808 380876 35860 380928
rect 39856 380876 39908 380928
rect 35624 379924 35676 379976
rect 41052 379924 41104 379976
rect 35808 379652 35860 379704
rect 39764 379652 39816 379704
rect 35440 379516 35492 379568
rect 41512 379516 41564 379568
rect 35808 378292 35860 378344
rect 39580 378292 39632 378344
rect 651656 378156 651708 378208
rect 661684 378156 661736 378208
rect 673368 377816 673420 377868
rect 675300 377816 675352 377868
rect 35624 377000 35676 377052
rect 41512 376932 41564 376984
rect 42064 376796 42116 376848
rect 35808 376728 35860 376780
rect 41696 376728 41748 376780
rect 53472 376728 53524 376780
rect 672908 376456 672960 376508
rect 675116 376456 675168 376508
rect 28816 375844 28868 375896
rect 33784 375844 33836 375896
rect 35808 375572 35860 375624
rect 41696 375572 41748 375624
rect 42064 375504 42116 375556
rect 52092 375504 52144 375556
rect 49332 375368 49384 375420
rect 62120 375368 62172 375420
rect 674472 375300 674524 375352
rect 675116 375300 675168 375352
rect 33784 373260 33836 373312
rect 41696 373260 41748 373312
rect 32404 371832 32456 371884
rect 41696 371832 41748 371884
rect 42064 371696 42116 371748
rect 42616 371696 42668 371748
rect 651656 364352 651708 364404
rect 664628 364352 664680 364404
rect 42248 364284 42300 364336
rect 52276 364284 52328 364336
rect 42340 364080 42392 364132
rect 43628 364080 43680 364132
rect 42432 360136 42484 360188
rect 44548 360136 44600 360188
rect 42156 359932 42208 359984
rect 43444 359932 43496 359984
rect 664996 357688 665048 357740
rect 675484 357688 675536 357740
rect 661868 357552 661920 357604
rect 675300 357552 675352 357604
rect 659108 357416 659160 357468
rect 675116 357416 675168 357468
rect 673920 357280 673972 357332
rect 674748 357280 674800 357332
rect 673920 357008 673972 357060
rect 675484 357008 675536 357060
rect 42432 355988 42484 356040
rect 45376 355988 45428 356040
rect 672724 355172 672776 355224
rect 675484 355172 675536 355224
rect 673092 354832 673144 354884
rect 675484 354832 675536 354884
rect 673092 354696 673144 354748
rect 675300 354696 675352 354748
rect 673368 353540 673420 353592
rect 675484 353540 675536 353592
rect 672816 353404 672868 353456
rect 675116 353404 675168 353456
rect 669780 353268 669832 353320
rect 675300 353268 675352 353320
rect 671896 351908 671948 351960
rect 675484 351908 675536 351960
rect 669596 350684 669648 350736
rect 675484 350684 675536 350736
rect 651656 350548 651708 350600
rect 661868 350548 661920 350600
rect 671804 350548 671856 350600
rect 675300 350548 675352 350600
rect 673552 349256 673604 349308
rect 675484 349256 675536 349308
rect 672632 348848 672684 348900
rect 675484 348848 675536 348900
rect 45376 347012 45428 347064
rect 62948 347012 63000 347064
rect 675852 346400 675904 346452
rect 683120 346400 683172 346452
rect 671712 344972 671764 345024
rect 675484 344972 675536 345024
rect 35808 344020 35860 344072
rect 39580 344020 39632 344072
rect 35624 343748 35676 343800
rect 40408 343816 40460 343868
rect 35348 343612 35400 343664
rect 41696 343612 41748 343664
rect 42064 343612 42116 343664
rect 56232 343612 56284 343664
rect 35808 342660 35860 342712
rect 39948 342660 40000 342712
rect 35348 342388 35400 342440
rect 39580 342456 39632 342508
rect 35532 342252 35584 342304
rect 40316 342252 40368 342304
rect 35808 341436 35860 341488
rect 39764 341436 39816 341488
rect 35624 341164 35676 341216
rect 40316 341232 40368 341284
rect 35624 341028 35676 341080
rect 41696 341028 41748 341080
rect 42064 341028 42116 341080
rect 45192 341028 45244 341080
rect 35808 340892 35860 340944
rect 41696 340892 41748 340944
rect 42064 340892 42116 340944
rect 44180 340892 44232 340944
rect 673368 340688 673420 340740
rect 675116 340688 675168 340740
rect 35624 339600 35676 339652
rect 39580 339600 39632 339652
rect 35808 338308 35860 338360
rect 41512 338308 41564 338360
rect 35624 338104 35676 338156
rect 41696 338104 41748 338156
rect 42064 338104 42116 338156
rect 47216 338104 47268 338156
rect 651656 338104 651708 338156
rect 667112 338104 667164 338156
rect 673276 337968 673328 338020
rect 675116 337968 675168 338020
rect 35808 337152 35860 337204
rect 40040 337152 40092 337204
rect 35532 336880 35584 336932
rect 41696 336948 41748 337000
rect 42064 336948 42116 337000
rect 43076 336948 43128 337000
rect 35808 336744 35860 336796
rect 41696 336744 41748 336796
rect 42064 336744 42116 336796
rect 43812 336744 43864 336796
rect 46756 336744 46808 336796
rect 62120 336744 62172 336796
rect 674472 336676 674524 336728
rect 675116 336676 675168 336728
rect 35624 335588 35676 335640
rect 40316 335588 40368 335640
rect 669596 335588 669648 335640
rect 674472 335588 674524 335640
rect 673552 335452 673604 335504
rect 675116 335452 675168 335504
rect 35808 335316 35860 335368
rect 39672 335316 39724 335368
rect 674472 335112 674524 335164
rect 674840 335112 674892 335164
rect 35808 334364 35860 334416
rect 40316 334364 40368 334416
rect 35440 334092 35492 334144
rect 39580 334092 39632 334144
rect 42064 334092 42116 334144
rect 35624 333956 35676 334008
rect 41696 333956 41748 334008
rect 54852 333956 54904 334008
rect 671896 333888 671948 333940
rect 675300 333888 675352 333940
rect 35624 332732 35676 332784
rect 39580 332732 39632 332784
rect 35808 332596 35860 332648
rect 41696 332596 41748 332648
rect 42064 332596 42116 332648
rect 56232 332596 56284 332648
rect 672632 332392 672684 332444
rect 675116 332392 675168 332444
rect 42432 327020 42484 327072
rect 43444 327020 43496 327072
rect 42432 325592 42484 325644
rect 45560 325592 45612 325644
rect 669780 325592 669832 325644
rect 674932 325592 674984 325644
rect 669228 325456 669280 325508
rect 675116 325456 675168 325508
rect 651656 324300 651708 324352
rect 673552 324300 673604 324352
rect 42432 324232 42484 324284
rect 46572 324232 46624 324284
rect 49516 322940 49568 322992
rect 62120 322940 62172 322992
rect 42432 321512 42484 321564
rect 43628 321512 43680 321564
rect 42248 321240 42300 321292
rect 44456 321240 44508 321292
rect 42432 320084 42484 320136
rect 44640 320084 44692 320136
rect 42432 318792 42484 318844
rect 47032 318792 47084 318844
rect 43628 318044 43680 318096
rect 62764 318044 62816 318096
rect 42432 317364 42484 317416
rect 43812 317364 43864 317416
rect 42248 317228 42300 317280
rect 43996 317228 44048 317280
rect 42432 315868 42484 315920
rect 43076 315868 43128 315920
rect 666376 313556 666428 313608
rect 663248 313420 663300 313472
rect 663432 313284 663484 313336
rect 666376 313284 666428 313336
rect 675484 313420 675536 313472
rect 675484 313284 675536 313336
rect 673920 312468 673972 312520
rect 675484 312468 675536 312520
rect 660672 311992 660724 312044
rect 675300 311992 675352 312044
rect 666192 311856 666244 311908
rect 675484 311856 675536 311908
rect 673092 310836 673144 310888
rect 675300 310836 675352 310888
rect 43444 310496 43496 310548
rect 62120 310496 62172 310548
rect 666376 310496 666428 310548
rect 675484 310496 675536 310548
rect 42432 310360 42484 310412
rect 47216 310360 47268 310412
rect 672816 310020 672868 310072
rect 675484 310020 675536 310072
rect 664260 309340 664312 309392
rect 675484 309340 675536 309392
rect 665088 309136 665140 309188
rect 675300 309136 675352 309188
rect 673092 305464 673144 305516
rect 675484 305464 675536 305516
rect 673368 303832 673420 303884
rect 675484 303832 675536 303884
rect 672540 303424 672592 303476
rect 675484 303424 675536 303476
rect 680360 302200 680412 302252
rect 683120 302200 683172 302252
rect 43812 301180 43864 301232
rect 49332 301180 49384 301232
rect 669780 300772 669832 300824
rect 675484 300772 675536 300824
rect 674794 298460 674846 298512
rect 675024 298460 675076 298512
rect 40960 298256 41012 298308
rect 41144 298256 41196 298308
rect 41696 298324 41748 298376
rect 42064 298324 42116 298376
rect 42892 298324 42944 298376
rect 42064 298188 42116 298240
rect 45192 298188 45244 298240
rect 41696 298120 41748 298172
rect 47952 298120 48004 298172
rect 62120 298120 62172 298172
rect 672356 297712 672408 297764
rect 672724 297712 672776 297764
rect 675852 297168 675904 297220
rect 681004 297168 681056 297220
rect 40960 296692 41012 296744
rect 41696 296692 41748 296744
rect 42064 296692 42116 296744
rect 45192 296692 45244 296744
rect 675484 296216 675536 296268
rect 675484 295876 675536 295928
rect 40500 292544 40552 292596
rect 41604 292544 41656 292596
rect 674472 292272 674524 292324
rect 675116 292272 675168 292324
rect 42892 289960 42944 290012
rect 64144 289960 64196 290012
rect 41144 289824 41196 289876
rect 41696 289824 41748 289876
rect 42064 289824 42116 289876
rect 61384 289824 61436 289876
rect 672356 289824 672408 289876
rect 672724 289824 672776 289876
rect 40960 289076 41012 289128
rect 41696 289076 41748 289128
rect 35164 284928 35216 284980
rect 41696 284928 41748 284980
rect 651656 284316 651708 284368
rect 662052 284316 662104 284368
rect 42248 280100 42300 280152
rect 43996 280100 44048 280152
rect 406936 278672 406988 278724
rect 499580 278672 499632 278724
rect 42432 278536 42484 278588
rect 50712 278536 50764 278588
rect 467564 278536 467616 278588
rect 476488 278536 476540 278588
rect 482284 278536 482336 278588
rect 590568 278536 590620 278588
rect 42432 278400 42484 278452
rect 44364 278400 44416 278452
rect 64144 278400 64196 278452
rect 661040 278400 661092 278452
rect 61384 278264 61436 278316
rect 659660 278264 659712 278316
rect 53288 278128 53340 278180
rect 654140 278128 654192 278180
rect 56232 277992 56284 278044
rect 658280 277992 658332 278044
rect 437204 277788 437256 277840
rect 546684 277788 546736 277840
rect 421932 277652 421984 277704
rect 524328 277652 524380 277704
rect 413652 277516 413704 277568
rect 510344 277516 510396 277568
rect 466092 277312 466144 277364
rect 471244 277312 471296 277364
rect 471428 277312 471480 277364
rect 475936 277380 475988 277432
rect 476488 277380 476540 277432
rect 596640 277380 596692 277432
rect 442540 277176 442592 277228
rect 557632 277176 557684 277228
rect 409328 277040 409380 277092
rect 475568 277040 475620 277092
rect 476396 277040 476448 277092
rect 502340 277040 502392 277092
rect 502524 277040 502576 277092
rect 509056 277040 509108 277092
rect 509240 277040 509292 277092
rect 512000 277040 512052 277092
rect 512184 277040 512236 277092
rect 571984 277040 572036 277092
rect 380716 276904 380768 276956
rect 457168 276904 457220 276956
rect 471244 276904 471296 276956
rect 475752 276904 475804 276956
rect 476672 276904 476724 276956
rect 587164 277040 587216 277092
rect 581644 276904 581696 276956
rect 606116 276904 606168 276956
rect 387340 276768 387392 276820
rect 467840 276768 467892 276820
rect 469036 276768 469088 276820
rect 471428 276768 471480 276820
rect 472900 276768 472952 276820
rect 475752 276768 475804 276820
rect 475936 276768 475988 276820
rect 599032 276768 599084 276820
rect 43812 276632 43864 276684
rect 509056 276632 509108 276684
rect 509240 276632 509292 276684
rect 659844 276632 659896 276684
rect 446312 276496 446364 276548
rect 451280 276496 451332 276548
rect 456984 276496 457036 276548
rect 570696 276496 570748 276548
rect 571984 276496 572036 276548
rect 581644 276496 581696 276548
rect 420368 276360 420420 276412
rect 521016 276360 521068 276412
rect 446956 276224 447008 276276
rect 531228 276224 531280 276276
rect 402796 276088 402848 276140
rect 485734 276088 485786 276140
rect 485872 276088 485924 276140
rect 499396 276088 499448 276140
rect 499534 276088 499586 276140
rect 110788 275952 110840 276004
rect 156420 275952 156472 276004
rect 171048 275952 171100 276004
rect 175648 275952 175700 276004
rect 175832 275952 175884 276004
rect 177396 275952 177448 276004
rect 344008 275952 344060 276004
rect 354312 275952 354364 276004
rect 356980 275952 357032 276004
rect 388628 275952 388680 276004
rect 388996 275952 389048 276004
rect 418160 275952 418212 276004
rect 418344 275952 418396 276004
rect 427636 275952 427688 276004
rect 217140 275884 217192 275936
rect 218520 275884 218572 275936
rect 103704 275816 103756 275868
rect 160652 275816 160704 275868
rect 174636 275816 174688 275868
rect 197544 275816 197596 275868
rect 316776 275816 316828 275868
rect 327080 275816 327132 275868
rect 331220 275816 331272 275868
rect 340144 275816 340196 275868
rect 343824 275816 343876 275868
rect 370872 275816 370924 275868
rect 371056 275816 371108 275868
rect 407488 275816 407540 275868
rect 410064 275816 410116 275868
rect 421656 275816 421708 275868
rect 426072 275816 426124 275868
rect 436744 275952 436796 276004
rect 436928 275952 436980 276004
rect 471244 275952 471296 276004
rect 471428 275952 471480 276004
rect 473728 275952 473780 276004
rect 473912 275952 473964 276004
rect 477224 275952 477276 276004
rect 477408 275952 477460 276004
rect 485228 275952 485280 276004
rect 428004 275816 428056 275868
rect 465540 275816 465592 275868
rect 465724 275816 465776 275868
rect 470876 275816 470928 275868
rect 471060 275816 471112 275868
rect 480812 275816 480864 275868
rect 480996 275816 481048 275868
rect 484308 275816 484360 275868
rect 484492 275816 484544 275868
rect 487896 275952 487948 276004
rect 490564 275952 490616 276004
rect 498568 275952 498620 276004
rect 498752 275952 498804 276004
rect 501788 275952 501840 276004
rect 501972 275952 502024 276004
rect 511540 275952 511592 276004
rect 561036 275952 561088 276004
rect 565912 275952 565964 276004
rect 635648 275952 635700 276004
rect 485872 275816 485924 275868
rect 612004 275816 612056 275868
rect 96620 275680 96672 275732
rect 153844 275680 153896 275732
rect 160468 275680 160520 275732
rect 174452 275680 174504 275732
rect 181720 275680 181772 275732
rect 207020 275680 207072 275732
rect 298008 275680 298060 275732
rect 85948 275544 86000 275596
rect 149060 275544 149112 275596
rect 153292 275544 153344 275596
rect 185768 275544 185820 275596
rect 199476 275544 199528 275596
rect 210976 275544 211028 275596
rect 218336 275544 218388 275596
rect 68192 275408 68244 275460
rect 135260 275408 135312 275460
rect 156880 275408 156932 275460
rect 166172 275408 166224 275460
rect 167552 275408 167604 275460
rect 200028 275408 200080 275460
rect 207756 275408 207808 275460
rect 216680 275408 216732 275460
rect 221924 275544 221976 275596
rect 228456 275544 228508 275596
rect 282920 275544 282972 275596
rect 285772 275544 285824 275596
rect 299020 275544 299072 275596
rect 302332 275544 302384 275596
rect 305092 275680 305144 275732
rect 316500 275680 316552 275732
rect 317328 275680 317380 275732
rect 329472 275680 329524 275732
rect 311716 275544 311768 275596
rect 313280 275544 313332 275596
rect 325976 275544 326028 275596
rect 329196 275544 329248 275596
rect 374368 275680 374420 275732
rect 380900 275680 380952 275732
rect 411076 275680 411128 275732
rect 414204 275680 414256 275732
rect 508688 275680 508740 275732
rect 511356 275680 511408 275732
rect 633348 275680 633400 275732
rect 333612 275544 333664 275596
rect 381544 275544 381596 275596
rect 394608 275544 394660 275596
rect 470508 275544 470560 275596
rect 471244 275544 471296 275596
rect 222844 275408 222896 275460
rect 236092 275408 236144 275460
rect 242256 275408 242308 275460
rect 285864 275408 285916 275460
rect 303436 275408 303488 275460
rect 70584 275272 70636 275324
rect 139768 275272 139820 275324
rect 149796 275272 149848 275324
rect 184756 275272 184808 275324
rect 188804 275272 188856 275324
rect 107200 275136 107252 275188
rect 151176 275136 151228 275188
rect 152188 275136 152240 275188
rect 162584 275136 162636 275188
rect 227812 275272 227864 275324
rect 237380 275272 237432 275324
rect 238484 275272 238536 275324
rect 243728 275272 243780 275324
rect 265900 275272 265952 275324
rect 271512 275272 271564 275324
rect 278412 275272 278464 275324
rect 292856 275272 292908 275324
rect 302240 275272 302292 275324
rect 318800 275408 318852 275460
rect 320088 275408 320140 275460
rect 336556 275408 336608 275460
rect 340236 275408 340288 275460
rect 392124 275408 392176 275460
rect 392308 275408 392360 275460
rect 396908 275408 396960 275460
rect 397092 275408 397144 275460
rect 471060 275408 471112 275460
rect 471244 275408 471296 275460
rect 484860 275408 484912 275460
rect 485228 275544 485280 275596
rect 490564 275544 490616 275596
rect 490748 275544 490800 275596
rect 494980 275544 495032 275596
rect 495164 275544 495216 275596
rect 604920 275544 604972 275596
rect 499396 275408 499448 275460
rect 211252 275204 211304 275256
rect 212448 275204 212500 275256
rect 245568 275136 245620 275188
rect 246304 275136 246356 275188
rect 301504 275136 301556 275188
rect 322388 275272 322440 275324
rect 322572 275272 322624 275324
rect 333060 275272 333112 275324
rect 342260 275272 342312 275324
rect 350724 275272 350776 275324
rect 350908 275272 350960 275324
rect 399208 275272 399260 275324
rect 399852 275272 399904 275324
rect 484492 275272 484544 275324
rect 336464 275136 336516 275188
rect 343640 275136 343692 275188
rect 350540 275136 350592 275188
rect 357900 275136 357952 275188
rect 365628 275136 365680 275188
rect 375564 275136 375616 275188
rect 376024 275136 376076 275188
rect 403992 275136 404044 275188
rect 404268 275136 404320 275188
rect 425244 275136 425296 275188
rect 425428 275136 425480 275188
rect 428004 275136 428056 275188
rect 430580 275136 430632 275188
rect 436560 275136 436612 275188
rect 436744 275136 436796 275188
rect 465724 275136 465776 275188
rect 465908 275136 465960 275188
rect 466414 275136 466466 275188
rect 466552 275136 466604 275188
rect 487344 275272 487396 275324
rect 487528 275272 487580 275324
rect 491484 275272 491536 275324
rect 491668 275272 491720 275324
rect 498752 275272 498804 275324
rect 498936 275272 498988 275324
rect 616788 275408 616840 275460
rect 499672 275272 499724 275324
rect 640432 275272 640484 275324
rect 485228 275136 485280 275188
rect 213920 275068 213972 275120
rect 81256 274932 81308 274984
rect 86224 274932 86276 274984
rect 116676 274864 116728 274916
rect 135628 274864 135680 274916
rect 142712 275000 142764 275052
rect 169760 275000 169812 275052
rect 249064 275000 249116 275052
rect 250352 275000 250404 275052
rect 347044 275000 347096 275052
rect 350908 275000 350960 275052
rect 375288 275000 375340 275052
rect 178132 274932 178184 274984
rect 180064 274932 180116 274984
rect 214840 274932 214892 274984
rect 221464 274932 221516 274984
rect 365260 274932 365312 274984
rect 369676 274932 369728 274984
rect 140320 274728 140372 274780
rect 140780 274728 140832 274780
rect 142988 274864 143040 274916
rect 150992 274864 151044 274916
rect 152648 274864 152700 274916
rect 374552 274864 374604 274916
rect 379152 274864 379204 274916
rect 382372 275000 382424 275052
rect 408684 275000 408736 275052
rect 408868 275000 408920 275052
rect 412456 275000 412508 275052
rect 414020 275000 414072 275052
rect 415768 275000 415820 275052
rect 422116 275000 422168 275052
rect 523408 275000 523460 275052
rect 523868 275136 523920 275188
rect 537576 275136 537628 275188
rect 537760 275136 537812 275188
rect 552940 275136 552992 275188
rect 556160 275136 556212 275188
rect 561220 275136 561272 275188
rect 530492 275000 530544 275052
rect 393320 274864 393372 274916
rect 397368 274864 397420 274916
rect 414572 274864 414624 274916
rect 418068 274864 418120 274916
rect 516232 274864 516284 274916
rect 186412 274796 186464 274848
rect 188436 274796 188488 274848
rect 358728 274796 358780 274848
rect 364984 274796 365036 274848
rect 156604 274728 156656 274780
rect 378784 274728 378836 274780
rect 386236 274728 386288 274780
rect 408500 274728 408552 274780
rect 412272 274728 412324 274780
rect 412456 274728 412508 274780
rect 491668 274728 491720 274780
rect 491852 274728 491904 274780
rect 494152 274728 494204 274780
rect 494336 274728 494388 274780
rect 499396 274728 499448 274780
rect 500132 274728 500184 274780
rect 523868 274864 523920 274916
rect 523684 274728 523736 274780
rect 549352 275000 549404 275052
rect 563060 275000 563112 275052
rect 577780 275000 577832 275052
rect 531228 274864 531280 274916
rect 563520 274864 563572 274916
rect 552664 274728 552716 274780
rect 556436 274728 556488 274780
rect 619456 274728 619508 274780
rect 623872 274728 623924 274780
rect 89536 274660 89588 274712
rect 92480 274660 92532 274712
rect 161572 274660 161624 274712
rect 163688 274660 163740 274712
rect 163964 274660 164016 274712
rect 167828 274660 167880 274712
rect 185216 274660 185268 274712
rect 186964 274660 187016 274712
rect 241980 274660 242032 274712
rect 246028 274660 246080 274712
rect 246764 274660 246816 274712
rect 248880 274660 248932 274712
rect 271144 274660 271196 274712
rect 276296 274660 276348 274712
rect 276664 274660 276716 274712
rect 278688 274660 278740 274712
rect 280712 274660 280764 274712
rect 283380 274660 283432 274712
rect 293224 274660 293276 274712
rect 294052 274660 294104 274712
rect 295524 274660 295576 274712
rect 298744 274660 298796 274712
rect 339224 274660 339276 274712
rect 344836 274660 344888 274712
rect 355692 274660 355744 274712
rect 356704 274660 356756 274712
rect 643744 274660 643796 274712
rect 645124 274660 645176 274712
rect 93032 274456 93084 274508
rect 119344 274592 119396 274644
rect 120264 274592 120316 274644
rect 161434 274592 161486 274644
rect 359464 274592 359516 274644
rect 400404 274592 400456 274644
rect 401324 274592 401376 274644
rect 489828 274592 489880 274644
rect 490012 274592 490064 274644
rect 495256 274592 495308 274644
rect 495394 274592 495446 274644
rect 497004 274592 497056 274644
rect 497188 274592 497240 274644
rect 621480 274592 621532 274644
rect 119068 274456 119120 274508
rect 168472 274456 168524 274508
rect 169760 274456 169812 274508
rect 184940 274456 184992 274508
rect 306196 274456 306248 274508
rect 320088 274456 320140 274508
rect 329656 274456 329708 274508
rect 365628 274456 365680 274508
rect 366364 274456 366416 274508
rect 111984 274320 112036 274372
rect 164240 274320 164292 274372
rect 177396 274320 177448 274372
rect 204260 274320 204312 274372
rect 299204 274320 299256 274372
rect 313280 274320 313332 274372
rect 322756 274320 322808 274372
rect 358728 274320 358780 274372
rect 358912 274320 358964 274372
rect 368020 274320 368072 274372
rect 102508 274184 102560 274236
rect 159088 274184 159140 274236
rect 166356 274184 166408 274236
rect 198924 274184 198976 274236
rect 200580 274184 200632 274236
rect 213184 274184 213236 274236
rect 274364 274184 274416 274236
rect 286876 274184 286928 274236
rect 290464 274184 290516 274236
rect 305828 274184 305880 274236
rect 310060 274184 310112 274236
rect 336464 274184 336516 274236
rect 234896 274116 234948 274168
rect 239496 274116 239548 274168
rect 77668 274048 77720 274100
rect 143632 274048 143684 274100
rect 158076 274048 158128 274100
rect 193220 274048 193272 274100
rect 198280 274048 198332 274100
rect 217968 274048 218020 274100
rect 283932 274048 283984 274100
rect 299020 274048 299072 274100
rect 307576 274048 307628 274100
rect 331220 274048 331272 274100
rect 336556 274048 336608 274100
rect 378784 274184 378836 274236
rect 353944 274048 353996 274100
rect 382648 274048 382700 274100
rect 390284 274456 390336 274508
rect 466414 274456 466466 274508
rect 466552 274456 466604 274508
rect 471060 274456 471112 274508
rect 471244 274456 471296 274508
rect 479616 274456 479668 274508
rect 480352 274456 480404 274508
rect 610808 274456 610860 274508
rect 393228 274320 393280 274372
rect 476212 274320 476264 274372
rect 478604 274320 478656 274372
rect 614396 274320 614448 274372
rect 394332 274184 394384 274236
rect 471244 274184 471296 274236
rect 471428 274184 471480 274236
rect 484860 274184 484912 274236
rect 485228 274184 485280 274236
rect 395712 274048 395764 274100
rect 397184 274048 397236 274100
rect 483204 274048 483256 274100
rect 486424 274184 486476 274236
rect 617984 274184 618036 274236
rect 625068 274048 625120 274100
rect 72976 273912 73028 273964
rect 140964 273912 141016 273964
rect 141792 273912 141844 273964
rect 183744 273912 183796 273964
rect 184480 273912 184532 273964
rect 206284 273912 206336 273964
rect 206560 273912 206612 273964
rect 223856 273912 223908 273964
rect 224224 273912 224276 273964
rect 234896 273912 234948 273964
rect 279884 273912 279936 273964
rect 295156 273912 295208 273964
rect 130844 273776 130896 273828
rect 176752 273776 176804 273828
rect 294604 273776 294656 273828
rect 314108 273912 314160 273964
rect 314476 273912 314528 273964
rect 342260 273912 342312 273964
rect 351184 273912 351236 273964
rect 359464 273912 359516 273964
rect 368020 273912 368072 273964
rect 389732 273912 389784 273964
rect 391848 273912 391900 273964
rect 394608 273912 394660 273964
rect 396724 273912 396776 273964
rect 435180 273912 435232 273964
rect 435364 273912 435416 273964
rect 451234 273912 451286 273964
rect 451372 273912 451424 273964
rect 561036 273912 561088 273964
rect 632704 273912 632756 273964
rect 643928 273912 643980 273964
rect 318708 273776 318760 273828
rect 350540 273776 350592 273828
rect 354220 273776 354272 273828
rect 397368 273776 397420 273828
rect 398748 273776 398800 273828
rect 484308 273776 484360 273828
rect 484860 273776 484912 273828
rect 488724 273776 488776 273828
rect 628564 273776 628616 273828
rect 124956 273640 125008 273692
rect 157984 273640 158036 273692
rect 161480 273640 161532 273692
rect 169944 273640 169996 273692
rect 361212 273640 361264 273692
rect 404268 273640 404320 273692
rect 405556 273640 405608 273692
rect 486884 273640 486936 273692
rect 543464 273640 543516 273692
rect 332508 273504 332560 273556
rect 374552 273504 374604 273556
rect 378784 273504 378836 273556
rect 420552 273504 420604 273556
rect 426256 273504 426308 273556
rect 529296 273504 529348 273556
rect 343548 273368 343600 273420
rect 392308 273368 392360 273420
rect 416136 273368 416188 273420
rect 515128 273368 515180 273420
rect 395436 273300 395488 273352
rect 396908 273300 396960 273352
rect 358176 273232 358228 273284
rect 358728 273232 358780 273284
rect 451096 273232 451148 273284
rect 451234 273232 451286 273284
rect 451372 273232 451424 273284
rect 460756 273232 460808 273284
rect 42432 273164 42484 273216
rect 43076 273164 43128 273216
rect 127348 273164 127400 273216
rect 174268 273164 174320 273216
rect 326896 273164 326948 273216
rect 343824 273164 343876 273216
rect 364340 273164 364392 273216
rect 430764 273164 430816 273216
rect 430948 273164 431000 273216
rect 121368 273028 121420 273080
rect 171600 273028 171652 273080
rect 174452 273028 174504 273080
rect 196164 273028 196216 273080
rect 295156 273028 295208 273080
rect 302240 273028 302292 273080
rect 317144 273028 317196 273080
rect 344008 273028 344060 273080
rect 357992 273028 358044 273080
rect 361396 273028 361448 273080
rect 368848 273028 368900 273080
rect 436928 273028 436980 273080
rect 437434 273164 437486 273216
rect 445484 273164 445536 273216
rect 441620 273028 441672 273080
rect 442080 273028 442132 273080
rect 447692 273164 447744 273216
rect 460940 273164 460992 273216
rect 568304 273164 568356 273216
rect 446128 273028 446180 273080
rect 555240 273028 555292 273080
rect 572168 273028 572220 273080
rect 608508 273028 608560 273080
rect 71780 272892 71832 272944
rect 109684 272892 109736 272944
rect 109960 272892 110012 272944
rect 163320 272892 163372 272944
rect 180800 272892 180852 272944
rect 207480 272892 207532 272944
rect 302884 272892 302936 272944
rect 317696 272892 317748 272944
rect 325516 272892 325568 272944
rect 368480 272892 368532 272944
rect 381360 272892 381412 272944
rect 384488 272892 384540 272944
rect 387800 272892 387852 272944
rect 97724 272756 97776 272808
rect 155408 272756 155460 272808
rect 168656 272756 168708 272808
rect 198740 272756 198792 272808
rect 91836 272620 91888 272672
rect 152372 272620 152424 272672
rect 159272 272620 159324 272672
rect 194784 272620 194836 272672
rect 195704 272620 195756 272672
rect 210608 272756 210660 272808
rect 300676 272756 300728 272808
rect 317328 272756 317380 272808
rect 321468 272756 321520 272808
rect 357992 272756 358044 272808
rect 359464 272756 359516 272808
rect 365260 272756 365312 272808
rect 376576 272756 376628 272808
rect 446312 272756 446364 272808
rect 447416 272892 447468 272944
rect 451096 272892 451148 272944
rect 451924 272892 451976 272944
rect 456616 272892 456668 272944
rect 452108 272756 452160 272808
rect 453856 272756 453908 272808
rect 575388 272892 575440 272944
rect 457444 272756 457496 272808
rect 571800 272756 571852 272808
rect 578884 272756 578936 272808
rect 636844 272756 636896 272808
rect 210056 272620 210108 272672
rect 226432 272620 226484 272672
rect 289084 272620 289136 272672
rect 299940 272620 299992 272672
rect 300124 272620 300176 272672
rect 319628 272620 319680 272672
rect 333244 272620 333296 272672
rect 377956 272620 378008 272672
rect 378140 272620 378192 272672
rect 239680 272552 239732 272604
rect 244556 272552 244608 272604
rect 74080 272484 74132 272536
rect 142160 272484 142212 272536
rect 154488 272484 154540 272536
rect 190736 272484 190788 272536
rect 197084 272484 197136 272536
rect 137928 272348 137980 272400
rect 181168 272348 181220 272400
rect 218520 272484 218572 272536
rect 230572 272484 230624 272536
rect 231400 272484 231452 272536
rect 239312 272484 239364 272536
rect 271696 272484 271748 272536
rect 280988 272484 281040 272536
rect 282184 272484 282236 272536
rect 297548 272484 297600 272536
rect 303436 272484 303488 272536
rect 322572 272484 322624 272536
rect 326712 272484 326764 272536
rect 218244 272348 218296 272400
rect 280988 272348 281040 272400
rect 289268 272348 289320 272400
rect 345664 272484 345716 272536
rect 372068 272484 372120 272536
rect 374460 272484 374512 272536
rect 380900 272484 380952 272536
rect 384488 272620 384540 272672
rect 458364 272620 458416 272672
rect 460480 272620 460532 272672
rect 466276 272620 466328 272672
rect 466460 272620 466512 272672
rect 582472 272620 582524 272672
rect 442080 272484 442132 272536
rect 359464 272348 359516 272400
rect 361856 272348 361908 272400
rect 417240 272348 417292 272400
rect 447416 272484 447468 272536
rect 455880 272484 455932 272536
rect 456064 272484 456116 272536
rect 113180 272212 113232 272264
rect 142804 272212 142856 272264
rect 142988 272212 143040 272264
rect 167460 272212 167512 272264
rect 348424 272212 348476 272264
rect 374644 272212 374696 272264
rect 374828 272212 374880 272264
rect 378140 272212 378192 272264
rect 379152 272212 379204 272264
rect 442724 272348 442776 272400
rect 446772 272348 446824 272400
rect 454224 272348 454276 272400
rect 454408 272348 454460 272400
rect 564716 272348 564768 272400
rect 571984 272484 572036 272536
rect 585600 272484 585652 272536
rect 585784 272484 585836 272536
rect 622676 272484 622728 272536
rect 578516 272348 578568 272400
rect 340696 272076 340748 272128
rect 375288 272076 375340 272128
rect 376760 272076 376812 272128
rect 409880 272076 409932 272128
rect 412272 272076 412324 272128
rect 485734 272212 485786 272264
rect 485872 272212 485924 272264
rect 571984 272212 572036 272264
rect 417700 272076 417752 272128
rect 418344 272076 418396 272128
rect 351736 271940 351788 271992
rect 374460 271940 374512 271992
rect 374644 271940 374696 271992
rect 385040 271940 385092 271992
rect 410708 271940 410760 271992
rect 427774 272076 427826 272128
rect 427912 272076 427964 272128
rect 442724 272076 442776 272128
rect 443368 272076 443420 272128
rect 446128 272076 446180 272128
rect 451280 272076 451332 272128
rect 556160 272076 556212 272128
rect 423496 271940 423548 271992
rect 427084 271940 427136 271992
rect 427268 271940 427320 271992
rect 532792 271940 532844 271992
rect 101312 271804 101364 271856
rect 157616 271804 157668 271856
rect 165160 271804 165212 271856
rect 197360 271804 197412 271856
rect 297364 271804 297416 271856
rect 309416 271804 309468 271856
rect 312544 271804 312596 271856
rect 338580 271804 338632 271856
rect 338948 271804 339000 271856
rect 363788 271804 363840 271856
rect 263416 271736 263468 271788
rect 269212 271736 269264 271788
rect 88616 271668 88668 271720
rect 145564 271668 145616 271720
rect 179328 271668 179380 271720
rect 204904 271668 204956 271720
rect 296628 271668 296680 271720
rect 301504 271668 301556 271720
rect 304908 271668 304960 271720
rect 334164 271668 334216 271720
rect 338028 271668 338080 271720
rect 356980 271668 357032 271720
rect 363696 271668 363748 271720
rect 98920 271532 98972 271584
rect 156236 271532 156288 271584
rect 170128 271532 170180 271584
rect 201040 271532 201092 271584
rect 213644 271532 213696 271584
rect 228272 271532 228324 271584
rect 229008 271532 229060 271584
rect 237840 271532 237892 271584
rect 289636 271532 289688 271584
rect 298008 271532 298060 271584
rect 309048 271532 309100 271584
rect 342444 271532 342496 271584
rect 345848 271532 345900 271584
rect 362592 271532 362644 271584
rect 92480 271396 92532 271448
rect 150440 271396 150492 271448
rect 156604 271396 156656 271448
rect 180800 271396 180852 271448
rect 201776 271396 201828 271448
rect 221004 271396 221056 271448
rect 233700 271396 233752 271448
rect 240784 271396 240836 271448
rect 268844 271396 268896 271448
rect 277492 271396 277544 271448
rect 285588 271396 285640 271448
rect 304632 271396 304684 271448
rect 311716 271396 311768 271448
rect 347228 271396 347280 271448
rect 361488 271396 361540 271448
rect 422760 271668 422812 271720
rect 365536 271532 365588 271584
rect 428188 271668 428240 271720
rect 428556 271804 428608 271856
rect 440608 271804 440660 271856
rect 440976 271804 441028 271856
rect 444564 271804 444616 271856
rect 444748 271804 444800 271856
rect 551744 271804 551796 271856
rect 551928 271804 551980 271856
rect 553860 271804 553912 271856
rect 429200 271668 429252 271720
rect 429384 271668 429436 271720
rect 433340 271668 433392 271720
rect 433524 271668 433576 271720
rect 535184 271668 535236 271720
rect 543004 271668 543056 271720
rect 423128 271532 423180 271584
rect 432604 271532 432656 271584
rect 432788 271532 432840 271584
rect 442264 271532 442316 271584
rect 442724 271532 442776 271584
rect 551928 271532 551980 271584
rect 554044 271668 554096 271720
rect 615592 271668 615644 271720
rect 562324 271532 562376 271584
rect 383200 271396 383252 271448
rect 456800 271396 456852 271448
rect 457444 271396 457496 271448
rect 84752 271260 84804 271312
rect 147680 271260 147732 271312
rect 155684 271260 155736 271312
rect 192392 271260 192444 271312
rect 193496 271260 193548 271312
rect 215760 271260 215812 271312
rect 223120 271260 223172 271312
rect 234160 271260 234212 271312
rect 273076 271260 273128 271312
rect 284576 271260 284628 271312
rect 291844 271260 291896 271312
rect 310520 271260 310572 271312
rect 315948 271260 316000 271312
rect 353116 271260 353168 271312
rect 65892 271124 65944 271176
rect 136640 271124 136692 271176
rect 139124 271124 139176 271176
rect 140044 271124 140096 271176
rect 145012 271124 145064 271176
rect 185584 271124 185636 271176
rect 192208 271124 192260 271176
rect 215300 271124 215352 271176
rect 215944 271124 215996 271176
rect 229744 271124 229796 271176
rect 277308 271124 277360 271176
rect 291660 271124 291712 271176
rect 292396 271124 292448 271176
rect 315304 271124 315356 271176
rect 322204 271124 322256 271176
rect 360200 271260 360252 271312
rect 369952 271260 370004 271312
rect 428556 271260 428608 271312
rect 432604 271260 432656 271312
rect 440976 271260 441028 271312
rect 442264 271260 442316 271312
rect 461860 271396 461912 271448
rect 465172 271396 465224 271448
rect 465632 271396 465684 271448
rect 466414 271396 466466 271448
rect 466552 271396 466604 271448
rect 580080 271396 580132 271448
rect 114284 270988 114336 271040
rect 164884 270988 164936 271040
rect 185768 270988 185820 271040
rect 192208 270988 192260 271040
rect 319444 270988 319496 271040
rect 346032 270988 346084 271040
rect 350448 270988 350500 271040
rect 382372 271124 382424 271176
rect 389824 271124 389876 271176
rect 456800 271124 456852 271176
rect 456984 271124 457036 271176
rect 461400 271124 461452 271176
rect 562140 271260 562192 271312
rect 562324 271260 562376 271312
rect 594340 271260 594392 271312
rect 485734 271124 485786 271176
rect 485872 271124 485924 271176
rect 495440 271124 495492 271176
rect 495624 271124 495676 271176
rect 360108 270988 360160 271040
rect 422484 270988 422536 271040
rect 123760 270852 123812 270904
rect 172704 270852 172756 270904
rect 334624 270852 334676 270904
rect 349620 270852 349672 270904
rect 357164 270852 357216 270904
rect 412594 270852 412646 270904
rect 412732 270852 412784 270904
rect 414020 270852 414072 270904
rect 414664 270852 414716 270904
rect 417240 270852 417292 270904
rect 432788 270988 432840 271040
rect 432972 270988 433024 271040
rect 495624 270988 495676 271040
rect 496544 271124 496596 271176
rect 639236 271124 639288 271176
rect 538404 270988 538456 271040
rect 538864 270988 538916 271040
rect 597836 270988 597888 271040
rect 134432 270716 134484 270768
rect 178960 270716 179012 270768
rect 342536 270716 342588 270768
rect 348148 270716 348200 270768
rect 354496 270716 354548 270768
rect 412088 270716 412140 270768
rect 412456 270716 412508 270768
rect 423312 270852 423364 270904
rect 426440 270852 426492 270904
rect 418252 270716 418304 270768
rect 423128 270716 423180 270768
rect 423312 270716 423364 270768
rect 495072 270852 495124 270904
rect 495808 270852 495860 270904
rect 513840 270852 513892 270904
rect 514024 270852 514076 270904
rect 543004 270852 543056 270904
rect 426992 270716 427044 270768
rect 495072 270716 495124 270768
rect 136824 270580 136876 270632
rect 174636 270580 174688 270632
rect 108948 270444 109000 270496
rect 162400 270444 162452 270496
rect 173808 270444 173860 270496
rect 176936 270444 176988 270496
rect 353208 270580 353260 270632
rect 403992 270580 404044 270632
rect 404176 270580 404228 270632
rect 409512 270580 409564 270632
rect 409696 270580 409748 270632
rect 495440 270580 495492 270632
rect 495900 270580 495952 270632
rect 531596 270716 531648 270768
rect 496360 270580 496412 270632
rect 514024 270580 514076 270632
rect 514208 270580 514260 270632
rect 518624 270580 518676 270632
rect 78864 270308 78916 270360
rect 132592 270308 132644 270360
rect 133788 270308 133840 270360
rect 177580 270308 177632 270360
rect 203616 270444 203668 270496
rect 207020 270444 207072 270496
rect 209504 270444 209556 270496
rect 216680 270444 216732 270496
rect 224960 270444 225012 270496
rect 244372 270444 244424 270496
rect 247776 270444 247828 270496
rect 250168 270444 250220 270496
rect 251456 270444 251508 270496
rect 258816 270444 258868 270496
rect 261300 270444 261352 270496
rect 292672 270444 292724 270496
rect 305092 270444 305144 270496
rect 323584 270444 323636 270496
rect 365812 270444 365864 270496
rect 367744 270444 367796 270496
rect 436100 270444 436152 270496
rect 438400 270444 438452 270496
rect 543004 270444 543056 270496
rect 543188 270444 543240 270496
rect 557816 270444 557868 270496
rect 205824 270308 205876 270360
rect 212264 270308 212316 270360
rect 219440 270308 219492 270360
rect 243176 270308 243228 270360
rect 247040 270308 247092 270360
rect 261024 270308 261076 270360
rect 264980 270308 265032 270360
rect 301964 270308 302016 270360
rect 320272 270308 320324 270360
rect 334992 270308 335044 270360
rect 383660 270308 383712 270360
rect 383844 270308 383896 270360
rect 386420 270308 386472 270360
rect 386604 270308 386656 270360
rect 456616 270308 456668 270360
rect 456754 270308 456806 270360
rect 475936 270308 475988 270360
rect 476488 270308 476540 270360
rect 599400 270308 599452 270360
rect 94228 270172 94280 270224
rect 153568 270172 153620 270224
rect 163688 270172 163740 270224
rect 195520 270172 195572 270224
rect 197544 270172 197596 270224
rect 205088 270172 205140 270224
rect 205548 270172 205600 270224
rect 223488 270172 223540 270224
rect 290832 270172 290884 270224
rect 311900 270172 311952 270224
rect 312820 270172 312872 270224
rect 331404 270172 331456 270224
rect 346400 270172 346452 270224
rect 393504 270172 393556 270224
rect 393872 270172 393924 270224
rect 67548 270036 67600 270088
rect 78220 270036 78272 270088
rect 80060 270036 80112 270088
rect 144460 270036 144512 270088
rect 152648 270036 152700 270088
rect 188896 270036 188948 270088
rect 202972 270036 203024 270088
rect 222016 270036 222068 270088
rect 226616 270036 226668 270088
rect 236736 270036 236788 270088
rect 266176 270036 266228 270088
rect 273260 270036 273312 270088
rect 276480 270036 276532 270088
rect 289820 270036 289872 270088
rect 301228 270036 301280 270088
rect 324320 270036 324372 270088
rect 337200 270036 337252 270088
rect 383844 270036 383896 270088
rect 384120 270036 384172 270088
rect 393688 270036 393740 270088
rect 395988 270036 396040 270088
rect 398472 270172 398524 270224
rect 401876 270172 401928 270224
rect 402244 270172 402296 270224
rect 412594 270172 412646 270224
rect 412732 270172 412784 270224
rect 475752 270172 475804 270224
rect 476212 270172 476264 270224
rect 490288 270172 490340 270224
rect 500224 270172 500276 270224
rect 500408 270172 500460 270224
rect 501972 270172 502024 270224
rect 502156 270172 502208 270224
rect 633624 270172 633676 270224
rect 75828 269900 75880 269952
rect 141792 269900 141844 269952
rect 143908 269900 143960 269952
rect 184480 269900 184532 269952
rect 184756 269900 184808 269952
rect 189632 269900 189684 269952
rect 194600 269900 194652 269952
rect 216864 269900 216916 269952
rect 221464 269900 221516 269952
rect 229376 269900 229428 269952
rect 230388 269900 230440 269952
rect 238944 269900 238996 269952
rect 266912 269900 266964 269952
rect 274640 269900 274692 269952
rect 275008 269900 275060 269952
rect 287060 269900 287112 269952
rect 287520 269900 287572 269952
rect 307760 269900 307812 269952
rect 310336 269900 310388 269952
rect 339224 269900 339276 269952
rect 339408 269900 339460 269952
rect 390560 269900 390612 269952
rect 390744 269900 390796 269952
rect 475752 270036 475804 270088
rect 475936 270036 475988 270088
rect 619456 270036 619508 270088
rect 69388 269764 69440 269816
rect 138848 269764 138900 269816
rect 140780 269764 140832 269816
rect 182272 269764 182324 269816
rect 191748 269764 191800 269816
rect 214656 269764 214708 269816
rect 219624 269764 219676 269816
rect 232320 269764 232372 269816
rect 237196 269764 237248 269816
rect 243360 269764 243412 269816
rect 261760 269764 261812 269816
rect 263600 269764 263652 269816
rect 265440 269764 265492 269816
rect 271880 269764 271932 269816
rect 283104 269764 283156 269816
rect 300860 269764 300912 269816
rect 305552 269764 305604 269816
rect 335360 269764 335412 269816
rect 341248 269764 341300 269816
rect 384120 269764 384172 269816
rect 122748 269628 122800 269680
rect 171232 269628 171284 269680
rect 172428 269628 172480 269680
rect 202144 269628 202196 269680
rect 271880 269628 271932 269680
rect 281540 269628 281592 269680
rect 311532 269628 311584 269680
rect 327264 269628 327316 269680
rect 332324 269628 332376 269680
rect 84108 269492 84160 269544
rect 126704 269492 126756 269544
rect 126888 269492 126940 269544
rect 173440 269492 173492 269544
rect 183468 269492 183520 269544
rect 194508 269492 194560 269544
rect 259644 269492 259696 269544
rect 260840 269492 260892 269544
rect 330208 269492 330260 269544
rect 374460 269492 374512 269544
rect 374828 269628 374880 269680
rect 397552 269764 397604 269816
rect 481640 269900 481692 269952
rect 484308 269900 484360 269952
rect 407948 269764 408000 269816
rect 408132 269764 408184 269816
rect 484676 269764 484728 269816
rect 485044 269900 485096 269952
rect 490196 269900 490248 269952
rect 490840 269900 490892 269952
rect 495256 269900 495308 269952
rect 490840 269764 490892 269816
rect 491392 269764 491444 269816
rect 491576 269764 491628 269816
rect 626540 269900 626592 269952
rect 495532 269764 495584 269816
rect 637580 269764 637632 269816
rect 638316 269764 638368 269816
rect 647240 269764 647292 269816
rect 384488 269628 384540 269680
rect 412732 269628 412784 269680
rect 413100 269628 413152 269680
rect 427820 269628 427872 269680
rect 428004 269628 428056 269680
rect 527180 269628 527232 269680
rect 543004 269628 543056 269680
rect 549904 269628 549956 269680
rect 379520 269492 379572 269544
rect 379704 269492 379756 269544
rect 129372 269356 129424 269408
rect 175648 269356 175700 269408
rect 328000 269356 328052 269408
rect 264704 269288 264756 269340
rect 265900 269288 265952 269340
rect 128544 269220 128596 269272
rect 162952 269220 163004 269272
rect 365720 269356 365772 269408
rect 374828 269356 374880 269408
rect 375012 269356 375064 269408
rect 393412 269356 393464 269408
rect 393596 269356 393648 269408
rect 398288 269356 398340 269408
rect 398472 269356 398524 269408
rect 407948 269492 408000 269544
rect 422576 269492 422628 269544
rect 500040 269492 500092 269544
rect 500224 269492 500276 269544
rect 543188 269492 543240 269544
rect 248328 269084 248380 269136
rect 249984 269084 250036 269136
rect 274640 269084 274692 269136
rect 278964 269084 279016 269136
rect 372528 269220 372580 269272
rect 406108 269220 406160 269272
rect 412916 269356 412968 269408
rect 413100 269356 413152 269408
rect 413928 269356 413980 269408
rect 414112 269356 414164 269408
rect 423128 269356 423180 269408
rect 423680 269356 423732 269408
rect 424416 269356 424468 269408
rect 427636 269356 427688 269408
rect 427820 269356 427872 269408
rect 521660 269356 521712 269408
rect 408132 269220 408184 269272
rect 408316 269220 408368 269272
rect 412456 269220 412508 269272
rect 412732 269220 412784 269272
rect 416412 269220 416464 269272
rect 416688 269152 416740 269204
rect 513380 269220 513432 269272
rect 372712 269084 372764 269136
rect 373908 269084 373960 269136
rect 375012 269084 375064 269136
rect 42340 269016 42392 269068
rect 45560 269016 45612 269068
rect 118608 269016 118660 269068
rect 169760 269016 169812 269068
rect 225420 269016 225472 269068
rect 227628 269016 227680 269068
rect 324320 269016 324372 269068
rect 336740 269016 336792 269068
rect 338488 269016 338540 269068
rect 359096 269016 359148 269068
rect 269120 268948 269172 269000
rect 276664 268948 276716 269000
rect 374460 268948 374512 269000
rect 376944 269084 376996 269136
rect 378048 269016 378100 269068
rect 384304 269016 384356 269068
rect 384488 269016 384540 269068
rect 398104 269016 398156 269068
rect 398288 269016 398340 269068
rect 466276 269016 466328 269068
rect 466460 269016 466512 269068
rect 468116 269016 468168 269068
rect 471244 269016 471296 269068
rect 587900 269016 587952 269068
rect 104900 268880 104952 268932
rect 160192 268880 160244 268932
rect 187516 268880 187568 268932
rect 208492 268880 208544 268932
rect 304172 268880 304224 268932
rect 329840 268880 329892 268932
rect 347412 268880 347464 268932
rect 77208 268744 77260 268796
rect 104900 268744 104952 268796
rect 106280 268744 106332 268796
rect 161664 268744 161716 268796
rect 166172 268744 166224 268796
rect 194048 268744 194100 268796
rect 203892 268744 203944 268796
rect 211160 268744 211212 268796
rect 284576 268744 284628 268796
rect 285864 268744 285916 268796
rect 314752 268744 314804 268796
rect 352104 268744 352156 268796
rect 375840 268880 375892 268932
rect 449900 268880 449952 268932
rect 455328 268880 455380 268932
rect 461400 268880 461452 268932
rect 462504 268880 462556 268932
rect 581000 268880 581052 268932
rect 376024 268744 376076 268796
rect 384304 268744 384356 268796
rect 440424 268744 440476 268796
rect 95424 268608 95476 268660
rect 155040 268608 155092 268660
rect 162584 268608 162636 268660
rect 190092 268608 190144 268660
rect 190368 268608 190420 268660
rect 204076 268608 204128 268660
rect 285772 268608 285824 268660
rect 295340 268608 295392 268660
rect 299296 268608 299348 268660
rect 316776 268608 316828 268660
rect 317696 268608 317748 268660
rect 355692 268608 355744 268660
rect 369216 268608 369268 268660
rect 437296 268608 437348 268660
rect 437434 268608 437486 268660
rect 460112 268744 460164 268796
rect 87144 268472 87196 268524
rect 149888 268472 149940 268524
rect 162768 268472 162820 268524
rect 196992 268472 197044 268524
rect 208860 268472 208912 268524
rect 225696 268472 225748 268524
rect 281632 268472 281684 268524
rect 295524 268472 295576 268524
rect 297088 268472 297140 268524
rect 322940 268472 322992 268524
rect 329472 268472 329524 268524
rect 340880 268472 340932 268524
rect 349344 268472 349396 268524
rect 371056 268472 371108 268524
rect 371424 268472 371476 268524
rect 432604 268472 432656 268524
rect 434720 268472 434772 268524
rect 456432 268608 456484 268660
rect 460296 268608 460348 268660
rect 583852 268744 583904 268796
rect 461952 268608 462004 268660
rect 440884 268472 440936 268524
rect 442816 268472 442868 268524
rect 443000 268472 443052 268524
rect 456432 268472 456484 268524
rect 456984 268472 457036 268524
rect 466414 268472 466466 268524
rect 467104 268608 467156 268660
rect 594800 268608 594852 268660
rect 594984 268608 595036 268660
rect 645860 268608 645912 268660
rect 471244 268472 471296 268524
rect 471428 268472 471480 268524
rect 474740 268472 474792 268524
rect 475200 268472 475252 268524
rect 608692 268472 608744 268524
rect 669320 268472 669372 268524
rect 675484 268472 675536 268524
rect 82728 268336 82780 268388
rect 146944 268336 146996 268388
rect 148876 268336 148928 268388
rect 188160 268336 188212 268388
rect 188436 268336 188488 268388
rect 115756 268200 115808 268252
rect 166816 268200 166868 268252
rect 210976 268336 211028 268388
rect 219808 268336 219860 268388
rect 220728 268336 220780 268388
rect 230756 268336 230808 268388
rect 273536 268336 273588 268388
rect 282920 268336 282972 268388
rect 286784 268336 286836 268388
rect 306380 268336 306432 268388
rect 316960 268336 317012 268388
rect 354680 268336 354732 268388
rect 358544 268336 358596 268388
rect 407396 268336 407448 268388
rect 210976 268200 211028 268252
rect 324688 268200 324740 268252
rect 367100 268200 367152 268252
rect 382464 268200 382516 268252
rect 384488 268200 384540 268252
rect 387616 268200 387668 268252
rect 397920 268200 397972 268252
rect 398104 268200 398156 268252
rect 417424 268336 417476 268388
rect 417608 268336 417660 268388
rect 456616 268336 456668 268388
rect 456800 268336 456852 268388
rect 495072 268336 495124 268388
rect 495532 268336 495584 268388
rect 504916 268336 504968 268388
rect 505054 268336 505106 268388
rect 607220 268336 607272 268388
rect 407948 268200 408000 268252
rect 446772 268200 446824 268252
rect 452384 268200 452436 268252
rect 456616 268200 456668 268252
rect 461584 268200 461636 268252
rect 480904 268200 480956 268252
rect 481088 268200 481140 268252
rect 484860 268200 484912 268252
rect 485688 268200 485740 268252
rect 485872 268200 485924 268252
rect 486056 268200 486108 268252
rect 572720 268200 572772 268252
rect 135260 268064 135312 268116
rect 138112 268064 138164 268116
rect 147496 268064 147548 268116
rect 186688 268064 186740 268116
rect 365352 268064 365404 268116
rect 432052 268064 432104 268116
rect 432604 268064 432656 268116
rect 440240 268064 440292 268116
rect 440424 268064 440476 268116
rect 452660 268064 452712 268116
rect 457536 268064 457588 268116
rect 461032 268064 461084 268116
rect 461400 268064 461452 268116
rect 484676 268064 484728 268116
rect 486424 268064 486476 268116
rect 563060 268064 563112 268116
rect 658924 267996 658976 268048
rect 675484 268268 675536 268320
rect 354680 267928 354732 267980
rect 42524 267656 42576 267708
rect 45928 267656 45980 267708
rect 104900 267656 104952 267708
rect 137560 267724 137612 267776
rect 140044 267656 140096 267708
rect 143448 267792 143500 267844
rect 355968 267792 356020 267844
rect 388996 267792 389048 267844
rect 402612 267928 402664 267980
rect 407948 267928 408000 267980
rect 411168 267928 411220 267980
rect 404452 267792 404504 267844
rect 407396 267792 407448 267844
rect 410064 267792 410116 267844
rect 410248 267792 410300 267844
rect 263968 267724 264020 267776
rect 269580 267724 269632 267776
rect 344192 267724 344244 267776
rect 347044 267724 347096 267776
rect 142804 267656 142856 267708
rect 166080 267656 166132 267708
rect 213184 267656 213236 267708
rect 220544 267656 220596 267708
rect 288256 267656 288308 267708
rect 297364 267656 297416 267708
rect 305920 267656 305972 267708
rect 324320 267656 324372 267708
rect 343364 267588 343416 267640
rect 132408 267520 132460 267572
rect 178592 267520 178644 267572
rect 180064 267520 180116 267572
rect 207296 267520 207348 267572
rect 286048 267520 286100 267572
rect 290464 267520 290516 267572
rect 294880 267520 294932 267572
rect 300124 267520 300176 267572
rect 319168 267520 319220 267572
rect 338488 267520 338540 267572
rect 350264 267520 350316 267572
rect 364156 267520 364208 267572
rect 364800 267656 364852 267708
rect 372528 267656 372580 267708
rect 372896 267656 372948 267708
rect 365720 267520 365772 267572
rect 366272 267520 366324 267572
rect 374460 267520 374512 267572
rect 375012 267656 375064 267708
rect 410708 267656 410760 267708
rect 415308 267792 415360 267844
rect 417424 267928 417476 267980
rect 427636 267928 427688 267980
rect 427820 267928 427872 267980
rect 437296 267928 437348 267980
rect 437434 267928 437486 267980
rect 541348 267928 541400 267980
rect 660304 267860 660356 267912
rect 669320 267860 669372 267912
rect 417608 267792 417660 267844
rect 417792 267792 417844 267844
rect 422300 267792 422352 267844
rect 422944 267792 422996 267844
rect 475752 267792 475804 267844
rect 476212 267792 476264 267844
rect 480720 267792 480772 267844
rect 480904 267792 480956 267844
rect 485044 267792 485096 267844
rect 486240 267792 486292 267844
rect 494520 267792 494572 267844
rect 415308 267656 415360 267708
rect 417884 267656 417936 267708
rect 418344 267656 418396 267708
rect 490196 267656 490248 267708
rect 491392 267656 491444 267708
rect 492588 267656 492640 267708
rect 492772 267656 492824 267708
rect 524696 267792 524748 267844
rect 664812 267724 664864 267776
rect 494888 267656 494940 267708
rect 525984 267656 526036 267708
rect 675484 267792 675536 267844
rect 411996 267520 412048 267572
rect 412180 267520 412232 267572
rect 412594 267520 412646 267572
rect 412732 267520 412784 267572
rect 414664 267520 414716 267572
rect 415308 267520 415360 267572
rect 100668 267384 100720 267436
rect 158720 267384 158772 267436
rect 162952 267384 163004 267436
rect 78220 267248 78272 267300
rect 137376 267248 137428 267300
rect 137560 267248 137612 267300
rect 143264 267248 143316 267300
rect 143448 267248 143500 267300
rect 173900 267248 173952 267300
rect 175924 267384 175976 267436
rect 202880 267384 202932 267436
rect 204076 267384 204128 267436
rect 213184 267384 213236 267436
rect 222844 267384 222896 267436
rect 231584 267384 231636 267436
rect 295616 267384 295668 267436
rect 301964 267384 302016 267436
rect 308128 267384 308180 267436
rect 329472 267384 329524 267436
rect 176384 267248 176436 267300
rect 86224 267112 86276 267164
rect 145932 267112 145984 267164
rect 146208 267112 146260 267164
rect 187424 267248 187476 267300
rect 194508 267248 194560 267300
rect 208768 267248 208820 267300
rect 228456 267248 228508 267300
rect 233792 267248 233844 267300
rect 262864 267248 262916 267300
rect 267924 267248 267976 267300
rect 275744 267248 275796 267300
rect 280988 267248 281040 267300
rect 282368 267248 282420 267300
rect 289084 267248 289136 267300
rect 257344 267180 257396 267232
rect 259460 267180 259512 267232
rect 186964 267112 187016 267164
rect 91008 266976 91060 267028
rect 152096 266976 152148 267028
rect 156512 266976 156564 267028
rect 165344 266976 165396 267028
rect 167920 266976 167972 267028
rect 198464 266976 198516 267028
rect 211160 267112 211212 267164
rect 222752 267112 222804 267164
rect 233240 267112 233292 267164
rect 240416 267112 240468 267164
rect 267648 267112 267700 267164
rect 271144 267112 271196 267164
rect 272064 267112 272116 267164
rect 280712 267112 280764 267164
rect 293408 267112 293460 267164
rect 302884 267248 302936 267300
rect 306656 267248 306708 267300
rect 312544 267248 312596 267300
rect 302240 267112 302292 267164
rect 312820 267112 312872 267164
rect 313280 267112 313332 267164
rect 334624 267248 334676 267300
rect 330484 267112 330536 267164
rect 345848 267384 345900 267436
rect 347688 267384 347740 267436
rect 353944 267384 353996 267436
rect 335728 267248 335780 267300
rect 348424 267248 348476 267300
rect 350080 267248 350132 267300
rect 364984 267384 365036 267436
rect 365168 267384 365220 267436
rect 370504 267384 370556 267436
rect 370688 267384 370740 267436
rect 374828 267384 374880 267436
rect 355232 267248 355284 267300
rect 363236 267248 363288 267300
rect 376760 267384 376812 267436
rect 341984 267112 342036 267164
rect 350264 267112 350316 267164
rect 350816 267112 350868 267164
rect 375472 267248 375524 267300
rect 384304 267384 384356 267436
rect 384488 267384 384540 267436
rect 379520 267248 379572 267300
rect 383660 267248 383712 267300
rect 383936 267248 383988 267300
rect 388996 267248 389048 267300
rect 392032 267384 392084 267436
rect 393228 267384 393280 267436
rect 393412 267384 393464 267436
rect 421104 267384 421156 267436
rect 421472 267520 421524 267572
rect 422116 267520 422168 267572
rect 422300 267520 422352 267572
rect 423496 267520 423548 267572
rect 423680 267520 423732 267572
rect 424968 267520 425020 267572
rect 425152 267520 425204 267572
rect 426256 267520 426308 267572
rect 426440 267520 426492 267572
rect 427774 267520 427826 267572
rect 427912 267520 427964 267572
rect 442264 267384 442316 267436
rect 442724 267384 442776 267436
rect 446588 267384 446640 267436
rect 447232 267384 447284 267436
rect 461584 267384 461636 267436
rect 461768 267384 461820 267436
rect 466092 267384 466144 267436
rect 467840 267520 467892 267572
rect 475752 267520 475804 267572
rect 476120 267520 476172 267572
rect 538864 267520 538916 267572
rect 415492 267248 415544 267300
rect 364984 267112 365036 267164
rect 373908 267112 373960 267164
rect 374460 267112 374512 267164
rect 402244 267112 402296 267164
rect 402980 267112 403032 267164
rect 446772 267248 446824 267300
rect 447416 267248 447468 267300
rect 477132 267248 477184 267300
rect 480352 267384 480404 267436
rect 481456 267384 481508 267436
rect 481640 267384 481692 267436
rect 490564 267384 490616 267436
rect 490840 267384 490892 267436
rect 572168 267384 572220 267436
rect 490564 267248 490616 267300
rect 490840 267248 490892 267300
rect 494888 267248 494940 267300
rect 416320 267112 416372 267164
rect 426440 267112 426492 267164
rect 426624 267112 426676 267164
rect 431224 267112 431276 267164
rect 434720 267112 434772 267164
rect 436192 267112 436244 267164
rect 437112 267112 437164 267164
rect 437296 267112 437348 267164
rect 442080 267112 442132 267164
rect 442264 267112 442316 267164
rect 211712 266976 211764 267028
rect 212448 266976 212500 267028
rect 227168 266976 227220 267028
rect 227628 266976 227680 267028
rect 236000 266976 236052 267028
rect 278688 266976 278740 267028
rect 293224 266976 293276 267028
rect 300032 266976 300084 267028
rect 311532 266976 311584 267028
rect 312544 266976 312596 267028
rect 342536 266976 342588 267028
rect 344928 266976 344980 267028
rect 351184 266976 351236 267028
rect 353024 266976 353076 267028
rect 379704 266976 379756 267028
rect 379888 266976 379940 267028
rect 384488 266976 384540 267028
rect 384672 266976 384724 267028
rect 387800 266976 387852 267028
rect 388352 266976 388404 267028
rect 393136 266976 393188 267028
rect 393320 266976 393372 267028
rect 430672 266976 430724 267028
rect 436744 266976 436796 267028
rect 437112 266976 437164 267028
rect 446772 266976 446824 267028
rect 451924 267112 451976 267164
rect 466414 267112 466466 267164
rect 466552 267112 466604 267164
rect 475752 267112 475804 267164
rect 461400 266976 461452 267028
rect 461584 266976 461636 267028
rect 490840 267112 490892 267164
rect 496544 267248 496596 267300
rect 504916 267248 504968 267300
rect 505054 267248 505106 267300
rect 550364 267248 550416 267300
rect 497464 267112 497516 267164
rect 498752 267112 498804 267164
rect 490564 267044 490616 267096
rect 638316 267112 638368 267164
rect 476396 266976 476448 267028
rect 476948 266976 477000 267028
rect 477132 266976 477184 267028
rect 487528 266976 487580 267028
rect 487712 266976 487764 267028
rect 489828 266976 489880 267028
rect 504548 266976 504600 267028
rect 505192 266976 505244 267028
rect 632704 266976 632756 267028
rect 119344 266840 119396 266892
rect 109684 266704 109736 266756
rect 140320 266704 140372 266756
rect 145564 266840 145616 266892
rect 151360 266840 151412 266892
rect 157984 266840 158036 266892
rect 174176 266840 174228 266892
rect 256516 266840 256568 266892
rect 258080 266840 258132 266892
rect 311072 266840 311124 266892
rect 319444 266840 319496 266892
rect 321284 266840 321336 266892
rect 330484 266840 330536 266892
rect 154304 266704 154356 266756
rect 173900 266704 173952 266756
rect 183008 266704 183060 266756
rect 206284 266704 206336 266756
rect 210240 266704 210292 266756
rect 327264 266704 327316 266756
rect 330944 266704 330996 266756
rect 333244 266704 333296 266756
rect 126704 266568 126756 266620
rect 148416 266568 148468 266620
rect 151176 266568 151228 266620
rect 163136 266568 163188 266620
rect 210608 266568 210660 266620
rect 217600 266568 217652 266620
rect 246304 266568 246356 266620
rect 248512 266568 248564 266620
rect 325792 266568 325844 266620
rect 326712 266568 326764 266620
rect 331680 266568 331732 266620
rect 332508 266568 332560 266620
rect 333888 266840 333940 266892
rect 347688 266840 347740 266892
rect 347872 266840 347924 266892
rect 353576 266840 353628 266892
rect 359648 266840 359700 266892
rect 390744 266840 390796 266892
rect 391296 266840 391348 266892
rect 392216 266840 392268 266892
rect 392768 266840 392820 266892
rect 466276 266840 466328 266892
rect 338304 266704 338356 266756
rect 358176 266704 358228 266756
rect 345664 266568 345716 266620
rect 353576 266568 353628 266620
rect 354680 266568 354732 266620
rect 357440 266568 357492 266620
rect 365168 266704 365220 266756
rect 367008 266704 367060 266756
rect 396724 266704 396776 266756
rect 397184 266704 397236 266756
rect 402796 266704 402848 266756
rect 403072 266704 403124 266756
rect 404176 266704 404228 266756
rect 406016 266704 406068 266756
rect 410248 266704 410300 266756
rect 410432 266704 410484 266756
rect 412088 266704 412140 266756
rect 412456 266704 412508 266756
rect 415308 266704 415360 266756
rect 415584 266704 415636 266756
rect 416688 266704 416740 266756
rect 418252 266704 418304 266756
rect 426624 266704 426676 266756
rect 358912 266568 358964 266620
rect 360108 266568 360160 266620
rect 360384 266568 360436 266620
rect 361212 266568 361264 266620
rect 363236 266568 363288 266620
rect 382188 266568 382240 266620
rect 241336 266500 241388 266552
rect 245568 266500 245620 266552
rect 259920 266500 259972 266552
rect 262588 266500 262640 266552
rect 269856 266500 269908 266552
rect 274640 266500 274692 266552
rect 280160 266500 280212 266552
rect 285772 266500 285824 266552
rect 291200 266500 291252 266552
rect 294604 266500 294656 266552
rect 301504 266500 301556 266552
rect 304172 266500 304224 266552
rect 304448 266500 304500 266552
rect 305552 266500 305604 266552
rect 319904 266500 319956 266552
rect 322204 266500 322256 266552
rect 348608 266500 348660 266552
rect 132592 266432 132644 266484
rect 145472 266432 145524 266484
rect 208492 266432 208544 266484
rect 212448 266432 212500 266484
rect 322480 266432 322532 266484
rect 338948 266432 339000 266484
rect 364800 266432 364852 266484
rect 370504 266432 370556 266484
rect 378784 266432 378836 266484
rect 381728 266432 381780 266484
rect 384948 266568 385000 266620
rect 385408 266568 385460 266620
rect 389824 266568 389876 266620
rect 390560 266568 390612 266620
rect 391848 266568 391900 266620
rect 392216 266568 392268 266620
rect 436560 266704 436612 266756
rect 437940 266704 437992 266756
rect 451924 266704 451976 266756
rect 452108 266704 452160 266756
rect 454592 266704 454644 266756
rect 454776 266704 454828 266756
rect 491208 266840 491260 266892
rect 629300 266840 629352 266892
rect 666192 266772 666244 266824
rect 675484 266772 675536 266824
rect 466736 266704 466788 266756
rect 469864 266704 469916 266756
rect 470048 266704 470100 266756
rect 504732 266704 504784 266756
rect 504916 266704 504968 266756
rect 543740 266704 543792 266756
rect 550364 266704 550416 266756
rect 594984 266704 595036 266756
rect 427912 266568 427964 266620
rect 437112 266568 437164 266620
rect 384304 266432 384356 266484
rect 401140 266432 401192 266484
rect 401600 266432 401652 266484
rect 402612 266432 402664 266484
rect 402796 266432 402848 266484
rect 466552 266568 466604 266620
rect 466920 266568 466972 266620
rect 476028 266568 476080 266620
rect 476212 266568 476264 266620
rect 481640 266568 481692 266620
rect 482560 266568 482612 266620
rect 485596 266568 485648 266620
rect 485780 266568 485832 266620
rect 554044 266568 554096 266620
rect 666376 266500 666428 266552
rect 675484 266568 675536 266620
rect 437756 266432 437808 266484
rect 153844 266364 153896 266416
rect 156144 266364 156196 266416
rect 164884 266364 164936 266416
rect 167552 266364 167604 266416
rect 174728 266364 174780 266416
rect 180064 266364 180116 266416
rect 204904 266364 204956 266416
rect 206560 266364 206612 266416
rect 219440 266364 219492 266416
rect 227904 266364 227956 266416
rect 230756 266364 230808 266416
rect 233056 266364 233108 266416
rect 239496 266364 239548 266416
rect 241888 266364 241940 266416
rect 251180 266364 251232 266416
rect 252192 266364 252244 266416
rect 255872 266364 255924 266416
rect 256700 266364 256752 266416
rect 258080 266364 258132 266416
rect 259644 266364 259696 266416
rect 260288 266364 260340 266416
rect 261760 266364 261812 266416
rect 262128 266364 262180 266416
rect 266360 266364 266412 266416
rect 270592 266364 270644 266416
rect 271604 266364 271656 266416
rect 280896 266364 280948 266416
rect 282184 266364 282236 266416
rect 288992 266364 289044 266416
rect 291844 266364 291896 266416
rect 294144 266364 294196 266416
rect 295156 266364 295208 266416
rect 297824 266364 297876 266416
rect 301228 266364 301280 266416
rect 303712 266364 303764 266416
rect 304908 266364 304960 266416
rect 305184 266364 305236 266416
rect 306196 266364 306248 266416
rect 316224 266364 316276 266416
rect 317144 266364 317196 266416
rect 320640 266364 320692 266416
rect 321468 266364 321520 266416
rect 342720 266364 342772 266416
rect 343548 266364 343600 266416
rect 346400 266364 346452 266416
rect 350080 266364 350132 266416
rect 352288 266364 352340 266416
rect 353208 266364 353260 266416
rect 372160 266296 372212 266348
rect 432604 266296 432656 266348
rect 373632 266160 373684 266212
rect 441712 266296 441764 266348
rect 442080 266432 442132 266484
rect 532976 266432 533028 266484
rect 664812 266364 664864 266416
rect 675300 266364 675352 266416
rect 442724 266296 442776 266348
rect 442908 266296 442960 266348
rect 445944 266296 445996 266348
rect 450544 266296 450596 266348
rect 452108 266296 452160 266348
rect 404176 266024 404228 266076
rect 412456 266024 412508 266076
rect 432604 266024 432656 266076
rect 443184 266160 443236 266212
rect 443920 266160 443972 266212
rect 448520 266160 448572 266212
rect 448704 266160 448756 266212
rect 566280 266296 566332 266348
rect 454592 266160 454644 266212
rect 575756 266160 575808 266212
rect 442264 266024 442316 266076
rect 461584 266024 461636 266076
rect 462136 266024 462188 266076
rect 463976 266024 464028 266076
rect 464160 266024 464212 266076
rect 591028 266024 591080 266076
rect 198740 265888 198792 265940
rect 199660 265888 199712 265940
rect 218060 265888 218112 265940
rect 218796 265888 218848 265940
rect 389088 265888 389140 265940
rect 470600 265888 470652 265940
rect 470784 265888 470836 265940
rect 601700 265888 601752 265940
rect 362592 265752 362644 265804
rect 428280 265752 428332 265804
rect 437664 265752 437716 265804
rect 523684 265752 523736 265804
rect 384672 265616 384724 265668
rect 461400 265616 461452 265668
rect 461584 265616 461636 265668
rect 495900 265616 495952 265668
rect 499488 265616 499540 265668
rect 648620 265616 648672 265668
rect 669320 265548 669372 265600
rect 675484 265548 675536 265600
rect 404544 265480 404596 265532
rect 442264 265480 442316 265532
rect 444288 265480 444340 265532
rect 559288 265480 559340 265532
rect 665272 265412 665324 265464
rect 675484 265412 675536 265464
rect 442080 265344 442132 265396
rect 552664 265344 552716 265396
rect 417792 265208 417844 265260
rect 516416 265208 516468 265260
rect 665088 265208 665140 265260
rect 675300 265208 675352 265260
rect 439872 265072 439924 265124
rect 537760 265072 537812 265124
rect 664260 265072 664312 265124
rect 675484 265004 675536 265056
rect 386144 264936 386196 264988
rect 467288 264936 467340 264988
rect 477408 264936 477460 264988
rect 612740 264936 612792 264988
rect 664260 264936 664312 264988
rect 669320 264868 669372 264920
rect 435456 264732 435508 264784
rect 545120 264732 545172 264784
rect 453120 264596 453172 264648
rect 574100 264596 574152 264648
rect 471888 264460 471940 264512
rect 603080 264460 603132 264512
rect 491024 264324 491076 264376
rect 491576 264324 491628 264376
rect 497648 264324 497700 264376
rect 643744 264324 643796 264376
rect 51908 264188 51960 264240
rect 655520 264188 655572 264240
rect 507124 264052 507176 264104
rect 600596 264052 600648 264104
rect 666192 263576 666244 263628
rect 675484 263576 675536 263628
rect 666376 262488 666428 262540
rect 675484 262488 675536 262540
rect 669412 262080 669464 262132
rect 675484 262080 675536 262132
rect 511540 261468 511592 261520
rect 568580 261468 568632 261520
rect 675852 260992 675904 261044
rect 676404 260992 676456 261044
rect 673368 260448 673420 260500
rect 675484 260448 675536 260500
rect 669136 259836 669188 259888
rect 675484 259836 675536 259888
rect 671896 259632 671948 259684
rect 675484 259632 675536 259684
rect 510988 259428 511040 259480
rect 514024 259428 514076 259480
rect 673092 258816 673144 258868
rect 675484 258816 675536 258868
rect 672724 258408 672776 258460
rect 675484 258408 675536 258460
rect 35808 258204 35860 258256
rect 40040 258204 40092 258256
rect 35808 257116 35860 257168
rect 39580 257116 39632 257168
rect 35808 256844 35860 256896
rect 40408 256912 40460 256964
rect 42064 256844 42116 256896
rect 49516 256844 49568 256896
rect 35624 256708 35676 256760
rect 41696 256776 41748 256828
rect 510804 256708 510856 256760
rect 567200 256708 567252 256760
rect 675852 256708 675904 256760
rect 683120 256708 683172 256760
rect 35808 255688 35860 255740
rect 41420 255688 41472 255740
rect 35624 255416 35676 255468
rect 41696 255484 41748 255536
rect 42064 255484 42116 255536
rect 42892 255484 42944 255536
rect 35808 255280 35860 255332
rect 41696 255280 41748 255332
rect 42064 255280 42116 255332
rect 45560 255280 45612 255332
rect 35532 254532 35584 254584
rect 39304 254532 39356 254584
rect 35808 254260 35860 254312
rect 39948 254328 40000 254380
rect 35348 254056 35400 254108
rect 40316 254124 40368 254176
rect 35164 253920 35216 253972
rect 41696 253920 41748 253972
rect 42064 253920 42116 253972
rect 43812 253920 43864 253972
rect 669596 253172 669648 253224
rect 675484 253172 675536 253224
rect 35808 252832 35860 252884
rect 41696 252832 41748 252884
rect 42064 252832 42116 252884
rect 42708 252832 42760 252884
rect 35624 252696 35676 252748
rect 41696 252696 41748 252748
rect 35808 252560 35860 252612
rect 41512 252560 41564 252612
rect 511908 252560 511960 252612
rect 559564 252560 559616 252612
rect 35808 251608 35860 251660
rect 40592 251608 40644 251660
rect 35808 251336 35860 251388
rect 41328 251336 41380 251388
rect 35624 251200 35676 251252
rect 41512 251200 41564 251252
rect 511540 250452 511592 250504
rect 571340 250452 571392 250504
rect 669412 250384 669464 250436
rect 672908 250384 672960 250436
rect 35808 250180 35860 250232
rect 39396 250180 39448 250232
rect 35624 249908 35676 249960
rect 40132 249976 40184 250028
rect 35440 249772 35492 249824
rect 39580 249772 39632 249824
rect 35532 248684 35584 248736
rect 39948 248684 40000 248736
rect 35808 248412 35860 248464
rect 40132 248412 40184 248464
rect 674840 247868 674892 247920
rect 675392 247868 675444 247920
rect 35808 247528 35860 247580
rect 41512 247528 41564 247580
rect 42156 247460 42208 247512
rect 129096 247460 129148 247512
rect 35624 247324 35676 247376
rect 40132 247324 40184 247376
rect 35624 247188 35676 247240
rect 41052 247188 41104 247240
rect 510988 247120 511040 247172
rect 512644 247120 512696 247172
rect 35440 247052 35492 247104
rect 41512 247052 41564 247104
rect 42064 247052 42116 247104
rect 129004 247052 129056 247104
rect 674472 246984 674524 247036
rect 675392 246984 675444 247036
rect 510804 246304 510856 246356
rect 570052 246304 570104 246356
rect 663708 244876 663760 244928
rect 669320 244876 669372 244928
rect 511264 242156 511316 242208
rect 632704 242156 632756 242208
rect 673092 241680 673144 241732
rect 675300 241680 675352 241732
rect 673368 241544 673420 241596
rect 666376 241408 666428 241460
rect 674932 241408 674984 241460
rect 675300 241068 675352 241120
rect 511908 240728 511960 240780
rect 629944 240728 629996 240780
rect 42248 240048 42300 240100
rect 45192 240048 45244 240100
rect 514024 238144 514076 238196
rect 568764 238144 568816 238196
rect 674840 238076 674892 238128
rect 675300 238076 675352 238128
rect 512644 238008 512696 238060
rect 633440 238008 633492 238060
rect 42340 235900 42392 235952
rect 44364 235900 44416 235952
rect 42340 234540 42392 234592
rect 44548 234540 44600 234592
rect 510896 233996 510948 234048
rect 577504 233996 577556 234048
rect 511080 233860 511132 233912
rect 631324 233860 631376 233912
rect 42340 232024 42392 232076
rect 45836 232024 45888 232076
rect 157340 231888 157392 231940
rect 164884 231888 164936 231940
rect 190460 231888 190512 231940
rect 191380 231888 191432 231940
rect 42340 231752 42392 231804
rect 43628 231752 43680 231804
rect 54484 231752 54536 231804
rect 641904 231752 641956 231804
rect 53104 231616 53156 231668
rect 641720 231616 641772 231668
rect 46204 231480 46256 231532
rect 643100 231480 643152 231532
rect 47584 231344 47636 231396
rect 645860 231344 645912 231396
rect 51724 231208 51776 231260
rect 650368 231208 650420 231260
rect 44824 231072 44876 231124
rect 644480 231072 644532 231124
rect 129188 230936 129240 230988
rect 661316 230936 661368 230988
rect 120724 230868 120776 230920
rect 123300 230868 123352 230920
rect 99288 230732 99340 230784
rect 176016 230732 176068 230784
rect 176476 230732 176528 230784
rect 176752 230800 176804 230852
rect 178316 230800 178368 230852
rect 185032 230800 185084 230852
rect 475200 230732 475252 230784
rect 479984 230732 480036 230784
rect 481272 230732 481324 230784
rect 489828 230732 489880 230784
rect 113088 230596 113140 230648
rect 186688 230596 186740 230648
rect 194784 230596 194836 230648
rect 195980 230596 196032 230648
rect 450544 230596 450596 230648
rect 510620 230596 510672 230648
rect 123300 230460 123352 230512
rect 147128 230460 147180 230512
rect 42156 230392 42208 230444
rect 43076 230392 43128 230444
rect 107568 230392 107620 230444
rect 42340 230256 42392 230308
rect 43260 230256 43312 230308
rect 90364 230256 90416 230308
rect 117872 230392 117924 230444
rect 123116 230392 123168 230444
rect 206008 230460 206060 230512
rect 147496 230324 147548 230376
rect 213552 230392 213604 230444
rect 253480 230392 253532 230444
rect 339592 230392 339644 230444
rect 341064 230392 341116 230444
rect 407212 230392 407264 230444
rect 412824 230392 412876 230444
rect 421288 230392 421340 230444
rect 422208 230392 422260 230444
rect 427912 230392 427964 230444
rect 429016 230392 429068 230444
rect 429200 230392 429252 230444
rect 441896 230460 441948 230512
rect 442816 230460 442868 230512
rect 451096 230460 451148 230512
rect 512736 230460 512788 230512
rect 450728 230392 450780 230444
rect 159548 230324 159600 230376
rect 167184 230324 167236 230376
rect 167828 230324 167880 230376
rect 171600 230324 171652 230376
rect 200672 230324 200724 230376
rect 147036 230256 147088 230308
rect 149336 230256 149388 230308
rect 156328 230256 156380 230308
rect 171784 230256 171836 230308
rect 200488 230256 200540 230308
rect 204168 230324 204220 230376
rect 205456 230324 205508 230376
rect 205732 230324 205784 230376
rect 207664 230324 207716 230376
rect 298744 230324 298796 230376
rect 299848 230324 299900 230376
rect 313464 230324 313516 230376
rect 313924 230324 313976 230376
rect 319444 230324 319496 230376
rect 321376 230324 321428 230376
rect 328828 230324 328880 230376
rect 329656 230324 329708 230376
rect 331864 230324 331916 230376
rect 333060 230324 333112 230376
rect 333520 230324 333572 230376
rect 334532 230324 334584 230376
rect 335728 230324 335780 230376
rect 337200 230324 337252 230376
rect 337384 230324 337436 230376
rect 338304 230324 338356 230376
rect 342352 230324 342404 230376
rect 343272 230324 343324 230376
rect 344008 230324 344060 230376
rect 344928 230324 344980 230376
rect 348976 230324 349028 230376
rect 352564 230324 352616 230376
rect 356152 230324 356204 230376
rect 357256 230324 357308 230376
rect 360568 230324 360620 230376
rect 362684 230324 362736 230376
rect 364432 230324 364484 230376
rect 365444 230324 365496 230376
rect 367192 230324 367244 230376
rect 368296 230324 368348 230376
rect 368848 230324 368900 230376
rect 369768 230324 369820 230376
rect 371056 230324 371108 230376
rect 372068 230324 372120 230376
rect 378232 230324 378284 230376
rect 379336 230324 379388 230376
rect 385408 230324 385460 230376
rect 386328 230324 386380 230376
rect 387064 230324 387116 230376
rect 388444 230324 388496 230376
rect 403072 230324 403124 230376
rect 404268 230324 404320 230376
rect 405832 230324 405884 230376
rect 407028 230324 407080 230376
rect 413560 230324 413612 230376
rect 418804 230324 418856 230376
rect 441712 230324 441764 230376
rect 442908 230324 442960 230376
rect 443368 230324 443420 230376
rect 444196 230324 444248 230376
rect 208032 230256 208084 230308
rect 240232 230256 240284 230308
rect 244924 230256 244976 230308
rect 246856 230256 246908 230308
rect 255964 230256 256016 230308
rect 279976 230256 280028 230308
rect 285312 230256 285364 230308
rect 291016 230256 291068 230308
rect 339040 230256 339092 230308
rect 339868 230256 339920 230308
rect 390376 230256 390428 230308
rect 399392 230256 399444 230308
rect 122932 230120 122984 230172
rect 123116 230120 123168 230172
rect 204904 230188 204956 230240
rect 186136 230120 186188 230172
rect 186274 230120 186326 230172
rect 187792 230120 187844 230172
rect 189908 230120 189960 230172
rect 83464 229984 83516 230036
rect 157294 229984 157346 230036
rect 162124 229984 162176 230036
rect 171784 229984 171836 230036
rect 171968 229984 172020 230036
rect 174544 229984 174596 230036
rect 174912 229984 174964 230036
rect 176384 229984 176436 230036
rect 176568 229984 176620 230036
rect 190368 229984 190420 230036
rect 191380 230120 191432 230172
rect 194416 230120 194468 230172
rect 194600 230120 194652 230172
rect 198832 230120 198884 230172
rect 199200 230120 199252 230172
rect 203248 230120 203300 230172
rect 205548 230120 205600 230172
rect 244648 230120 244700 230172
rect 247776 230120 247828 230172
rect 275560 230120 275612 230172
rect 279792 230120 279844 230172
rect 297640 230188 297692 230240
rect 313924 230188 313976 230240
rect 315304 230188 315356 230240
rect 341248 230188 341300 230240
rect 343824 230188 343876 230240
rect 355048 230188 355100 230240
rect 360844 230188 360896 230240
rect 378784 230188 378836 230240
rect 380164 230188 380216 230240
rect 380992 230188 381044 230240
rect 389732 230188 389784 230240
rect 404728 230188 404780 230240
rect 413284 230256 413336 230308
rect 420184 230256 420236 230308
rect 434904 230256 434956 230308
rect 435088 230256 435140 230308
rect 436008 230256 436060 230308
rect 446128 230256 446180 230308
rect 505744 230256 505796 230308
rect 344560 230120 344612 230172
rect 349804 230120 349856 230172
rect 369400 230120 369452 230172
rect 371884 230120 371936 230172
rect 372712 230120 372764 230172
rect 297364 230052 297416 230104
rect 299296 230052 299348 230104
rect 320824 230052 320876 230104
rect 321928 230052 321980 230104
rect 340696 230052 340748 230104
rect 344284 230052 344336 230104
rect 357440 230052 357492 230104
rect 363604 230052 363656 230104
rect 196624 229984 196676 230036
rect 196808 229984 196860 230036
rect 235816 229984 235868 230036
rect 241612 229984 241664 230036
rect 271144 229984 271196 230036
rect 275652 229984 275704 230036
rect 293224 229984 293276 230036
rect 367744 229984 367796 230036
rect 370872 229984 370924 230036
rect 77944 229848 77996 229900
rect 133052 229848 133104 229900
rect 133236 229848 133288 229900
rect 182824 229848 182876 229900
rect 183468 229848 183520 229900
rect 231400 229848 231452 229900
rect 233240 229848 233292 229900
rect 266728 229848 266780 229900
rect 267004 229848 267056 229900
rect 288808 229848 288860 229900
rect 338488 229848 338540 229900
rect 339316 229848 339368 229900
rect 359464 229848 359516 229900
rect 369124 229848 369176 229900
rect 374368 229984 374420 230036
rect 377404 229984 377456 230036
rect 379152 229984 379204 230036
rect 392216 230120 392268 230172
rect 392400 230120 392452 230172
rect 394976 230120 395028 230172
rect 411352 230120 411404 230172
rect 414848 230120 414900 230172
rect 415216 230120 415268 230172
rect 441712 230120 441764 230172
rect 441896 230120 441948 230172
rect 447508 230120 447560 230172
rect 455512 230120 455564 230172
rect 456708 230120 456760 230172
rect 457168 230120 457220 230172
rect 458088 230120 458140 230172
rect 458456 230120 458508 230172
rect 475200 230120 475252 230172
rect 476488 230120 476540 230172
rect 479524 230120 479576 230172
rect 479984 230120 480036 230172
rect 481364 230120 481416 230172
rect 482560 230120 482612 230172
rect 541992 230120 542044 230172
rect 392032 229984 392084 230036
rect 396724 229984 396776 230036
rect 398748 229984 398800 230036
rect 382280 229848 382332 229900
rect 300584 229780 300636 229832
rect 301504 229780 301556 229832
rect 67548 229712 67600 229764
rect 149336 229712 149388 229764
rect 150992 229712 151044 229764
rect 154120 229712 154172 229764
rect 154580 229712 154632 229764
rect 157984 229712 158036 229764
rect 158168 229712 158220 229764
rect 160744 229712 160796 229764
rect 161112 229712 161164 229764
rect 163504 229712 163556 229764
rect 163964 229712 164016 229764
rect 171784 229712 171836 229764
rect 171968 229712 172020 229764
rect 218152 229712 218204 229764
rect 220544 229712 220596 229764
rect 257896 229712 257948 229764
rect 261576 229712 261628 229764
rect 284392 229712 284444 229764
rect 289728 229712 289780 229764
rect 305644 229712 305696 229764
rect 313096 229712 313148 229764
rect 342904 229712 342956 229764
rect 348424 229712 348476 229764
rect 361672 229712 361724 229764
rect 374000 229712 374052 229764
rect 377128 229712 377180 229764
rect 391204 229848 391256 229900
rect 391480 229848 391532 229900
rect 392584 229848 392636 229900
rect 400864 229848 400916 229900
rect 414112 229984 414164 230036
rect 415308 229984 415360 230036
rect 416320 229984 416372 230036
rect 304264 229644 304316 229696
rect 122932 229576 122984 229628
rect 132868 229576 132920 229628
rect 130108 229440 130160 229492
rect 133236 229440 133288 229492
rect 126888 229304 126940 229356
rect 194784 229576 194836 229628
rect 195244 229576 195296 229628
rect 200488 229576 200540 229628
rect 201224 229576 201276 229628
rect 226984 229576 227036 229628
rect 230664 229576 230716 229628
rect 262312 229576 262364 229628
rect 313188 229576 313240 229628
rect 319720 229576 319772 229628
rect 374920 229576 374972 229628
rect 391664 229712 391716 229764
rect 392952 229712 393004 229764
rect 399576 229712 399628 229764
rect 416044 229848 416096 229900
rect 419080 229848 419132 229900
rect 424048 229984 424100 230036
rect 429200 229984 429252 230036
rect 429384 229984 429436 230036
rect 446772 229984 446824 230036
rect 448152 229984 448204 230036
rect 507124 229984 507176 230036
rect 420184 229712 420236 229764
rect 427084 229848 427136 229900
rect 428464 229848 428516 229900
rect 473452 229848 473504 229900
rect 475200 229848 475252 229900
rect 484032 229848 484084 229900
rect 484216 229848 484268 229900
rect 487344 229848 487396 229900
rect 487528 229848 487580 229900
rect 428096 229712 428148 229764
rect 438952 229712 439004 229764
rect 484860 229712 484912 229764
rect 485044 229712 485096 229764
rect 495394 229712 495446 229764
rect 499488 229848 499540 229900
rect 551928 229848 551980 229900
rect 558184 229712 558236 229764
rect 389272 229576 389324 229628
rect 390468 229576 390520 229628
rect 394240 229576 394292 229628
rect 400864 229576 400916 229628
rect 407488 229576 407540 229628
rect 424324 229576 424376 229628
rect 425704 229576 425756 229628
rect 133052 229168 133104 229220
rect 133696 229304 133748 229356
rect 152556 229304 152608 229356
rect 153016 229440 153068 229492
rect 162124 229440 162176 229492
rect 163596 229440 163648 229492
rect 165712 229440 165764 229492
rect 167000 229440 167052 229492
rect 171600 229440 171652 229492
rect 171784 229440 171836 229492
rect 200672 229440 200724 229492
rect 200856 229440 200908 229492
rect 208032 229440 208084 229492
rect 208216 229440 208268 229492
rect 209320 229440 209372 229492
rect 211160 229440 211212 229492
rect 220912 229440 220964 229492
rect 225972 229440 226024 229492
rect 229744 229440 229796 229492
rect 156328 229304 156380 229356
rect 156880 229304 156932 229356
rect 200074 229304 200126 229356
rect 200488 229304 200540 229356
rect 213736 229304 213788 229356
rect 220820 229304 220872 229356
rect 225328 229304 225380 229356
rect 226984 229304 227036 229356
rect 236368 229304 236420 229356
rect 133880 229168 133932 229220
rect 147312 229168 147364 229220
rect 147680 229168 147732 229220
rect 157294 229168 157346 229220
rect 157616 229168 157668 229220
rect 195244 229168 195296 229220
rect 196532 229168 196584 229220
rect 201040 229168 201092 229220
rect 201408 229168 201460 229220
rect 208216 229168 208268 229220
rect 208400 229168 208452 229220
rect 216496 229168 216548 229220
rect 222936 229168 222988 229220
rect 249064 229440 249116 229492
rect 385960 229440 386012 229492
rect 392400 229440 392452 229492
rect 397000 229440 397052 229492
rect 290464 229372 290516 229424
rect 295432 229372 295484 229424
rect 372528 229372 372580 229424
rect 374552 229372 374604 229424
rect 405280 229440 405332 229492
rect 428464 229440 428516 229492
rect 428832 229576 428884 229628
rect 441896 229576 441948 229628
rect 444472 229576 444524 229628
rect 495440 229576 495492 229628
rect 429752 229440 429804 229492
rect 434904 229440 434956 229492
rect 439504 229440 439556 229492
rect 441712 229440 441764 229492
rect 450544 229440 450596 229492
rect 450728 229440 450780 229492
rect 499120 229644 499172 229696
rect 499856 229576 499908 229628
rect 495900 229440 495952 229492
rect 499488 229440 499540 229492
rect 499672 229440 499724 229492
rect 502524 229440 502576 229492
rect 502984 229576 503036 229628
rect 511264 229576 511316 229628
rect 504180 229440 504232 229492
rect 504364 229440 504416 229492
rect 507492 229440 507544 229492
rect 404636 229372 404688 229424
rect 396448 229304 396500 229356
rect 397368 229304 397420 229356
rect 412824 229304 412876 229356
rect 421564 229304 421616 229356
rect 421840 229304 421892 229356
rect 451188 229304 451240 229356
rect 453304 229304 453356 229356
rect 455880 229304 455932 229356
rect 456064 229304 456116 229356
rect 458456 229304 458508 229356
rect 458824 229304 458876 229356
rect 480168 229304 480220 229356
rect 480536 229304 480588 229356
rect 481732 229304 481784 229356
rect 484860 229304 484912 229356
rect 489552 229304 489604 229356
rect 334072 229236 334124 229288
rect 335728 229236 335780 229288
rect 350632 229236 350684 229288
rect 355324 229236 355376 229288
rect 390192 229236 390244 229288
rect 393964 229236 394016 229288
rect 399208 229236 399260 229288
rect 405004 229236 405056 229288
rect 422944 229168 422996 229220
rect 429384 229168 429436 229220
rect 429752 229168 429804 229220
rect 446956 229168 447008 229220
rect 448336 229168 448388 229220
rect 463700 229168 463752 229220
rect 464160 229168 464212 229220
rect 466368 229168 466420 229220
rect 466552 229168 466604 229220
rect 470784 229168 470836 229220
rect 473452 229168 473504 229220
rect 476396 229168 476448 229220
rect 479248 229168 479300 229220
rect 485044 229168 485096 229220
rect 485872 229168 485924 229220
rect 490012 229304 490064 229356
rect 490196 229304 490248 229356
rect 536840 229304 536892 229356
rect 489920 229168 489972 229220
rect 533344 229168 533396 229220
rect 304080 229100 304132 229152
rect 308680 229100 308732 229152
rect 322756 229100 322808 229152
rect 326344 229100 326396 229152
rect 335176 229100 335228 229152
rect 335912 229100 335964 229152
rect 87604 229032 87656 229084
rect 147496 229032 147548 229084
rect 147634 229032 147686 229084
rect 152464 229032 152516 229084
rect 152924 229032 152976 229084
rect 185860 229032 185912 229084
rect 188988 229032 189040 229084
rect 195244 229032 195296 229084
rect 195704 229032 195756 229084
rect 119988 228896 120040 228948
rect 189724 228896 189776 228948
rect 194232 228896 194284 228948
rect 196808 228896 196860 228948
rect 198648 229032 198700 229084
rect 201224 229032 201276 229084
rect 212264 229032 212316 229084
rect 251824 229032 251876 229084
rect 262036 229032 262088 229084
rect 284944 229032 284996 229084
rect 361120 229032 361172 229084
rect 373540 229032 373592 229084
rect 382280 229032 382332 229084
rect 202420 228896 202472 228948
rect 202604 228896 202656 228948
rect 245200 228896 245252 228948
rect 245476 228896 245528 228948
rect 273904 228896 273956 228948
rect 286692 228896 286744 228948
rect 300952 228896 301004 228948
rect 373264 228896 373316 228948
rect 388444 228896 388496 228948
rect 391204 229032 391256 229084
rect 397736 229032 397788 229084
rect 407764 229032 407816 229084
rect 429936 229032 429988 229084
rect 430120 229032 430172 229084
rect 457444 229032 457496 229084
rect 459928 229032 459980 229084
rect 525984 229032 526036 229084
rect 391848 228896 391900 228948
rect 110328 228760 110380 228812
rect 183100 228760 183152 228812
rect 183284 228760 183336 228812
rect 225972 228760 226024 228812
rect 238576 228760 238628 228812
rect 269488 228760 269540 228812
rect 275836 228760 275888 228812
rect 293776 228760 293828 228812
rect 295156 228760 295208 228812
rect 307024 228760 307076 228812
rect 352840 228760 352892 228812
rect 361028 228760 361080 228812
rect 362224 228760 362276 228812
rect 376760 228760 376812 228812
rect 377680 228760 377732 228812
rect 400680 228896 400732 228948
rect 401968 228896 402020 228948
rect 437112 228896 437164 228948
rect 439504 228896 439556 228948
rect 465264 228896 465316 228948
rect 477592 228896 477644 228948
rect 495394 228896 495446 228948
rect 495992 228896 496044 228948
rect 507952 228896 508004 228948
rect 508136 228896 508188 228948
rect 552204 228896 552256 228948
rect 397552 228760 397604 228812
rect 407764 228760 407816 228812
rect 423496 228760 423548 228812
rect 468024 228760 468076 228812
rect 468208 228760 468260 228812
rect 538404 228760 538456 228812
rect 85488 228624 85540 228676
rect 100668 228488 100720 228540
rect 166908 228488 166960 228540
rect 167828 228624 167880 228676
rect 171968 228624 172020 228676
rect 172428 228624 172480 228676
rect 213828 228624 213880 228676
rect 169024 228488 169076 228540
rect 171600 228488 171652 228540
rect 193036 228488 193088 228540
rect 195244 228488 195296 228540
rect 226984 228624 227036 228676
rect 231676 228624 231728 228676
rect 266176 228624 266228 228676
rect 266360 228624 266412 228676
rect 287152 228624 287204 228676
rect 292488 228624 292540 228676
rect 304816 228624 304868 228676
rect 315672 228624 315724 228676
rect 320272 228624 320324 228676
rect 349528 228624 349580 228676
rect 359464 228624 359516 228676
rect 370504 228624 370556 228676
rect 387064 228624 387116 228676
rect 393136 228624 393188 228676
rect 424048 228624 424100 228676
rect 426808 228624 426860 228676
rect 475200 228624 475252 228676
rect 475384 228624 475436 228676
rect 495624 228624 495676 228676
rect 495808 228624 495860 228676
rect 214748 228488 214800 228540
rect 248512 228488 248564 228540
rect 253572 228488 253624 228540
rect 278872 228488 278924 228540
rect 285588 228488 285640 228540
rect 300400 228488 300452 228540
rect 300768 228488 300820 228540
rect 309784 228488 309836 228540
rect 325608 228488 325660 228540
rect 328368 228488 328420 228540
rect 353392 228488 353444 228540
rect 364432 228488 364484 228540
rect 364984 228488 365036 228540
rect 376392 228488 376444 228540
rect 376760 228488 376812 228540
rect 377680 228488 377732 228540
rect 386512 228488 386564 228540
rect 414204 228488 414256 228540
rect 414848 228488 414900 228540
rect 451464 228488 451516 228540
rect 451648 228488 451700 228540
rect 505054 228488 505106 228540
rect 505192 228488 505244 228540
rect 507492 228488 507544 228540
rect 507952 228624 508004 228676
rect 548340 228624 548392 228676
rect 548524 228488 548576 228540
rect 49148 228352 49200 228404
rect 653220 228352 653272 228404
rect 96436 228216 96488 228268
rect 69572 228080 69624 228132
rect 147956 228080 148008 228132
rect 149244 228080 149296 228132
rect 151360 228080 151412 228132
rect 152464 228216 152516 228268
rect 171600 228216 171652 228268
rect 159824 228080 159876 228132
rect 160008 228080 160060 228132
rect 208400 228216 208452 228268
rect 213828 228216 213880 228268
rect 220820 228216 220872 228268
rect 222016 228216 222068 228268
rect 258448 228216 258500 228268
rect 376392 228216 376444 228268
rect 382648 228216 382700 228268
rect 388444 228216 388496 228268
rect 394240 228216 394292 228268
rect 400312 228216 400364 228268
rect 432604 228216 432656 228268
rect 434536 228216 434588 228268
rect 442448 228216 442500 228268
rect 446772 228216 446824 228268
rect 466184 228216 466236 228268
rect 466368 228216 466420 228268
rect 531688 228216 531740 228268
rect 171968 228080 172020 228132
rect 211160 228080 211212 228132
rect 456524 228080 456576 228132
rect 520924 228080 520976 228132
rect 133512 227944 133564 227996
rect 147496 227944 147548 227996
rect 147680 227944 147732 227996
rect 204168 227944 204220 227996
rect 205272 227944 205324 227996
rect 214748 227944 214800 227996
rect 454960 227944 455012 227996
rect 517796 227944 517848 227996
rect 310336 227876 310388 227928
rect 316408 227876 316460 227928
rect 136548 227808 136600 227860
rect 196532 227808 196584 227860
rect 201040 227808 201092 227860
rect 222568 227808 222620 227860
rect 226248 227808 226300 227860
rect 230664 227808 230716 227860
rect 236644 227808 236696 227860
rect 238024 227808 238076 227860
rect 240048 227808 240100 227860
rect 241612 227808 241664 227860
rect 259276 227808 259328 227860
rect 261576 227808 261628 227860
rect 436744 227808 436796 227860
rect 249064 227740 249116 227792
rect 251272 227740 251324 227792
rect 251732 227740 251784 227792
rect 255688 227740 255740 227792
rect 308772 227740 308824 227792
rect 315488 227740 315540 227792
rect 317052 227740 317104 227792
rect 320548 227740 320600 227792
rect 321468 227740 321520 227792
rect 324688 227740 324740 227792
rect 345112 227740 345164 227792
rect 352840 227740 352892 227792
rect 394792 227740 394844 227792
rect 402244 227740 402296 227792
rect 111708 227672 111760 227724
rect 183928 227672 183980 227724
rect 196624 227672 196676 227724
rect 207112 227672 207164 227724
rect 209596 227672 209648 227724
rect 249616 227604 249668 227656
rect 251088 227604 251140 227656
rect 276664 227672 276716 227724
rect 429568 227672 429620 227724
rect 476212 227672 476264 227724
rect 481364 227808 481416 227860
rect 489874 227808 489926 227860
rect 487620 227672 487672 227724
rect 489552 227672 489604 227724
rect 630680 227740 630732 227792
rect 93768 227536 93820 227588
rect 173992 227536 174044 227588
rect 184204 227536 184256 227588
rect 198280 227536 198332 227588
rect 199476 227536 199528 227588
rect 205548 227536 205600 227588
rect 205916 227536 205968 227588
rect 247408 227536 247460 227588
rect 256516 227536 256568 227588
rect 276112 227536 276164 227588
rect 395344 227536 395396 227588
rect 427360 227536 427412 227588
rect 461584 227536 461636 227588
rect 527824 227536 527876 227588
rect 68928 227400 68980 227452
rect 154580 227400 154632 227452
rect 155684 227400 155736 227452
rect 73712 227264 73764 227316
rect 160192 227264 160244 227316
rect 166724 227400 166776 227452
rect 167828 227400 167880 227452
rect 176568 227400 176620 227452
rect 182824 227400 182876 227452
rect 233056 227400 233108 227452
rect 234436 227400 234488 227452
rect 268292 227400 268344 227452
rect 374552 227400 374604 227452
rect 390100 227400 390152 227452
rect 392216 227400 392268 227452
rect 401692 227400 401744 227452
rect 404084 227400 404136 227452
rect 440608 227400 440660 227452
rect 446956 227400 447008 227452
rect 471244 227400 471296 227452
rect 473728 227400 473780 227452
rect 546592 227400 546644 227452
rect 66168 227128 66220 227180
rect 149520 227128 149572 227180
rect 63408 226992 63460 227044
rect 151728 227128 151780 227180
rect 156696 227128 156748 227180
rect 163964 227128 164016 227180
rect 227536 227264 227588 227316
rect 228824 227264 228876 227316
rect 262864 227264 262916 227316
rect 272432 227264 272484 227316
rect 282184 227264 282236 227316
rect 293776 227264 293828 227316
rect 305368 227264 305420 227316
rect 376576 227264 376628 227316
rect 396724 227264 396776 227316
rect 417976 227264 418028 227316
rect 462136 227264 462188 227316
rect 471520 227264 471572 227316
rect 543464 227264 543516 227316
rect 214288 227128 214340 227180
rect 215208 227128 215260 227180
rect 255136 227128 255188 227180
rect 277216 227128 277268 227180
rect 294328 227128 294380 227180
rect 363880 227128 363932 227180
rect 374644 227128 374696 227180
rect 384304 227128 384356 227180
rect 410616 227128 410668 227180
rect 424600 227128 424652 227180
rect 472164 227128 472216 227180
rect 474280 227128 474332 227180
rect 547512 227128 547564 227180
rect 149888 226992 149940 227044
rect 117228 226856 117280 226908
rect 184848 226856 184900 226908
rect 205456 226992 205508 227044
rect 205916 226992 205968 227044
rect 210976 226992 211028 227044
rect 250168 226992 250220 227044
rect 256148 226992 256200 227044
rect 281632 226992 281684 227044
rect 282736 226992 282788 227044
rect 298192 226992 298244 227044
rect 304632 226992 304684 227044
rect 314752 226992 314804 227044
rect 351736 226992 351788 227044
rect 361580 226992 361632 227044
rect 366640 226992 366692 227044
rect 384304 226992 384356 227044
rect 388168 226992 388220 227044
rect 414940 226992 414992 227044
rect 426256 226992 426308 227044
rect 473728 226992 473780 227044
rect 479800 226992 479852 227044
rect 555700 226992 555752 227044
rect 210700 226856 210752 226908
rect 249616 226856 249668 226908
rect 256516 226856 256568 226908
rect 470784 226856 470836 226908
rect 535920 226856 535972 226908
rect 146116 226720 146168 226772
rect 205732 226720 205784 226772
rect 458640 226720 458692 226772
rect 523500 226720 523552 226772
rect 129556 226584 129608 226636
rect 189908 226584 189960 226636
rect 441896 226584 441948 226636
rect 477592 226584 477644 226636
rect 481732 226584 481784 226636
rect 515956 226584 516008 226636
rect 139308 226448 139360 226500
rect 199292 226448 199344 226500
rect 391664 226380 391716 226432
rect 395068 226380 395120 226432
rect 484032 226380 484084 226432
rect 206100 226312 206152 226364
rect 211528 226312 211580 226364
rect 64788 226244 64840 226296
rect 125692 226244 125744 226296
rect 125876 226244 125928 226296
rect 118608 226108 118660 226160
rect 129372 226244 129424 226296
rect 122748 225972 122800 226024
rect 125876 225972 125928 226024
rect 137100 226108 137152 226160
rect 137468 226244 137520 226296
rect 147956 226244 148008 226296
rect 148508 226108 148560 226160
rect 156512 226108 156564 226160
rect 157294 226244 157346 226296
rect 202144 226244 202196 226296
rect 214380 226244 214432 226296
rect 245752 226244 245804 226296
rect 393688 226244 393740 226296
rect 425704 226244 425756 226296
rect 428096 226244 428148 226296
rect 461308 226244 461360 226296
rect 462688 226244 462740 226296
rect 489874 226244 489926 226296
rect 509608 226380 509660 226432
rect 510160 226380 510212 226432
rect 197728 226108 197780 226160
rect 197912 226108 197964 226160
rect 181996 225972 182048 226024
rect 193312 225972 193364 226024
rect 193680 225972 193732 226024
rect 195704 225972 195756 226024
rect 195888 225972 195940 226024
rect 199292 225972 199344 226024
rect 200120 226108 200172 226160
rect 242992 226108 243044 226160
rect 270132 226108 270184 226160
rect 289912 226108 289964 226160
rect 382096 226108 382148 226160
rect 407488 226108 407540 226160
rect 415768 226108 415820 226160
rect 449164 226108 449216 226160
rect 453856 226108 453908 226160
rect 514576 226244 514628 226296
rect 530584 226244 530636 226296
rect 533344 226244 533396 226296
rect 556712 226244 556764 226296
rect 238300 225972 238352 226024
rect 246856 225972 246908 226024
rect 274456 225972 274508 226024
rect 399760 225972 399812 226024
rect 433984 225972 434036 226024
rect 436560 225972 436612 226024
rect 467288 225972 467340 226024
rect 469312 225972 469364 226024
rect 489874 225972 489926 226024
rect 490012 225972 490064 226024
rect 505054 225972 505106 226024
rect 505192 225972 505244 226024
rect 509608 225972 509660 226024
rect 518900 226108 518952 226160
rect 536840 226108 536892 226160
rect 561772 226108 561824 226160
rect 514576 225972 514628 226024
rect 514714 225972 514766 226024
rect 540244 225972 540296 226024
rect 57888 225836 57940 225888
rect 107568 225836 107620 225888
rect 115296 225836 115348 225888
rect 190184 225836 190236 225888
rect 190368 225836 190420 225888
rect 204536 225836 204588 225888
rect 204720 225836 204772 225888
rect 214564 225836 214616 225888
rect 244188 225836 244240 225888
rect 272248 225836 272300 225888
rect 390928 225836 390980 225888
rect 419724 225836 419776 225888
rect 422392 225836 422444 225888
rect 458640 225836 458692 225888
rect 467656 225836 467708 225888
rect 536840 225836 536892 225888
rect 93584 225700 93636 225752
rect 166356 225700 166408 225752
rect 181260 225700 181312 225752
rect 188620 225700 188672 225752
rect 190414 225700 190466 225752
rect 234160 225700 234212 225752
rect 235908 225700 235960 225752
rect 267280 225700 267332 225752
rect 267648 225700 267700 225752
rect 290188 225700 290240 225752
rect 291016 225700 291068 225752
rect 303160 225700 303212 225752
rect 363328 225700 363380 225752
rect 376852 225700 376904 225752
rect 402520 225700 402572 225752
rect 439044 225700 439096 225752
rect 447508 225700 447560 225752
rect 469312 225700 469364 225752
rect 472624 225700 472676 225752
rect 543740 225700 543792 225752
rect 75736 225564 75788 225616
rect 147772 225564 147824 225616
rect 147956 225564 148008 225616
rect 156972 225564 157024 225616
rect 157156 225564 157208 225616
rect 157294 225564 157346 225616
rect 157432 225564 157484 225616
rect 169024 225564 169076 225616
rect 214196 225564 214248 225616
rect 214564 225564 214616 225616
rect 240784 225564 240836 225616
rect 241152 225564 241204 225616
rect 272800 225564 272852 225616
rect 274548 225564 274600 225616
rect 292120 225564 292172 225616
rect 294972 225564 295024 225616
rect 308128 225564 308180 225616
rect 308956 225564 309008 225616
rect 317512 225564 317564 225616
rect 359280 225564 359332 225616
rect 370228 225564 370280 225616
rect 371608 225564 371660 225616
rect 392584 225564 392636 225616
rect 438400 225564 438452 225616
rect 472624 225564 472676 225616
rect 475936 225564 475988 225616
rect 504732 225564 504784 225616
rect 505192 225564 505244 225616
rect 549904 225564 549956 225616
rect 125232 225428 125284 225480
rect 195520 225428 195572 225480
rect 195704 225428 195756 225480
rect 197728 225428 197780 225480
rect 197912 225428 197964 225480
rect 204720 225428 204772 225480
rect 204904 225428 204956 225480
rect 241888 225428 241940 225480
rect 432880 225428 432932 225480
rect 464528 225428 464580 225480
rect 464712 225428 464764 225480
rect 531964 225428 532016 225480
rect 125692 225292 125744 225344
rect 133880 225292 133932 225344
rect 137100 225292 137152 225344
rect 141608 225292 141660 225344
rect 141792 225292 141844 225344
rect 206560 225292 206612 225344
rect 208032 225292 208084 225344
rect 250720 225292 250772 225344
rect 418528 225292 418580 225344
rect 446404 225292 446456 225344
rect 459376 225292 459428 225344
rect 525064 225292 525116 225344
rect 107568 225156 107620 225208
rect 130108 225156 130160 225208
rect 132408 225156 132460 225208
rect 199660 225156 199712 225208
rect 199844 225156 199896 225208
rect 204904 225156 204956 225208
rect 205088 225156 205140 225208
rect 214380 225156 214432 225208
rect 217324 225156 217376 225208
rect 229192 225156 229244 225208
rect 406384 225156 406436 225208
rect 443920 225156 443972 225208
rect 461124 225156 461176 225208
rect 528468 225156 528520 225208
rect 116952 225020 117004 225072
rect 117872 225020 117924 225072
rect 135076 225020 135128 225072
rect 137468 225020 137520 225072
rect 139124 225020 139176 225072
rect 204352 225020 204404 225072
rect 204536 225020 204588 225072
rect 212080 225020 212132 225072
rect 214196 225020 214248 225072
rect 218704 225020 218756 225072
rect 466000 225020 466052 225072
rect 535000 225020 535052 225072
rect 273168 224952 273220 225004
rect 275652 224952 275704 225004
rect 42432 224884 42484 224936
rect 47124 224884 47176 224936
rect 96252 224884 96304 224936
rect 171600 224884 171652 224936
rect 106188 224748 106240 224800
rect 182272 224884 182324 224936
rect 185400 224884 185452 224936
rect 171968 224748 172020 224800
rect 173440 224748 173492 224800
rect 175096 224748 175148 224800
rect 185584 224748 185636 224800
rect 191472 224884 191524 224936
rect 239680 224884 239732 224936
rect 420000 224884 420052 224936
rect 454868 224884 454920 224936
rect 470968 224884 471020 224936
rect 542360 224884 542412 224936
rect 543740 224884 543792 224936
rect 545028 224884 545080 224936
rect 553400 225020 553452 225072
rect 552756 224884 552808 224936
rect 559012 224884 559064 224936
rect 194784 224748 194836 224800
rect 195244 224748 195296 224800
rect 237472 224748 237524 224800
rect 255228 224748 255280 224800
rect 280528 224748 280580 224800
rect 408592 224748 408644 224800
rect 447232 224748 447284 224800
rect 480352 224748 480404 224800
rect 483664 224748 483716 224800
rect 485872 224748 485924 224800
rect 85304 224612 85356 224664
rect 165988 224612 166040 224664
rect 166264 224612 166316 224664
rect 221648 224612 221700 224664
rect 89628 224476 89680 224528
rect 171232 224476 171284 224528
rect 171600 224476 171652 224528
rect 175648 224476 175700 224528
rect 82728 224340 82780 224392
rect 166540 224340 166592 224392
rect 168196 224340 168248 224392
rect 171968 224340 172020 224392
rect 173256 224340 173308 224392
rect 185400 224476 185452 224528
rect 185584 224476 185636 224528
rect 221280 224476 221332 224528
rect 221464 224476 221516 224528
rect 257344 224612 257396 224664
rect 379888 224612 379940 224664
rect 402980 224612 403032 224664
rect 413008 224612 413060 224664
rect 453856 224612 453908 224664
rect 457720 224612 457772 224664
rect 486240 224748 486292 224800
rect 556528 224748 556580 224800
rect 556712 224748 556764 224800
rect 557356 224748 557408 224800
rect 557816 224748 557868 224800
rect 561496 224748 561548 224800
rect 250904 224476 250956 224528
rect 279424 224476 279476 224528
rect 279976 224476 280028 224528
rect 296536 224476 296588 224528
rect 370872 224476 370924 224528
rect 383476 224476 383528 224528
rect 387616 224476 387668 224528
rect 413284 224476 413336 224528
rect 414664 224476 414716 224528
rect 425888 224476 425940 224528
rect 434168 224476 434220 224528
rect 481824 224476 481876 224528
rect 482008 224476 482060 224528
rect 484860 224476 484912 224528
rect 552756 224612 552808 224664
rect 552940 224612 552992 224664
rect 487988 224476 488040 224528
rect 491944 224476 491996 224528
rect 557816 224476 557868 224528
rect 558000 224476 558052 224528
rect 566464 224476 566516 224528
rect 176016 224340 176068 224392
rect 224224 224340 224276 224392
rect 226064 224340 226116 224392
rect 260380 224340 260432 224392
rect 57244 224204 57296 224256
rect 142114 224204 142166 224256
rect 142252 224204 142304 224256
rect 156696 224204 156748 224256
rect 156972 224204 157024 224256
rect 158536 224204 158588 224256
rect 158720 224204 158772 224256
rect 217600 224204 217652 224256
rect 224592 224204 224644 224256
rect 261760 224204 261812 224256
rect 262680 224204 262732 224256
rect 264520 224204 264572 224256
rect 101404 224068 101456 224120
rect 168380 224068 168432 224120
rect 168564 224068 168616 224120
rect 172244 224068 172296 224120
rect 172612 224068 172664 224120
rect 92112 223932 92164 223984
rect 173072 223932 173124 223984
rect 173440 224068 173492 224120
rect 176016 224068 176068 224120
rect 176384 224068 176436 224120
rect 193864 224068 193916 224120
rect 194784 224068 194836 224120
rect 198648 224068 198700 224120
rect 216496 224068 216548 224120
rect 254032 224068 254084 224120
rect 260196 224068 260248 224120
rect 283288 224340 283340 224392
rect 296628 224340 296680 224392
rect 304080 224340 304132 224392
rect 358452 224340 358504 224392
rect 372712 224340 372764 224392
rect 383016 224340 383068 224392
rect 403440 224340 403492 224392
rect 403624 224340 403676 224392
rect 405372 224340 405424 224392
rect 410800 224340 410852 224392
rect 434168 224340 434220 224392
rect 275284 224204 275336 224256
rect 294788 224204 294840 224256
rect 296444 224204 296496 224256
rect 307300 224204 307352 224256
rect 307484 224204 307536 224256
rect 316684 224204 316736 224256
rect 331220 224204 331272 224256
rect 332140 224204 332192 224256
rect 335728 224204 335780 224256
rect 336280 224204 336332 224256
rect 352288 224204 352340 224256
rect 358084 224204 358136 224256
rect 370412 224204 370464 224256
rect 386788 224204 386840 224256
rect 388812 224204 388864 224256
rect 417424 224204 417476 224256
rect 432328 224204 432380 224256
rect 435364 224204 435416 224256
rect 403440 224068 403492 224120
rect 409144 224068 409196 224120
rect 409696 224068 409748 224120
rect 421840 224068 421892 224120
rect 433800 224068 433852 224120
rect 485044 224340 485096 224392
rect 490748 224340 490800 224392
rect 563980 224340 564032 224392
rect 438216 224204 438268 224256
rect 484676 224204 484728 224256
rect 442632 224068 442684 224120
rect 486792 224272 486844 224324
rect 590936 224408 590988 224460
rect 597560 224408 597612 224460
rect 486976 224204 487028 224256
rect 558000 224204 558052 224256
rect 487988 224068 488040 224120
rect 522580 224068 522632 224120
rect 536840 224000 536892 224052
rect 537484 224000 537536 224052
rect 210424 223932 210476 223984
rect 113824 223796 113876 223848
rect 161848 223796 161900 223848
rect 162492 223796 162544 223848
rect 219348 223932 219400 223984
rect 221280 223932 221332 223984
rect 228640 223932 228692 223984
rect 417608 223932 417660 223984
rect 431224 223932 431276 223984
rect 431776 223932 431828 223984
rect 438308 223932 438360 223984
rect 454408 223932 454460 223984
rect 485688 223932 485740 223984
rect 485872 223932 485924 223984
rect 517612 223932 517664 223984
rect 544016 223864 544068 223916
rect 544384 224000 544436 224052
rect 591120 224136 591172 224188
rect 610440 224272 610492 224324
rect 610808 224136 610860 224188
rect 617708 224136 617760 224188
rect 558552 224000 558604 224052
rect 626724 224000 626776 224052
rect 552940 223864 552992 223916
rect 553400 223864 553452 223916
rect 623780 223864 623832 223916
rect 219348 223796 219400 223848
rect 256332 223796 256384 223848
rect 452752 223796 452804 223848
rect 485688 223796 485740 223848
rect 485872 223796 485924 223848
rect 515128 223796 515180 223848
rect 317236 223728 317288 223780
rect 323584 223728 323636 223780
rect 129740 223660 129792 223712
rect 187240 223660 187292 223712
rect 188804 223660 188856 223712
rect 195244 223660 195296 223712
rect 210424 223660 210476 223712
rect 221096 223660 221148 223712
rect 440056 223660 440108 223712
rect 496084 223660 496136 223712
rect 505008 223660 505060 223712
rect 590936 223592 590988 223644
rect 591120 223592 591172 223644
rect 610440 223592 610492 223644
rect 610808 223728 610860 223780
rect 622584 223728 622636 223780
rect 617064 223592 617116 223644
rect 42248 223524 42300 223576
rect 46940 223524 46992 223576
rect 121092 223524 121144 223576
rect 190552 223524 190604 223576
rect 194416 223524 194468 223576
rect 239128 223524 239180 223576
rect 246672 223524 246724 223576
rect 271696 223524 271748 223576
rect 305920 223524 305972 223576
rect 306472 223524 306524 223576
rect 347872 223524 347924 223576
rect 353668 223524 353720 223576
rect 399392 223524 399444 223576
rect 418252 223524 418304 223576
rect 435640 223524 435692 223576
rect 474648 223524 474700 223576
rect 477040 223524 477092 223576
rect 484124 223524 484176 223576
rect 487068 223524 487120 223576
rect 511264 223524 511316 223576
rect 108672 223388 108724 223440
rect 133144 223388 133196 223440
rect 133788 223388 133840 223440
rect 197176 223388 197228 223440
rect 198096 223388 198148 223440
rect 243820 223456 243872 223508
rect 245292 223456 245344 223508
rect 529388 223456 529440 223508
rect 536104 223456 536156 223508
rect 242164 223320 242216 223372
rect 246304 223320 246356 223372
rect 97908 223252 97960 223304
rect 171416 223252 171468 223304
rect 171600 223252 171652 223304
rect 180616 223252 180668 223304
rect 187332 223252 187384 223304
rect 234712 223252 234764 223304
rect 267464 223388 267516 223440
rect 287704 223388 287756 223440
rect 410248 223388 410300 223440
rect 448060 223388 448112 223440
rect 451280 223388 451332 223440
rect 467104 223388 467156 223440
rect 468760 223388 468812 223440
rect 529204 223388 529256 223440
rect 551928 223388 551980 223440
rect 564808 223388 564860 223440
rect 275008 223252 275060 223304
rect 375472 223252 375524 223304
rect 397828 223252 397880 223304
rect 399576 223252 399628 223304
rect 421564 223252 421616 223304
rect 431592 223252 431644 223304
rect 469864 223252 469916 223304
rect 470416 223252 470468 223304
rect 541624 223252 541676 223304
rect 541992 223252 542044 223304
rect 558000 223252 558052 223304
rect 81348 223116 81400 223168
rect 160468 223116 160520 223168
rect 184480 223116 184532 223168
rect 184848 223116 184900 223168
rect 232504 223116 232556 223168
rect 237012 223116 237064 223168
rect 268108 223116 268160 223168
rect 284208 223116 284260 223168
rect 300584 223116 300636 223168
rect 365720 223116 365772 223168
rect 380164 223116 380216 223168
rect 384120 223116 384172 223168
rect 408316 223116 408368 223168
rect 417240 223116 417292 223168
rect 456892 223116 456944 223168
rect 460480 223116 460532 223168
rect 523224 223116 523276 223168
rect 523684 223116 523736 223168
rect 529020 223116 529072 223168
rect 529204 223116 529256 223168
rect 539232 223116 539284 223168
rect 548340 223116 548392 223168
rect 549076 223116 549128 223168
rect 550640 223116 550692 223168
rect 42616 222980 42668 223032
rect 62764 222980 62816 223032
rect 75552 222980 75604 223032
rect 152280 222980 152332 223032
rect 152464 222980 152516 223032
rect 156420 222980 156472 223032
rect 62028 222844 62080 222896
rect 146668 222844 146720 222896
rect 146944 222844 146996 222896
rect 161480 222980 161532 223032
rect 171600 222980 171652 223032
rect 171784 222980 171836 223032
rect 176200 222980 176252 223032
rect 177948 222980 178000 223032
rect 228088 222980 228140 223032
rect 233056 222980 233108 223032
rect 265072 222980 265124 223032
rect 271788 222980 271840 223032
rect 292672 222980 292724 223032
rect 300584 222980 300636 223032
rect 312544 222980 312596 223032
rect 353944 222980 353996 223032
rect 366088 222980 366140 223032
rect 376024 222980 376076 223032
rect 399208 222980 399260 223032
rect 404636 222980 404688 223032
rect 428188 222980 428240 223032
rect 430672 222980 430724 223032
rect 471428 222980 471480 223032
rect 478696 222980 478748 223032
rect 483020 222980 483072 223032
rect 484124 222980 484176 223032
rect 551560 222980 551612 223032
rect 551744 222980 551796 223032
rect 558552 222980 558604 223032
rect 567752 222980 567804 223032
rect 156788 222844 156840 222896
rect 213184 222844 213236 222896
rect 215944 222844 215996 222896
rect 220268 222844 220320 222896
rect 221280 222844 221332 222896
rect 259552 222844 259604 222896
rect 261852 222844 261904 222896
rect 286048 222844 286100 222896
rect 293224 222844 293276 222896
rect 306104 222844 306156 222896
rect 362684 222844 362736 222896
rect 376024 222844 376076 222896
rect 380440 222844 380492 222896
rect 405832 222844 405884 222896
rect 412456 222844 412508 222896
rect 451464 222844 451516 222896
rect 471980 222844 472032 222896
rect 544200 222844 544252 222896
rect 128268 222708 128320 222760
rect 194968 222708 195020 222760
rect 197268 222708 197320 222760
rect 133144 222572 133196 222624
rect 146944 222572 146996 222624
rect 147128 222572 147180 222624
rect 151268 222572 151320 222624
rect 151452 222572 151504 222624
rect 156420 222572 156472 222624
rect 156604 222572 156656 222624
rect 208768 222572 208820 222624
rect 210332 222572 210384 222624
rect 231952 222572 232004 222624
rect 239312 222708 239364 222760
rect 242440 222708 242492 222760
rect 242808 222708 242860 222760
rect 246672 222708 246724 222760
rect 408040 222708 408092 222760
rect 444748 222708 444800 222760
rect 465816 222708 465868 222760
rect 533528 222708 533580 222760
rect 533804 222708 533856 222760
rect 534172 222708 534224 222760
rect 554044 222844 554096 222896
rect 554688 222844 554740 222896
rect 240968 222572 241020 222624
rect 395252 222572 395304 222624
rect 411628 222572 411680 222624
rect 425336 222572 425388 222624
rect 459008 222572 459060 222624
rect 467472 222572 467524 222624
rect 131028 222436 131080 222488
rect 133788 222436 133840 222488
rect 137652 222436 137704 222488
rect 201592 222436 201644 222488
rect 205640 222436 205692 222488
rect 215668 222436 215720 222488
rect 427728 222436 427780 222488
rect 460204 222436 460256 222488
rect 461952 222436 462004 222488
rect 524880 222436 524932 222488
rect 529020 222572 529072 222624
rect 555424 222708 555476 222760
rect 559564 222844 559616 222896
rect 571432 222980 571484 223032
rect 568120 222844 568172 222896
rect 596824 222844 596876 222896
rect 620468 222980 620520 223032
rect 619180 222844 619232 222896
rect 620284 222844 620336 222896
rect 625344 222844 625396 222896
rect 664628 222844 664680 222896
rect 675484 222844 675536 222896
rect 630956 222708 631008 222760
rect 664812 222708 664864 222760
rect 675300 222708 675352 222760
rect 536104 222504 536156 222556
rect 533528 222436 533580 222488
rect 88984 222300 89036 222352
rect 148876 222300 148928 222352
rect 151774 222300 151826 222352
rect 156604 222300 156656 222352
rect 158996 222300 159048 222352
rect 161296 222300 161348 222352
rect 161434 222300 161486 222352
rect 209872 222300 209924 222352
rect 459192 222300 459244 222352
rect 523040 222300 523092 222352
rect 523224 222300 523276 222352
rect 526720 222368 526772 222420
rect 527640 222368 527692 222420
rect 528468 222368 528520 222420
rect 533988 222368 534040 222420
rect 596640 222572 596692 222624
rect 596824 222572 596876 222624
rect 618720 222572 618772 222624
rect 619180 222572 619232 222624
rect 629300 222572 629352 222624
rect 661684 222572 661736 222624
rect 549904 222368 549956 222420
rect 620284 222436 620336 222488
rect 620468 222436 620520 222488
rect 631232 222436 631284 222488
rect 668400 222572 668452 222624
rect 675116 222572 675168 222624
rect 597008 222300 597060 222352
rect 619732 222300 619784 222352
rect 416044 222232 416096 222284
rect 91284 222096 91336 222148
rect 161572 222096 161624 222148
rect 161756 222096 161808 222148
rect 167644 222096 167696 222148
rect 171600 222096 171652 222148
rect 179696 222096 179748 222148
rect 184664 222096 184716 222148
rect 234988 222096 235040 222148
rect 258172 222096 258224 222148
rect 261024 222096 261076 222148
rect 265992 222096 266044 222148
rect 267004 222096 267056 222148
rect 377404 222096 377456 222148
rect 393412 222096 393464 222148
rect 393964 222096 394016 222148
rect 416596 222096 416648 222148
rect 429752 222096 429804 222148
rect 452568 222096 452620 222148
rect 79692 222028 79744 222080
rect 511264 222164 511316 222216
rect 523684 222164 523736 222216
rect 523868 222164 523920 222216
rect 618352 222164 618404 222216
rect 618720 222164 618772 222216
rect 619916 222164 619968 222216
rect 663064 222164 663116 222216
rect 668400 222164 668452 222216
rect 675484 222164 675536 222216
rect 529388 222096 529440 222148
rect 553308 222096 553360 222148
rect 555976 222096 556028 222148
rect 565728 222096 565780 222148
rect 567660 222096 567712 222148
rect 567844 222096 567896 222148
rect 591304 222096 591356 222148
rect 591488 222096 591540 222148
rect 80520 221892 80572 221944
rect 83464 221892 83516 221944
rect 514300 222028 514352 222080
rect 517796 222028 517848 222080
rect 518440 222028 518492 222080
rect 88800 221960 88852 222012
rect 156604 221960 156656 222012
rect 156788 221960 156840 222012
rect 178132 221960 178184 222012
rect 180064 221960 180116 222012
rect 230480 221960 230532 222012
rect 251916 221960 251968 222012
rect 278044 221960 278096 222012
rect 280896 221960 280948 222012
rect 297364 221960 297416 222012
rect 369768 221960 369820 222012
rect 387616 221960 387668 222012
rect 396908 221960 396960 222012
rect 419908 221960 419960 222012
rect 424324 221960 424376 222012
rect 443092 221960 443144 222012
rect 449900 221960 449952 222012
rect 509194 221960 509246 222012
rect 597836 222028 597888 222080
rect 591994 221960 592046 222012
rect 73896 221688 73948 221740
rect 77944 221688 77996 221740
rect 60648 221552 60700 221604
rect 79324 221688 79376 221740
rect 83004 221688 83056 221740
rect 88800 221688 88852 221740
rect 89260 221824 89312 221876
rect 161434 221824 161486 221876
rect 161572 221824 161624 221876
rect 164424 221824 164476 221876
rect 164608 221824 164660 221876
rect 170404 221824 170456 221876
rect 170772 221824 170824 221876
rect 173716 221824 173768 221876
rect 173900 221824 173952 221876
rect 174728 221824 174780 221876
rect 174912 221824 174964 221876
rect 223948 221824 224000 221876
rect 227076 221824 227128 221876
rect 258172 221824 258224 221876
rect 151912 221688 151964 221740
rect 152280 221688 152332 221740
rect 156420 221688 156472 221740
rect 156604 221688 156656 221740
rect 163596 221688 163648 221740
rect 164056 221688 164108 221740
rect 218888 221688 218940 221740
rect 223764 221688 223816 221740
rect 258632 221824 258684 221876
rect 263508 221824 263560 221876
rect 285128 221824 285180 221876
rect 351552 221824 351604 221876
rect 361212 221824 361264 221876
rect 372068 221824 372120 221876
rect 390928 221824 390980 221876
rect 397368 221824 397420 221876
rect 426532 221824 426584 221876
rect 427084 221824 427136 221876
rect 456340 221824 456392 221876
rect 456708 221824 456760 221876
rect 519268 221824 519320 221876
rect 520924 221824 520976 221876
rect 258540 221688 258592 221740
rect 282460 221688 282512 221740
rect 78864 221552 78916 221604
rect 161434 221552 161486 221604
rect 161572 221552 161624 221604
rect 171784 221552 171836 221604
rect 171968 221552 172020 221604
rect 226432 221552 226484 221604
rect 227904 221552 227956 221604
rect 263784 221552 263836 221604
rect 278412 221552 278464 221604
rect 295708 221552 295760 221604
rect 59360 221416 59412 221468
rect 147036 221416 147088 221468
rect 147220 221416 147272 221468
rect 150716 221416 150768 221468
rect 150900 221416 150952 221468
rect 197728 221416 197780 221468
rect 214012 221416 214064 221468
rect 220636 221416 220688 221468
rect 256792 221416 256844 221468
rect 257712 221416 257764 221468
rect 283196 221416 283248 221468
rect 283380 221416 283432 221468
rect 298468 221688 298520 221740
rect 303252 221688 303304 221740
rect 311992 221688 312044 221740
rect 357348 221688 357400 221740
rect 369400 221688 369452 221740
rect 379980 221688 380032 221740
rect 400036 221688 400088 221740
rect 404268 221688 404320 221740
rect 436468 221688 436520 221740
rect 441528 221688 441580 221740
rect 449900 221688 449952 221740
rect 458088 221688 458140 221740
rect 521752 221688 521804 221740
rect 522580 221824 522632 221876
rect 523868 221824 523920 221876
rect 600320 221824 600372 221876
rect 529756 221688 529808 221740
rect 602252 221688 602304 221740
rect 317420 221620 317472 221672
rect 318800 221620 318852 221672
rect 296904 221552 296956 221604
rect 301780 221552 301832 221604
rect 297456 221416 297508 221468
rect 310060 221552 310112 221604
rect 344928 221552 344980 221604
rect 348700 221552 348752 221604
rect 360016 221552 360068 221604
rect 374368 221552 374420 221604
rect 383200 221552 383252 221604
rect 406660 221552 406712 221604
rect 412272 221552 412324 221604
rect 446956 221552 447008 221604
rect 486608 221552 486660 221604
rect 555976 221552 556028 221604
rect 304908 221416 304960 221468
rect 313648 221416 313700 221468
rect 315764 221416 315816 221468
rect 320824 221416 320876 221468
rect 347596 221416 347648 221468
rect 356152 221416 356204 221468
rect 368296 221416 368348 221468
rect 385960 221416 386012 221468
rect 386328 221416 386380 221468
rect 409972 221416 410024 221468
rect 422208 221416 422260 221468
rect 464620 221416 464672 221468
rect 484492 221416 484544 221468
rect 563244 221552 563296 221604
rect 556344 221416 556396 221468
rect 567844 221416 567896 221468
rect 568304 221552 568356 221604
rect 611360 221552 611412 221604
rect 609980 221416 610032 221468
rect 87144 221280 87196 221332
rect 90364 221280 90416 221332
rect 102048 221280 102100 221332
rect 171600 221280 171652 221332
rect 171784 221280 171836 221332
rect 195612 221280 195664 221332
rect 210056 221280 210108 221332
rect 211344 221280 211396 221332
rect 252652 221280 252704 221332
rect 400864 221280 400916 221332
rect 423220 221280 423272 221332
rect 428464 221280 428516 221332
rect 439780 221280 439832 221332
rect 444932 221280 444984 221332
rect 503536 221280 503588 221332
rect 504548 221280 504600 221332
rect 529388 221280 529440 221332
rect 529572 221280 529624 221332
rect 593972 221280 594024 221332
rect 86316 221144 86368 221196
rect 89260 221144 89312 221196
rect 97724 221144 97776 221196
rect 173716 221144 173768 221196
rect 173900 221144 173952 221196
rect 594156 221212 594208 221264
rect 601056 221212 601108 221264
rect 664260 221212 664312 221264
rect 675484 221212 675536 221264
rect 222752 221144 222804 221196
rect 389732 221144 389784 221196
rect 403348 221144 403400 221196
rect 409512 221144 409564 221196
rect 422300 221144 422352 221196
rect 444288 221144 444340 221196
rect 501052 221144 501104 221196
rect 509240 221144 509292 221196
rect 511080 221144 511132 221196
rect 515956 221076 516008 221128
rect 600872 221076 600924 221128
rect 104532 221008 104584 221060
rect 179420 221008 179472 221060
rect 179880 221008 179932 221060
rect 183468 221008 183520 221060
rect 186504 221008 186556 221060
rect 194232 221008 194284 221060
rect 195612 221008 195664 221060
rect 197728 221008 197780 221060
rect 213368 221008 213420 221060
rect 252100 221008 252152 221060
rect 420184 221008 420236 221060
rect 433156 221008 433208 221060
rect 439964 221008 440016 221060
rect 491208 221008 491260 221060
rect 669044 221008 669096 221060
rect 675484 221008 675536 221060
rect 513564 220940 513616 220992
rect 598940 220940 598992 220992
rect 117780 220872 117832 220924
rect 187976 220872 188028 220924
rect 253848 220872 253900 220924
rect 259828 220872 259880 220924
rect 343456 220872 343508 220924
rect 347044 220872 347096 220924
rect 463700 220872 463752 220924
rect 508596 220872 508648 220924
rect 313004 220804 313056 220856
rect 318248 220804 318300 220856
rect 320640 220804 320692 220856
rect 325792 220804 325844 220856
rect 591120 220804 591172 220856
rect 591304 220804 591356 220856
rect 607220 220804 607272 220856
rect 667480 220804 667532 220856
rect 675300 220804 675352 220856
rect 83188 220736 83240 220788
rect 152096 220736 152148 220788
rect 155868 220736 155920 220788
rect 215392 220736 215444 220788
rect 240324 220736 240376 220788
rect 269764 220736 269816 220788
rect 310520 220736 310572 220788
rect 311164 220736 311216 220788
rect 337936 220736 337988 220788
rect 341248 220736 341300 220788
rect 345848 220736 345900 220788
rect 346400 220736 346452 220788
rect 348424 220736 348476 220788
rect 349528 220736 349580 220788
rect 349804 220736 349856 220788
rect 351184 220736 351236 220788
rect 369124 220736 369176 220788
rect 371884 220736 371936 220788
rect 379336 220736 379388 220788
rect 402520 220736 402572 220788
rect 413468 220736 413520 220788
rect 442264 220736 442316 220788
rect 446220 220736 446272 220788
rect 505008 220736 505060 220788
rect 506020 220736 506072 220788
rect 318156 220668 318208 220720
rect 322204 220668 322256 220720
rect 107844 220600 107896 220652
rect 181536 220600 181588 220652
rect 190644 220600 190696 220652
rect 236460 220600 236512 220652
rect 247868 220600 247920 220652
rect 276940 220600 276992 220652
rect 288348 220600 288400 220652
rect 302424 220600 302476 220652
rect 340604 220600 340656 220652
rect 344560 220600 344612 220652
rect 347228 220600 347280 220652
rect 354496 220600 354548 220652
rect 392768 220600 392820 220652
rect 422484 220600 422536 220652
rect 437296 220600 437348 220652
rect 478788 220600 478840 220652
rect 479524 220600 479576 220652
rect 543556 220600 543608 220652
rect 103428 220464 103480 220516
rect 177028 220464 177080 220516
rect 180708 220464 180760 220516
rect 229928 220464 229980 220516
rect 233700 220464 233752 220516
rect 265348 220464 265400 220516
rect 268476 220464 268528 220516
rect 288992 220464 289044 220516
rect 352564 220464 352616 220516
rect 357808 220464 357860 220516
rect 362868 220464 362920 220516
rect 379336 220464 379388 220516
rect 384672 220464 384724 220516
rect 412456 220464 412508 220516
rect 415308 220464 415360 220516
rect 453028 220464 453080 220516
rect 473176 220464 473228 220516
rect 539048 220464 539100 220516
rect 540796 220464 540848 220516
rect 94596 220328 94648 220380
rect 172888 220328 172940 220380
rect 174084 220328 174136 220380
rect 225512 220328 225564 220380
rect 230388 220328 230440 220380
rect 263048 220328 263100 220380
rect 264336 220328 264388 220380
rect 287888 220328 287940 220380
rect 288532 220328 288584 220380
rect 303712 220328 303764 220380
rect 354312 220328 354364 220380
rect 361764 220328 361816 220380
rect 365444 220328 365496 220380
rect 380992 220328 381044 220380
rect 390468 220328 390520 220380
rect 419080 220328 419132 220380
rect 420552 220328 420604 220380
rect 459836 220328 459888 220380
rect 477776 220328 477828 220380
rect 543832 220328 543884 220380
rect 553354 220668 553406 220720
rect 544384 220600 544436 220652
rect 553124 220600 553176 220652
rect 558000 220464 558052 220516
rect 558368 220668 558420 220720
rect 562784 220668 562836 220720
rect 562968 220668 563020 220720
rect 572536 220668 572588 220720
rect 572674 220600 572726 220652
rect 574560 220600 574612 220652
rect 574744 220600 574796 220652
rect 597008 220600 597060 220652
rect 607772 220464 607824 220516
rect 545764 220328 545816 220380
rect 76380 220192 76432 220244
rect 153936 220192 153988 220244
rect 69756 220056 69808 220108
rect 156052 220192 156104 220244
rect 156236 220192 156288 220244
rect 160652 220192 160704 220244
rect 160836 220192 160888 220244
rect 216864 220192 216916 220244
rect 226892 220192 226944 220244
rect 233424 220192 233476 220244
rect 237840 220192 237892 220244
rect 270592 220192 270644 220244
rect 271604 220192 271656 220244
rect 291384 220192 291436 220244
rect 303436 220192 303488 220244
rect 310796 220192 310848 220244
rect 343272 220192 343324 220244
rect 347872 220192 347924 220244
rect 358268 220192 358320 220244
rect 371056 220192 371108 220244
rect 372068 220192 372120 220244
rect 389272 220192 389324 220244
rect 395712 220192 395764 220244
rect 429016 220192 429068 220244
rect 436008 220192 436060 220244
rect 480260 220192 480312 220244
rect 481548 220192 481600 220244
rect 552940 220192 552992 220244
rect 553860 220328 553912 220380
rect 608876 220328 608928 220380
rect 557816 220192 557868 220244
rect 558000 220192 558052 220244
rect 564624 220192 564676 220244
rect 596640 220192 596692 220244
rect 605012 220192 605064 220244
rect 154304 220056 154356 220108
rect 212632 220056 212684 220108
rect 217140 220056 217192 220108
rect 254308 220056 254360 220108
rect 256884 220056 256936 220108
rect 280712 220056 280764 220108
rect 281264 220056 281316 220108
rect 297088 220056 297140 220108
rect 298284 220056 298336 220108
rect 309232 220056 309284 220108
rect 355968 220056 356020 220108
rect 367744 220056 367796 220108
rect 373724 220056 373776 220108
rect 395896 220056 395948 220108
rect 398564 220056 398616 220108
rect 432328 220056 432380 220108
rect 442908 220056 442960 220108
rect 485734 220056 485786 220108
rect 485872 220056 485924 220108
rect 553400 220056 553452 220108
rect 596456 220124 596508 220176
rect 124404 219920 124456 219972
rect 192484 219920 192536 219972
rect 200580 219920 200632 219972
rect 243268 219920 243320 219972
rect 388628 219920 388680 219972
rect 415768 219920 415820 219972
rect 418804 219920 418856 219972
rect 455512 219920 455564 219972
rect 469496 219920 469548 219972
rect 526444 219920 526496 219972
rect 126060 219784 126112 219836
rect 191288 219784 191340 219836
rect 193036 219784 193088 219836
rect 200856 219784 200908 219836
rect 207204 219784 207256 219836
rect 247500 219784 247552 219836
rect 428832 219784 428884 219836
rect 462320 219784 462372 219836
rect 464988 219784 465040 219836
rect 533344 219852 533396 219904
rect 48964 219648 49016 219700
rect 54208 219648 54260 219700
rect 138296 219648 138348 219700
rect 143632 219648 143684 219700
rect 128452 219580 128504 219632
rect 129740 219580 129792 219632
rect 140964 219512 141016 219564
rect 203524 219648 203576 219700
rect 205364 219648 205416 219700
rect 205824 219648 205876 219700
rect 213920 219648 213972 219700
rect 224408 219648 224460 219700
rect 421380 219648 421432 219700
rect 445576 219648 445628 219700
rect 463516 219648 463568 219700
rect 530860 219716 530912 219768
rect 538680 219852 538732 219904
rect 540796 219852 540848 219904
rect 540980 219852 541032 219904
rect 565360 219988 565412 220040
rect 574744 219988 574796 220040
rect 574928 219988 574980 220040
rect 610164 219988 610216 220040
rect 557816 219852 557868 219904
rect 350264 219580 350316 219632
rect 145012 219512 145064 219564
rect 147404 219512 147456 219564
rect 147588 219512 147640 219564
rect 207848 219512 207900 219564
rect 63132 219376 63184 219428
rect 83188 219444 83240 219496
rect 97080 219376 97132 219428
rect 98000 219376 98052 219428
rect 108304 219376 108356 219428
rect 113824 219376 113876 219428
rect 114468 219376 114520 219428
rect 144460 219444 144512 219496
rect 131672 219376 131724 219428
rect 131856 219376 131908 219428
rect 132408 219376 132460 219428
rect 132684 219376 132736 219428
rect 133420 219376 133472 219428
rect 135996 219376 136048 219428
rect 136548 219376 136600 219428
rect 136824 219376 136876 219428
rect 138296 219376 138348 219428
rect 138480 219376 138532 219428
rect 141148 219376 141200 219428
rect 169208 219376 169260 219428
rect 169944 219376 169996 219428
rect 178592 219376 178644 219428
rect 184020 219376 184072 219428
rect 184940 219376 184992 219428
rect 185308 219376 185360 219428
rect 189724 219376 189776 219428
rect 189908 219376 189960 219428
rect 226892 219444 226944 219496
rect 236184 219376 236236 219428
rect 311532 219444 311584 219496
rect 317696 219444 317748 219496
rect 267924 219376 267976 219428
rect 269304 219376 269356 219428
rect 284944 219376 284996 219428
rect 299940 219376 299992 219428
rect 300860 219376 300912 219428
rect 319812 219376 319864 219428
rect 323032 219444 323084 219496
rect 324044 219444 324096 219496
rect 327816 219444 327868 219496
rect 344284 219444 344336 219496
rect 346216 219444 346268 219496
rect 529388 219580 529440 219632
rect 538680 219580 538732 219632
rect 539048 219716 539100 219768
rect 543832 219716 543884 219768
rect 545212 219716 545264 219768
rect 596640 219716 596692 219768
rect 597008 219852 597060 219904
rect 605932 219852 605984 219904
rect 606116 219716 606168 219768
rect 666192 219716 666244 219768
rect 675484 219784 675536 219836
rect 603908 219580 603960 219632
rect 665088 219580 665140 219632
rect 675300 219580 675352 219632
rect 447692 219512 447744 219564
rect 506848 219512 506900 219564
rect 511080 219444 511132 219496
rect 422300 219376 422352 219428
rect 448888 219376 448940 219428
rect 449164 219376 449216 219428
rect 64604 219104 64656 219156
rect 88984 219240 89036 219292
rect 100392 219240 100444 219292
rect 356980 219308 357032 219360
rect 147220 219240 147272 219292
rect 147404 219240 147456 219292
rect 192484 219240 192536 219292
rect 195612 219240 195664 219292
rect 197912 219240 197964 219292
rect 198924 219240 198976 219292
rect 200028 219240 200080 219292
rect 200212 219240 200264 219292
rect 201040 219240 201092 219292
rect 208860 219240 208912 219292
rect 209596 219240 209648 219292
rect 209780 219240 209832 219292
rect 210332 219240 210384 219292
rect 210516 219240 210568 219292
rect 210976 219240 211028 219292
rect 213000 219240 213052 219292
rect 213552 219240 213604 219292
rect 213736 219240 213788 219292
rect 239312 219240 239364 219292
rect 249432 219240 249484 219292
rect 59820 218968 59872 219020
rect 87604 219104 87656 219156
rect 87972 219104 88024 219156
rect 101404 219104 101456 219156
rect 113640 219104 113692 219156
rect 120908 219104 120960 219156
rect 121920 219104 121972 219156
rect 122748 219104 122800 219156
rect 123576 219104 123628 219156
rect 126428 219104 126480 219156
rect 126612 219104 126664 219156
rect 128498 219104 128550 219156
rect 128636 219104 128688 219156
rect 164424 219104 164476 219156
rect 164608 219104 164660 219156
rect 171600 219104 171652 219156
rect 83832 218968 83884 219020
rect 70584 218832 70636 218884
rect 156420 218832 156472 218884
rect 157524 218832 157576 218884
rect 161388 218832 161440 218884
rect 161756 218968 161808 219020
rect 178408 219104 178460 219156
rect 178592 219104 178644 219156
rect 213920 219104 213972 219156
rect 214656 219104 214708 219156
rect 215208 219104 215260 219156
rect 224224 219104 224276 219156
rect 251732 219104 251784 219156
rect 252744 219104 252796 219156
rect 255964 219104 256016 219156
rect 262864 219104 262916 219156
rect 272432 219104 272484 219156
rect 178592 218968 178644 219020
rect 180064 218968 180116 219020
rect 180248 218968 180300 219020
rect 185768 218968 185820 219020
rect 185952 218968 186004 219020
rect 209136 218968 209188 219020
rect 167368 218832 167420 218884
rect 167552 218832 167604 218884
rect 170128 218832 170180 218884
rect 171600 218832 171652 218884
rect 215944 218968 215996 219020
rect 217968 218968 218020 219020
rect 221464 218968 221516 219020
rect 242624 218968 242676 219020
rect 273444 218968 273496 219020
rect 209688 218832 209740 218884
rect 56508 218696 56560 218748
rect 144920 218696 144972 218748
rect 78036 218560 78088 218612
rect 108304 218560 108356 218612
rect 111984 218560 112036 218612
rect 113088 218560 113140 218612
rect 110144 218424 110196 218476
rect 116124 218424 116176 218476
rect 117228 218424 117280 218476
rect 119436 218424 119488 218476
rect 119988 218424 120040 218476
rect 120356 218560 120408 218612
rect 125508 218560 125560 218612
rect 125692 218560 125744 218612
rect 120724 218424 120776 218476
rect 120908 218424 120960 218476
rect 126612 218424 126664 218476
rect 127716 218424 127768 218476
rect 128268 218424 128320 218476
rect 128544 218424 128596 218476
rect 129280 218424 129332 218476
rect 131672 218424 131724 218476
rect 137928 218424 137980 218476
rect 138480 218424 138532 218476
rect 139124 218424 139176 218476
rect 140136 218424 140188 218476
rect 140688 218424 140740 218476
rect 141148 218560 141200 218612
rect 142252 218560 142304 218612
rect 144460 218560 144512 218612
rect 147404 218696 147456 218748
rect 149244 218696 149296 218748
rect 142620 218424 142672 218476
rect 143448 218424 143500 218476
rect 143632 218424 143684 218476
rect 146760 218560 146812 218612
rect 151084 218560 151136 218612
rect 145104 218424 145156 218476
rect 145932 218424 145984 218476
rect 148416 218424 148468 218476
rect 149888 218424 149940 218476
rect 151912 218696 151964 218748
rect 151452 218560 151504 218612
rect 191932 218560 191984 218612
rect 192300 218560 192352 218612
rect 193772 218560 193824 218612
rect 193956 218560 194008 218612
rect 194416 218560 194468 218612
rect 194784 218560 194836 218612
rect 195888 218560 195940 218612
rect 196256 218560 196308 218612
rect 199844 218560 199896 218612
rect 200212 218696 200264 218748
rect 202880 218696 202932 218748
rect 205502 218696 205554 218748
rect 213736 218696 213788 218748
rect 214104 218832 214156 218884
rect 222844 218832 222896 218884
rect 229560 218832 229612 218884
rect 262680 218832 262732 218884
rect 295800 219240 295852 219292
rect 296720 219240 296772 219292
rect 342260 219240 342312 219292
rect 345388 219240 345440 219292
rect 402244 219240 402296 219292
rect 424876 219240 424928 219292
rect 285864 219104 285916 219156
rect 296904 219104 296956 219156
rect 302424 219104 302476 219156
rect 305644 219104 305696 219156
rect 405004 219104 405056 219156
rect 430856 219240 430908 219292
rect 431224 219240 431276 219292
rect 425888 219104 425940 219156
rect 436928 219240 436980 219292
rect 454684 219240 454736 219292
rect 457444 219376 457496 219428
rect 458824 219240 458876 219292
rect 462320 219376 462372 219428
rect 474556 219376 474608 219428
rect 474740 219376 474792 219428
rect 489368 219376 489420 219428
rect 471060 219240 471112 219292
rect 471428 219240 471480 219292
rect 475752 219240 475804 219292
rect 480260 219240 480312 219292
rect 483572 219240 483624 219292
rect 483756 219240 483808 219292
rect 484308 219240 484360 219292
rect 490196 219308 490248 219360
rect 490380 219308 490432 219360
rect 275652 218968 275704 219020
rect 290464 218968 290516 219020
rect 301596 218968 301648 219020
rect 310520 218968 310572 219020
rect 314016 218968 314068 219020
rect 319444 218968 319496 219020
rect 363604 218968 363656 219020
rect 368572 218968 368624 219020
rect 407028 218968 407080 219020
rect 436284 218968 436336 219020
rect 436928 218968 436980 219020
rect 446404 218968 446456 219020
rect 459652 218968 459704 219020
rect 460204 219104 460256 219156
rect 472900 219104 472952 219156
rect 475108 219104 475160 219156
rect 482836 219104 482888 219156
rect 489828 219172 489880 219224
rect 547512 219308 547564 219360
rect 549444 219308 549496 219360
rect 559840 219308 559892 219360
rect 568028 219308 568080 219360
rect 568212 219308 568264 219360
rect 596456 219444 596508 219496
rect 604552 219444 604604 219496
rect 671896 219444 671948 219496
rect 675484 219444 675536 219496
rect 599124 219308 599176 219360
rect 574744 219240 574796 219292
rect 460480 218968 460532 219020
rect 467288 218968 467340 219020
rect 485044 219104 485096 219156
rect 486148 219104 486200 219156
rect 491484 219036 491536 219088
rect 495256 219036 495308 219088
rect 526444 219036 526496 219088
rect 529388 219036 529440 219088
rect 530124 219036 530176 219088
rect 530584 219036 530636 219088
rect 531964 219036 532016 219088
rect 532516 219036 532568 219088
rect 535920 219036 535972 219088
rect 540980 219036 541032 219088
rect 551744 219172 551796 219224
rect 554872 219104 554924 219156
rect 550640 219036 550692 219088
rect 485412 218968 485464 219020
rect 277584 218832 277636 218884
rect 282552 218832 282604 218884
rect 298744 218832 298796 218884
rect 305736 218832 305788 218884
rect 313832 218832 313884 218884
rect 366732 218832 366784 218884
rect 381820 218832 381872 218884
rect 382188 218832 382240 218884
rect 405004 218832 405056 218884
rect 405372 218832 405424 218884
rect 438124 218832 438176 218884
rect 454868 218832 454920 218884
rect 463792 218832 463844 218884
rect 469864 218832 469916 218884
rect 474924 218832 474976 218884
rect 243544 218696 243596 218748
rect 262680 218696 262732 218748
rect 286048 218696 286100 218748
rect 292304 218696 292356 218748
rect 305920 218696 305972 218748
rect 310704 218696 310756 218748
rect 317420 218696 317472 218748
rect 323124 218696 323176 218748
rect 324688 218696 324740 218748
rect 355324 218696 355376 218748
rect 358636 218696 358688 218748
rect 360844 218696 360896 218748
rect 365260 218696 365312 218748
rect 368112 218696 368164 218748
rect 385132 218696 385184 218748
rect 401324 218696 401376 218748
rect 434812 218696 434864 218748
rect 438308 218696 438360 218748
rect 475108 218696 475160 218748
rect 485412 218832 485464 218884
rect 485872 218968 485924 219020
rect 491300 218968 491352 219020
rect 498384 218968 498436 219020
rect 524328 218968 524380 219020
rect 552204 218968 552256 219020
rect 552388 218968 552440 219020
rect 558184 218968 558236 219020
rect 561772 219104 561824 219156
rect 562324 219104 562376 219156
rect 567476 219104 567528 219156
rect 567660 219104 567712 219156
rect 574928 219104 574980 219156
rect 567844 218968 567896 219020
rect 568028 218968 568080 219020
rect 575296 218968 575348 219020
rect 529572 218832 529624 218884
rect 530584 218832 530636 218884
rect 596088 218832 596140 218884
rect 254400 218628 254452 218680
rect 256148 218628 256200 218680
rect 207848 218560 207900 218612
rect 244924 218560 244976 218612
rect 324780 218560 324832 218612
rect 326068 218560 326120 218612
rect 349160 218560 349212 218612
rect 355324 218560 355376 218612
rect 357164 218560 357216 218612
rect 366916 218560 366968 218612
rect 421840 218560 421892 218612
rect 446404 218560 446456 218612
rect 450544 218560 450596 218612
rect 457168 218560 457220 218612
rect 459008 218560 459060 218612
rect 469588 218560 469640 218612
rect 206100 218492 206152 218544
rect 256056 218492 256108 218544
rect 262864 218492 262916 218544
rect 152464 218424 152516 218476
rect 89444 218288 89496 218340
rect 55680 218152 55732 218204
rect 57244 218152 57296 218204
rect 66444 218152 66496 218204
rect 69572 218152 69624 218204
rect 90456 218152 90508 218204
rect 95424 218288 95476 218340
rect 96252 218288 96304 218340
rect 103704 218288 103756 218340
rect 153384 218288 153436 218340
rect 154120 218288 154172 218340
rect 155040 218288 155092 218340
rect 155960 218288 156012 218340
rect 156696 218424 156748 218476
rect 161296 218424 161348 218476
rect 161480 218424 161532 218476
rect 183560 218424 183612 218476
rect 158996 218288 159048 218340
rect 159180 218288 159232 218340
rect 160008 218288 160060 218340
rect 160192 218288 160244 218340
rect 164792 218288 164844 218340
rect 166632 218288 166684 218340
rect 164976 218220 165028 218272
rect 166264 218220 166316 218272
rect 57336 218016 57388 218068
rect 57888 218016 57940 218068
rect 58164 218016 58216 218068
rect 59360 218016 59412 218068
rect 61476 218016 61528 218068
rect 62028 218016 62080 218068
rect 62304 218016 62356 218068
rect 63408 218016 63460 218068
rect 63960 218016 64012 218068
rect 64788 218016 64840 218068
rect 65616 218016 65668 218068
rect 66168 218016 66220 218068
rect 68100 218016 68152 218068
rect 68744 218016 68796 218068
rect 72240 218016 72292 218068
rect 73712 218016 73764 218068
rect 74724 218016 74776 218068
rect 75552 218016 75604 218068
rect 82176 218016 82228 218068
rect 82728 218016 82780 218068
rect 84660 218016 84712 218068
rect 85304 218016 85356 218068
rect 88800 218016 88852 218068
rect 89628 218016 89680 218068
rect 92940 218016 92992 218068
rect 93584 218016 93636 218068
rect 161480 218152 161532 218204
rect 163320 218152 163372 218204
rect 164608 218152 164660 218204
rect 169116 218152 169168 218204
rect 173900 218152 173952 218204
rect 175740 218152 175792 218204
rect 176568 218152 176620 218204
rect 178408 218288 178460 218340
rect 205456 218424 205508 218476
rect 206376 218424 206428 218476
rect 214104 218424 214156 218476
rect 216312 218424 216364 218476
rect 224224 218424 224276 218476
rect 224408 218424 224460 218476
rect 253848 218424 253900 218476
rect 434168 218424 434220 218476
rect 450544 218424 450596 218476
rect 458640 218424 458692 218476
rect 468760 218424 468812 218476
rect 196256 218288 196308 218340
rect 196440 218288 196492 218340
rect 200212 218288 200264 218340
rect 201408 218288 201460 218340
rect 205456 218288 205508 218340
rect 205640 218288 205692 218340
rect 242164 218288 242216 218340
rect 243544 218288 243596 218340
rect 249064 218288 249116 218340
rect 436284 218288 436336 218340
rect 441436 218288 441488 218340
rect 459836 218288 459888 218340
rect 462964 218288 463016 218340
rect 464804 218288 464856 218340
rect 475752 218560 475804 218612
rect 481180 218696 481232 218748
rect 482652 218696 482704 218748
rect 486976 218696 487028 218748
rect 487896 218696 487948 218748
rect 490380 218696 490432 218748
rect 491300 218696 491352 218748
rect 498384 218696 498436 218748
rect 498752 218696 498804 218748
rect 554688 218696 554740 218748
rect 558184 218696 558236 218748
rect 567660 218696 567712 218748
rect 567844 218696 567896 218748
rect 625068 218696 625120 218748
rect 480444 218560 480496 218612
rect 502984 218560 503036 218612
rect 542360 218560 542412 218612
rect 623320 218560 623372 218612
rect 472624 218424 472676 218476
rect 490334 218424 490386 218476
rect 491300 218424 491352 218476
rect 497740 218424 497792 218476
rect 498752 218424 498804 218476
rect 540060 218424 540112 218476
rect 601700 218424 601752 218476
rect 474924 218288 474976 218340
rect 482008 218288 482060 218340
rect 482192 218288 482244 218340
rect 491944 218288 491996 218340
rect 503352 218288 503404 218340
rect 535000 218288 535052 218340
rect 608508 218288 608560 218340
rect 185768 218152 185820 218204
rect 215208 218152 215260 218204
rect 215484 218152 215536 218204
rect 216496 218152 216548 218204
rect 218796 218152 218848 218204
rect 219348 218152 219400 218204
rect 219624 218152 219676 218204
rect 220360 218152 220412 218204
rect 222936 218152 222988 218204
rect 224408 218152 224460 218204
rect 225420 218152 225472 218204
rect 226064 218152 226116 218204
rect 161664 218084 161716 218136
rect 162492 218084 162544 218136
rect 165804 218084 165856 218136
rect 166816 218084 166868 218136
rect 177396 218084 177448 218136
rect 177948 218084 178000 218136
rect 98736 218016 98788 218068
rect 99288 218016 99340 218068
rect 99564 218016 99616 218068
rect 100668 218016 100720 218068
rect 101220 218016 101272 218068
rect 103428 218016 103480 218068
rect 105360 218016 105412 218068
rect 106188 218016 106240 218068
rect 107016 218016 107068 218068
rect 107568 218016 107620 218068
rect 109500 218016 109552 218068
rect 110328 218016 110380 218068
rect 111156 218016 111208 218068
rect 111708 218016 111760 218068
rect 112812 218016 112864 218068
rect 181536 218016 181588 218068
rect 182824 218016 182876 218068
rect 183008 218016 183060 218068
rect 185124 217880 185176 217932
rect 185676 218016 185728 218068
rect 186136 218016 186188 218068
rect 188160 218016 188212 218068
rect 188804 218016 188856 218068
rect 189816 218016 189868 218068
rect 236644 218152 236696 218204
rect 274272 218152 274324 218204
rect 275284 218152 275336 218204
rect 277584 218152 277636 218204
rect 281264 218152 281316 218204
rect 290832 218152 290884 218204
rect 293224 218152 293276 218204
rect 306564 218152 306616 218204
rect 313464 218152 313516 218204
rect 318984 218152 319036 218204
rect 323308 218152 323360 218204
rect 327264 218152 327316 218204
rect 329932 218152 329984 218204
rect 339316 218152 339368 218204
rect 342904 218152 342956 218204
rect 346032 218152 346084 218204
rect 352012 218152 352064 218204
rect 361028 218152 361080 218204
rect 361948 218152 362000 218204
rect 449900 218152 449952 218204
rect 490564 218152 490616 218204
rect 490932 218152 490984 218204
rect 493692 218152 493744 218204
rect 493876 218152 493928 218204
rect 496912 218152 496964 218204
rect 532516 218152 532568 218204
rect 597192 218152 597244 218204
rect 231216 218016 231268 218068
rect 231676 218016 231728 218068
rect 232044 218016 232096 218068
rect 233056 218016 233108 218068
rect 235356 218016 235408 218068
rect 235908 218016 235960 218068
rect 239496 218016 239548 218068
rect 240048 218016 240100 218068
rect 241980 218016 242032 218068
rect 242808 218016 242860 218068
rect 243636 218016 243688 218068
rect 244188 218016 244240 218068
rect 244464 218016 244516 218068
rect 245292 218016 245344 218068
rect 246120 218016 246172 218068
rect 247592 218016 247644 218068
rect 248604 218016 248656 218068
rect 249616 218016 249668 218068
rect 250260 218016 250312 218068
rect 251180 218016 251232 218068
rect 261024 218016 261076 218068
rect 261852 218016 261904 218068
rect 265164 218016 265216 218068
rect 266268 218016 266320 218068
rect 266820 218016 266872 218068
rect 267464 218016 267516 218068
rect 270960 218016 271012 218068
rect 271880 218016 271932 218068
rect 272616 218016 272668 218068
rect 273168 218016 273220 218068
rect 273444 218016 273496 218068
rect 274548 218016 274600 218068
rect 275100 218016 275152 218068
rect 275836 218016 275888 218068
rect 276756 218016 276808 218068
rect 277216 218016 277268 218068
rect 279240 218016 279292 218068
rect 279792 218016 279844 218068
rect 281724 218016 281776 218068
rect 282736 218016 282788 218068
rect 285036 218016 285088 218068
rect 285588 218016 285640 218068
rect 287520 218016 287572 218068
rect 288532 218016 288584 218068
rect 289176 218016 289228 218068
rect 289728 218016 289780 218068
rect 290004 218016 290056 218068
rect 291016 218016 291068 218068
rect 291660 218016 291712 218068
rect 292488 218016 292540 218068
rect 293316 218016 293368 218068
rect 293776 218016 293828 218068
rect 294144 218016 294196 218068
rect 294972 218016 295024 218068
rect 299112 218016 299164 218068
rect 303436 218016 303488 218068
rect 304080 218016 304132 218068
rect 304632 218016 304684 218068
rect 308220 218016 308272 218068
rect 308772 218016 308824 218068
rect 309876 218016 309928 218068
rect 310336 218016 310388 218068
rect 312360 218016 312412 218068
rect 313280 218016 313332 218068
rect 314844 218016 314896 218068
rect 315580 218016 315632 218068
rect 316500 218016 316552 218068
rect 317052 218016 317104 218068
rect 322296 218016 322348 218068
rect 322756 218016 322808 218068
rect 326436 218016 326488 218068
rect 327632 218016 327684 218068
rect 328092 218016 328144 218068
rect 328552 218016 328604 218068
rect 328920 218016 328972 218068
rect 330116 218016 330168 218068
rect 330576 218016 330628 218068
rect 331220 218016 331272 218068
rect 332232 218016 332284 218068
rect 332692 218016 332744 218068
rect 336556 218016 336608 218068
rect 339592 218016 339644 218068
rect 346400 218016 346452 218068
rect 350356 218016 350408 218068
rect 358084 218016 358136 218068
rect 360292 218016 360344 218068
rect 361764 218016 361816 218068
rect 363604 218016 363656 218068
rect 374644 218016 374696 218068
rect 378508 218016 378560 218068
rect 387064 218016 387116 218068
rect 388444 218016 388496 218068
rect 429936 218016 429988 218068
rect 430672 218016 430724 218068
rect 430856 218016 430908 218068
rect 431500 218016 431552 218068
rect 432604 218016 432656 218068
rect 435640 218016 435692 218068
rect 446956 218016 447008 218068
rect 449716 218016 449768 218068
rect 471060 218016 471112 218068
rect 477868 218016 477920 218068
rect 479616 218016 479668 218068
rect 504364 218016 504416 218068
rect 549444 218016 549496 218068
rect 567660 218016 567712 218068
rect 574192 218016 574244 218068
rect 614120 218016 614172 218068
rect 527824 217948 527876 218000
rect 528376 217948 528428 218000
rect 543832 217948 543884 218000
rect 545856 217948 545908 218000
rect 185952 217880 186004 217932
rect 205456 217880 205508 217932
rect 205640 217880 205692 217932
rect 486516 217880 486568 217932
rect 492772 217880 492824 217932
rect 567844 217948 567896 218000
rect 570144 217948 570196 218000
rect 167276 217812 167328 217864
rect 167460 217812 167512 217864
rect 172612 217812 172664 217864
rect 176568 217812 176620 217864
rect 180248 217812 180300 217864
rect 397644 217812 397696 217864
rect 398380 217812 398432 217864
rect 530860 217812 530912 217864
rect 548156 217812 548208 217864
rect 601976 217812 602028 217864
rect 134340 217676 134392 217728
rect 199108 217676 199160 217728
rect 445392 217676 445444 217728
rect 456064 217676 456116 217728
rect 528376 217676 528428 217728
rect 596640 217676 596692 217728
rect 596824 217676 596876 217728
rect 608324 217676 608376 217728
rect 608508 217676 608560 217728
rect 621664 217676 621716 217728
rect 122748 217540 122800 217592
rect 192116 217540 192168 217592
rect 444104 217540 444156 217592
rect 501880 217540 501932 217592
rect 548156 217540 548208 217592
rect 601516 217540 601568 217592
rect 601700 217540 601752 217592
rect 622768 217540 622820 217592
rect 106188 217404 106240 217456
rect 181168 217404 181220 217456
rect 456064 217404 456116 217456
rect 504364 217404 504416 217456
rect 555700 217404 555752 217456
rect 449532 217336 449584 217388
rect 102830 217200 102882 217252
rect 178040 217268 178092 217320
rect 203018 217200 203070 217252
rect 207848 217200 207900 217252
rect 361580 217200 361632 217252
rect 362822 217200 362874 217252
rect 374000 217200 374052 217252
rect 375242 217200 375294 217252
rect 402980 217200 403032 217252
rect 404222 217200 404274 217252
rect 419724 217200 419776 217252
rect 420782 217200 420834 217252
rect 509378 217200 509430 217252
rect 510620 217200 510672 217252
rect 511862 217200 511914 217252
rect 518900 217200 518952 217252
rect 520142 217200 520194 217252
rect 523040 217200 523092 217252
rect 524282 217200 524334 217252
rect 524880 217200 524932 217252
rect 529250 217200 529302 217252
rect 544154 217200 544206 217252
rect 544568 217200 544620 217252
rect 552940 217200 552992 217252
rect 558230 217200 558282 217252
rect 567844 217200 567896 217252
rect 568580 217200 568632 217252
rect 569822 217200 569874 217252
rect 570144 217404 570196 217456
rect 596824 217404 596876 217456
rect 597008 217404 597060 217456
rect 601332 217404 601384 217456
rect 601654 217404 601706 217456
rect 620560 217404 620612 217456
rect 672356 217336 672408 217388
rect 672908 217336 672960 217388
rect 609060 217268 609112 217320
rect 167276 217132 167328 217184
rect 171232 217132 171284 217184
rect 451280 217132 451332 217184
rect 452246 217132 452298 217184
rect 456892 217132 456944 217184
rect 458042 217132 458094 217184
rect 469312 217132 469364 217184
rect 470462 217132 470514 217184
rect 477592 217132 477644 217184
rect 478742 217132 478794 217184
rect 498200 217132 498252 217184
rect 499442 217132 499494 217184
rect 597008 217132 597060 217184
rect 628840 217268 628892 217320
rect 483572 217064 483624 217116
rect 488678 217064 488730 217116
rect 491392 217064 491444 217116
rect 523454 217064 523506 217116
rect 523684 217064 523736 217116
rect 601792 216996 601844 217048
rect 574284 216928 574336 216980
rect 597008 216860 597060 216912
rect 597192 216792 597244 216844
rect 621112 216928 621164 216980
rect 670608 216928 670660 216980
rect 675392 216928 675444 216980
rect 609612 216792 609664 216844
rect 615684 216792 615736 216844
rect 596088 216656 596140 216708
rect 601608 216656 601660 216708
rect 601976 216656 602028 216708
rect 606760 216656 606812 216708
rect 574928 216316 574980 216368
rect 625528 216316 625580 216368
rect 575296 216180 575348 216232
rect 627184 216180 627236 216232
rect 673368 216112 673420 216164
rect 675392 216112 675444 216164
rect 574928 216044 574980 216096
rect 628288 216044 628340 216096
rect 671988 215976 672040 216028
rect 574560 215908 574612 215960
rect 627920 215908 627972 215960
rect 672264 215568 672316 215620
rect 672172 215432 672224 215484
rect 672264 215228 672316 215280
rect 672356 215092 672408 215144
rect 672908 215092 672960 215144
rect 35532 214684 35584 214736
rect 39764 214684 39816 214736
rect 575112 214684 575164 214736
rect 612280 214684 612332 214736
rect 574744 214548 574796 214600
rect 597836 214412 597888 214464
rect 598480 214412 598532 214464
rect 598940 214412 598992 214464
rect 599584 214412 599636 214464
rect 600320 214412 600372 214464
rect 601240 214412 601292 214464
rect 609980 214548 610032 214600
rect 610624 214548 610676 214600
rect 618352 214548 618404 214600
rect 618904 214548 618956 214600
rect 624424 214412 624476 214464
rect 35808 214276 35860 214328
rect 40684 214276 40736 214328
rect 35348 213936 35400 213988
rect 40224 213936 40276 213988
rect 625160 213936 625212 213988
rect 626080 213936 626132 213988
rect 632704 213868 632756 213920
rect 633440 213868 633492 213920
rect 637212 213868 637264 213920
rect 650920 213868 650972 213920
rect 608324 213732 608376 213784
rect 609520 213732 609572 213784
rect 638868 213732 638920 213784
rect 652484 213732 652536 213784
rect 673092 213664 673144 213716
rect 675484 213664 675536 213716
rect 639972 213596 640024 213648
rect 652760 213596 652812 213648
rect 638316 213460 638368 213512
rect 651472 213460 651524 213512
rect 629944 213392 629996 213444
rect 633808 213392 633860 213444
rect 575480 213324 575532 213376
rect 594800 213324 594852 213376
rect 636660 213324 636712 213376
rect 650828 213324 650880 213376
rect 672908 213256 672960 213308
rect 675484 213256 675536 213308
rect 574376 213188 574428 213240
rect 629944 213188 629996 213240
rect 635556 213188 635608 213240
rect 650092 213188 650144 213240
rect 641536 213052 641588 213104
rect 651840 213052 651892 213104
rect 35808 212916 35860 212968
rect 39304 212984 39356 213036
rect 640248 212916 640300 212968
rect 651104 212916 651156 212968
rect 631416 212712 631468 212764
rect 632704 212712 632756 212764
rect 35808 212644 35860 212696
rect 39764 212644 39816 212696
rect 42156 212644 42208 212696
rect 50988 212644 51040 212696
rect 35624 212508 35676 212560
rect 41236 212576 41288 212628
rect 647240 212372 647292 212424
rect 648160 212372 648212 212424
rect 659660 212372 659712 212424
rect 660304 212372 660356 212424
rect 661316 212372 661368 212424
rect 661960 212372 662012 212424
rect 662420 212372 662472 212424
rect 663064 212372 663116 212424
rect 670976 212032 671028 212084
rect 675484 212032 675536 212084
rect 35808 211556 35860 211608
rect 41236 211556 41288 211608
rect 35808 211284 35860 211336
rect 39672 211352 39724 211404
rect 578332 211284 578384 211336
rect 580632 211284 580684 211336
rect 35624 211148 35676 211200
rect 41052 211216 41104 211268
rect 644480 211012 644532 211064
rect 644848 211012 644900 211064
rect 663800 211012 663852 211064
rect 664168 211012 664220 211064
rect 661776 210672 661828 210724
rect 672540 210672 672592 210724
rect 652208 210536 652260 210588
rect 667296 210536 667348 210588
rect 652024 210400 652076 210452
rect 673920 210400 673972 210452
rect 662144 210264 662196 210316
rect 667480 210264 667532 210316
rect 579528 210060 579580 210112
rect 582288 210060 582340 210112
rect 597560 210060 597612 210112
rect 597928 210060 597980 210112
rect 35624 209924 35676 209976
rect 41696 209924 41748 209976
rect 35808 209788 35860 209840
rect 40040 209788 40092 209840
rect 591304 209788 591356 209840
rect 632152 209788 632204 209840
rect 672264 209380 672316 209432
rect 672264 208904 672316 208956
rect 35808 208632 35860 208684
rect 39672 208564 39724 208616
rect 35624 208360 35676 208412
rect 39580 208360 39632 208412
rect 578884 208224 578936 208276
rect 589464 208224 589516 208276
rect 35808 207272 35860 207324
rect 39764 207272 39816 207324
rect 35532 207000 35584 207052
rect 40316 207000 40368 207052
rect 580632 206932 580684 206984
rect 589556 206932 589608 206984
rect 671712 206728 671764 206780
rect 671712 206592 671764 206644
rect 35808 205912 35860 205964
rect 39396 205912 39448 205964
rect 579528 205776 579580 205828
rect 581000 205776 581052 205828
rect 35624 205640 35676 205692
rect 41144 205640 41196 205692
rect 582288 205504 582340 205556
rect 589464 205504 589516 205556
rect 35808 204824 35860 204876
rect 39948 204824 40000 204876
rect 35624 204620 35676 204672
rect 41696 204552 41748 204604
rect 42064 204552 42116 204604
rect 44364 204552 44416 204604
rect 35532 204416 35584 204468
rect 41696 204416 41748 204468
rect 42064 204416 42116 204468
rect 47584 204416 47636 204468
rect 35808 204280 35860 204332
rect 41696 204280 41748 204332
rect 42064 204280 42116 204332
rect 48964 204280 49016 204332
rect 579712 204212 579764 204264
rect 589464 204212 589516 204264
rect 35624 203124 35676 203176
rect 41236 203192 41288 203244
rect 42064 202988 42116 203040
rect 50344 202988 50396 203040
rect 35808 202852 35860 202904
rect 41696 202852 41748 202904
rect 578332 202852 578384 202904
rect 580264 202852 580316 202904
rect 581000 202784 581052 202836
rect 589464 202784 589516 202836
rect 673368 201832 673420 201884
rect 675392 201832 675444 201884
rect 671988 201288 672040 201340
rect 675208 201288 675260 201340
rect 674840 200880 674892 200932
rect 675300 200880 675352 200932
rect 673092 200472 673144 200524
rect 675024 200472 675076 200524
rect 579160 200132 579212 200184
rect 590568 200132 590620 200184
rect 580264 199996 580316 200048
rect 589464 199996 589516 200048
rect 578884 197344 578936 197396
rect 589464 197344 589516 197396
rect 666928 196664 666980 196716
rect 667848 196664 667900 196716
rect 667664 196528 667716 196580
rect 667848 196324 667900 196376
rect 579528 195984 579580 196036
rect 589556 195984 589608 196036
rect 42432 195644 42484 195696
rect 43812 195644 43864 195696
rect 674472 194488 674524 194540
rect 675116 194488 675168 194540
rect 579528 193808 579580 193860
rect 589556 193808 589608 193860
rect 42432 193128 42484 193180
rect 43628 193128 43680 193180
rect 666928 192244 666980 192296
rect 669320 192244 669372 192296
rect 42432 191768 42484 191820
rect 44548 191768 44600 191820
rect 42432 191632 42484 191684
rect 44364 191632 44416 191684
rect 579528 191088 579580 191140
rect 589464 191088 589516 191140
rect 42432 190340 42484 190392
rect 42984 190340 43036 190392
rect 675852 189728 675904 189780
rect 683120 189728 683172 189780
rect 579528 188980 579580 189032
rect 589464 188980 589516 189032
rect 42432 187620 42484 187672
rect 43444 187620 43496 187672
rect 579528 186940 579580 186992
rect 589464 186940 589516 186992
rect 579436 184900 579488 184952
rect 589464 184900 589516 184952
rect 578516 184764 578568 184816
rect 589648 184764 589700 184816
rect 42432 183472 42484 183524
rect 44180 183472 44232 183524
rect 668216 183472 668268 183524
rect 670976 183472 671028 183524
rect 669228 182860 669280 182912
rect 672356 182860 672408 182912
rect 580908 182180 580960 182232
rect 589464 182180 589516 182232
rect 583116 180820 583168 180872
rect 589464 180820 589516 180872
rect 581736 179392 581788 179444
rect 589464 179392 589516 179444
rect 578332 179324 578384 179376
rect 580908 179324 580960 179376
rect 672540 178236 672592 178288
rect 675484 178236 675536 178288
rect 579712 178032 579764 178084
rect 589464 178032 589516 178084
rect 667112 178032 667164 178084
rect 675300 178032 675352 178084
rect 667940 177896 667992 177948
rect 673184 177896 673236 177948
rect 667756 176808 667808 176860
rect 675300 176808 675352 176860
rect 673276 176672 673328 176724
rect 675484 176672 675536 176724
rect 579528 176604 579580 176656
rect 583116 176604 583168 176656
rect 587164 175312 587216 175364
rect 589280 175312 589332 175364
rect 673092 175176 673144 175228
rect 675484 175176 675536 175228
rect 578700 174836 578752 174888
rect 581736 174836 581788 174888
rect 667940 174700 667992 174752
rect 669964 174700 670016 174752
rect 581736 173136 581788 173188
rect 589464 173136 589516 173188
rect 669412 171912 669464 171964
rect 675484 171912 675536 171964
rect 673368 171164 673420 171216
rect 675484 171164 675536 171216
rect 579804 171096 579856 171148
rect 589464 171096 589516 171148
rect 578884 170348 578936 170400
rect 587164 170348 587216 170400
rect 670608 170280 670660 170332
rect 675484 170280 675536 170332
rect 667940 169668 667992 169720
rect 670148 169668 670200 169720
rect 579252 169532 579304 169584
rect 581736 169532 581788 169584
rect 672356 169056 672408 169108
rect 675484 169056 675536 169108
rect 671988 168648 672040 168700
rect 675484 168648 675536 168700
rect 583024 168376 583076 168428
rect 589464 168376 589516 168428
rect 672540 168240 672592 168292
rect 675484 168240 675536 168292
rect 669964 167832 670016 167884
rect 675484 167832 675536 167884
rect 581644 167016 581696 167068
rect 589464 167016 589516 167068
rect 670976 166880 671028 166932
rect 675392 166880 675444 166932
rect 579528 166268 579580 166320
rect 589740 166268 589792 166320
rect 668032 164908 668084 164960
rect 670332 164908 670384 164960
rect 580264 164228 580316 164280
rect 589464 164228 589516 164280
rect 587348 162868 587400 162920
rect 589740 162868 589792 162920
rect 675852 162664 675904 162716
rect 678244 162664 678296 162716
rect 585968 160080 586020 160132
rect 589464 160080 589516 160132
rect 579528 159944 579580 159996
rect 588544 159944 588596 159996
rect 668584 158312 668636 158364
rect 674104 158312 674156 158364
rect 584404 157360 584456 157412
rect 589464 157360 589516 157412
rect 579252 157292 579304 157344
rect 583024 157292 583076 157344
rect 673368 156952 673420 157004
rect 675116 156952 675168 157004
rect 578700 155456 578752 155508
rect 581644 155456 581696 155508
rect 583208 154572 583260 154624
rect 589372 154572 589424 154624
rect 578332 153416 578384 153468
rect 580264 153416 580316 153468
rect 581828 153212 581880 153264
rect 589464 153212 589516 153264
rect 672356 153144 672408 153196
rect 675116 153144 675168 153196
rect 578424 152464 578476 152516
rect 590108 152464 590160 152516
rect 671988 151716 672040 151768
rect 675116 151716 675168 151768
rect 580632 151036 580684 151088
rect 589740 151036 589792 151088
rect 579528 150356 579580 150408
rect 587348 150356 587400 150408
rect 668768 150220 668820 150272
rect 671252 150220 671304 150272
rect 587164 149064 587216 149116
rect 589280 149064 589332 149116
rect 669412 148996 669464 149048
rect 675300 148996 675352 149048
rect 670608 147568 670660 147620
rect 675116 147568 675168 147620
rect 586888 146276 586940 146328
rect 589464 146276 589516 146328
rect 668768 145528 668820 145580
rect 671436 145528 671488 145580
rect 578792 145392 578844 145444
rect 585968 145392 586020 145444
rect 585784 144916 585836 144968
rect 589464 144916 589516 144968
rect 578884 144168 578936 144220
rect 586888 144168 586940 144220
rect 579252 143420 579304 143472
rect 588728 143420 588780 143472
rect 583760 140768 583812 140820
rect 589464 140768 589516 140820
rect 579528 140564 579580 140616
rect 584404 140564 584456 140616
rect 668676 140428 668728 140480
rect 671620 140428 671672 140480
rect 580264 140020 580316 140072
rect 590292 140020 590344 140072
rect 579068 138660 579120 138712
rect 589924 138660 589976 138712
rect 668768 138388 668820 138440
rect 674288 138388 674340 138440
rect 578332 137844 578384 137896
rect 583208 137844 583260 137896
rect 583024 137232 583076 137284
rect 589464 137232 589516 137284
rect 668768 136484 668820 136536
rect 671804 136484 671856 136536
rect 581644 135260 581696 135312
rect 589464 135260 589516 135312
rect 579344 135124 579396 135176
rect 581828 135124 581880 135176
rect 580448 133900 580500 133952
rect 589464 133900 589516 133952
rect 578332 133764 578384 133816
rect 580632 133764 580684 133816
rect 579252 133424 579304 133476
rect 583760 133424 583812 133476
rect 673920 132948 673972 133000
rect 675484 132948 675536 133000
rect 667480 132744 667532 132796
rect 675484 132744 675536 132796
rect 584772 132472 584824 132524
rect 589464 132472 589516 132524
rect 667296 132472 667348 132524
rect 675300 132472 675352 132524
rect 673368 131248 673420 131300
rect 675300 131248 675352 131300
rect 668768 131112 668820 131164
rect 675484 131112 675536 131164
rect 667940 130908 667992 130960
rect 669780 130908 669832 130960
rect 674104 130840 674156 130892
rect 675484 130840 675536 130892
rect 673092 130228 673144 130280
rect 675484 130228 675536 130280
rect 669136 129888 669188 129940
rect 675484 129888 675536 129940
rect 668584 129752 668636 129804
rect 669136 129752 669188 129804
rect 669228 129004 669280 129056
rect 672724 129004 672776 129056
rect 585968 128324 586020 128376
rect 589464 128324 589516 128376
rect 668952 128324 669004 128376
rect 675484 128324 675536 128376
rect 579528 128188 579580 128240
rect 587164 128188 587216 128240
rect 667940 126148 667992 126200
rect 669596 126148 669648 126200
rect 673184 125944 673236 125996
rect 675484 125944 675536 125996
rect 587348 125604 587400 125656
rect 589280 125604 589332 125656
rect 672724 125604 672776 125656
rect 675484 125604 675536 125656
rect 578424 124856 578476 124908
rect 588544 124856 588596 124908
rect 673920 124720 673972 124772
rect 675484 124720 675536 124772
rect 669228 124108 669280 124160
rect 672908 124108 672960 124160
rect 673368 122952 673420 123004
rect 675300 122952 675352 123004
rect 671344 122816 671396 122868
rect 675484 122816 675536 122868
rect 578884 122612 578936 122664
rect 585784 122612 585836 122664
rect 581828 121456 581880 121508
rect 589464 121456 589516 121508
rect 670148 121456 670200 121508
rect 675300 121456 675352 121508
rect 586152 120708 586204 120760
rect 589924 120708 589976 120760
rect 671528 120708 671580 120760
rect 675484 120708 675536 120760
rect 669136 119212 669188 119264
rect 672540 119212 672592 119264
rect 584588 118668 584640 118720
rect 589464 118668 589516 118720
rect 578516 118260 578568 118312
rect 580264 118260 580316 118312
rect 667940 117784 667992 117836
rect 669964 117784 670016 117836
rect 579068 117308 579120 117360
rect 589464 117308 589516 117360
rect 675852 117240 675904 117292
rect 679624 117240 679676 117292
rect 578884 115948 578936 116000
rect 589464 115948 589516 116000
rect 668400 115812 668452 115864
rect 670976 115812 671028 115864
rect 580632 115200 580684 115252
rect 590292 115200 590344 115252
rect 668400 114316 668452 114368
rect 671344 114316 671396 114368
rect 585784 113160 585836 113212
rect 589464 113160 589516 113212
rect 579528 113092 579580 113144
rect 583024 113092 583076 113144
rect 668032 112888 668084 112940
rect 670148 112888 670200 112940
rect 673184 111732 673236 111784
rect 675116 111732 675168 111784
rect 668768 111596 668820 111648
rect 671528 111596 671580 111648
rect 579528 111188 579580 111240
rect 586152 111188 586204 111240
rect 672724 111120 672776 111172
rect 675392 111120 675444 111172
rect 587164 110440 587216 110492
rect 589648 110440 589700 110492
rect 584404 109012 584456 109064
rect 589464 109012 589516 109064
rect 579252 108740 579304 108792
rect 581644 108740 581696 108792
rect 583208 107652 583260 107704
rect 589464 107652 589516 107704
rect 669228 107652 669280 107704
rect 674104 107652 674156 107704
rect 579252 107176 579304 107228
rect 584772 107176 584824 107228
rect 673920 106972 673972 107024
rect 675300 106972 675352 107024
rect 578332 106768 578384 106820
rect 580448 106768 580500 106820
rect 580264 106292 580316 106344
rect 589464 106292 589516 106344
rect 583024 104864 583076 104916
rect 589464 104864 589516 104916
rect 581644 103504 581696 103556
rect 589464 103504 589516 103556
rect 579528 103368 579580 103420
rect 591304 103368 591356 103420
rect 579528 99288 579580 99340
rect 588912 99288 588964 99340
rect 625068 99152 625120 99204
rect 634452 99152 634504 99204
rect 623688 99016 623740 99068
rect 632152 99016 632204 99068
rect 629760 98880 629812 98932
rect 640984 98880 641036 98932
rect 621664 98744 621716 98796
rect 628380 98744 628432 98796
rect 629024 98744 629076 98796
rect 640248 98744 640300 98796
rect 622308 98608 622360 98660
rect 629484 98608 629536 98660
rect 630496 98608 630548 98660
rect 642088 98608 642140 98660
rect 588544 97996 588596 98048
rect 589372 97996 589424 98048
rect 577504 97928 577556 97980
rect 594064 97928 594116 97980
rect 596180 97928 596232 97980
rect 620192 97928 620244 97980
rect 626080 97928 626132 97980
rect 626816 97928 626868 97980
rect 636384 97928 636436 97980
rect 592684 97792 592736 97844
rect 597560 97792 597612 97844
rect 625896 97792 625948 97844
rect 635280 97792 635332 97844
rect 643008 97792 643060 97844
rect 659752 97928 659804 97980
rect 659936 97928 659988 97980
rect 665732 97928 665784 97980
rect 647148 97792 647200 97844
rect 661960 97792 662012 97844
rect 595260 97656 595312 97708
rect 595628 97656 595680 97708
rect 623136 97656 623188 97708
rect 630680 97656 630732 97708
rect 632704 97656 632756 97708
rect 595444 97520 595496 97572
rect 598940 97520 598992 97572
rect 624608 97520 624660 97572
rect 632980 97520 633032 97572
rect 633348 97656 633400 97708
rect 643928 97656 643980 97708
rect 655428 97656 655480 97708
rect 662512 97656 662564 97708
rect 644756 97520 644808 97572
rect 627552 97384 627604 97436
rect 637580 97384 637632 97436
rect 639328 97384 639380 97436
rect 646504 97384 646556 97436
rect 658832 97520 658884 97572
rect 591304 97248 591356 97300
rect 600412 97248 600464 97300
rect 605472 97248 605524 97300
rect 611912 97248 611964 97300
rect 628196 97248 628248 97300
rect 639052 97248 639104 97300
rect 641536 97248 641588 97300
rect 643008 97248 643060 97300
rect 644296 97248 644348 97300
rect 658188 97384 658240 97436
rect 663064 97384 663116 97436
rect 656808 97248 656860 97300
rect 661408 97248 661460 97300
rect 654784 97180 654836 97232
rect 655244 97180 655296 97232
rect 634176 97112 634228 97164
rect 643468 97112 643520 97164
rect 656716 97044 656768 97096
rect 612648 96976 612700 97028
rect 613384 96976 613436 97028
rect 601700 96908 601752 96960
rect 602620 96908 602672 96960
rect 606208 96908 606260 96960
rect 606944 96908 606996 96960
rect 614028 96908 614080 96960
rect 614764 96908 614816 96960
rect 615776 96908 615828 96960
rect 616788 96908 616840 96960
rect 617248 96908 617300 96960
rect 617892 96908 617944 96960
rect 646688 96908 646740 96960
rect 647148 96908 647200 96960
rect 650368 96908 650420 96960
rect 658280 96908 658332 96960
rect 660120 96908 660172 96960
rect 609152 96840 609204 96892
rect 609704 96840 609756 96892
rect 612096 96840 612148 96892
rect 612648 96840 612700 96892
rect 618720 96840 618772 96892
rect 626264 96840 626316 96892
rect 613568 96772 613620 96824
rect 614028 96772 614080 96824
rect 651840 96772 651892 96824
rect 659568 96772 659620 96824
rect 578608 96568 578660 96620
rect 587348 96568 587400 96620
rect 635648 96568 635700 96620
rect 642824 96704 642876 96756
rect 645216 96704 645268 96756
rect 645768 96704 645820 96756
rect 651104 96636 651156 96688
rect 654324 96636 654376 96688
rect 642272 96568 642324 96620
rect 643284 96568 643336 96620
rect 638592 96432 638644 96484
rect 650920 96568 650972 96620
rect 653312 96432 653364 96484
rect 663984 96432 664036 96484
rect 631232 96296 631284 96348
rect 642640 96296 642692 96348
rect 642824 96296 642876 96348
rect 648804 96296 648856 96348
rect 652576 96296 652628 96348
rect 665364 96296 665416 96348
rect 620928 96228 620980 96280
rect 626448 96228 626500 96280
rect 631876 96160 631928 96212
rect 644480 96160 644532 96212
rect 648620 96160 648672 96212
rect 663800 96160 663852 96212
rect 586520 96024 586572 96076
rect 590108 96024 590160 96076
rect 610624 96024 610676 96076
rect 621664 96024 621716 96076
rect 637856 96024 637908 96076
rect 660672 96024 660724 96076
rect 608416 95888 608468 95940
rect 620284 95888 620336 95940
rect 640800 95888 640852 95940
rect 665180 95888 665232 95940
rect 640064 95752 640116 95804
rect 652024 95752 652076 95804
rect 634728 95616 634780 95668
rect 643100 95616 643152 95668
rect 645584 95616 645636 95668
rect 656164 95616 656216 95668
rect 659200 95616 659252 95668
rect 664168 95616 664220 95668
rect 616512 95140 616564 95192
rect 622676 95140 622728 95192
rect 643744 94596 643796 94648
rect 653404 94596 653456 94648
rect 607680 94460 607732 94512
rect 624976 94460 625028 94512
rect 642916 94460 642968 94512
rect 663248 94460 663300 94512
rect 649632 93984 649684 94036
rect 650644 93984 650696 94036
rect 579528 93780 579580 93832
rect 586520 93780 586572 93832
rect 619548 93780 619600 93832
rect 626448 93780 626500 93832
rect 643284 93780 643336 93832
rect 654140 93712 654192 93764
rect 609704 93100 609756 93152
rect 618904 93100 618956 93152
rect 618076 92420 618128 92472
rect 625436 92420 625488 92472
rect 650920 92420 650972 92472
rect 654324 92420 654376 92472
rect 579528 90992 579580 91044
rect 585968 90992 586020 91044
rect 611268 90992 611320 91044
rect 617340 90992 617392 91044
rect 617892 90992 617944 91044
rect 626448 90992 626500 91044
rect 646504 90992 646556 91044
rect 654140 90992 654192 91044
rect 622676 89632 622728 89684
rect 626448 89632 626500 89684
rect 578516 89564 578568 89616
rect 580632 89564 580684 89616
rect 647148 88952 647200 89004
rect 656900 88952 656952 89004
rect 656164 88748 656216 88800
rect 657452 88748 657504 88800
rect 662328 88748 662380 88800
rect 664168 88748 664220 88800
rect 607312 88272 607364 88324
rect 626448 88272 626500 88324
rect 655244 88272 655296 88324
rect 658464 88272 658516 88324
rect 617340 88136 617392 88188
rect 625620 88136 625672 88188
rect 656532 87252 656584 87304
rect 662512 87252 662564 87304
rect 645768 87116 645820 87168
rect 660672 87116 660724 87168
rect 648344 86980 648396 87032
rect 656532 86980 656584 87032
rect 579528 86912 579580 86964
rect 588728 86912 588780 86964
rect 656716 86912 656768 86964
rect 659568 86912 659620 86964
rect 653404 86708 653456 86760
rect 661408 86708 661460 86760
rect 652024 86572 652076 86624
rect 660120 86572 660172 86624
rect 650644 86436 650696 86488
rect 658832 86436 658884 86488
rect 621664 86232 621716 86284
rect 626448 86232 626500 86284
rect 609888 85484 609940 85536
rect 626448 85484 626500 85536
rect 620284 84124 620336 84176
rect 626264 84124 626316 84176
rect 579344 83988 579396 84040
rect 581828 83988 581880 84040
rect 618904 83988 618956 84040
rect 626448 83920 626500 83972
rect 579528 81336 579580 81388
rect 584588 81336 584640 81388
rect 628564 80928 628616 80980
rect 642456 80928 642508 80980
rect 612648 80792 612700 80844
rect 645860 80792 645912 80844
rect 595628 80656 595680 80708
rect 636108 80656 636160 80708
rect 579252 80044 579304 80096
rect 583208 80044 583260 80096
rect 629208 79432 629260 79484
rect 637488 79432 637540 79484
rect 616788 79296 616840 79348
rect 647424 79296 647476 79348
rect 637488 78208 637540 78260
rect 645308 78208 645360 78260
rect 631048 78072 631100 78124
rect 638960 78072 639012 78124
rect 614028 77936 614080 77988
rect 647608 77936 647660 77988
rect 624424 77392 624476 77444
rect 631048 77664 631100 77716
rect 628288 77528 628340 77580
rect 631508 77528 631560 77580
rect 625804 77392 625856 77444
rect 633900 77392 633952 77444
rect 577504 77256 577556 77308
rect 637120 77256 637172 77308
rect 639604 77256 639656 77308
rect 614764 76644 614816 76696
rect 646320 76644 646372 76696
rect 613384 76508 613436 76560
rect 648988 76508 649040 76560
rect 584588 75896 584640 75948
rect 628288 75896 628340 75948
rect 615408 75284 615460 75336
rect 646136 75284 646188 75336
rect 607128 75148 607180 75200
rect 646872 75148 646924 75200
rect 579528 74468 579580 74520
rect 589924 74468 589976 74520
rect 579528 71476 579580 71528
rect 584404 71476 584456 71528
rect 578516 68960 578568 69012
rect 587164 68960 587216 69012
rect 579528 67464 579580 67516
rect 585784 67464 585836 67516
rect 578516 61956 578568 62008
rect 580264 61956 580316 62008
rect 579528 58964 579580 59016
rect 583024 58964 583076 59016
rect 579068 57876 579120 57928
rect 581644 57876 581696 57928
rect 612004 57196 612056 57248
rect 662420 57196 662472 57248
rect 578516 55156 578568 55208
rect 588544 55156 588596 55208
rect 145380 53048 145432 53100
rect 584588 53048 584640 53100
rect 391940 52436 391992 52488
rect 392584 52436 392636 52488
rect 577504 52436 577556 52488
rect 288164 52300 288216 52352
rect 625804 52300 625856 52352
rect 405096 51688 405148 51740
rect 595444 51688 595496 51740
rect 235816 51008 235868 51060
rect 288164 51008 288216 51060
rect 340512 51008 340564 51060
rect 391940 51008 391992 51060
rect 445208 50464 445260 50516
rect 498108 50464 498160 50516
rect 183468 50328 183520 50380
rect 445024 50328 445076 50380
rect 498108 47268 498160 47320
rect 499580 47268 499632 47320
rect 194048 44820 194100 44872
rect 662604 44820 662656 44872
rect 315948 43392 316000 43444
rect 663800 43392 663852 43444
rect 409604 42340 409656 42392
rect 464896 42328 464948 42380
rect 315948 42173 316000 42225
<< metal2 >>
rect 110170 1029098 110262 1029126
rect 212934 1029098 213026 1029126
rect 264362 1029098 264454 1029126
rect 315974 1029098 316066 1029126
rect 366390 1029098 366482 1029126
rect 433734 1029098 433826 1029126
rect 510738 1029098 510830 1029126
rect 562166 1029098 562258 1029126
rect 110170 1028622 110262 1028650
rect 212934 1028622 213026 1028650
rect 264362 1028622 264454 1028650
rect 315974 1028622 316066 1028650
rect 366390 1028622 366482 1028650
rect 433734 1028622 433826 1028650
rect 510738 1028622 510830 1028650
rect 562166 1028622 562258 1028650
rect 110170 1028177 110262 1028205
rect 212934 1028177 213026 1028205
rect 264362 1028177 264454 1028205
rect 315974 1028177 316066 1028205
rect 366390 1028177 366482 1028205
rect 433734 1028177 433826 1028205
rect 510738 1028177 510830 1028205
rect 562166 1028177 562258 1028205
rect 366180 1027880 366232 1027886
rect 366180 1027822 366232 1027828
rect 366548 1027880 366600 1027886
rect 366548 1027822 366600 1027828
rect 110170 1027738 110262 1027766
rect 212934 1027738 213026 1027766
rect 264362 1027738 264454 1027766
rect 315974 1027738 316066 1027766
rect 366192 1027752 366220 1027822
rect 366560 1027752 366588 1027822
rect 433734 1027738 433826 1027766
rect 510738 1027738 510830 1027766
rect 562166 1027738 562258 1027766
rect 110170 1027262 110262 1027290
rect 212934 1027262 213026 1027290
rect 264362 1027262 264454 1027290
rect 315974 1027262 316066 1027290
rect 366390 1027262 366482 1027290
rect 433734 1027262 433826 1027290
rect 510738 1027262 510830 1027290
rect 562166 1027262 562258 1027290
rect 110170 1026786 110262 1026814
rect 212934 1026786 213026 1026814
rect 264362 1026786 264454 1026814
rect 315974 1026786 316066 1026814
rect 366390 1026786 366482 1026814
rect 433734 1026786 433826 1026814
rect 510738 1026786 510830 1026814
rect 562166 1026786 562258 1026814
rect 110170 1026310 110262 1026338
rect 212934 1026310 213026 1026338
rect 264362 1026310 264454 1026338
rect 315974 1026310 316066 1026338
rect 366284 1026202 366312 1026324
rect 366468 1026202 366496 1026324
rect 433734 1026310 433826 1026338
rect 510738 1026310 510830 1026338
rect 562166 1026310 562258 1026338
rect 366284 1026174 366496 1026202
rect 366284 1026038 366496 1026066
rect 110170 1025902 110262 1025930
rect 212934 1025902 213026 1025930
rect 264362 1025902 264454 1025930
rect 315974 1025902 316066 1025930
rect 366284 1025916 366312 1026038
rect 366468 1025916 366496 1026038
rect 433734 1025902 433826 1025930
rect 510738 1025902 510830 1025930
rect 562166 1025902 562258 1025930
rect 110170 1025426 110262 1025454
rect 212934 1025426 213026 1025454
rect 264362 1025426 264454 1025454
rect 315974 1025426 316066 1025454
rect 366390 1025426 366482 1025454
rect 433734 1025426 433826 1025454
rect 510738 1025426 510830 1025454
rect 562166 1025426 562258 1025454
rect 110170 1024950 110262 1024978
rect 212934 1024950 213026 1024978
rect 264362 1024950 264454 1024978
rect 315974 1024950 316066 1024978
rect 366390 1024950 366482 1024978
rect 433734 1024950 433826 1024978
rect 510738 1024950 510830 1024978
rect 562166 1024950 562258 1024978
rect 110170 1024474 110262 1024502
rect 212934 1024474 213026 1024502
rect 264362 1024474 264454 1024502
rect 315974 1024474 316066 1024502
rect 366192 1024418 366220 1024488
rect 366560 1024418 366588 1024488
rect 433734 1024474 433826 1024502
rect 510738 1024474 510830 1024502
rect 562166 1024474 562258 1024502
rect 366180 1024412 366232 1024418
rect 366180 1024354 366232 1024360
rect 366548 1024412 366600 1024418
rect 366548 1024354 366600 1024360
rect 110170 1024037 110262 1024065
rect 212934 1024037 213026 1024065
rect 264362 1024037 264454 1024065
rect 315974 1024037 316066 1024065
rect 366390 1024037 366482 1024065
rect 433734 1024037 433826 1024065
rect 510738 1024037 510830 1024065
rect 562166 1024037 562258 1024065
rect 110170 1023590 110262 1023618
rect 212934 1023590 213026 1023618
rect 264362 1023590 264454 1023618
rect 315974 1023590 316066 1023618
rect 366390 1023590 366482 1023618
rect 433734 1023590 433826 1023618
rect 510738 1023590 510830 1023618
rect 562166 1023590 562258 1023618
rect 504548 1007072 504600 1007078
rect 504546 1007040 504548 1007049
rect 514208 1007072 514260 1007078
rect 504600 1007040 504602 1007049
rect 514208 1007014 514260 1007020
rect 559654 1007040 559710 1007049
rect 504546 1006975 504602 1006984
rect 506204 1006936 506256 1006942
rect 151726 1006904 151782 1006913
rect 145748 1006868 145800 1006874
rect 151726 1006839 151728 1006848
rect 145748 1006810 145800 1006816
rect 151780 1006839 151782 1006848
rect 428002 1006904 428058 1006913
rect 506202 1006904 506204 1006913
rect 514024 1006936 514076 1006942
rect 506256 1006904 506258 1006913
rect 428002 1006839 428004 1006848
rect 151728 1006810 151780 1006816
rect 428056 1006839 428058 1006848
rect 439504 1006868 439556 1006874
rect 428004 1006810 428056 1006816
rect 514024 1006878 514076 1006884
rect 506202 1006839 506258 1006848
rect 439504 1006810 439556 1006816
rect 144552 1006596 144604 1006602
rect 144552 1006538 144604 1006544
rect 101126 1006496 101182 1006505
rect 94688 1006460 94740 1006466
rect 101126 1006431 101128 1006440
rect 94688 1006402 94740 1006408
rect 101180 1006431 101182 1006440
rect 101128 1006402 101180 1006408
rect 94504 1006324 94556 1006330
rect 94504 1006266 94556 1006272
rect 93124 1006188 93176 1006194
rect 93124 1006130 93176 1006136
rect 92664 999796 92716 999802
rect 92664 999738 92716 999744
rect 92296 998300 92348 998306
rect 92296 998242 92348 998248
rect 82266 995752 82322 995761
rect 82018 995710 82266 995738
rect 82266 995687 82322 995696
rect 81070 995480 81126 995489
rect 77036 995042 77064 995452
rect 77680 995178 77708 995452
rect 77668 995172 77720 995178
rect 77668 995114 77720 995120
rect 77024 995036 77076 995042
rect 77024 994978 77076 994984
rect 78324 994906 78352 995452
rect 78312 994900 78364 994906
rect 78312 994842 78364 994848
rect 80164 994809 80192 995452
rect 80730 995438 81070 995466
rect 86590 995480 86646 995489
rect 81070 995415 81126 995424
rect 80150 994800 80206 994809
rect 81360 994770 81388 995452
rect 84488 995217 84516 995452
rect 84474 995208 84530 995217
rect 84474 995143 84530 995152
rect 80150 994735 80206 994744
rect 81348 994764 81400 994770
rect 81348 994706 81400 994712
rect 85040 994265 85068 995452
rect 85684 994537 85712 995452
rect 86342 995438 86590 995466
rect 87538 995438 87828 995466
rect 86590 995415 86646 995424
rect 87800 995017 87828 995438
rect 87786 995008 87842 995017
rect 87786 994943 87842 994952
rect 85670 994528 85726 994537
rect 85670 994463 85726 994472
rect 88720 994294 88748 995452
rect 89378 995438 89668 995466
rect 90022 995438 90312 995466
rect 91218 995438 91692 995466
rect 89640 995382 89668 995438
rect 89628 995376 89680 995382
rect 89628 995318 89680 995324
rect 90284 994634 90312 995438
rect 91664 995330 91692 995438
rect 92308 995330 92336 998242
rect 92480 997756 92532 997762
rect 92480 997698 92532 997704
rect 92492 997642 92520 997698
rect 92400 997614 92520 997642
rect 92400 996418 92428 997614
rect 92676 997257 92704 999738
rect 92662 997248 92718 997257
rect 92662 997183 92718 997192
rect 92400 996390 92520 996418
rect 92492 995382 92520 996390
rect 93136 995489 93164 1006130
rect 93308 1006052 93360 1006058
rect 93308 1005994 93360 1006000
rect 93122 995480 93178 995489
rect 93122 995415 93178 995424
rect 91664 995302 92336 995330
rect 92480 995376 92532 995382
rect 92480 995318 92532 995324
rect 93320 994634 93348 1005994
rect 93674 995888 93730 995897
rect 93674 995823 93730 995832
rect 93688 995081 93716 995823
rect 93674 995072 93730 995081
rect 93674 995007 93730 995016
rect 90272 994628 90324 994634
rect 90272 994570 90324 994576
rect 93308 994628 93360 994634
rect 93308 994570 93360 994576
rect 88708 994288 88760 994294
rect 85026 994256 85082 994265
rect 94516 994265 94544 1006266
rect 94700 994537 94728 1006402
rect 100298 1006360 100354 1006369
rect 100298 1006295 100300 1006304
rect 100352 1006295 100354 1006304
rect 144184 1006324 144236 1006330
rect 100300 1006266 100352 1006272
rect 144184 1006266 144236 1006272
rect 99470 1006224 99526 1006233
rect 103978 1006224 104034 1006233
rect 99470 1006159 99472 1006168
rect 99524 1006159 99526 1006168
rect 102784 1006188 102836 1006194
rect 99472 1006130 99524 1006136
rect 103978 1006159 103980 1006168
rect 102784 1006130 102836 1006136
rect 104032 1006159 104034 1006168
rect 106830 1006224 106886 1006233
rect 106830 1006159 106832 1006168
rect 103980 1006130 104032 1006136
rect 106884 1006159 106886 1006168
rect 124864 1006188 124916 1006194
rect 106832 1006130 106884 1006136
rect 124864 1006130 124916 1006136
rect 98274 1006088 98330 1006097
rect 98274 1006023 98276 1006032
rect 98328 1006023 98330 1006032
rect 101404 1006052 101456 1006058
rect 98276 1005994 98328 1006000
rect 101404 1005994 101456 1006000
rect 94872 1004692 94924 1004698
rect 94872 1004634 94924 1004640
rect 94884 998306 94912 1004634
rect 97264 1002652 97316 1002658
rect 97264 1002594 97316 1002600
rect 96528 1002108 96580 1002114
rect 96528 1002050 96580 1002056
rect 96344 1001972 96396 1001978
rect 96344 1001914 96396 1001920
rect 94872 998300 94924 998306
rect 94872 998242 94924 998248
rect 94686 994528 94742 994537
rect 94686 994463 94742 994472
rect 88708 994230 88760 994236
rect 94502 994256 94558 994265
rect 85026 994191 85082 994200
rect 94502 994191 94558 994200
rect 51724 993064 51776 993070
rect 51724 993006 51776 993012
rect 46204 992928 46256 992934
rect 46204 992870 46256 992876
rect 42524 969468 42576 969474
rect 42524 969410 42576 969416
rect 41800 968833 41828 969272
rect 41786 968824 41842 968833
rect 41786 968759 41842 968768
rect 42182 968034 42288 968062
rect 41984 967201 42012 967405
rect 41970 967192 42026 967201
rect 41970 967127 42026 967136
rect 42260 966890 42288 968034
rect 42248 966884 42300 966890
rect 42248 966826 42300 966832
rect 42536 966770 42564 969410
rect 42708 966884 42760 966890
rect 42708 966826 42760 966832
rect 42182 966742 42564 966770
rect 42182 965551 42472 965579
rect 42444 964714 42472 965551
rect 42432 964708 42484 964714
rect 42432 964650 42484 964656
rect 42182 964362 42472 964390
rect 42444 963898 42472 964362
rect 42432 963892 42484 963898
rect 42432 963834 42484 963840
rect 42182 963711 42472 963739
rect 42444 963490 42472 963711
rect 42432 963484 42484 963490
rect 42432 963426 42484 963432
rect 42182 963070 42472 963098
rect 41800 962169 41828 962540
rect 41786 962160 41842 962169
rect 41786 962095 41842 962104
rect 42444 961926 42472 963070
rect 42432 961920 42484 961926
rect 42432 961862 42484 961868
rect 42168 960078 42288 960106
rect 42168 960024 42196 960078
rect 42260 960038 42288 960078
rect 42260 960010 42472 960038
rect 41800 959177 41828 959412
rect 41786 959168 41842 959177
rect 42444 959138 42472 960010
rect 41786 959103 41842 959112
rect 42432 959132 42484 959138
rect 42432 959074 42484 959080
rect 42168 958854 42288 958882
rect 42168 958732 42196 958854
rect 42260 958746 42288 958854
rect 42260 958718 42472 958746
rect 42168 958310 42288 958338
rect 42444 958322 42472 958718
rect 42168 958188 42196 958310
rect 42260 958202 42288 958310
rect 42432 958316 42484 958322
rect 42432 958258 42484 958264
rect 42260 958174 42380 958202
rect 41786 956584 41842 956593
rect 41786 956519 41842 956528
rect 41800 956352 41828 956519
rect 41800 955505 41828 955740
rect 41786 955496 41842 955505
rect 41786 955431 41842 955440
rect 42168 955182 42288 955210
rect 42168 955060 42196 955182
rect 42260 954122 42288 955182
rect 41708 954094 42288 954122
rect 35162 952912 35218 952921
rect 35162 952847 35218 952856
rect 8588 944180 8616 944316
rect 9048 944180 9076 944316
rect 9508 944180 9536 944316
rect 9968 944180 9996 944316
rect 10428 944180 10456 944316
rect 10888 944180 10916 944316
rect 11348 944180 11376 944316
rect 11808 944180 11836 944316
rect 12268 944180 12296 944316
rect 12728 944180 12756 944316
rect 13188 944180 13216 944316
rect 13648 944180 13676 944316
rect 14108 944180 14136 944316
rect 35176 937009 35204 952847
rect 41708 952270 41736 954094
rect 42352 953986 42380 958174
rect 42260 953958 42380 953986
rect 37924 952264 37976 952270
rect 41696 952264 41748 952270
rect 37924 952206 37976 952212
rect 39302 952232 39358 952241
rect 37936 938471 37964 952206
rect 41696 952206 41748 952212
rect 39302 952167 39358 952176
rect 37922 938462 37978 938471
rect 37922 938397 37978 938406
rect 39316 937417 39344 952167
rect 40038 951824 40094 951833
rect 40038 951759 40094 951768
rect 39302 937408 39358 937417
rect 39302 937343 39358 937352
rect 35162 937000 35218 937009
rect 35162 936935 35218 936944
rect 40052 935785 40080 951759
rect 41418 951688 41474 951697
rect 41418 951623 41474 951632
rect 41234 941896 41290 941905
rect 41234 941831 41290 941840
rect 41248 941526 41276 941831
rect 41236 941520 41288 941526
rect 41236 941462 41288 941468
rect 41234 941080 41290 941089
rect 41234 941015 41290 941024
rect 41248 940438 41276 941015
rect 41236 940432 41288 940438
rect 41236 940374 41288 940380
rect 41234 940264 41290 940273
rect 41234 940199 41290 940208
rect 41248 940030 41276 940199
rect 41236 940024 41288 940030
rect 41236 939966 41288 939972
rect 41050 939448 41106 939457
rect 41050 939383 41106 939392
rect 41064 938466 41092 939383
rect 41432 938602 41460 951623
rect 41696 941520 41748 941526
rect 41748 941468 42012 941474
rect 41696 941462 42012 941468
rect 41708 941446 42012 941462
rect 41604 940432 41656 940438
rect 41524 940380 41604 940386
rect 41524 940374 41656 940380
rect 41524 940358 41644 940374
rect 41524 939794 41552 940358
rect 41696 940024 41748 940030
rect 41696 939966 41748 939972
rect 41708 939794 41736 939966
rect 41984 939794 42012 941446
rect 41524 939766 41644 939794
rect 41708 939766 41920 939794
rect 41984 939766 42104 939794
rect 41236 938596 41288 938602
rect 41236 938538 41288 938544
rect 41420 938596 41472 938602
rect 41420 938538 41472 938544
rect 41248 938471 41276 938538
rect 41052 938460 41104 938466
rect 41052 938402 41104 938408
rect 41234 938462 41290 938471
rect 41234 938397 41290 938406
rect 41420 938460 41472 938466
rect 41420 938402 41472 938408
rect 40038 935776 40094 935785
rect 40038 935711 40094 935720
rect 40682 881920 40738 881929
rect 40682 881855 40738 881864
rect 40222 819088 40278 819097
rect 40222 819023 40278 819032
rect 39578 818680 39634 818689
rect 39578 818615 39634 818624
rect 8588 818380 8616 818516
rect 9048 818380 9076 818516
rect 9508 818380 9536 818516
rect 9968 818380 9996 818516
rect 10428 818380 10456 818516
rect 10888 818380 10916 818516
rect 11348 818380 11376 818516
rect 11808 818380 11836 818516
rect 12268 818380 12296 818516
rect 12728 818380 12756 818516
rect 13188 818380 13216 818516
rect 13648 818380 13676 818516
rect 14108 818380 14136 818516
rect 35622 818000 35678 818009
rect 35622 817935 35678 817944
rect 35636 817018 35664 817935
rect 35806 817320 35862 817329
rect 35806 817255 35862 817264
rect 35820 817154 35848 817255
rect 35808 817148 35860 817154
rect 35808 817090 35860 817096
rect 35624 817012 35676 817018
rect 35624 816954 35676 816960
rect 35438 816912 35494 816921
rect 35438 816847 35494 816856
rect 35452 815658 35480 816847
rect 35806 816504 35862 816513
rect 35806 816439 35862 816448
rect 35820 816270 35848 816439
rect 39592 816270 39620 818615
rect 39762 818000 39818 818009
rect 39762 817935 39818 817944
rect 35808 816264 35860 816270
rect 35808 816206 35860 816212
rect 39580 816264 39632 816270
rect 39580 816206 39632 816212
rect 35806 816096 35862 816105
rect 35806 816031 35862 816040
rect 35624 815992 35676 815998
rect 35624 815934 35676 815940
rect 35636 815697 35664 815934
rect 35820 815862 35848 816031
rect 35808 815856 35860 815862
rect 35808 815798 35860 815804
rect 35622 815688 35678 815697
rect 35440 815652 35492 815658
rect 35622 815623 35678 815632
rect 35440 815594 35492 815600
rect 35622 815280 35678 815289
rect 35622 815215 35678 815224
rect 35636 814298 35664 815215
rect 35806 814872 35862 814881
rect 35806 814807 35862 814816
rect 35820 814638 35848 814807
rect 35808 814632 35860 814638
rect 35808 814574 35860 814580
rect 39776 814570 39804 817935
rect 40236 817018 40264 819023
rect 40696 817154 40724 881855
rect 40684 817148 40736 817154
rect 40684 817090 40736 817096
rect 40224 817012 40276 817018
rect 40224 816954 40276 816960
rect 39764 814564 39816 814570
rect 39764 814506 39816 814512
rect 35806 814464 35862 814473
rect 35806 814399 35808 814408
rect 35860 814399 35862 814408
rect 35808 814370 35860 814376
rect 35624 814292 35676 814298
rect 35624 814234 35676 814240
rect 41050 814056 41106 814065
rect 41050 813991 41106 814000
rect 41064 813006 41092 813991
rect 41432 813006 41460 938402
rect 41616 930134 41644 939766
rect 41616 930106 41736 930134
rect 41708 815998 41736 930106
rect 41892 818009 41920 939766
rect 42076 818689 42104 939766
rect 42260 937825 42288 953958
rect 42720 953594 42748 966826
rect 42892 964708 42944 964714
rect 42892 964650 42944 964656
rect 42904 953594 42932 964650
rect 44180 963892 44232 963898
rect 44180 963834 44232 963840
rect 43076 963484 43128 963490
rect 43076 963426 43128 963432
rect 42352 953566 42748 953594
rect 42812 953566 42932 953594
rect 42352 939794 42380 953566
rect 42352 939766 42472 939794
rect 42246 937816 42302 937825
rect 42246 937751 42302 937760
rect 42444 932929 42472 939766
rect 42812 935377 42840 953566
rect 42798 935368 42854 935377
rect 42798 935303 42854 935312
rect 43088 934969 43116 963426
rect 43260 959132 43312 959138
rect 43260 959074 43312 959080
rect 43074 934960 43130 934969
rect 43074 934895 43130 934904
rect 43272 934561 43300 959074
rect 43536 946008 43588 946014
rect 43536 945950 43588 945956
rect 43548 943537 43576 945950
rect 43534 943528 43590 943537
rect 43534 943463 43590 943472
rect 43626 942304 43682 942313
rect 43626 942239 43682 942248
rect 43444 941384 43496 941390
rect 43442 941352 43444 941361
rect 43496 941352 43498 941361
rect 43442 941287 43498 941296
rect 43640 941254 43668 942239
rect 43628 941248 43680 941254
rect 43628 941190 43680 941196
rect 43442 939856 43498 939865
rect 43442 939791 43444 939800
rect 43496 939791 43498 939800
rect 43444 939762 43496 939768
rect 43258 934552 43314 934561
rect 43258 934487 43314 934496
rect 44192 933745 44220 963834
rect 44456 961920 44508 961926
rect 44456 961862 44508 961868
rect 44468 934153 44496 961862
rect 44640 958316 44692 958322
rect 44640 958258 44692 958264
rect 44652 949454 44680 958258
rect 44652 949426 44864 949454
rect 44638 943120 44694 943129
rect 44638 943055 44694 943064
rect 44652 937038 44680 943055
rect 44640 937032 44692 937038
rect 44640 936974 44692 936980
rect 44836 936193 44864 949426
rect 46216 940681 46244 992870
rect 50344 991500 50396 991506
rect 50344 991442 50396 991448
rect 48964 990140 49016 990146
rect 48964 990082 49016 990088
rect 47584 961920 47636 961926
rect 47584 961862 47636 961868
rect 47596 942721 47624 961862
rect 47582 942712 47638 942721
rect 47582 942647 47638 942656
rect 48976 941390 49004 990082
rect 48964 941384 49016 941390
rect 48964 941326 49016 941332
rect 50356 941254 50384 991442
rect 50344 941248 50396 941254
rect 50344 941190 50396 941196
rect 46202 940672 46258 940681
rect 46202 940607 46258 940616
rect 51736 939826 51764 993006
rect 73436 991636 73488 991642
rect 73436 991578 73488 991584
rect 73448 983620 73476 991578
rect 96356 987426 96384 1001914
rect 96344 987420 96396 987426
rect 96344 987362 96396 987368
rect 89628 985992 89680 985998
rect 89628 985934 89680 985940
rect 89640 983620 89668 985934
rect 96540 984638 96568 1002050
rect 97276 995178 97304 1002594
rect 98644 1002516 98696 1002522
rect 98644 1002458 98696 1002464
rect 97448 1002380 97500 1002386
rect 97448 1002322 97500 1002328
rect 97460 996033 97488 1002322
rect 98274 1002008 98330 1002017
rect 98274 1001943 98276 1001952
rect 98328 1001943 98330 1001952
rect 98276 1001914 98328 1001920
rect 97446 996024 97502 996033
rect 97446 995959 97502 995968
rect 97264 995172 97316 995178
rect 97264 995114 97316 995120
rect 98656 994770 98684 1002458
rect 100298 1002416 100354 1002425
rect 100298 1002351 100300 1002360
rect 100352 1002351 100354 1002360
rect 100300 1002322 100352 1002328
rect 101126 1002280 101182 1002289
rect 98828 1002244 98880 1002250
rect 101126 1002215 101128 1002224
rect 98828 1002186 98880 1002192
rect 101180 1002215 101182 1002224
rect 101128 1002186 101180 1002192
rect 98840 999802 98868 1002186
rect 99102 1002144 99158 1002153
rect 99102 1002079 99104 1002088
rect 99156 1002079 99158 1002088
rect 100208 1002108 100260 1002114
rect 99104 1002050 99156 1002056
rect 100208 1002050 100260 1002056
rect 100024 1001972 100076 1001978
rect 100024 1001914 100076 1001920
rect 98828 999796 98880 999802
rect 98828 999738 98880 999744
rect 100036 995081 100064 1001914
rect 100220 995353 100248 1002050
rect 100206 995344 100262 995353
rect 100206 995279 100262 995288
rect 100022 995072 100078 995081
rect 100022 995007 100078 995016
rect 101416 994906 101444 1005994
rect 102322 1002688 102378 1002697
rect 102322 1002623 102324 1002632
rect 102376 1002623 102378 1002632
rect 102324 1002594 102376 1002600
rect 101954 1002552 102010 1002561
rect 101954 1002487 101956 1002496
rect 102008 1002487 102010 1002496
rect 101956 1002458 102008 1002464
rect 101954 1002008 102010 1002017
rect 101954 1001943 101956 1001952
rect 102008 1001943 102010 1001952
rect 101956 1001914 102008 1001920
rect 102796 995042 102824 1006130
rect 104806 1006088 104862 1006097
rect 104806 1006023 104808 1006032
rect 104860 1006023 104862 1006032
rect 107658 1006088 107714 1006097
rect 107658 1006023 107660 1006032
rect 104808 1005994 104860 1006000
rect 107712 1006023 107714 1006032
rect 107660 1005994 107712 1006000
rect 103150 1004728 103206 1004737
rect 108486 1004728 108542 1004737
rect 103150 1004663 103152 1004672
rect 103204 1004663 103206 1004672
rect 106188 1004692 106240 1004698
rect 103152 1004634 103204 1004640
rect 108486 1004663 108488 1004672
rect 106188 1004634 106240 1004640
rect 108540 1004663 108542 1004672
rect 108488 1004634 108540 1004640
rect 106004 1002584 106056 1002590
rect 106002 1002552 106004 1002561
rect 106056 1002552 106058 1002561
rect 106002 1002487 106058 1002496
rect 105636 1002312 105688 1002318
rect 105634 1002280 105636 1002289
rect 105688 1002280 105690 1002289
rect 105634 1002215 105690 1002224
rect 104808 1002176 104860 1002182
rect 103150 1002144 103206 1002153
rect 103150 1002079 103152 1002088
rect 103204 1002079 103206 1002088
rect 104806 1002144 104808 1002153
rect 104860 1002144 104862 1002153
rect 104806 1002079 104862 1002088
rect 103152 1002050 103204 1002056
rect 106004 1002040 106056 1002046
rect 103978 1002008 104034 1002017
rect 103532 1001966 103978 1001994
rect 102784 995036 102836 995042
rect 102784 994978 102836 994984
rect 101404 994900 101456 994906
rect 101404 994842 101456 994848
rect 103532 994809 103560 1001966
rect 103978 1001943 104034 1001952
rect 106002 1002008 106004 1002017
rect 106056 1002008 106058 1002017
rect 106002 1001943 106058 1001952
rect 103518 994800 103574 994809
rect 98644 994764 98696 994770
rect 103518 994735 103574 994744
rect 98644 994706 98696 994712
rect 106200 992234 106228 1004634
rect 109500 1002584 109552 1002590
rect 109500 1002526 109552 1002532
rect 108028 1002448 108080 1002454
rect 108026 1002416 108028 1002425
rect 108080 1002416 108082 1002425
rect 108026 1002351 108082 1002360
rect 107844 1002312 107896 1002318
rect 108488 1002312 108540 1002318
rect 107844 1002254 107896 1002260
rect 108486 1002280 108488 1002289
rect 108540 1002280 108542 1002289
rect 106372 1002176 106424 1002182
rect 106832 1002176 106884 1002182
rect 106372 1002118 106424 1002124
rect 106830 1002144 106832 1002153
rect 106884 1002144 106886 1002153
rect 106384 997762 106412 1002118
rect 107856 1002130 107884 1002254
rect 108486 1002215 108542 1002224
rect 109040 1002176 109092 1002182
rect 107856 1002102 107976 1002130
rect 109040 1002118 109092 1002124
rect 106830 1002079 106886 1002088
rect 107752 1002040 107804 1002046
rect 107752 1001982 107804 1001988
rect 106372 997756 106424 997762
rect 106372 997698 106424 997704
rect 106924 996940 106976 996946
rect 106924 996882 106976 996888
rect 106108 992206 106228 992234
rect 96528 984632 96580 984638
rect 96528 984574 96580 984580
rect 106108 983634 106136 992206
rect 106936 985998 106964 996882
rect 107764 992934 107792 1001982
rect 107948 993070 107976 1002102
rect 108854 1002008 108910 1002017
rect 108854 1001943 108856 1001952
rect 108908 1001943 108910 1001952
rect 108856 1001914 108908 1001920
rect 107936 993064 107988 993070
rect 107936 993006 107988 993012
rect 107752 992928 107804 992934
rect 107752 992870 107804 992876
rect 109052 990146 109080 1002118
rect 109512 996130 109540 1002526
rect 110420 1002448 110472 1002454
rect 110420 1002390 110472 1002396
rect 109682 1002144 109738 1002153
rect 109682 1002079 109684 1002088
rect 109736 1002079 109738 1002088
rect 109684 1002050 109736 1002056
rect 109500 996124 109552 996130
rect 109500 996066 109552 996072
rect 110432 991506 110460 1002390
rect 111064 1002312 111116 1002318
rect 111064 1002254 111116 1002260
rect 111076 995450 111104 1002254
rect 111892 1002108 111944 1002114
rect 111892 1002050 111944 1002056
rect 111904 996946 111932 1002050
rect 112076 1001972 112128 1001978
rect 112076 1001914 112128 1001920
rect 111892 996940 111944 996946
rect 111892 996882 111944 996888
rect 111064 995444 111116 995450
rect 111064 995386 111116 995392
rect 112088 991642 112116 1001914
rect 124876 995858 124904 1006130
rect 126244 1006052 126296 1006058
rect 126244 1005994 126296 1006000
rect 126256 995994 126284 1005994
rect 126244 995988 126296 995994
rect 126244 995930 126296 995936
rect 124864 995852 124916 995858
rect 124864 995794 124916 995800
rect 133602 995752 133658 995761
rect 133446 995710 133602 995738
rect 139122 995752 139178 995761
rect 138966 995710 139122 995738
rect 133602 995687 133658 995696
rect 140962 995752 141018 995761
rect 140806 995710 140962 995738
rect 139122 995687 139178 995696
rect 142894 995752 142950 995761
rect 142646 995710 142894 995738
rect 140962 995687 141018 995696
rect 142894 995687 142950 995696
rect 143448 995580 143500 995586
rect 143448 995522 143500 995528
rect 128464 994838 128492 995452
rect 128452 994832 128504 994838
rect 128452 994774 128504 994780
rect 129108 994702 129136 995452
rect 129752 994974 129780 995452
rect 129740 994968 129792 994974
rect 129740 994910 129792 994916
rect 131592 994809 131620 995452
rect 131578 994800 131634 994809
rect 131578 994735 131634 994744
rect 129096 994696 129148 994702
rect 129096 994638 129148 994644
rect 132144 994430 132172 995452
rect 132788 994537 132816 995452
rect 135916 994566 135944 995452
rect 135904 994560 135956 994566
rect 132774 994528 132830 994537
rect 135904 994502 135956 994508
rect 132774 994463 132830 994472
rect 132132 994424 132184 994430
rect 132132 994366 132184 994372
rect 121736 994288 121788 994294
rect 136468 994265 136496 995452
rect 137112 995081 137140 995452
rect 137770 995438 137968 995466
rect 137940 995178 137968 995438
rect 137928 995172 137980 995178
rect 137928 995114 137980 995120
rect 137098 995072 137154 995081
rect 137098 995007 137154 995016
rect 140148 994294 140176 995452
rect 141450 995438 141832 995466
rect 141804 995353 141832 995438
rect 141790 995344 141846 995353
rect 141790 995279 141846 995288
rect 142068 995308 142120 995314
rect 142068 995250 142120 995256
rect 142080 994566 142108 995250
rect 142068 994560 142120 994566
rect 142068 994502 142120 994508
rect 143460 994430 143488 995522
rect 144196 995178 144224 1006266
rect 144368 997348 144420 997354
rect 144368 997290 144420 997296
rect 144380 996713 144408 997290
rect 144366 996704 144422 996713
rect 144366 996639 144422 996648
rect 144564 995450 144592 1006538
rect 145564 1006188 145616 1006194
rect 145564 1006130 145616 1006136
rect 144828 997756 144880 997762
rect 144828 997698 144880 997704
rect 144840 996441 144868 997698
rect 144826 996432 144882 996441
rect 144826 996367 144882 996376
rect 144552 995444 144604 995450
rect 144552 995386 144604 995392
rect 144184 995172 144236 995178
rect 144184 995114 144236 995120
rect 143448 994424 143500 994430
rect 143448 994366 143500 994372
rect 140136 994288 140188 994294
rect 121736 994230 121788 994236
rect 136454 994256 136510 994265
rect 112076 991636 112128 991642
rect 112076 991578 112128 991584
rect 110420 991500 110472 991506
rect 110420 991442 110472 991448
rect 109040 990140 109092 990146
rect 109040 990082 109092 990088
rect 106924 985992 106976 985998
rect 106924 985934 106976 985940
rect 105846 983606 106136 983634
rect 121748 983634 121776 994230
rect 145576 994265 145604 1006130
rect 145760 996985 145788 1006810
rect 307758 1006768 307814 1006777
rect 300124 1006732 300176 1006738
rect 307758 1006703 307760 1006712
rect 300124 1006674 300176 1006680
rect 307812 1006703 307814 1006712
rect 357714 1006768 357770 1006777
rect 430854 1006768 430910 1006777
rect 357714 1006703 357716 1006712
rect 307760 1006674 307812 1006680
rect 357768 1006703 357770 1006712
rect 374000 1006732 374052 1006738
rect 357716 1006674 357768 1006680
rect 374000 1006674 374052 1006680
rect 400864 1006732 400916 1006738
rect 430854 1006703 430856 1006712
rect 400864 1006674 400916 1006680
rect 430908 1006703 430910 1006712
rect 430856 1006674 430908 1006680
rect 151452 1006596 151504 1006602
rect 151452 1006538 151504 1006544
rect 298744 1006596 298796 1006602
rect 298744 1006538 298796 1006544
rect 148324 1006460 148376 1006466
rect 148324 1006402 148376 1006408
rect 146942 1006088 146998 1006097
rect 146942 1006023 146998 1006032
rect 146956 1001894 146984 1006023
rect 147588 1001972 147640 1001978
rect 147588 1001914 147640 1001920
rect 146772 1001866 146984 1001894
rect 145746 996976 145802 996985
rect 145746 996911 145802 996920
rect 146772 995353 146800 1001866
rect 146944 995580 146996 995586
rect 146944 995522 146996 995528
rect 146758 995344 146814 995353
rect 146956 995314 146984 995522
rect 146758 995279 146814 995288
rect 146944 995308 146996 995314
rect 146944 995250 146996 995256
rect 140136 994230 140188 994236
rect 145562 994256 145618 994265
rect 136454 994191 136510 994200
rect 145562 994191 145618 994200
rect 147600 992934 147628 1001914
rect 148336 995081 148364 1006402
rect 150898 1006360 150954 1006369
rect 150898 1006295 150900 1006304
rect 150952 1006295 150954 1006304
rect 150900 1006266 150952 1006272
rect 151266 1006224 151322 1006233
rect 151464 1006194 151492 1006538
rect 255318 1006496 255374 1006505
rect 249064 1006460 249116 1006466
rect 255318 1006431 255320 1006440
rect 249064 1006402 249116 1006408
rect 255372 1006431 255374 1006440
rect 255320 1006402 255372 1006408
rect 152096 1006392 152148 1006398
rect 152094 1006360 152096 1006369
rect 210424 1006392 210476 1006398
rect 152148 1006360 152150 1006369
rect 152094 1006295 152150 1006304
rect 158258 1006360 158314 1006369
rect 158258 1006295 158260 1006304
rect 158312 1006295 158314 1006304
rect 210422 1006360 210424 1006369
rect 228364 1006392 228416 1006398
rect 210476 1006360 210478 1006369
rect 228364 1006334 228416 1006340
rect 210422 1006295 210478 1006304
rect 158260 1006266 158312 1006272
rect 208400 1006256 208452 1006262
rect 159454 1006224 159510 1006233
rect 151266 1006159 151268 1006168
rect 151320 1006159 151322 1006168
rect 151452 1006188 151504 1006194
rect 151268 1006130 151320 1006136
rect 159454 1006159 159456 1006168
rect 151452 1006130 151504 1006136
rect 159508 1006159 159510 1006168
rect 160282 1006224 160338 1006233
rect 208398 1006224 208400 1006233
rect 208452 1006224 208454 1006233
rect 160282 1006159 160284 1006168
rect 159456 1006130 159508 1006136
rect 160336 1006159 160338 1006168
rect 164884 1006188 164936 1006194
rect 160284 1006130 160336 1006136
rect 164884 1006130 164936 1006136
rect 175924 1006188 175976 1006194
rect 208398 1006159 208454 1006168
rect 175924 1006130 175976 1006136
rect 148874 1006088 148930 1006097
rect 148874 1006023 148876 1006032
rect 148928 1006023 148930 1006032
rect 150070 1006088 150126 1006097
rect 150070 1006023 150072 1006032
rect 148876 1005994 148928 1006000
rect 150124 1006023 150126 1006032
rect 158626 1006088 158682 1006097
rect 158626 1006023 158628 1006032
rect 150072 1005994 150124 1006000
rect 158680 1006023 158682 1006032
rect 158628 1005994 158680 1006000
rect 152922 1005272 152978 1005281
rect 149704 1005236 149756 1005242
rect 152922 1005207 152924 1005216
rect 149704 1005178 149756 1005184
rect 152976 1005207 152978 1005216
rect 152924 1005178 152976 1005184
rect 148968 1002108 149020 1002114
rect 148968 1002050 149020 1002056
rect 148322 995072 148378 995081
rect 148322 995007 148378 995016
rect 148980 993070 149008 1002050
rect 149242 1002008 149298 1002017
rect 149242 1001943 149244 1001952
rect 149296 1001943 149298 1001952
rect 149244 1001914 149296 1001920
rect 149716 994537 149744 1005178
rect 153750 1005136 153806 1005145
rect 151084 1005100 151136 1005106
rect 153750 1005071 153752 1005080
rect 151084 1005042 151136 1005048
rect 153804 1005071 153806 1005080
rect 153752 1005042 153804 1005048
rect 149888 1004964 149940 1004970
rect 149888 1004906 149940 1004912
rect 149900 997354 149928 1004906
rect 150898 1002144 150954 1002153
rect 150898 1002079 150900 1002088
rect 150952 1002079 150954 1002088
rect 150900 1002050 150952 1002056
rect 149888 997348 149940 997354
rect 149888 997290 149940 997296
rect 151096 994702 151124 1005042
rect 152922 1005000 152978 1005009
rect 160650 1005000 160706 1005009
rect 152922 1004935 152924 1004944
rect 152976 1004935 152978 1004944
rect 154396 1004964 154448 1004970
rect 152924 1004906 152976 1004912
rect 160650 1004935 160652 1004944
rect 154396 1004906 154448 1004912
rect 160704 1004935 160706 1004944
rect 160652 1004906 160704 1004912
rect 154118 1004864 154174 1004873
rect 151268 1004828 151320 1004834
rect 154118 1004799 154120 1004808
rect 151268 1004770 151320 1004776
rect 154172 1004799 154174 1004808
rect 154120 1004770 154172 1004776
rect 151280 995761 151308 1004770
rect 153936 1002312 153988 1002318
rect 153936 1002254 153988 1002260
rect 152648 1002176 152700 1002182
rect 152648 1002118 152700 1002124
rect 152464 1002040 152516 1002046
rect 152464 1001982 152516 1001988
rect 151266 995752 151322 995761
rect 151266 995687 151322 995696
rect 152476 995314 152504 1001982
rect 152660 995450 152688 1002118
rect 153752 1002040 153804 1002046
rect 153750 1002008 153752 1002017
rect 153804 1002008 153806 1002017
rect 153750 1001943 153806 1001952
rect 153948 997762 153976 1002254
rect 153936 997756 153988 997762
rect 153936 997698 153988 997704
rect 152648 995444 152700 995450
rect 152648 995386 152700 995392
rect 152464 995308 152516 995314
rect 152464 995250 152516 995256
rect 151084 994696 151136 994702
rect 151084 994638 151136 994644
rect 149702 994528 149758 994537
rect 149702 994463 149758 994472
rect 148968 993064 149020 993070
rect 148968 993006 149020 993012
rect 147588 992928 147640 992934
rect 147588 992870 147640 992876
rect 154408 992234 154436 1004906
rect 159454 1004864 159510 1004873
rect 159454 1004799 159456 1004808
rect 159508 1004799 159510 1004808
rect 162124 1004828 162176 1004834
rect 159456 1004770 159508 1004776
rect 162124 1004770 162176 1004776
rect 160650 1004728 160706 1004737
rect 160650 1004663 160652 1004672
rect 160704 1004663 160706 1004672
rect 160652 1004634 160704 1004640
rect 157430 1002552 157486 1002561
rect 157430 1002487 157432 1002496
rect 157484 1002487 157486 1002496
rect 159364 1002516 159416 1002522
rect 157432 1002458 157484 1002464
rect 159364 1002458 159416 1002464
rect 158626 1002416 158682 1002425
rect 158626 1002351 158628 1002360
rect 158680 1002351 158682 1002360
rect 158628 1002322 158680 1002328
rect 155776 1002312 155828 1002318
rect 155774 1002280 155776 1002289
rect 155828 1002280 155830 1002289
rect 155774 1002215 155830 1002224
rect 156602 1002280 156658 1002289
rect 156602 1002215 156604 1002224
rect 156656 1002215 156658 1002224
rect 158720 1002244 158772 1002250
rect 156604 1002186 156656 1002192
rect 158720 1002186 158772 1002192
rect 154580 1002176 154632 1002182
rect 154578 1002144 154580 1002153
rect 154632 1002144 154634 1002153
rect 154578 1002079 154634 1002088
rect 154946 1002144 155002 1002153
rect 154946 1002079 154948 1002088
rect 155000 1002079 155002 1002088
rect 157340 1002108 157392 1002114
rect 154948 1002050 155000 1002056
rect 157340 1002050 157392 1002056
rect 155774 1002008 155830 1002017
rect 154580 1001972 154632 1001978
rect 156602 1002008 156658 1002017
rect 155774 1001943 155776 1001952
rect 154580 1001914 154632 1001920
rect 155828 1001943 155830 1001952
rect 155972 1001966 156602 1001994
rect 155776 1001914 155828 1001920
rect 154592 994838 154620 1001914
rect 155972 994974 156000 1001966
rect 156602 1001943 156658 1001952
rect 155960 994968 156012 994974
rect 155960 994910 156012 994916
rect 154580 994832 154632 994838
rect 157352 994809 157380 1002050
rect 157798 1002008 157854 1002017
rect 157798 1001943 157800 1001952
rect 157852 1001943 157854 1001952
rect 157800 1001914 157852 1001920
rect 158732 996130 158760 1002186
rect 159376 996130 159404 1002458
rect 160376 1002380 160428 1002386
rect 160376 1002322 160428 1002328
rect 160192 1001972 160244 1001978
rect 160192 1001914 160244 1001920
rect 158720 996124 158772 996130
rect 158720 996066 158772 996072
rect 159364 996124 159416 996130
rect 159364 996066 159416 996072
rect 160204 995858 160232 1001914
rect 160388 995994 160416 1002322
rect 162136 995994 162164 1004770
rect 162860 1004692 162912 1004698
rect 162860 1004634 162912 1004640
rect 160376 995988 160428 995994
rect 160376 995930 160428 995936
rect 162124 995988 162176 995994
rect 162124 995930 162176 995936
rect 160192 995852 160244 995858
rect 160192 995794 160244 995800
rect 154580 994774 154632 994780
rect 157338 994800 157394 994809
rect 157338 994735 157394 994744
rect 154408 992206 154528 992234
rect 138296 991500 138348 991506
rect 138296 991442 138348 991448
rect 121748 983606 122130 983634
rect 138308 983620 138336 991442
rect 154500 983620 154528 992206
rect 162872 991506 162900 1004634
rect 164896 997694 164924 1006130
rect 164884 997688 164936 997694
rect 164884 997630 164936 997636
rect 170312 997688 170364 997694
rect 170312 997630 170364 997636
rect 162860 991500 162912 991506
rect 162860 991442 162912 991448
rect 170324 983634 170352 997630
rect 175936 995858 175964 1006130
rect 201038 1006088 201094 1006097
rect 177304 1006052 177356 1006058
rect 177304 1005994 177356 1006000
rect 198004 1006052 198056 1006058
rect 201038 1006023 201040 1006032
rect 198004 1005994 198056 1006000
rect 201092 1006023 201094 1006032
rect 201040 1005994 201092 1006000
rect 175924 995852 175976 995858
rect 175924 995794 175976 995800
rect 177316 995081 177344 1005994
rect 195336 1001972 195388 1001978
rect 195336 1001914 195388 1001920
rect 195152 997824 195204 997830
rect 195152 997766 195204 997772
rect 195164 997665 195192 997766
rect 195150 997656 195206 997665
rect 195150 997591 195206 997600
rect 195348 995761 195376 1001914
rect 195980 999184 196032 999190
rect 195980 999126 196032 999132
rect 195520 998436 195572 998442
rect 195520 998378 195572 998384
rect 184478 995752 184534 995761
rect 187514 995752 187570 995761
rect 184534 995710 184828 995738
rect 187312 995710 187514 995738
rect 184478 995687 184534 995696
rect 189538 995752 189594 995761
rect 189152 995710 189538 995738
rect 187514 995687 187570 995696
rect 190458 995752 190514 995761
rect 190348 995710 190458 995738
rect 189538 995687 189594 995696
rect 190458 995687 190514 995696
rect 195334 995752 195390 995761
rect 195334 995687 195390 995696
rect 195244 995580 195296 995586
rect 195244 995522 195296 995528
rect 183834 995480 183890 995489
rect 179860 995438 180196 995466
rect 180504 995438 180656 995466
rect 181148 995438 181484 995466
rect 182988 995438 183324 995466
rect 183540 995438 183834 995466
rect 177302 995072 177358 995081
rect 177302 995007 177358 995016
rect 180168 994906 180196 995438
rect 180156 994900 180208 994906
rect 180156 994842 180208 994848
rect 180628 994770 180656 995438
rect 181456 995042 181484 995438
rect 181444 995036 181496 995042
rect 181444 994978 181496 994984
rect 180616 994764 180668 994770
rect 180616 994706 180668 994712
rect 180614 994528 180670 994537
rect 183296 994498 183324 995438
rect 192482 995480 192538 995489
rect 184184 995438 184520 995466
rect 187864 995438 188200 995466
rect 188508 995438 188844 995466
rect 191544 995438 191788 995466
rect 192188 995438 192482 995466
rect 183834 995415 183890 995424
rect 184492 994809 184520 995438
rect 184478 994800 184534 994809
rect 184478 994735 184534 994744
rect 180614 994463 180616 994472
rect 180668 994463 180670 994472
rect 183284 994492 183336 994498
rect 180616 994434 180668 994440
rect 183284 994434 183336 994440
rect 186504 994288 186556 994294
rect 186504 994230 186556 994236
rect 186516 983634 186544 994230
rect 188172 993993 188200 995438
rect 188816 994537 188844 995438
rect 188802 994528 188858 994537
rect 188802 994463 188858 994472
rect 188158 993984 188214 993993
rect 188158 993919 188214 993928
rect 191760 993177 191788 995438
rect 192832 995438 193168 995466
rect 194028 995438 194364 995466
rect 192482 995415 192538 995424
rect 193140 994809 193168 995438
rect 194336 995382 194364 995438
rect 194324 995376 194376 995382
rect 194324 995318 194376 995324
rect 192942 994800 192998 994809
rect 192942 994735 192998 994744
rect 193126 994800 193182 994809
rect 193126 994735 193182 994744
rect 192956 994265 192984 994735
rect 195256 994498 195284 995522
rect 195532 995382 195560 998378
rect 195520 995376 195572 995382
rect 195520 995318 195572 995324
rect 195992 994634 196020 999126
rect 196624 998572 196676 998578
rect 196624 998514 196676 998520
rect 195980 994628 196032 994634
rect 195980 994570 196032 994576
rect 195244 994492 195296 994498
rect 195244 994434 195296 994440
rect 192942 994256 192998 994265
rect 192942 994191 192998 994200
rect 196636 993993 196664 998514
rect 198016 994809 198044 1005994
rect 209226 1005000 209282 1005009
rect 209226 1004935 209228 1004944
rect 209280 1004935 209282 1004944
rect 211804 1004964 211856 1004970
rect 209228 1004906 209280 1004912
rect 211804 1004906 211856 1004912
rect 207202 1004864 207258 1004873
rect 207202 1004799 207204 1004808
rect 207256 1004799 207258 1004808
rect 209872 1004828 209924 1004834
rect 207204 1004770 207256 1004776
rect 209872 1004770 209924 1004776
rect 209226 1004728 209282 1004737
rect 209226 1004663 209228 1004672
rect 209280 1004663 209282 1004672
rect 209228 1004634 209280 1004640
rect 206374 1002552 206430 1002561
rect 203340 1002516 203392 1002522
rect 206374 1002487 206376 1002496
rect 203340 1002458 203392 1002464
rect 206428 1002487 206430 1002496
rect 206376 1002458 206428 1002464
rect 199844 998844 199896 998850
rect 199844 998786 199896 998792
rect 199384 998708 199436 998714
rect 199384 998650 199436 998656
rect 198648 997960 198700 997966
rect 198648 997902 198700 997908
rect 198002 994800 198058 994809
rect 198002 994735 198058 994744
rect 196622 993984 196678 993993
rect 196622 993919 196678 993928
rect 191746 993168 191802 993177
rect 191746 993103 191802 993112
rect 198660 991642 198688 997902
rect 199396 994265 199424 998650
rect 199856 996441 199884 998786
rect 202694 998608 202750 998617
rect 202694 998543 202696 998552
rect 202748 998543 202750 998552
rect 202696 998514 202748 998520
rect 202144 998232 202196 998238
rect 202144 998174 202196 998180
rect 200672 997960 200724 997966
rect 200670 997928 200672 997937
rect 200856 997960 200908 997966
rect 200724 997928 200726 997937
rect 200856 997902 200908 997908
rect 200670 997863 200726 997872
rect 200028 997824 200080 997830
rect 200028 997766 200080 997772
rect 199842 996432 199898 996441
rect 199842 996367 199898 996376
rect 199382 994256 199438 994265
rect 199382 994191 199438 994200
rect 198648 991636 198700 991642
rect 198648 991578 198700 991584
rect 200040 991506 200068 997766
rect 200868 997754 200896 997902
rect 201868 997824 201920 997830
rect 200776 997726 200896 997754
rect 201866 997792 201868 997801
rect 201920 997792 201922 997801
rect 201866 997727 201922 997736
rect 200212 997280 200264 997286
rect 200210 997248 200212 997257
rect 200264 997248 200266 997257
rect 200210 997183 200266 997192
rect 200776 994537 200804 997726
rect 202156 994770 202184 998174
rect 202696 998096 202748 998102
rect 202694 998064 202696 998073
rect 202748 998064 202750 998073
rect 202694 997999 202750 998008
rect 202328 997824 202380 997830
rect 202328 997766 202380 997772
rect 202340 995489 202368 997766
rect 203352 997286 203380 1002458
rect 206374 1002280 206430 1002289
rect 204904 1002244 204956 1002250
rect 206374 1002215 206376 1002224
rect 204904 1002186 204956 1002192
rect 206428 1002215 206430 1002224
rect 206376 1002186 206428 1002192
rect 203890 1002008 203946 1002017
rect 203890 1001943 203892 1001952
rect 203944 1001943 203946 1001952
rect 204168 1001972 204220 1001978
rect 203892 1001914 203944 1001920
rect 204168 1001914 204220 1001920
rect 203524 999184 203576 999190
rect 203522 999152 203524 999161
rect 203576 999152 203578 999161
rect 203522 999087 203578 999096
rect 204180 998442 204208 1001914
rect 204350 998744 204406 998753
rect 204350 998679 204352 998688
rect 204404 998679 204406 998688
rect 204352 998650 204404 998656
rect 204168 998436 204220 998442
rect 204168 998378 204220 998384
rect 203524 997960 203576 997966
rect 203522 997928 203524 997937
rect 203576 997928 203578 997937
rect 203522 997863 203578 997872
rect 204720 997824 204772 997830
rect 204718 997792 204720 997801
rect 204772 997792 204774 997801
rect 204718 997727 204774 997736
rect 203340 997280 203392 997286
rect 203340 997222 203392 997228
rect 204916 995586 204944 1002186
rect 207202 1002144 207258 1002153
rect 206296 1002102 207202 1002130
rect 205546 1002008 205602 1002017
rect 205546 1001943 205548 1001952
rect 205600 1001943 205602 1001952
rect 205548 1001914 205600 1001920
rect 206296 998578 206324 1002102
rect 207202 1002079 207258 1002088
rect 207570 1002008 207626 1002017
rect 207032 1001966 207570 1001994
rect 206284 998572 206336 998578
rect 206284 998514 206336 998520
rect 205548 998232 205600 998238
rect 205546 998200 205548 998209
rect 205600 998200 205602 998209
rect 205546 998135 205602 998144
rect 204904 995580 204956 995586
rect 204904 995522 204956 995528
rect 202326 995480 202382 995489
rect 202326 995415 202382 995424
rect 207032 995042 207060 1001966
rect 207570 1001943 207626 1001952
rect 208398 1002008 208454 1002017
rect 208398 1001943 208454 1001952
rect 208412 996130 208440 1001943
rect 208400 996124 208452 996130
rect 208400 996066 208452 996072
rect 207020 995036 207072 995042
rect 207020 994978 207072 994984
rect 209884 994906 209912 1004770
rect 211160 1004692 211212 1004698
rect 211160 1004634 211212 1004640
rect 211172 1002538 211200 1004634
rect 211080 1002510 211200 1002538
rect 210422 1002008 210478 1002017
rect 210068 1001966 210422 1001994
rect 210068 995994 210096 1001966
rect 211080 1001994 211108 1002510
rect 211250 1002416 211306 1002425
rect 211250 1002351 211252 1002360
rect 211304 1002351 211306 1002360
rect 211252 1002322 211304 1002328
rect 211250 1002144 211306 1002153
rect 211250 1002079 211252 1002088
rect 211304 1002079 211306 1002088
rect 211252 1002050 211304 1002056
rect 211080 1001966 211200 1001994
rect 210422 1001943 210478 1001952
rect 210056 995988 210108 995994
rect 210056 995930 210108 995936
rect 211172 995858 211200 1001966
rect 211160 995852 211212 995858
rect 211160 995794 211212 995800
rect 211816 995450 211844 1004906
rect 212538 1004728 212594 1004737
rect 212538 1004663 212540 1004672
rect 212592 1004663 212594 1004672
rect 217324 1004692 217376 1004698
rect 212540 1004634 212592 1004640
rect 217324 1004634 217376 1004640
rect 215944 1002380 215996 1002386
rect 215944 1002322 215996 1002328
rect 213184 1002108 213236 1002114
rect 213184 1002050 213236 1002056
rect 212078 1002008 212134 1002017
rect 212078 1001943 212080 1001952
rect 212132 1001943 212134 1001952
rect 212080 1001914 212132 1001920
rect 213196 995994 213224 1002050
rect 213920 1001972 213972 1001978
rect 213920 1001914 213972 1001920
rect 213184 995988 213236 995994
rect 213184 995930 213236 995936
rect 211804 995444 211856 995450
rect 211804 995386 211856 995392
rect 209872 994900 209924 994906
rect 209872 994842 209924 994848
rect 202144 994764 202196 994770
rect 202144 994706 202196 994712
rect 200762 994528 200818 994537
rect 200762 994463 200818 994472
rect 213932 994294 213960 1001914
rect 207756 994288 207808 994294
rect 207756 994230 207808 994236
rect 213920 994288 213972 994294
rect 213920 994230 213972 994236
rect 200028 991500 200080 991506
rect 200028 991442 200080 991448
rect 207768 986678 207796 994230
rect 203156 986672 203208 986678
rect 203156 986614 203208 986620
rect 207756 986672 207808 986678
rect 207756 986614 207808 986620
rect 170324 983606 170798 983634
rect 186516 983606 186990 983634
rect 203168 983620 203196 986614
rect 215956 985998 215984 1002322
rect 217336 986678 217364 1004634
rect 228376 995858 228404 1006334
rect 247868 1006188 247920 1006194
rect 247868 1006130 247920 1006136
rect 229744 1006052 229796 1006058
rect 229744 1005994 229796 1006000
rect 247684 1006052 247736 1006058
rect 247684 1005994 247736 1006000
rect 229756 996130 229784 1005994
rect 246856 997892 246908 997898
rect 246856 997834 246908 997840
rect 246672 997756 246724 997762
rect 246672 997698 246724 997704
rect 246684 996441 246712 997698
rect 246670 996432 246726 996441
rect 246670 996367 246726 996376
rect 229744 996124 229796 996130
rect 229744 996066 229796 996072
rect 228364 995852 228416 995858
rect 228364 995794 228416 995800
rect 240874 995752 240930 995761
rect 240580 995710 240874 995738
rect 245566 995752 245622 995761
rect 245456 995710 245566 995738
rect 240874 995687 240930 995696
rect 245566 995687 245622 995696
rect 243910 995480 243966 995489
rect 231288 995438 231624 995466
rect 231932 995438 232268 995466
rect 232576 995438 232912 995466
rect 234416 995438 234568 995466
rect 234968 995438 235304 995466
rect 235612 995438 235948 995466
rect 236256 995438 236592 995466
rect 231596 994634 231624 995438
rect 232240 994906 232268 995438
rect 232884 995042 232912 995438
rect 232872 995036 232924 995042
rect 232872 994978 232924 994984
rect 232228 994900 232280 994906
rect 232228 994842 232280 994848
rect 231584 994628 231636 994634
rect 231584 994570 231636 994576
rect 234540 994498 234568 995438
rect 234528 994492 234580 994498
rect 234528 994434 234580 994440
rect 235276 994362 235304 995438
rect 235920 994770 235948 995438
rect 235908 994764 235960 994770
rect 235908 994706 235960 994712
rect 235264 994356 235316 994362
rect 235264 994298 235316 994304
rect 236564 994265 236592 995438
rect 238680 995438 238740 995466
rect 239292 995438 239628 995466
rect 239936 995438 240088 995466
rect 241776 995438 242112 995466
rect 238680 994537 238708 995438
rect 239600 994945 239628 995438
rect 239586 994936 239642 994945
rect 239586 994871 239642 994880
rect 238666 994528 238722 994537
rect 238666 994463 238722 994472
rect 236550 994256 236606 994265
rect 236550 994191 236606 994200
rect 240060 994106 240088 995438
rect 242084 995314 242112 995438
rect 242072 995308 242124 995314
rect 242072 995250 242124 995256
rect 242958 995217 242986 995452
rect 243616 995438 243910 995466
rect 243910 995415 243966 995424
rect 244246 995217 244274 995452
rect 246868 995314 246896 997834
rect 246856 995308 246908 995314
rect 246856 995250 246908 995256
rect 242944 995208 243000 995217
rect 242716 995172 242768 995178
rect 242944 995143 243000 995152
rect 244232 995208 244288 995217
rect 244232 995143 244288 995152
rect 242716 995114 242768 995120
rect 242728 994770 242756 995114
rect 247696 994945 247724 1005994
rect 247880 996713 247908 1006130
rect 249076 997898 249104 1006402
rect 254122 1006360 254178 1006369
rect 250260 1006324 250312 1006330
rect 254122 1006295 254124 1006304
rect 250260 1006266 250312 1006272
rect 254176 1006295 254178 1006304
rect 254124 1006266 254176 1006272
rect 250272 1006058 250300 1006266
rect 253662 1006224 253718 1006233
rect 253662 1006159 253664 1006168
rect 253716 1006159 253718 1006168
rect 262678 1006224 262734 1006233
rect 262678 1006159 262680 1006168
rect 253664 1006130 253716 1006136
rect 262732 1006159 262734 1006168
rect 278044 1006188 278096 1006194
rect 262680 1006130 262732 1006136
rect 278044 1006130 278096 1006136
rect 252466 1006088 252522 1006097
rect 250260 1006052 250312 1006058
rect 250260 1005994 250312 1006000
rect 250444 1006052 250496 1006058
rect 252466 1006023 252468 1006032
rect 250444 1005994 250496 1006000
rect 252520 1006023 252522 1006032
rect 261850 1006088 261906 1006097
rect 261850 1006023 261852 1006032
rect 252468 1005994 252520 1006000
rect 261904 1006023 261906 1006032
rect 261852 1005994 261904 1006000
rect 249708 1001972 249760 1001978
rect 249708 1001914 249760 1001920
rect 249340 999184 249392 999190
rect 249340 999126 249392 999132
rect 249064 997892 249116 997898
rect 249064 997834 249116 997840
rect 247866 996704 247922 996713
rect 247866 996639 247922 996648
rect 249352 995217 249380 999126
rect 249338 995208 249394 995217
rect 249338 995143 249394 995152
rect 247682 994936 247738 994945
rect 242900 994900 242952 994906
rect 242900 994842 242952 994848
rect 244556 994900 244608 994906
rect 247682 994871 247738 994880
rect 244556 994842 244608 994848
rect 242912 994786 242940 994842
rect 242912 994770 243124 994786
rect 242716 994764 242768 994770
rect 242912 994764 243136 994770
rect 242912 994758 243084 994764
rect 242716 994706 242768 994712
rect 243084 994706 243136 994712
rect 243728 994628 243780 994634
rect 243728 994570 243780 994576
rect 243360 994492 243412 994498
rect 243360 994434 243412 994440
rect 243372 994226 243400 994434
rect 243740 994362 243768 994570
rect 243728 994356 243780 994362
rect 243728 994298 243780 994304
rect 244568 994226 244596 994842
rect 243360 994220 243412 994226
rect 243360 994162 243412 994168
rect 244556 994220 244608 994226
rect 244556 994162 244608 994168
rect 240060 994078 240180 994106
rect 240152 993993 240180 994078
rect 240138 993984 240194 993993
rect 240138 993919 240194 993928
rect 249720 990146 249748 1001914
rect 250456 999190 250484 1005994
rect 263048 1005304 263100 1005310
rect 263046 1005272 263048 1005281
rect 263100 1005272 263102 1005281
rect 263046 1005207 263102 1005216
rect 255318 1002552 255374 1002561
rect 251824 1002516 251876 1002522
rect 255318 1002487 255320 1002496
rect 251824 1002458 251876 1002464
rect 255372 1002487 255374 1002496
rect 261022 1002552 261078 1002561
rect 261022 1002487 261024 1002496
rect 255320 1002458 255372 1002464
rect 261076 1002487 261078 1002496
rect 264244 1002516 264296 1002522
rect 261024 1002458 261076 1002464
rect 264244 1002458 264296 1002464
rect 250996 1002108 251048 1002114
rect 250996 1002050 251048 1002056
rect 250444 999184 250496 999190
rect 250444 999126 250496 999132
rect 249708 990140 249760 990146
rect 249708 990082 249760 990088
rect 251008 988786 251036 1002050
rect 251836 993993 251864 1002458
rect 256146 1002416 256202 1002425
rect 253112 1002380 253164 1002386
rect 256146 1002351 256148 1002360
rect 253112 1002322 253164 1002328
rect 256200 1002351 256202 1002360
rect 256148 1002322 256200 1002328
rect 252008 1002244 252060 1002250
rect 252008 1002186 252060 1002192
rect 252020 994265 252048 1002186
rect 252466 1002008 252522 1002017
rect 252466 1001943 252468 1001952
rect 252520 1001943 252522 1001952
rect 252468 1001914 252520 1001920
rect 253124 994634 253152 1002322
rect 254490 1002280 254546 1002289
rect 254490 1002215 254492 1002224
rect 254544 1002215 254546 1002224
rect 254492 1002186 254544 1002192
rect 253294 1002144 253350 1002153
rect 256146 1002144 256202 1002153
rect 253294 1002079 253296 1002088
rect 253348 1002079 253350 1002088
rect 253480 1002108 253532 1002114
rect 253296 1002050 253348 1002056
rect 256146 1002079 256148 1002088
rect 253480 1002050 253532 1002056
rect 256200 1002079 256202 1002088
rect 263506 1002144 263562 1002153
rect 263506 1002079 263508 1002088
rect 256148 1002050 256200 1002056
rect 263560 1002079 263562 1002088
rect 263508 1002050 263560 1002056
rect 253492 995178 253520 1002050
rect 261022 1002008 261078 1002017
rect 263874 1002008 263930 1002017
rect 261022 1001943 261024 1001952
rect 261076 1001943 261078 1001952
rect 263600 1001972 263652 1001978
rect 261024 1001914 261076 1001920
rect 263874 1001943 263876 1001952
rect 263600 1001914 263652 1001920
rect 263928 1001943 263930 1001952
rect 263876 1001914 263928 1001920
rect 258170 998200 258226 998209
rect 258170 998135 258172 998144
rect 258224 998135 258226 998144
rect 259460 998164 259512 998170
rect 258172 998106 258224 998112
rect 259460 998106 259512 998112
rect 257342 998064 257398 998073
rect 254584 998028 254636 998034
rect 257342 997999 257344 998008
rect 254584 997970 254636 997976
rect 257396 997999 257398 998008
rect 257344 997970 257396 997976
rect 253480 995172 253532 995178
rect 253480 995114 253532 995120
rect 253112 994628 253164 994634
rect 253112 994570 253164 994576
rect 254596 994537 254624 997970
rect 256974 997928 257030 997937
rect 254768 997892 254820 997898
rect 258170 997928 258226 997937
rect 256974 997863 256976 997872
rect 254768 997834 254820 997840
rect 257028 997863 257030 997872
rect 257356 997886 258170 997914
rect 256976 997834 257028 997840
rect 254780 997762 254808 997834
rect 256514 997792 256570 997801
rect 254768 997756 254820 997762
rect 254768 997698 254820 997704
rect 255976 997736 256514 997754
rect 255976 997727 256570 997736
rect 255976 997726 256556 997727
rect 255976 994770 256004 997726
rect 255964 994764 256016 994770
rect 255964 994706 256016 994712
rect 254582 994528 254638 994537
rect 257356 994498 257384 997886
rect 258170 997863 258226 997872
rect 258998 997792 259054 997801
rect 258092 997736 258998 997754
rect 258092 997727 259054 997736
rect 258092 997726 259040 997727
rect 258092 995042 258120 997726
rect 258080 995036 258132 995042
rect 258080 994978 258132 994984
rect 259472 994906 259500 998106
rect 260196 998096 260248 998102
rect 260194 998064 260196 998073
rect 262864 998096 262916 998102
rect 260248 998064 260250 998073
rect 262864 998038 262916 998044
rect 260194 997999 260250 998008
rect 259828 997960 259880 997966
rect 259826 997928 259828 997937
rect 262220 997960 262272 997966
rect 259880 997928 259882 997937
rect 262220 997902 262272 997908
rect 259826 997863 259882 997872
rect 260196 997824 260248 997830
rect 260194 997792 260196 997801
rect 260932 997824 260984 997830
rect 260248 997792 260250 997801
rect 260932 997766 260984 997772
rect 261850 997792 261906 997801
rect 260194 997727 260250 997736
rect 260944 995450 260972 997766
rect 261128 997736 261850 997754
rect 261128 997727 261906 997736
rect 261128 997726 261892 997727
rect 261128 995994 261156 997726
rect 262232 996130 262260 997902
rect 262876 996130 262904 998038
rect 262220 996124 262272 996130
rect 262220 996066 262272 996072
rect 262864 996124 262916 996130
rect 262864 996066 262916 996072
rect 261116 995988 261168 995994
rect 261116 995930 261168 995936
rect 263612 995858 263640 1001914
rect 264256 995994 264284 1002458
rect 265624 1002108 265676 1002114
rect 265624 1002050 265676 1002056
rect 264244 995988 264296 995994
rect 264244 995930 264296 995936
rect 263600 995852 263652 995858
rect 263600 995794 263652 995800
rect 260932 995444 260984 995450
rect 260932 995386 260984 995392
rect 259460 994900 259512 994906
rect 259460 994842 259512 994848
rect 254582 994463 254638 994472
rect 257344 994492 257396 994498
rect 257344 994434 257396 994440
rect 252006 994256 252062 994265
rect 252006 994191 252062 994200
rect 265636 994158 265664 1002050
rect 267004 1001972 267056 1001978
rect 267004 1001914 267056 1001920
rect 265624 994152 265676 994158
rect 265624 994094 265676 994100
rect 251822 993984 251878 993993
rect 251822 993919 251878 993928
rect 251454 993168 251510 993177
rect 251454 993103 251510 993112
rect 250996 988780 251048 988786
rect 250996 988722 251048 988728
rect 217324 986672 217376 986678
rect 217324 986614 217376 986620
rect 219440 986672 219492 986678
rect 219440 986614 219492 986620
rect 215944 985992 215996 985998
rect 215944 985934 215996 985940
rect 219452 983620 219480 986614
rect 235632 985992 235684 985998
rect 235632 985934 235684 985940
rect 235644 983620 235672 985934
rect 251468 983634 251496 993103
rect 267016 991778 267044 1001914
rect 278056 995858 278084 1006130
rect 280804 1006052 280856 1006058
rect 280804 1005994 280856 1006000
rect 279424 1005304 279476 1005310
rect 279424 1005246 279476 1005252
rect 278044 995852 278096 995858
rect 278044 995794 278096 995800
rect 267740 994152 267792 994158
rect 267740 994094 267792 994100
rect 267004 991772 267056 991778
rect 267004 991714 267056 991720
rect 267752 983634 267780 994094
rect 279436 985998 279464 1005246
rect 280816 995246 280844 1005994
rect 298468 1000476 298520 1000482
rect 298468 1000418 298520 1000424
rect 298100 997824 298152 997830
rect 298100 997766 298152 997772
rect 298282 997792 298338 997801
rect 281908 995988 281960 995994
rect 281908 995930 281960 995936
rect 281920 995450 281948 995930
rect 291750 995752 291806 995761
rect 291502 995710 291750 995738
rect 293498 995752 293554 995761
rect 293342 995710 293498 995738
rect 291750 995687 291806 995696
rect 297270 995752 297326 995761
rect 297022 995710 297270 995738
rect 293498 995687 293554 995696
rect 298112 995738 298140 997766
rect 298282 997727 298338 997736
rect 298296 995761 298324 997727
rect 297270 995687 297326 995696
rect 297928 995710 298140 995738
rect 298282 995752 298338 995761
rect 286690 995480 286746 995489
rect 281908 995444 281960 995450
rect 281908 995386 281960 995392
rect 280804 995240 280856 995246
rect 280804 995182 280856 995188
rect 282840 994974 282868 995452
rect 282828 994968 282880 994974
rect 282828 994910 282880 994916
rect 283484 994566 283512 995452
rect 284128 994838 284156 995452
rect 284116 994832 284168 994838
rect 284116 994774 284168 994780
rect 285968 994702 285996 995452
rect 286534 995438 286690 995466
rect 292486 995480 292542 995489
rect 287178 995438 287560 995466
rect 286690 995415 286746 995424
rect 285956 994696 286008 994702
rect 285956 994638 286008 994644
rect 283472 994560 283524 994566
rect 283472 994502 283524 994508
rect 287532 994265 287560 995438
rect 287808 994537 287836 995452
rect 287794 994528 287850 994537
rect 287794 994463 287850 994472
rect 287518 994256 287574 994265
rect 287518 994191 287574 994200
rect 290292 993993 290320 995452
rect 290844 994809 290872 995452
rect 292146 995438 292486 995466
rect 296166 995480 296222 995489
rect 294538 995438 294920 995466
rect 292486 995415 292542 995424
rect 294696 995376 294748 995382
rect 294696 995318 294748 995324
rect 294708 995110 294736 995318
rect 294696 995104 294748 995110
rect 294696 995046 294748 995052
rect 290830 994800 290886 994809
rect 290830 994735 290886 994744
rect 294892 994294 294920 995438
rect 295168 995330 295196 995452
rect 295826 995438 296166 995466
rect 296166 995415 296222 995424
rect 295168 995314 295288 995330
rect 295168 995308 295300 995314
rect 295168 995302 295248 995308
rect 295248 995250 295300 995256
rect 296628 995172 296680 995178
rect 296628 995114 296680 995120
rect 296444 995104 296496 995110
rect 296442 995072 296444 995081
rect 296496 995072 296498 995081
rect 296442 995007 296498 995016
rect 296640 994566 296668 995114
rect 297928 994809 297956 995710
rect 298282 995687 298338 995696
rect 298100 995580 298152 995586
rect 298100 995522 298152 995528
rect 298112 994838 298140 995522
rect 298480 995314 298508 1000418
rect 298756 997754 298784 1006538
rect 298928 1006324 298980 1006330
rect 298928 1006266 298980 1006272
rect 298940 997754 298968 1006266
rect 298756 997726 298876 997754
rect 298940 997726 299060 997754
rect 298652 995988 298704 995994
rect 298652 995930 298704 995936
rect 298664 995450 298692 995930
rect 298652 995444 298704 995450
rect 298652 995386 298704 995392
rect 298468 995308 298520 995314
rect 298468 995250 298520 995256
rect 298848 995081 298876 997726
rect 299032 996849 299060 997726
rect 299018 996840 299074 996849
rect 299018 996775 299074 996784
rect 300136 995761 300164 1006674
rect 306104 1006596 306156 1006602
rect 306104 1006538 306156 1006544
rect 304078 1006496 304134 1006505
rect 304078 1006431 304080 1006440
rect 304132 1006431 304134 1006440
rect 304080 1006402 304132 1006408
rect 305274 1006360 305330 1006369
rect 305274 1006295 305276 1006304
rect 305328 1006295 305330 1006304
rect 305276 1006266 305328 1006272
rect 306116 1006194 306144 1006538
rect 314658 1006496 314714 1006505
rect 361394 1006496 361450 1006505
rect 314658 1006431 314660 1006440
rect 314712 1006431 314714 1006440
rect 319444 1006460 319496 1006466
rect 314660 1006402 314712 1006408
rect 361394 1006431 361396 1006440
rect 319444 1006402 319496 1006408
rect 361448 1006431 361450 1006440
rect 371884 1006460 371936 1006466
rect 361396 1006402 361448 1006408
rect 371884 1006402 371936 1006408
rect 306930 1006360 306986 1006369
rect 306930 1006295 306932 1006304
rect 306984 1006295 306986 1006304
rect 306932 1006266 306984 1006272
rect 311806 1006224 311862 1006233
rect 300308 1006188 300360 1006194
rect 300308 1006130 300360 1006136
rect 306104 1006188 306156 1006194
rect 311806 1006159 311808 1006168
rect 306104 1006130 306156 1006136
rect 311860 1006159 311862 1006168
rect 314658 1006224 314714 1006233
rect 314658 1006159 314660 1006168
rect 311808 1006130 311860 1006136
rect 314712 1006159 314714 1006168
rect 314660 1006130 314712 1006136
rect 300320 996033 300348 1006130
rect 301502 1006088 301558 1006097
rect 301502 1006023 301558 1006032
rect 303250 1006088 303306 1006097
rect 303250 1006023 303252 1006032
rect 301044 999184 301096 999190
rect 301044 999126 301096 999132
rect 300860 999048 300912 999054
rect 300860 998990 300912 998996
rect 300872 996441 300900 998990
rect 300858 996432 300914 996441
rect 300858 996367 300914 996376
rect 300306 996024 300362 996033
rect 300306 995959 300362 995968
rect 300122 995752 300178 995761
rect 300122 995687 300178 995696
rect 298834 995072 298890 995081
rect 298834 995007 298890 995016
rect 298100 994832 298152 994838
rect 297914 994800 297970 994809
rect 298100 994774 298152 994780
rect 297914 994735 297970 994744
rect 296628 994560 296680 994566
rect 301056 994537 301084 999126
rect 301516 995489 301544 1006023
rect 303304 1006023 303306 1006032
rect 304078 1006088 304134 1006097
rect 304078 1006023 304080 1006032
rect 303252 1005994 303304 1006000
rect 304132 1006023 304134 1006032
rect 305274 1006088 305330 1006097
rect 305274 1006023 305276 1006032
rect 304080 1005994 304132 1006000
rect 305328 1006023 305330 1006032
rect 305276 1005994 305328 1006000
rect 307298 1005272 307354 1005281
rect 304264 1005236 304316 1005242
rect 307298 1005207 307300 1005216
rect 304264 1005178 304316 1005184
rect 307352 1005207 307354 1005216
rect 307300 1005178 307352 1005184
rect 303068 1002244 303120 1002250
rect 303068 1002186 303120 1002192
rect 302884 1001972 302936 1001978
rect 302884 1001914 302936 1001920
rect 302896 997830 302924 1001914
rect 303080 999190 303108 1002186
rect 303068 999184 303120 999190
rect 303068 999126 303120 999132
rect 302884 997824 302936 997830
rect 303252 997824 303304 997830
rect 302884 997766 302936 997772
rect 303250 997792 303252 997801
rect 303304 997792 303306 997801
rect 303250 997727 303306 997736
rect 301502 995480 301558 995489
rect 301502 995415 301558 995424
rect 296628 994502 296680 994508
rect 301042 994528 301098 994537
rect 301042 994463 301098 994472
rect 294880 994288 294932 994294
rect 304276 994265 304304 1005178
rect 308954 1005000 309010 1005009
rect 305828 1004964 305880 1004970
rect 308954 1004935 308956 1004944
rect 305828 1004906 305880 1004912
rect 309008 1004935 309010 1004944
rect 308956 1004906 309008 1004912
rect 304448 1004828 304500 1004834
rect 304448 1004770 304500 1004776
rect 304460 999054 304488 1004770
rect 305644 1004692 305696 1004698
rect 305644 1004634 305696 1004640
rect 304448 999048 304500 999054
rect 304448 998990 304500 998996
rect 305656 995246 305684 1004634
rect 305840 997830 305868 1004906
rect 306930 1004864 306986 1004873
rect 306930 1004799 306932 1004808
rect 306984 1004799 306986 1004808
rect 313830 1004864 313886 1004873
rect 313830 1004799 313832 1004808
rect 306932 1004770 306984 1004776
rect 313884 1004799 313886 1004808
rect 316040 1004828 316092 1004834
rect 313832 1004770 313884 1004776
rect 316040 1004770 316092 1004776
rect 308126 1004728 308182 1004737
rect 308126 1004663 308128 1004672
rect 308180 1004663 308182 1004672
rect 315486 1004728 315542 1004737
rect 315486 1004663 315488 1004672
rect 308128 1004634 308180 1004640
rect 315540 1004663 315542 1004672
rect 315488 1004634 315540 1004640
rect 310150 1002416 310206 1002425
rect 310150 1002351 310152 1002360
rect 310204 1002351 310206 1002360
rect 311900 1002380 311952 1002386
rect 310152 1002322 310204 1002328
rect 311900 1002322 311952 1002328
rect 306102 1002280 306158 1002289
rect 306102 1002215 306104 1002224
rect 306156 1002215 306158 1002224
rect 306104 1002186 306156 1002192
rect 308954 1002144 309010 1002153
rect 307024 1002108 307076 1002114
rect 310150 1002144 310206 1002153
rect 308954 1002079 308956 1002088
rect 307024 1002050 307076 1002056
rect 309008 1002079 309010 1002088
rect 309152 1002102 310150 1002130
rect 308956 1002050 309008 1002056
rect 306102 1002008 306158 1002017
rect 306102 1001943 306104 1001952
rect 306156 1001943 306158 1001952
rect 306104 1001914 306156 1001920
rect 305828 997824 305880 997830
rect 305828 997766 305880 997772
rect 305644 995240 305696 995246
rect 305644 995182 305696 995188
rect 294880 994230 294932 994236
rect 304262 994256 304318 994265
rect 304262 994191 304318 994200
rect 307036 993993 307064 1002050
rect 308404 1001972 308456 1001978
rect 308404 1001914 308456 1001920
rect 308416 994702 308444 1001914
rect 309152 1000482 309180 1002102
rect 310150 1002079 310206 1002088
rect 310610 1002144 310666 1002153
rect 310610 1002079 310666 1002088
rect 310978 1002144 311034 1002153
rect 310978 1002079 310980 1002088
rect 309782 1002008 309838 1002017
rect 309782 1001943 309784 1001952
rect 309836 1001943 309838 1001952
rect 309784 1001914 309836 1001920
rect 309140 1000476 309192 1000482
rect 309140 1000418 309192 1000424
rect 310624 995586 310652 1002079
rect 311032 1002079 311034 1002088
rect 310980 1002050 311032 1002056
rect 310612 995580 310664 995586
rect 310612 995522 310664 995528
rect 311912 994974 311940 1002322
rect 313280 1002108 313332 1002114
rect 313280 1002050 313332 1002056
rect 312634 1002008 312690 1002017
rect 312634 1001943 312636 1001952
rect 312688 1001943 312690 1001952
rect 312636 1001914 312688 1001920
rect 313292 996130 313320 1002050
rect 314660 1001972 314712 1001978
rect 314660 1001914 314712 1001920
rect 313280 996124 313332 996130
rect 313280 996066 313332 996072
rect 314672 995994 314700 1001914
rect 314660 995988 314712 995994
rect 314660 995930 314712 995936
rect 316052 995858 316080 1004770
rect 318064 1004692 318116 1004698
rect 318064 1004634 318116 1004640
rect 318076 997082 318104 1004634
rect 319456 997218 319484 1006402
rect 331864 1006324 331916 1006330
rect 331864 1006266 331916 1006272
rect 324964 1006188 325016 1006194
rect 324964 1006130 325016 1006136
rect 319444 997212 319496 997218
rect 319444 997154 319496 997160
rect 318064 997076 318116 997082
rect 318064 997018 318116 997024
rect 316040 995852 316092 995858
rect 316040 995794 316092 995800
rect 324976 995586 325004 1006130
rect 324964 995580 325016 995586
rect 324964 995522 325016 995528
rect 311900 994968 311952 994974
rect 311900 994910 311952 994916
rect 308404 994696 308456 994702
rect 308404 994638 308456 994644
rect 290278 993984 290334 993993
rect 290278 993919 290334 993928
rect 307022 993984 307078 993993
rect 307022 993919 307078 993928
rect 316406 992896 316462 992905
rect 316406 992831 316462 992840
rect 284300 991772 284352 991778
rect 284300 991714 284352 991720
rect 279424 985992 279476 985998
rect 279424 985934 279476 985940
rect 251468 983606 251850 983634
rect 267752 983606 268134 983634
rect 284312 983620 284340 991714
rect 300492 985992 300544 985998
rect 300492 985934 300544 985940
rect 300504 983620 300532 985934
rect 316420 983634 316448 992831
rect 331876 984910 331904 1006266
rect 365074 1006224 365130 1006233
rect 365074 1006159 365076 1006168
rect 365128 1006159 365130 1006168
rect 367744 1006188 367796 1006194
rect 365076 1006130 365128 1006136
rect 367744 1006130 367796 1006136
rect 354862 1006088 354918 1006097
rect 332048 1006052 332100 1006058
rect 357346 1006088 357402 1006097
rect 354862 1006023 354864 1006032
rect 332048 1005994 332100 1006000
rect 354916 1006023 354918 1006032
rect 356704 1006052 356756 1006058
rect 354864 1005994 354916 1006000
rect 357346 1006023 357348 1006032
rect 356704 1005994 356756 1006000
rect 357400 1006023 357402 1006032
rect 357348 1005994 357400 1006000
rect 331864 984904 331916 984910
rect 331864 984846 331916 984852
rect 332060 984774 332088 1005994
rect 356520 1005440 356572 1005446
rect 356518 1005408 356520 1005417
rect 356572 1005408 356574 1005417
rect 356518 1005343 356574 1005352
rect 355690 1005000 355746 1005009
rect 353208 1004964 353260 1004970
rect 355690 1004935 355692 1004944
rect 353208 1004906 353260 1004912
rect 355744 1004935 355746 1004944
rect 355692 1004906 355744 1004912
rect 351828 1001972 351880 1001978
rect 351828 1001914 351880 1001920
rect 332600 997212 332652 997218
rect 332600 997154 332652 997160
rect 332048 984768 332100 984774
rect 332048 984710 332100 984716
rect 332612 983634 332640 997154
rect 349160 997076 349212 997082
rect 349160 997018 349212 997024
rect 316420 983606 316802 983634
rect 332612 983606 332994 983634
rect 349172 983620 349200 997018
rect 351840 993206 351868 1001914
rect 353220 998714 353248 1004906
rect 355690 1004728 355746 1004737
rect 354588 1004692 354640 1004698
rect 355690 1004663 355692 1004672
rect 354588 1004634 354640 1004640
rect 355744 1004663 355746 1004672
rect 355692 1004634 355744 1004640
rect 354034 1002008 354090 1002017
rect 354034 1001943 354036 1001952
rect 354088 1001943 354090 1001952
rect 354036 1001914 354088 1001920
rect 353208 998708 353260 998714
rect 353208 998650 353260 998656
rect 351828 993200 351880 993206
rect 351828 993142 351880 993148
rect 354600 987562 354628 1004634
rect 355968 1001972 356020 1001978
rect 355968 1001914 356020 1001920
rect 355980 998578 356008 1001914
rect 355968 998572 356020 998578
rect 355968 998514 356020 998520
rect 356716 994770 356744 1005994
rect 360568 1005712 360620 1005718
rect 360566 1005680 360568 1005689
rect 360620 1005680 360622 1005689
rect 360566 1005615 360622 1005624
rect 359740 1005576 359792 1005582
rect 359738 1005544 359740 1005553
rect 359792 1005544 359794 1005553
rect 359738 1005479 359794 1005488
rect 356888 1005304 356940 1005310
rect 356886 1005272 356888 1005281
rect 356940 1005272 356942 1005281
rect 356886 1005207 356942 1005216
rect 363418 1005136 363474 1005145
rect 365074 1005136 365130 1005145
rect 363418 1005071 363420 1005080
rect 363472 1005071 363474 1005080
rect 364524 1005100 364576 1005106
rect 363420 1005042 363472 1005048
rect 365074 1005071 365076 1005080
rect 364524 1005042 364576 1005048
rect 365128 1005071 365130 1005080
rect 365076 1005042 365128 1005048
rect 361394 1005000 361450 1005009
rect 361394 1004935 361396 1004944
rect 361448 1004935 361450 1004944
rect 361396 1004906 361448 1004912
rect 364246 1004864 364302 1004873
rect 364246 1004799 364248 1004808
rect 364300 1004799 364302 1004808
rect 364248 1004770 364300 1004776
rect 362590 1004728 362646 1004737
rect 362590 1004663 362592 1004672
rect 362644 1004663 362646 1004672
rect 362592 1004634 362644 1004640
rect 364536 1004562 364564 1005042
rect 365168 1004964 365220 1004970
rect 365168 1004906 365220 1004912
rect 364984 1004692 365036 1004698
rect 364984 1004634 365036 1004640
rect 364524 1004556 364576 1004562
rect 364524 1004498 364576 1004504
rect 358542 1002416 358598 1002425
rect 358542 1002351 358544 1002360
rect 358596 1002351 358598 1002360
rect 360844 1002380 360896 1002386
rect 358544 1002322 358596 1002328
rect 360844 1002322 360896 1002328
rect 359370 1002280 359426 1002289
rect 359370 1002215 359372 1002224
rect 359424 1002215 359426 1002224
rect 359372 1002186 359424 1002192
rect 358542 1002144 358598 1002153
rect 360566 1002144 360622 1002153
rect 358598 1002102 359504 1002130
rect 358542 1002079 358598 1002088
rect 358728 1002040 358780 1002046
rect 357346 1002008 357402 1002017
rect 358728 1001982 358780 1001988
rect 357346 1001943 357348 1001952
rect 357400 1001943 357402 1001952
rect 357348 1001914 357400 1001920
rect 358740 995042 358768 1001982
rect 359476 997626 359504 1002102
rect 360566 1002079 360568 1002088
rect 360620 1002079 360622 1002088
rect 360568 1002050 360620 1002056
rect 360198 1002008 360254 1002017
rect 360198 1001943 360200 1001952
rect 360252 1001943 360254 1001952
rect 360200 1001914 360252 1001920
rect 360856 998442 360884 1002322
rect 363604 1002108 363656 1002114
rect 363604 1002050 363656 1002056
rect 362224 1001972 362276 1001978
rect 362224 1001914 362276 1001920
rect 360844 998436 360896 998442
rect 360844 998378 360896 998384
rect 362236 997762 362264 1001914
rect 362224 997756 362276 997762
rect 362224 997698 362276 997704
rect 359464 997620 359516 997626
rect 359464 997562 359516 997568
rect 363616 997082 363644 1002050
rect 363604 997076 363656 997082
rect 363604 997018 363656 997024
rect 364996 996130 365024 1004634
rect 364984 996124 365036 996130
rect 364984 996066 365036 996072
rect 365180 995994 365208 1004906
rect 366364 1004828 366416 1004834
rect 366364 1004770 366416 1004776
rect 365902 1002008 365958 1002017
rect 365902 1001943 365904 1001952
rect 365956 1001943 365958 1001952
rect 365904 1001914 365956 1001920
rect 365168 995988 365220 995994
rect 365168 995930 365220 995936
rect 366376 995858 366404 1004770
rect 366548 1004556 366600 1004562
rect 366548 1004498 366600 1004504
rect 366560 996266 366588 1004498
rect 366548 996260 366600 996266
rect 366548 996202 366600 996208
rect 366364 995852 366416 995858
rect 366364 995794 366416 995800
rect 364984 995580 365036 995586
rect 364984 995522 365036 995528
rect 358728 995036 358780 995042
rect 358728 994978 358780 994984
rect 356704 994764 356756 994770
rect 356704 994706 356756 994712
rect 354588 987556 354640 987562
rect 354588 987498 354640 987504
rect 364996 983634 365024 995522
rect 367756 991778 367784 1006130
rect 370504 1005100 370556 1005106
rect 370504 1005042 370556 1005048
rect 369124 1001972 369176 1001978
rect 369124 1001914 369176 1001920
rect 367744 991772 367796 991778
rect 367744 991714 367796 991720
rect 369136 985998 369164 1001914
rect 370516 986134 370544 1005042
rect 371896 998850 371924 1006402
rect 373264 1005576 373316 1005582
rect 373264 1005518 373316 1005524
rect 371884 998844 371936 998850
rect 371884 998786 371936 998792
rect 372896 998708 372948 998714
rect 372896 998650 372948 998656
rect 372528 997756 372580 997762
rect 372528 997698 372580 997704
rect 372344 997620 372396 997626
rect 372344 997562 372396 997568
rect 372356 996713 372384 997562
rect 372342 996704 372398 996713
rect 372342 996639 372398 996648
rect 372540 996441 372568 997698
rect 372712 997076 372764 997082
rect 372712 997018 372764 997024
rect 372526 996432 372582 996441
rect 372526 996367 372582 996376
rect 372724 994906 372752 997018
rect 372712 994900 372764 994906
rect 372712 994842 372764 994848
rect 372908 994634 372936 998650
rect 373276 995081 373304 1005518
rect 374012 999190 374040 1006674
rect 376024 1006052 376076 1006058
rect 376024 1005994 376076 1006000
rect 374000 999184 374052 999190
rect 374000 999126 374052 999132
rect 376036 998102 376064 1005994
rect 377404 1005712 377456 1005718
rect 377404 1005654 377456 1005660
rect 376300 998572 376352 998578
rect 376300 998514 376352 998520
rect 376024 998096 376076 998102
rect 376024 998038 376076 998044
rect 375472 996260 375524 996266
rect 375472 996202 375524 996208
rect 375484 995586 375512 996202
rect 375472 995580 375524 995586
rect 375472 995522 375524 995528
rect 373262 995072 373318 995081
rect 373262 995007 373318 995016
rect 376312 994809 376340 998514
rect 377416 995178 377444 1005654
rect 378784 1005440 378836 1005446
rect 378784 1005382 378836 1005388
rect 378796 998170 378824 1005382
rect 381544 1005304 381596 1005310
rect 381544 1005246 381596 1005252
rect 378784 998164 378836 998170
rect 378784 998106 378836 998112
rect 381268 998164 381320 998170
rect 381268 998106 381320 998112
rect 378416 998096 378468 998102
rect 378416 998038 378468 998044
rect 377404 995172 377456 995178
rect 377404 995114 377456 995120
rect 376298 994800 376354 994809
rect 376298 994735 376354 994744
rect 372896 994628 372948 994634
rect 372896 994570 372948 994576
rect 378428 994265 378456 998038
rect 378600 994764 378652 994770
rect 378600 994706 378652 994712
rect 378612 994498 378640 994706
rect 381280 994537 381308 998106
rect 381556 995353 381584 1005246
rect 381728 999184 381780 999190
rect 381728 999126 381780 999132
rect 381740 995450 381768 999126
rect 383108 998844 383160 998850
rect 383108 998786 383160 998792
rect 383120 995761 383148 998786
rect 383292 998436 383344 998442
rect 383292 998378 383344 998384
rect 383106 995752 383162 995761
rect 383106 995687 383162 995696
rect 383304 995586 383332 998378
rect 385682 995752 385738 995761
rect 387890 995752 387946 995761
rect 385738 995710 385986 995738
rect 387826 995710 387890 995738
rect 385682 995687 385738 995696
rect 387890 995687 387946 995696
rect 388166 995752 388222 995761
rect 396538 995752 396594 995761
rect 388222 995710 388378 995738
rect 396382 995710 396538 995738
rect 388166 995687 388222 995696
rect 396538 995687 396594 995696
rect 385052 995586 385342 995602
rect 383292 995580 383344 995586
rect 383292 995522 383344 995528
rect 385040 995580 385342 995586
rect 385092 995574 385342 995580
rect 385040 995522 385092 995528
rect 381728 995444 381780 995450
rect 381728 995386 381780 995392
rect 381542 995344 381598 995353
rect 381542 995279 381598 995288
rect 384684 995178 384712 995452
rect 388640 995450 389022 995466
rect 388628 995444 389022 995450
rect 388680 995438 389022 995444
rect 389376 995438 389666 995466
rect 388628 995386 388680 995392
rect 389376 995353 389404 995438
rect 389362 995344 389418 995353
rect 389362 995279 389418 995288
rect 384672 995172 384724 995178
rect 384672 995114 384724 995120
rect 392136 995081 392164 995452
rect 392320 995438 392702 995466
rect 392122 995072 392178 995081
rect 392122 995007 392178 995016
rect 392320 994537 392348 995438
rect 393332 995217 393360 995452
rect 393318 995208 393374 995217
rect 393318 995143 393374 995152
rect 393226 995072 393282 995081
rect 393226 995007 393282 995016
rect 381266 994528 381322 994537
rect 378600 994492 378652 994498
rect 381266 994463 381322 994472
rect 392306 994528 392362 994537
rect 392306 994463 392362 994472
rect 378600 994434 378652 994440
rect 381176 994288 381228 994294
rect 378414 994256 378470 994265
rect 393240 994265 393268 995007
rect 393976 994770 394004 995452
rect 395172 994809 395200 995452
rect 397012 994906 397040 995452
rect 397000 994900 397052 994906
rect 397000 994842 397052 994848
rect 395158 994800 395214 994809
rect 393964 994764 394016 994770
rect 395158 994735 395214 994744
rect 393964 994706 394016 994712
rect 397656 994634 397684 995452
rect 398852 995042 398880 995452
rect 400876 995382 400904 1006674
rect 427174 1006632 427230 1006641
rect 427174 1006567 427176 1006576
rect 427228 1006567 427230 1006576
rect 427176 1006538 427228 1006544
rect 423494 1006496 423550 1006505
rect 423494 1006431 423496 1006440
rect 423548 1006431 423550 1006440
rect 423496 1006402 423548 1006408
rect 424322 1006360 424378 1006369
rect 424322 1006295 424324 1006304
rect 424376 1006295 424378 1006304
rect 438860 1006324 438912 1006330
rect 424324 1006266 424376 1006272
rect 438860 1006266 438912 1006272
rect 422666 1006088 422722 1006097
rect 422666 1006023 422722 1006032
rect 423494 1006088 423550 1006097
rect 429198 1006088 429254 1006097
rect 423494 1006023 423496 1006032
rect 422680 1004850 422708 1006023
rect 423548 1006023 423550 1006032
rect 427820 1006052 427872 1006058
rect 423496 1005994 423548 1006000
rect 429198 1006023 429200 1006032
rect 427820 1005994 427872 1006000
rect 429252 1006023 429254 1006032
rect 429200 1005994 429252 1006000
rect 427544 1005712 427596 1005718
rect 427542 1005680 427544 1005689
rect 427596 1005680 427598 1005689
rect 427542 1005615 427598 1005624
rect 425518 1005408 425574 1005417
rect 425518 1005343 425520 1005352
rect 425572 1005343 425574 1005352
rect 425520 1005314 425572 1005320
rect 424690 1005136 424746 1005145
rect 424690 1005071 424692 1005080
rect 424744 1005071 424746 1005080
rect 424692 1005042 424744 1005048
rect 422680 1004822 422984 1004850
rect 422666 1004728 422722 1004737
rect 422220 1004686 422666 1004714
rect 421470 1002008 421526 1002017
rect 419448 1001972 419500 1001978
rect 421470 1001943 421472 1001952
rect 419448 1001914 419500 1001920
rect 421524 1001943 421526 1001952
rect 421472 1001914 421524 1001920
rect 400864 995376 400916 995382
rect 400864 995318 400916 995324
rect 398840 995036 398892 995042
rect 398840 994978 398892 994984
rect 397644 994628 397696 994634
rect 397644 994570 397696 994576
rect 381176 994230 381228 994236
rect 393226 994256 393282 994265
rect 378414 994191 378470 994200
rect 370504 986128 370556 986134
rect 370504 986070 370556 986076
rect 369124 985992 369176 985998
rect 369124 985934 369176 985940
rect 381188 983634 381216 994230
rect 393226 994191 393282 994200
rect 419460 991778 419488 1001914
rect 421012 996464 421064 996470
rect 421010 996432 421012 996441
rect 421064 996432 421066 996441
rect 421010 996367 421066 996376
rect 415032 991772 415084 991778
rect 415032 991714 415084 991720
rect 419448 991772 419500 991778
rect 419448 991714 419500 991720
rect 397828 986128 397880 986134
rect 397828 986070 397880 986076
rect 364996 983606 365470 983634
rect 381188 983606 381662 983634
rect 397840 983620 397868 986070
rect 415044 985998 415072 991714
rect 422220 988922 422248 1004686
rect 422666 1004663 422722 1004672
rect 422956 994974 422984 1004822
rect 425520 1003944 425572 1003950
rect 425518 1003912 425520 1003921
rect 425572 1003912 425574 1003921
rect 425518 1003847 425574 1003856
rect 424692 1002720 424744 1002726
rect 424690 1002688 424692 1002697
rect 424744 1002688 424746 1002697
rect 424690 1002623 424746 1002632
rect 427832 1002590 427860 1005994
rect 428372 1005848 428424 1005854
rect 428370 1005816 428372 1005825
rect 428424 1005816 428426 1005825
rect 428370 1005751 428426 1005760
rect 438872 1005718 438900 1006266
rect 438860 1005712 438912 1005718
rect 438860 1005654 438912 1005660
rect 430856 1005576 430908 1005582
rect 430854 1005544 430856 1005553
rect 433984 1005576 434036 1005582
rect 430908 1005544 430910 1005553
rect 430854 1005479 430910 1005488
rect 431512 1005502 432000 1005530
rect 433984 1005518 434036 1005524
rect 430026 1005272 430082 1005281
rect 430026 1005207 430028 1005216
rect 430080 1005207 430082 1005216
rect 430028 1005178 430080 1005184
rect 431512 1005106 431540 1005502
rect 431972 1005446 432000 1005502
rect 431960 1005440 432012 1005446
rect 431960 1005382 432012 1005388
rect 431776 1005372 431828 1005378
rect 431776 1005314 431828 1005320
rect 431788 1005258 431816 1005314
rect 432420 1005304 432472 1005310
rect 432050 1005272 432106 1005281
rect 431788 1005230 431954 1005258
rect 431682 1005136 431738 1005145
rect 431500 1005100 431552 1005106
rect 431926 1005122 431954 1005230
rect 432106 1005252 432420 1005258
rect 432106 1005246 432472 1005252
rect 432106 1005230 432460 1005246
rect 432050 1005207 432106 1005216
rect 432604 1005168 432656 1005174
rect 431926 1005094 432000 1005122
rect 432604 1005110 432656 1005116
rect 431682 1005071 431684 1005080
rect 431500 1005042 431552 1005048
rect 431736 1005071 431738 1005080
rect 431972 1005088 432000 1005094
rect 431972 1005060 432460 1005088
rect 431684 1005042 431736 1005048
rect 429198 1005000 429254 1005009
rect 431926 1004970 432092 1004986
rect 429198 1004935 429200 1004944
rect 429252 1004935 429254 1004944
rect 431914 1004964 432092 1004970
rect 429200 1004906 429252 1004912
rect 431966 1004958 432092 1004964
rect 431914 1004906 431966 1004912
rect 430026 1004864 430082 1004873
rect 430026 1004799 430028 1004808
rect 430080 1004799 430082 1004808
rect 430028 1004770 430080 1004776
rect 431682 1004728 431738 1004737
rect 431682 1004663 431684 1004672
rect 431736 1004663 431738 1004672
rect 431684 1004634 431736 1004640
rect 427820 1002584 427872 1002590
rect 427820 1002526 427872 1002532
rect 426346 1002280 426402 1002289
rect 426402 1002238 426572 1002266
rect 426346 1002215 426402 1002224
rect 426346 1002008 426402 1002017
rect 425060 1001972 425112 1001978
rect 426544 1001978 426572 1002238
rect 428370 1002008 428426 1002017
rect 426346 1001943 426348 1001952
rect 425060 1001914 425112 1001920
rect 426400 1001943 426402 1001952
rect 426532 1001972 426584 1001978
rect 426348 1001914 426400 1001920
rect 426532 1001914 426584 1001920
rect 427820 1001972 427872 1001978
rect 428370 1001943 428372 1001952
rect 427820 1001914 427872 1001920
rect 428424 1001943 428426 1001952
rect 431224 1001972 431276 1001978
rect 428372 1001914 428424 1001920
rect 431224 1001914 431276 1001920
rect 425072 997626 425100 1001914
rect 427832 999802 427860 1001914
rect 427820 999796 427872 999802
rect 427820 999738 427872 999744
rect 431236 997762 431264 1001914
rect 431224 997756 431276 997762
rect 431224 997698 431276 997704
rect 425060 997620 425112 997626
rect 425060 997562 425112 997568
rect 425060 996464 425112 996470
rect 425060 996406 425112 996412
rect 422944 994968 422996 994974
rect 422944 994910 422996 994916
rect 425072 994294 425100 996406
rect 432064 995994 432092 1004958
rect 432432 1004902 432460 1005060
rect 432420 1004896 432472 1004902
rect 432420 1004838 432472 1004844
rect 432236 1004828 432288 1004834
rect 432236 1004770 432288 1004776
rect 432248 996130 432276 1004770
rect 432236 996124 432288 996130
rect 432236 996066 432288 996072
rect 432052 995988 432104 995994
rect 432052 995930 432104 995936
rect 432616 995450 432644 1005110
rect 433524 1004692 433576 1004698
rect 433524 1004634 433576 1004640
rect 432880 1004080 432932 1004086
rect 432878 1004048 432880 1004057
rect 432932 1004048 432934 1004057
rect 432878 1003983 432934 1003992
rect 433338 1002144 433394 1002153
rect 433338 1002079 433340 1002088
rect 433392 1002079 433394 1002088
rect 433340 1002050 433392 1002056
rect 433536 995858 433564 1004634
rect 433996 995858 434024 1005518
rect 434168 1005032 434220 1005038
rect 434168 1004974 434220 1004980
rect 434180 995994 434208 1004974
rect 438124 1004896 438176 1004902
rect 438124 1004838 438176 1004844
rect 436744 1002108 436796 1002114
rect 436744 1002050 436796 1002056
rect 434168 995988 434220 995994
rect 434168 995930 434220 995936
rect 433524 995852 433576 995858
rect 433524 995794 433576 995800
rect 433984 995852 434036 995858
rect 433984 995794 434036 995800
rect 432604 995444 432656 995450
rect 432604 995386 432656 995392
rect 425060 994288 425112 994294
rect 425060 994230 425112 994236
rect 422208 988916 422260 988922
rect 422208 988858 422260 988864
rect 436756 985998 436784 1002050
rect 437480 999796 437532 999802
rect 437480 999738 437532 999744
rect 437492 997082 437520 999738
rect 438136 999122 438164 1004838
rect 439516 1001230 439544 1006810
rect 445024 1006596 445076 1006602
rect 445024 1006538 445076 1006544
rect 440884 1005848 440936 1005854
rect 440884 1005790 440936 1005796
rect 439504 1001224 439556 1001230
rect 439504 1001166 439556 1001172
rect 438124 999116 438176 999122
rect 438124 999058 438176 999064
rect 439872 997756 439924 997762
rect 439872 997698 439924 997704
rect 439688 997620 439740 997626
rect 439688 997562 439740 997568
rect 437480 997076 437532 997082
rect 437480 997018 437532 997024
rect 439700 996713 439728 997562
rect 439686 996704 439742 996713
rect 439686 996639 439742 996648
rect 439884 996441 439912 997698
rect 439870 996432 439926 996441
rect 439870 996367 439926 996376
rect 440896 995586 440924 1005790
rect 443644 1005440 443696 1005446
rect 443644 1005382 443696 1005388
rect 443460 999116 443512 999122
rect 443460 999058 443512 999064
rect 440884 995580 440936 995586
rect 440884 995522 440936 995528
rect 443472 993993 443500 999058
rect 443656 998782 443684 1005382
rect 445036 1002862 445064 1006538
rect 501694 1006496 501750 1006505
rect 447140 1006460 447192 1006466
rect 501694 1006431 501696 1006440
rect 447140 1006402 447192 1006408
rect 501748 1006431 501750 1006440
rect 501696 1006402 501748 1006408
rect 447152 1005446 447180 1006402
rect 502154 1006360 502210 1006369
rect 502154 1006295 502156 1006304
rect 502208 1006295 502210 1006304
rect 502156 1006266 502208 1006272
rect 500498 1006224 500554 1006233
rect 500498 1006159 500500 1006168
rect 500552 1006159 500554 1006168
rect 505744 1006188 505796 1006194
rect 500500 1006130 500552 1006136
rect 505744 1006130 505796 1006136
rect 499670 1006088 499726 1006097
rect 471244 1006052 471296 1006058
rect 505374 1006088 505430 1006097
rect 499670 1006023 499672 1006032
rect 471244 1005994 471296 1006000
rect 499724 1006023 499726 1006032
rect 502984 1006052 503036 1006058
rect 499672 1005994 499724 1006000
rect 505374 1006023 505376 1006032
rect 502984 1005994 503036 1006000
rect 505428 1006023 505430 1006032
rect 505376 1005994 505428 1006000
rect 451924 1005712 451976 1005718
rect 451924 1005654 451976 1005660
rect 449164 1005576 449216 1005582
rect 449164 1005518 449216 1005524
rect 447140 1005440 447192 1005446
rect 447140 1005382 447192 1005388
rect 445024 1002856 445076 1002862
rect 445024 1002798 445076 1002804
rect 446220 1002720 446272 1002726
rect 446220 1002662 446272 1002668
rect 446232 999802 446260 1002662
rect 446404 1001224 446456 1001230
rect 446404 1001166 446456 1001172
rect 446220 999796 446272 999802
rect 446220 999738 446272 999744
rect 443644 998776 443696 998782
rect 443644 998718 443696 998724
rect 445760 998776 445812 998782
rect 445760 998718 445812 998724
rect 445772 994809 445800 998718
rect 446416 998442 446444 1001166
rect 449176 999122 449204 1005518
rect 449164 999116 449216 999122
rect 449164 999058 449216 999064
rect 451740 999116 451792 999122
rect 451740 999058 451792 999064
rect 446404 998436 446456 998442
rect 446404 998378 446456 998384
rect 448520 997076 448572 997082
rect 448520 997018 448572 997024
rect 448532 994838 448560 997018
rect 451752 995081 451780 999058
rect 451936 999054 451964 1005654
rect 457444 1005440 457496 1005446
rect 457444 1005382 457496 1005388
rect 454684 1002856 454736 1002862
rect 454684 1002798 454736 1002804
rect 451924 999048 451976 999054
rect 451924 998990 451976 998996
rect 451738 995072 451794 995081
rect 451738 995007 451794 995016
rect 448520 994832 448572 994838
rect 445758 994800 445814 994809
rect 448520 994774 448572 994780
rect 445758 994735 445814 994744
rect 446128 994288 446180 994294
rect 454696 994265 454724 1002798
rect 456800 999048 456852 999054
rect 456800 998990 456852 998996
rect 456812 996169 456840 998990
rect 457456 997082 457484 1005382
rect 465724 1005304 465776 1005310
rect 465724 1005246 465776 1005252
rect 462320 1004080 462372 1004086
rect 462320 1004022 462372 1004028
rect 459560 999796 459612 999802
rect 459560 999738 459612 999744
rect 457444 997076 457496 997082
rect 457444 997018 457496 997024
rect 456798 996160 456854 996169
rect 456798 996095 456854 996104
rect 459572 994702 459600 999738
rect 459560 994696 459612 994702
rect 459560 994638 459612 994644
rect 446128 994230 446180 994236
rect 454682 994256 454738 994265
rect 443458 993984 443514 993993
rect 443458 993919 443514 993928
rect 414112 985992 414164 985998
rect 414112 985934 414164 985940
rect 415032 985992 415084 985998
rect 415032 985934 415084 985940
rect 430304 985992 430356 985998
rect 430304 985934 430356 985940
rect 436744 985992 436796 985998
rect 436744 985934 436796 985940
rect 414124 983620 414152 985934
rect 430316 983620 430344 985934
rect 446140 983634 446168 994230
rect 454682 994191 454738 994200
rect 462332 983634 462360 1004022
rect 465736 986134 465764 1005246
rect 467840 1003944 467892 1003950
rect 467840 1003886 467892 1003892
rect 467852 1001978 467880 1003886
rect 468760 1002584 468812 1002590
rect 468760 1002526 468812 1002532
rect 467840 1001972 467892 1001978
rect 467840 1001914 467892 1001920
rect 468772 994566 468800 1002526
rect 471256 996130 471284 1005994
rect 500500 1005304 500552 1005310
rect 500498 1005272 500500 1005281
rect 500552 1005272 500554 1005281
rect 500498 1005207 500554 1005216
rect 499670 1004864 499726 1004873
rect 498108 1004828 498160 1004834
rect 499670 1004799 499672 1004808
rect 498108 1004770 498160 1004776
rect 499724 1004799 499726 1004808
rect 499672 1004770 499724 1004776
rect 472624 1001972 472676 1001978
rect 472624 1001914 472676 1001920
rect 496728 1001972 496780 1001978
rect 496728 1001914 496780 1001920
rect 472440 998436 472492 998442
rect 472440 998378 472492 998384
rect 471796 997076 471848 997082
rect 471796 997018 471848 997024
rect 471244 996124 471296 996130
rect 471244 996066 471296 996072
rect 468760 994560 468812 994566
rect 471808 994537 471836 997018
rect 472452 995586 472480 998378
rect 472636 995761 472664 1001914
rect 472622 995752 472678 995761
rect 472622 995687 472678 995696
rect 477038 995752 477094 995761
rect 478326 995752 478382 995761
rect 477094 995710 477342 995738
rect 477038 995687 477094 995696
rect 485594 995752 485650 995761
rect 478382 995710 478630 995738
rect 485346 995710 485594 995738
rect 478326 995687 478382 995696
rect 485594 995687 485650 995696
rect 473372 995586 473662 995602
rect 472256 995580 472308 995586
rect 472256 995522 472308 995528
rect 472440 995580 472492 995586
rect 472440 995522 472492 995528
rect 473360 995580 473662 995586
rect 473412 995574 473662 995580
rect 473360 995522 473412 995528
rect 468760 994502 468812 994508
rect 471794 994528 471850 994537
rect 471794 994463 471850 994472
rect 472268 994430 472296 995522
rect 474094 995480 474150 995489
rect 474738 995480 474794 995489
rect 474150 995438 474306 995466
rect 474094 995415 474150 995424
rect 480810 995480 480866 995489
rect 474794 995438 474950 995466
rect 474738 995415 474794 995424
rect 476776 995081 476804 995452
rect 476762 995072 476818 995081
rect 476762 995007 476818 995016
rect 472256 994424 472308 994430
rect 472256 994366 472308 994372
rect 477972 993993 478000 995452
rect 480866 995438 481114 995466
rect 480810 995415 480866 995424
rect 481652 995058 481680 995452
rect 481560 995030 481680 995058
rect 481560 994537 481588 995030
rect 482296 994809 482324 995452
rect 482282 994800 482338 994809
rect 482282 994735 482338 994744
rect 482940 994566 482968 995452
rect 484136 994702 484164 995452
rect 484124 994696 484176 994702
rect 484124 994638 484176 994644
rect 482928 994560 482980 994566
rect 481546 994528 481602 994537
rect 482928 994502 482980 994508
rect 481546 994463 481602 994472
rect 485976 994430 486004 995452
rect 486620 994838 486648 995452
rect 486608 994832 486660 994838
rect 486608 994774 486660 994780
rect 487816 994702 487844 995452
rect 489736 995240 489788 995246
rect 489736 995182 489788 995188
rect 489748 994838 489776 995182
rect 489736 994832 489788 994838
rect 489736 994774 489788 994780
rect 487804 994696 487856 994702
rect 487804 994638 487856 994644
rect 485964 994424 486016 994430
rect 485964 994366 486016 994372
rect 477958 993984 478014 993993
rect 477958 993919 478014 993928
rect 496740 993342 496768 1001914
rect 496728 993336 496780 993342
rect 496728 993278 496780 993284
rect 465724 986128 465776 986134
rect 465724 986070 465776 986076
rect 495164 986128 495216 986134
rect 495164 986070 495216 986076
rect 478972 985992 479024 985998
rect 478972 985934 479024 985940
rect 446140 983606 446522 983634
rect 462332 983606 462806 983634
rect 478984 983620 479012 985934
rect 495176 983620 495204 986070
rect 498120 985046 498148 1004770
rect 501326 1004728 501382 1004737
rect 499488 1004692 499540 1004698
rect 501326 1004663 501328 1004672
rect 499488 1004634 499540 1004640
rect 501380 1004663 501382 1004672
rect 501328 1004634 501380 1004640
rect 498474 1002008 498530 1002017
rect 498474 1001943 498476 1001952
rect 498528 1001943 498530 1001952
rect 498476 1001914 498528 1001920
rect 499500 995042 499528 1004634
rect 502524 1002584 502576 1002590
rect 502522 1002552 502524 1002561
rect 502576 1002552 502578 1002561
rect 502522 1002487 502578 1002496
rect 500684 1002244 500736 1002250
rect 500684 1002186 500736 1002192
rect 500696 1001230 500724 1002186
rect 502248 1002108 502300 1002114
rect 502248 1002050 502300 1002056
rect 500868 1001972 500920 1001978
rect 500868 1001914 500920 1001920
rect 500684 1001224 500736 1001230
rect 500684 1001166 500736 1001172
rect 500880 997762 500908 1001914
rect 502260 998442 502288 1002050
rect 502522 1002008 502578 1002017
rect 502522 1001943 502524 1001952
rect 502576 1001943 502578 1001952
rect 502524 1001914 502576 1001920
rect 502248 998436 502300 998442
rect 502248 998378 502300 998384
rect 500868 997756 500920 997762
rect 500868 997698 500920 997704
rect 499488 995036 499540 995042
rect 499488 994978 499540 994984
rect 502996 994906 503024 1005994
rect 505008 1005576 505060 1005582
rect 505006 1005544 505008 1005553
rect 505060 1005544 505062 1005553
rect 505006 1005479 505062 1005488
rect 505376 1003944 505428 1003950
rect 505374 1003912 505376 1003921
rect 505428 1003912 505430 1003921
rect 505374 1003847 505430 1003856
rect 503350 1002280 503406 1002289
rect 503350 1002215 503352 1002224
rect 503404 1002215 503406 1002224
rect 503352 1002186 503404 1002192
rect 504178 1002144 504234 1002153
rect 504178 1002079 504180 1002088
rect 504232 1002079 504234 1002088
rect 504180 1002050 504232 1002056
rect 503350 1002008 503406 1002017
rect 503350 1001943 503352 1001952
rect 503404 1001943 503406 1001952
rect 504364 1001972 504416 1001978
rect 503352 1001914 503404 1001920
rect 504364 1001914 504416 1001920
rect 504376 998322 504404 1001914
rect 504376 998294 504588 998322
rect 504364 996260 504416 996266
rect 504364 996202 504416 996208
rect 504376 995858 504404 996202
rect 504364 995852 504416 995858
rect 504364 995794 504416 995800
rect 502984 994900 503036 994906
rect 502984 994842 503036 994848
rect 504560 994634 504588 998294
rect 505756 994770 505784 1006130
rect 514036 1006058 514064 1006878
rect 514024 1006052 514076 1006058
rect 514024 1005994 514076 1006000
rect 509056 1005848 509108 1005854
rect 509054 1005816 509056 1005825
rect 514024 1005848 514076 1005854
rect 509108 1005816 509110 1005825
rect 514024 1005790 514076 1005796
rect 509054 1005751 509110 1005760
rect 508228 1005440 508280 1005446
rect 508226 1005408 508228 1005417
rect 510988 1005440 511040 1005446
rect 508280 1005408 508282 1005417
rect 510988 1005382 511040 1005388
rect 508226 1005343 508282 1005352
rect 507032 1005168 507084 1005174
rect 507030 1005136 507032 1005145
rect 509700 1005168 509752 1005174
rect 507084 1005136 507086 1005145
rect 509700 1005110 509752 1005116
rect 507030 1005071 507086 1005080
rect 508228 1005032 508280 1005038
rect 508226 1005000 508228 1005009
rect 508280 1005000 508282 1005009
rect 508226 1004935 508282 1004944
rect 507860 1004896 507912 1004902
rect 507858 1004864 507860 1004873
rect 507912 1004864 507914 1004873
rect 507858 1004799 507914 1004808
rect 509054 1004728 509110 1004737
rect 509054 1004663 509056 1004672
rect 509108 1004663 509110 1004672
rect 509056 1004634 509108 1004640
rect 506202 1002008 506258 1002017
rect 507030 1002008 507086 1002017
rect 506202 1001943 506204 1001952
rect 506256 1001943 506258 1001952
rect 506492 1001966 507030 1001994
rect 506204 1001914 506256 1001920
rect 506492 995450 506520 1001966
rect 507030 1001943 507086 1001952
rect 507860 1001972 507912 1001978
rect 507860 1001914 507912 1001920
rect 507872 996130 507900 1001914
rect 509712 996130 509740 1005110
rect 510068 1004896 510120 1004902
rect 510068 1004838 510120 1004844
rect 509882 1002144 509938 1002153
rect 509882 1002079 509884 1002088
rect 509936 1002079 509938 1002088
rect 509884 1002050 509936 1002056
rect 507860 996124 507912 996130
rect 507860 996066 507912 996072
rect 509700 996124 509752 996130
rect 509700 996066 509752 996072
rect 510080 995858 510108 1004838
rect 510342 1004728 510398 1004737
rect 510342 1004663 510344 1004672
rect 510396 1004663 510398 1004672
rect 510344 1004634 510396 1004640
rect 510804 1004556 510856 1004562
rect 510804 1004498 510856 1004504
rect 510816 995994 510844 1004498
rect 511000 996266 511028 1005382
rect 511264 1005032 511316 1005038
rect 511264 1004974 511316 1004980
rect 510988 996260 511040 996266
rect 510988 996202 511040 996208
rect 511276 995994 511304 1004974
rect 512644 1002108 512696 1002114
rect 512644 1002050 512696 1002056
rect 510804 995988 510856 995994
rect 510804 995930 510856 995936
rect 511264 995988 511316 995994
rect 511264 995930 511316 995936
rect 511078 995888 511134 995897
rect 510068 995852 510120 995858
rect 511078 995823 511134 995832
rect 510068 995794 510120 995800
rect 506480 995444 506532 995450
rect 506480 995386 506532 995392
rect 505744 994764 505796 994770
rect 505744 994706 505796 994712
rect 504548 994628 504600 994634
rect 504548 994570 504600 994576
rect 498108 985040 498160 985046
rect 498108 984982 498160 984988
rect 511092 983634 511120 995823
rect 512656 991914 512684 1002050
rect 512644 991908 512696 991914
rect 512644 991850 512696 991856
rect 514036 985998 514064 1005790
rect 514220 997626 514248 1007014
rect 554136 1007004 554188 1007010
rect 559654 1006975 559656 1006984
rect 554136 1006946 554188 1006952
rect 559708 1006975 559710 1006984
rect 559656 1006946 559708 1006952
rect 552294 1006496 552350 1006505
rect 518164 1006460 518216 1006466
rect 518164 1006402 518216 1006408
rect 520924 1006460 520976 1006466
rect 552294 1006431 552296 1006440
rect 520924 1006402 520976 1006408
rect 552348 1006431 552350 1006440
rect 552296 1006402 552348 1006408
rect 516784 1006188 516836 1006194
rect 516784 1006130 516836 1006136
rect 515404 1004692 515456 1004698
rect 515404 1004634 515456 1004640
rect 514208 997620 514260 997626
rect 514208 997562 514260 997568
rect 515416 986134 515444 1004634
rect 516600 1003944 516652 1003950
rect 516600 1003886 516652 1003892
rect 516048 1002584 516100 1002590
rect 516048 1002526 516100 1002532
rect 516060 996266 516088 1002526
rect 516612 999122 516640 1003886
rect 516600 999116 516652 999122
rect 516600 999058 516652 999064
rect 516796 998578 516824 1006130
rect 516784 998572 516836 998578
rect 516784 998514 516836 998520
rect 517060 998436 517112 998442
rect 517060 998378 517112 998384
rect 516692 997756 516744 997762
rect 516692 997698 516744 997704
rect 516704 996441 516732 997698
rect 516876 997620 516928 997626
rect 516876 997562 516928 997568
rect 516888 996849 516916 997562
rect 516874 996840 516930 996849
rect 516874 996775 516930 996784
rect 516690 996432 516746 996441
rect 516690 996367 516746 996376
rect 516048 996260 516100 996266
rect 516048 996202 516100 996208
rect 517072 995081 517100 998378
rect 517058 995072 517114 995081
rect 517058 995007 517114 995016
rect 518176 994265 518204 1006402
rect 519544 1005304 519596 1005310
rect 519544 1005246 519596 1005252
rect 519556 996305 519584 1005246
rect 520004 1001224 520056 1001230
rect 520004 1001166 520056 1001172
rect 520016 997966 520044 1001166
rect 520188 999116 520240 999122
rect 520188 999058 520240 999064
rect 520004 997960 520056 997966
rect 520004 997902 520056 997908
rect 519542 996296 519598 996305
rect 519542 996231 519598 996240
rect 520200 995761 520228 999058
rect 520186 995752 520242 995761
rect 520186 995687 520242 995696
rect 520936 994537 520964 1006402
rect 551466 1006224 551522 1006233
rect 551466 1006159 551468 1006168
rect 551520 1006159 551522 1006168
rect 551468 1006130 551520 1006136
rect 551098 1006088 551154 1006097
rect 522304 1006052 522356 1006058
rect 551098 1006023 551154 1006032
rect 553122 1006088 553178 1006097
rect 553122 1006023 553124 1006032
rect 522304 1005994 522356 1006000
rect 522316 995178 522344 1005994
rect 522488 1005440 522540 1005446
rect 522488 1005382 522540 1005388
rect 522500 997830 522528 1005382
rect 551112 1005310 551140 1006023
rect 553176 1006023 553178 1006032
rect 553124 1005994 553176 1006000
rect 551100 1005304 551152 1005310
rect 551100 1005246 551152 1005252
rect 551928 1002312 551980 1002318
rect 551928 1002254 551980 1002260
rect 522948 998572 523000 998578
rect 522948 998514 523000 998520
rect 522488 997824 522540 997830
rect 522488 997766 522540 997772
rect 522304 995172 522356 995178
rect 522304 995114 522356 995120
rect 520922 994528 520978 994537
rect 520922 994463 520978 994472
rect 518162 994256 518218 994265
rect 518162 994191 518218 994200
rect 522960 993993 522988 998514
rect 523868 997960 523920 997966
rect 523868 997902 523920 997908
rect 549168 997960 549220 997966
rect 551100 997960 551152 997966
rect 549168 997902 549220 997908
rect 551098 997928 551100 997937
rect 551152 997928 551154 997937
rect 523684 996260 523736 996266
rect 523684 996202 523736 996208
rect 523696 995314 523724 996202
rect 523880 995450 523908 997902
rect 524052 997824 524104 997830
rect 524052 997766 524104 997772
rect 547788 997824 547840 997830
rect 547788 997766 547840 997772
rect 524064 995586 524092 997766
rect 526074 995752 526130 995761
rect 528006 995752 528062 995761
rect 526130 995710 526378 995738
rect 526074 995687 526130 995696
rect 528558 995752 528614 995761
rect 528062 995710 528218 995738
rect 528006 995687 528062 995696
rect 532790 995752 532846 995761
rect 528614 995710 528770 995738
rect 528558 995687 528614 995696
rect 536562 995752 536618 995761
rect 532846 995710 533094 995738
rect 532790 995687 532846 995696
rect 536618 995710 536774 995738
rect 536562 995687 536618 995696
rect 524800 995586 525090 995602
rect 524052 995580 524104 995586
rect 524052 995522 524104 995528
rect 524788 995580 525090 995586
rect 524840 995574 525090 995580
rect 524788 995522 524840 995528
rect 525352 995450 525734 995466
rect 529032 995450 529414 995466
rect 523868 995444 523920 995450
rect 523868 995386 523920 995392
rect 525340 995444 525734 995450
rect 525392 995438 525734 995444
rect 529020 995444 529414 995450
rect 525340 995386 525392 995392
rect 529072 995438 529414 995444
rect 529020 995386 529072 995392
rect 523684 995308 523736 995314
rect 523684 995250 523736 995256
rect 530044 995042 530072 995452
rect 532528 995081 532556 995452
rect 532514 995072 532570 995081
rect 530032 995036 530084 995042
rect 532514 995007 532570 995016
rect 530032 994978 530084 994984
rect 533724 994265 533752 995452
rect 534092 995438 534382 995466
rect 534092 995058 534120 995438
rect 534000 995030 534120 995058
rect 534000 994770 534028 995030
rect 533988 994764 534040 994770
rect 533988 994706 534040 994712
rect 535564 994537 535592 995452
rect 536852 995438 537418 995466
rect 536852 995058 536880 995438
rect 536760 995030 536880 995058
rect 535550 994528 535606 994537
rect 535550 994463 535606 994472
rect 533710 994256 533766 994265
rect 533710 994191 533766 994200
rect 536760 993993 536788 995030
rect 538048 994906 538076 995452
rect 538036 994900 538088 994906
rect 538036 994842 538088 994848
rect 539244 994770 539272 995452
rect 539232 994764 539284 994770
rect 539232 994706 539284 994712
rect 547800 994294 547828 997766
rect 549180 994430 549208 997902
rect 551098 997863 551154 997872
rect 550272 997824 550324 997830
rect 550270 997792 550272 997801
rect 551284 997824 551336 997830
rect 550324 997792 550326 997801
rect 551284 997766 551336 997772
rect 550270 997727 550326 997736
rect 551296 997354 551324 997766
rect 551940 997694 551968 1002254
rect 553308 1002040 553360 1002046
rect 553952 1002040 554004 1002046
rect 553308 1001982 553360 1001988
rect 553950 1002008 553952 1002017
rect 554004 1002008 554006 1002017
rect 553320 998646 553348 1001982
rect 553950 1001943 554006 1001952
rect 553308 998640 553360 998646
rect 553308 998582 553360 998588
rect 553122 998472 553178 998481
rect 553122 998407 553124 998416
rect 553176 998407 553178 998416
rect 553124 998378 553176 998384
rect 552296 997824 552348 997830
rect 552294 997792 552296 997801
rect 552348 997792 552350 997801
rect 552294 997727 552350 997736
rect 551928 997688 551980 997694
rect 551928 997630 551980 997636
rect 551284 997348 551336 997354
rect 551284 997290 551336 997296
rect 554148 995858 554176 1006946
rect 555146 1006904 555202 1006913
rect 555146 1006839 555148 1006848
rect 555200 1006839 555202 1006848
rect 562324 1006868 562376 1006874
rect 555148 1006810 555200 1006816
rect 562324 1006810 562376 1006816
rect 557170 1006768 557226 1006777
rect 557170 1006703 557172 1006712
rect 557224 1006703 557226 1006712
rect 557172 1006674 557224 1006680
rect 556802 1006496 556858 1006505
rect 554780 1006460 554832 1006466
rect 556802 1006431 556804 1006440
rect 554780 1006402 554832 1006408
rect 556856 1006431 556858 1006440
rect 556804 1006402 556856 1006408
rect 554318 1006360 554374 1006369
rect 554318 1006295 554320 1006304
rect 554372 1006295 554374 1006304
rect 554320 1006266 554372 1006272
rect 554792 1005582 554820 1006402
rect 562336 1006330 562364 1006810
rect 566648 1006732 566700 1006738
rect 566648 1006674 566700 1006680
rect 562324 1006324 562376 1006330
rect 562324 1006266 562376 1006272
rect 560850 1006224 560906 1006233
rect 555424 1006188 555476 1006194
rect 560850 1006159 560852 1006168
rect 555424 1006130 555476 1006136
rect 560904 1006159 560906 1006168
rect 563980 1006188 564032 1006194
rect 560852 1006130 560904 1006136
rect 563980 1006130 564032 1006136
rect 554780 1005576 554832 1005582
rect 554780 1005518 554832 1005524
rect 555148 1005440 555200 1005446
rect 555146 1005408 555148 1005417
rect 555200 1005408 555202 1005417
rect 555146 1005343 555202 1005352
rect 554320 1002312 554372 1002318
rect 554318 1002280 554320 1002289
rect 554372 1002280 554374 1002289
rect 554318 1002215 554374 1002224
rect 555148 998640 555200 998646
rect 555148 998582 555200 998588
rect 554136 995852 554188 995858
rect 554136 995794 554188 995800
rect 555160 995042 555188 998582
rect 555436 998578 555464 1006130
rect 556804 1006052 556856 1006058
rect 556804 1005994 556856 1006000
rect 555976 1005712 556028 1005718
rect 555974 1005680 555976 1005689
rect 556028 1005680 556030 1005689
rect 555974 1005615 556030 1005624
rect 555974 1004864 556030 1004873
rect 555974 1004799 555976 1004808
rect 556028 1004799 556030 1004808
rect 555976 1004770 556028 1004776
rect 555424 998572 555476 998578
rect 555424 998514 555476 998520
rect 556816 997218 556844 1005994
rect 563992 1005718 564020 1006130
rect 563060 1005712 563112 1005718
rect 563060 1005654 563112 1005660
rect 563980 1005712 564032 1005718
rect 563980 1005654 564032 1005660
rect 558184 1004828 558236 1004834
rect 558184 1004770 558236 1004776
rect 557630 1004728 557686 1004737
rect 557630 1004663 557632 1004672
rect 557684 1004663 557686 1004672
rect 557632 1004634 557684 1004640
rect 557998 1002688 558054 1002697
rect 557998 1002623 558000 1002632
rect 558052 1002623 558054 1002632
rect 558000 1002594 558052 1002600
rect 558000 1002448 558052 1002454
rect 557998 1002416 558000 1002425
rect 558052 1002416 558054 1002425
rect 557998 1002351 558054 1002360
rect 558196 997558 558224 1004770
rect 561678 1004728 561734 1004737
rect 559564 1004692 559616 1004698
rect 561678 1004663 561680 1004672
rect 559564 1004634 559616 1004640
rect 561732 1004663 561734 1004672
rect 561680 1004634 561732 1004640
rect 558826 1002824 558882 1002833
rect 558826 1002759 558828 1002768
rect 558880 1002759 558882 1002768
rect 558828 1002730 558880 1002736
rect 558826 1002008 558882 1002017
rect 558826 1001943 558828 1001952
rect 558880 1001943 558882 1001952
rect 558828 1001914 558880 1001920
rect 558184 997552 558236 997558
rect 558184 997494 558236 997500
rect 556804 997212 556856 997218
rect 556804 997154 556856 997160
rect 555148 995036 555200 995042
rect 555148 994978 555200 994984
rect 549168 994424 549220 994430
rect 549168 994366 549220 994372
rect 547788 994288 547840 994294
rect 547788 994230 547840 994236
rect 522946 993984 523002 993993
rect 522946 993919 523002 993928
rect 536746 993984 536802 993993
rect 536746 993919 536802 993928
rect 527640 991908 527692 991914
rect 527640 991850 527692 991856
rect 515404 986128 515456 986134
rect 515404 986070 515456 986076
rect 514024 985992 514076 985998
rect 514024 985934 514076 985940
rect 511092 983606 511474 983634
rect 527652 983620 527680 991850
rect 559576 986134 559604 1004634
rect 562324 1002788 562376 1002794
rect 562324 1002730 562376 1002736
rect 560300 1002652 560352 1002658
rect 560300 1002594 560352 1002600
rect 560024 1002176 560076 1002182
rect 560022 1002144 560024 1002153
rect 560076 1002144 560078 1002153
rect 560312 1002130 560340 1002594
rect 561036 1002448 561088 1002454
rect 561036 1002390 561088 1002396
rect 560484 1002312 560536 1002318
rect 560482 1002280 560484 1002289
rect 560536 1002280 560538 1002289
rect 560482 1002215 560538 1002224
rect 560312 1002102 560616 1002130
rect 560022 1002079 560078 1002088
rect 560392 1001972 560444 1001978
rect 560392 1001914 560444 1001920
rect 560404 996130 560432 1001914
rect 560392 996124 560444 996130
rect 560392 996066 560444 996072
rect 560588 995450 560616 1002102
rect 560852 1002040 560904 1002046
rect 560850 1002008 560852 1002017
rect 560904 1002008 560906 1002017
rect 560850 1001943 560906 1001952
rect 560576 995444 560628 995450
rect 560576 995386 560628 995392
rect 561048 992234 561076 1002390
rect 560956 992206 561076 992234
rect 543832 986128 543884 986134
rect 543832 986070 543884 986076
rect 559564 986128 559616 986134
rect 559564 986070 559616 986076
rect 543844 983620 543872 986070
rect 560116 985992 560168 985998
rect 560116 985934 560168 985940
rect 560128 983620 560156 985934
rect 560956 985182 560984 992206
rect 562336 987698 562364 1002730
rect 563072 1002590 563100 1005654
rect 566464 1004692 566516 1004698
rect 566464 1004634 566516 1004640
rect 563060 1002584 563112 1002590
rect 563060 1002526 563112 1002532
rect 563060 1002312 563112 1002318
rect 563060 1002254 563112 1002260
rect 562508 1002176 562560 1002182
rect 562508 1002118 562560 1002124
rect 562520 990282 562548 1002118
rect 563072 995994 563100 1002254
rect 565084 1002040 565136 1002046
rect 565084 1001982 565136 1001988
rect 563060 995988 563112 995994
rect 563060 995930 563112 995936
rect 563702 995616 563758 995625
rect 563702 995551 563758 995560
rect 563716 991914 563744 995551
rect 565096 994566 565124 1001982
rect 565084 994560 565136 994566
rect 565084 994502 565136 994508
rect 563704 991908 563756 991914
rect 563704 991850 563756 991856
rect 562508 990276 562560 990282
rect 562508 990218 562560 990224
rect 562324 987692 562376 987698
rect 562324 987634 562376 987640
rect 566476 986270 566504 1004634
rect 566660 996946 566688 1006674
rect 569224 1006460 569276 1006466
rect 569224 1006402 569276 1006408
rect 567844 1005848 567896 1005854
rect 567844 1005790 567896 1005796
rect 567856 997082 567884 1005790
rect 568488 998572 568540 998578
rect 568488 998514 568540 998520
rect 567844 997076 567896 997082
rect 567844 997018 567896 997024
rect 566648 996940 566700 996946
rect 566648 996882 566700 996888
rect 568500 994158 568528 998514
rect 569236 994770 569264 1006402
rect 571984 1006324 572036 1006330
rect 571984 1006266 572036 1006272
rect 570604 1005712 570656 1005718
rect 570604 1005654 570656 1005660
rect 569868 998436 569920 998442
rect 569868 998378 569920 998384
rect 569880 995178 569908 998378
rect 570236 997212 570288 997218
rect 570236 997154 570288 997160
rect 569868 995172 569920 995178
rect 569868 995114 569920 995120
rect 570248 994809 570276 997154
rect 570234 994800 570290 994809
rect 569224 994764 569276 994770
rect 570234 994735 570290 994744
rect 569224 994706 569276 994712
rect 568488 994152 568540 994158
rect 568488 994094 568540 994100
rect 566464 986264 566516 986270
rect 566464 986206 566516 986212
rect 570616 986134 570644 1005654
rect 571248 1002584 571300 1002590
rect 571248 1002526 571300 1002532
rect 571260 996810 571288 1002526
rect 571248 996804 571300 996810
rect 571248 996746 571300 996752
rect 571996 995314 572024 1006266
rect 574744 1006052 574796 1006058
rect 574744 1005994 574796 1006000
rect 573548 1005440 573600 1005446
rect 573548 1005382 573600 1005388
rect 573364 1005304 573416 1005310
rect 573364 1005246 573416 1005252
rect 572720 997348 572772 997354
rect 572720 997290 572772 997296
rect 572732 996130 572760 997290
rect 572720 996124 572772 996130
rect 572720 996066 572772 996072
rect 571984 995308 572036 995314
rect 571984 995250 572036 995256
rect 573376 994906 573404 1005246
rect 573560 997218 573588 1005382
rect 574756 997422 574784 1005994
rect 591120 998096 591172 998102
rect 591120 998038 591172 998044
rect 625804 998096 625856 998102
rect 625804 998038 625856 998044
rect 590568 997552 590620 997558
rect 590396 997500 590568 997506
rect 590396 997494 590620 997500
rect 590396 997478 590608 997494
rect 574744 997416 574796 997422
rect 574744 997358 574796 997364
rect 573548 997212 573600 997218
rect 573548 997154 573600 997160
rect 590396 996418 590424 997478
rect 590568 996940 590620 996946
rect 590568 996882 590620 996888
rect 590580 996713 590608 996882
rect 591132 996810 591160 998038
rect 621020 997960 621072 997966
rect 621020 997902 621072 997908
rect 625620 997960 625672 997966
rect 625620 997902 625672 997908
rect 591304 997824 591356 997830
rect 591304 997766 591356 997772
rect 591316 997422 591344 997766
rect 621032 997694 621060 997902
rect 625252 997824 625304 997830
rect 625252 997766 625304 997772
rect 621020 997688 621072 997694
rect 621020 997630 621072 997636
rect 591304 997416 591356 997422
rect 591304 997358 591356 997364
rect 622400 997212 622452 997218
rect 622400 997154 622452 997160
rect 618168 997076 618220 997082
rect 618168 997018 618220 997024
rect 591120 996804 591172 996810
rect 591120 996746 591172 996752
rect 590566 996704 590622 996713
rect 590566 996639 590622 996648
rect 590566 996432 590622 996441
rect 590396 996390 590566 996418
rect 590566 996367 590622 996376
rect 618180 995858 618208 997018
rect 618168 995852 618220 995858
rect 618168 995794 618220 995800
rect 622412 995450 622440 997154
rect 625264 996033 625292 997766
rect 625436 996124 625488 996130
rect 625436 996066 625488 996072
rect 625250 996024 625306 996033
rect 625250 995959 625306 995968
rect 625252 995852 625304 995858
rect 625252 995794 625304 995800
rect 625264 995586 625292 995794
rect 625252 995580 625304 995586
rect 625252 995522 625304 995528
rect 622400 995444 622452 995450
rect 622400 995386 622452 995392
rect 625448 995314 625476 996066
rect 625632 995761 625660 997902
rect 625618 995752 625674 995761
rect 625618 995687 625674 995696
rect 625816 995586 625844 998038
rect 627182 995752 627238 995761
rect 627918 995752 627974 995761
rect 627238 995710 627532 995738
rect 627182 995687 627238 995696
rect 629758 995752 629814 995761
rect 627974 995710 628176 995738
rect 627918 995687 627974 995696
rect 629814 995710 630016 995738
rect 629758 995687 629814 995696
rect 626552 995586 626888 995602
rect 625620 995580 625672 995586
rect 625620 995522 625672 995528
rect 625804 995580 625856 995586
rect 625804 995522 625856 995528
rect 626540 995580 626888 995586
rect 626592 995574 626888 995580
rect 634740 995574 634892 995602
rect 626540 995522 626592 995528
rect 625252 995308 625304 995314
rect 625252 995250 625304 995256
rect 625436 995308 625488 995314
rect 625436 995250 625488 995256
rect 625264 995042 625292 995250
rect 625632 995217 625660 995522
rect 630310 995480 630366 995489
rect 630366 995438 630568 995466
rect 630876 995438 631212 995466
rect 631520 995438 631856 995466
rect 634004 995438 634340 995466
rect 630310 995415 630366 995424
rect 625618 995208 625674 995217
rect 630128 995172 630180 995178
rect 625618 995143 625674 995152
rect 629588 995132 630128 995160
rect 629588 995042 629616 995132
rect 630128 995114 630180 995120
rect 625114 995036 625166 995042
rect 625114 994978 625166 994984
rect 625252 995036 625304 995042
rect 625252 994978 625304 994984
rect 629576 995036 629628 995042
rect 629576 994978 629628 994984
rect 625126 994922 625154 994978
rect 573364 994900 573416 994906
rect 625126 994894 625200 994922
rect 573364 994842 573416 994848
rect 625172 994634 625200 994894
rect 630876 994634 630904 995438
rect 631520 995314 631548 995438
rect 631508 995308 631560 995314
rect 631508 995250 631560 995256
rect 634004 995178 634032 995438
rect 634740 995217 634768 995574
rect 635200 995438 635536 995466
rect 635844 995438 636180 995466
rect 637040 995438 637376 995466
rect 638572 995438 638908 995466
rect 634726 995208 634782 995217
rect 633992 995172 634044 995178
rect 634726 995143 634782 995152
rect 633992 995114 634044 995120
rect 635200 995042 635228 995438
rect 635188 995036 635240 995042
rect 635188 994978 635240 994984
rect 625160 994628 625212 994634
rect 625160 994570 625212 994576
rect 630864 994628 630916 994634
rect 630864 994570 630916 994576
rect 592040 994560 592092 994566
rect 592040 994502 592092 994508
rect 576308 991908 576360 991914
rect 576308 991850 576360 991856
rect 570604 986128 570656 986134
rect 570604 986070 570656 986076
rect 560944 985176 560996 985182
rect 560944 985118 560996 985124
rect 576320 983620 576348 991850
rect 592052 983634 592080 994502
rect 635844 994158 635872 995438
rect 637040 994809 637068 995438
rect 638880 994945 638908 995438
rect 639064 995438 639216 995466
rect 639524 995438 639860 995466
rect 640720 995438 641056 995466
rect 638866 994936 638922 994945
rect 638866 994871 638922 994880
rect 637026 994800 637082 994809
rect 639064 994770 639092 995438
rect 639524 994906 639552 995438
rect 640720 995382 640748 995438
rect 640708 995376 640760 995382
rect 640708 995318 640760 995324
rect 640798 994936 640854 994945
rect 639512 994900 639564 994906
rect 640798 994871 640854 994880
rect 639512 994842 639564 994848
rect 637026 994735 637082 994744
rect 639052 994764 639104 994770
rect 639052 994706 639104 994712
rect 635832 994152 635884 994158
rect 635832 994094 635884 994100
rect 608784 986264 608836 986270
rect 608784 986206 608836 986212
rect 592052 983606 592526 983634
rect 608796 983620 608824 986206
rect 624976 986128 625028 986134
rect 624976 986070 625028 986076
rect 624988 983620 625016 986070
rect 640812 983634 640840 994871
rect 667940 994424 667992 994430
rect 667940 994366 667992 994372
rect 666560 994288 666612 994294
rect 666560 994230 666612 994236
rect 652760 993064 652812 993070
rect 652760 993006 652812 993012
rect 652484 992928 652536 992934
rect 652484 992870 652536 992876
rect 650920 991636 650972 991642
rect 650920 991578 650972 991584
rect 650092 990140 650144 990146
rect 650092 990082 650144 990088
rect 640812 983606 641194 983634
rect 62118 976032 62174 976041
rect 62118 975967 62174 975976
rect 62132 975730 62160 975967
rect 55864 975724 55916 975730
rect 55864 975666 55916 975672
rect 62120 975724 62172 975730
rect 62120 975666 62172 975672
rect 55876 969474 55904 975666
rect 55864 969468 55916 969474
rect 55864 969410 55916 969416
rect 62118 962976 62174 962985
rect 62118 962911 62174 962920
rect 62132 961926 62160 962911
rect 62120 961920 62172 961926
rect 62120 961862 62172 961868
rect 62118 949920 62174 949929
rect 62118 949855 62174 949864
rect 62132 946014 62160 949855
rect 62120 946008 62172 946014
rect 62120 945950 62172 945956
rect 51724 939820 51776 939826
rect 51724 939762 51776 939768
rect 62120 937032 62172 937038
rect 62118 937000 62120 937009
rect 62172 937000 62174 937009
rect 62118 936935 62174 936944
rect 44822 936184 44878 936193
rect 44822 936119 44878 936128
rect 44454 934144 44510 934153
rect 44454 934079 44510 934088
rect 44178 933736 44234 933745
rect 44178 933671 44234 933680
rect 42982 933328 43038 933337
rect 42982 933263 43038 933272
rect 42996 932958 43024 933263
rect 42984 932952 43036 932958
rect 42430 932920 42486 932929
rect 42984 932894 43036 932900
rect 54484 932952 54536 932958
rect 54484 932894 54536 932900
rect 42430 932855 42486 932864
rect 42798 932104 42854 932113
rect 42798 932039 42854 932048
rect 42812 931598 42840 932039
rect 42800 931592 42852 931598
rect 42800 931534 42852 931540
rect 53104 931592 53156 931598
rect 53104 931534 53156 931540
rect 47584 923296 47636 923302
rect 47584 923238 47636 923244
rect 46204 897048 46256 897054
rect 46204 896990 46256 896996
rect 42432 884740 42484 884746
rect 42432 884682 42484 884688
rect 42444 881929 42472 884682
rect 42430 881920 42486 881929
rect 42430 881855 42486 881864
rect 43444 870868 43496 870874
rect 43444 870810 43496 870816
rect 42062 818680 42118 818689
rect 42062 818615 42118 818624
rect 41878 818000 41934 818009
rect 41878 817935 41934 817944
rect 41696 815992 41748 815998
rect 41696 815934 41748 815940
rect 41604 815856 41656 815862
rect 41524 815804 41604 815810
rect 41524 815798 41656 815804
rect 41524 815782 41644 815798
rect 41524 814042 41552 815782
rect 41708 815658 42104 815674
rect 41696 815652 42116 815658
rect 41748 815646 42064 815652
rect 41696 815594 41748 815600
rect 42064 815594 42116 815600
rect 41708 814434 42104 814450
rect 41696 814428 42116 814434
rect 41748 814422 42064 814428
rect 41696 814370 41748 814376
rect 42064 814370 42116 814376
rect 42892 814428 42944 814434
rect 42892 814370 42944 814376
rect 41708 814298 42104 814314
rect 41696 814292 42116 814298
rect 41748 814286 42064 814292
rect 41696 814234 41748 814240
rect 42064 814234 42116 814240
rect 41786 814056 41842 814065
rect 41524 814014 41786 814042
rect 41786 813991 41842 814000
rect 41052 813000 41104 813006
rect 41052 812942 41104 812948
rect 41420 813000 41472 813006
rect 41420 812942 41472 812948
rect 40774 812832 40830 812841
rect 40774 812767 40830 812776
rect 35162 812424 35218 812433
rect 35162 812359 35218 812368
rect 32402 811200 32458 811209
rect 32402 811135 32458 811144
rect 31666 809976 31722 809985
rect 31666 809911 31722 809920
rect 31680 802330 31708 809911
rect 32416 802602 32444 811135
rect 33782 809568 33838 809577
rect 33782 809503 33838 809512
rect 32404 802596 32456 802602
rect 32404 802538 32456 802544
rect 31668 802324 31720 802330
rect 31668 802266 31720 802272
rect 33796 801106 33824 809503
rect 35176 803865 35204 812359
rect 40788 810762 40816 812767
rect 40958 812016 41014 812025
rect 40958 811951 41014 811960
rect 40776 810756 40828 810762
rect 40776 810698 40828 810704
rect 40972 809282 41000 811951
rect 41328 811776 41380 811782
rect 41328 811718 41380 811724
rect 41696 811776 41748 811782
rect 41696 811718 41748 811724
rect 41340 811617 41368 811718
rect 41326 811608 41382 811617
rect 41708 811594 41736 811718
rect 41708 811566 42288 811594
rect 41326 811543 41382 811552
rect 41696 810756 41748 810762
rect 41696 810698 41748 810704
rect 41708 810642 41736 810698
rect 41708 810626 42104 810642
rect 41708 810620 42116 810626
rect 41708 810614 42064 810620
rect 42064 810562 42116 810568
rect 41786 809296 41842 809305
rect 40972 809254 41786 809282
rect 41786 809231 41842 809240
rect 36542 809160 36598 809169
rect 36542 809095 36598 809104
rect 35162 803856 35218 803865
rect 35162 803791 35218 803800
rect 36556 801650 36584 809095
rect 41786 808344 41842 808353
rect 41524 808302 41786 808330
rect 41326 807528 41382 807537
rect 41326 807463 41382 807472
rect 41340 807362 41368 807463
rect 41328 807356 41380 807362
rect 41328 807298 41380 807304
rect 41524 805089 41552 808302
rect 41786 808279 41842 808288
rect 41696 807356 41748 807362
rect 42064 807356 42116 807362
rect 41748 807316 42064 807344
rect 41696 807298 41748 807304
rect 42064 807298 42116 807304
rect 42062 806712 42118 806721
rect 42062 806647 42118 806656
rect 41510 805080 41566 805089
rect 41510 805015 41566 805024
rect 41696 802596 41748 802602
rect 41696 802538 41748 802544
rect 41708 802482 41736 802538
rect 41708 802454 41828 802482
rect 39764 802324 39816 802330
rect 39764 802266 39816 802272
rect 39776 802097 39804 802266
rect 39762 802088 39818 802097
rect 39762 802023 39818 802032
rect 36544 801644 36596 801650
rect 36544 801586 36596 801592
rect 40316 801644 40368 801650
rect 40316 801586 40368 801592
rect 33784 801100 33836 801106
rect 33784 801042 33836 801048
rect 40328 800737 40356 801586
rect 40592 801100 40644 801106
rect 40592 801042 40644 801048
rect 40604 800737 40632 801042
rect 40314 800728 40370 800737
rect 40314 800663 40370 800672
rect 40590 800728 40646 800737
rect 40590 800663 40646 800672
rect 41800 800329 41828 802454
rect 42076 801394 42104 806647
rect 42260 804554 42288 811566
rect 42616 810620 42668 810626
rect 42616 810562 42668 810568
rect 42628 804554 42656 810562
rect 42260 804526 42380 804554
rect 42076 801366 42288 801394
rect 41786 800320 41842 800329
rect 41786 800255 41842 800264
rect 41786 799912 41842 799921
rect 41786 799847 41842 799856
rect 41800 799445 41828 799847
rect 42260 798266 42288 801366
rect 42182 798238 42288 798266
rect 42352 798266 42380 804526
rect 42444 804526 42656 804554
rect 42444 801258 42472 804526
rect 42706 802088 42762 802097
rect 42706 802023 42762 802032
rect 42444 801230 42564 801258
rect 42536 798386 42564 801230
rect 42524 798380 42576 798386
rect 42524 798322 42576 798328
rect 42352 798238 42472 798266
rect 42248 798176 42300 798182
rect 42248 798118 42300 798124
rect 42444 798130 42472 798238
rect 42260 797619 42288 798118
rect 42444 798102 42564 798130
rect 42182 797591 42288 797619
rect 42062 797328 42118 797337
rect 42062 797263 42118 797272
rect 42076 796960 42104 797263
rect 41786 796240 41842 796249
rect 41786 796175 41842 796184
rect 41800 795765 41828 796175
rect 42248 795660 42300 795666
rect 42248 795602 42300 795608
rect 42260 794594 42288 795602
rect 42182 794566 42288 794594
rect 41786 794472 41842 794481
rect 41786 794407 41842 794416
rect 41800 793900 41828 794407
rect 41786 793520 41842 793529
rect 41786 793455 41842 793464
rect 41800 793288 41828 793455
rect 42536 792758 42564 798102
rect 42182 792730 42564 792758
rect 42720 792134 42748 802023
rect 42904 794894 42932 814370
rect 43258 813648 43314 813657
rect 43258 813583 43314 813592
rect 43074 808752 43130 808761
rect 43074 808687 43130 808696
rect 43088 794894 43116 808687
rect 42536 792106 42748 792134
rect 42812 794866 42932 794894
rect 42996 794866 43116 794894
rect 42536 791738 42564 792106
rect 42260 791710 42564 791738
rect 42062 790664 42118 790673
rect 42062 790599 42118 790608
rect 42076 790228 42104 790599
rect 42260 790106 42288 791710
rect 42430 791616 42486 791625
rect 42430 791551 42486 791560
rect 42076 790078 42288 790106
rect 42076 789616 42104 790078
rect 42246 789984 42302 789993
rect 42246 789919 42302 789928
rect 42260 789426 42288 789919
rect 42168 789398 42288 789426
rect 42168 788936 42196 789398
rect 42444 788406 42472 791551
rect 42614 790256 42670 790265
rect 42614 790191 42670 790200
rect 42182 788378 42472 788406
rect 42246 788216 42302 788225
rect 42246 788151 42302 788160
rect 42260 786570 42288 788151
rect 42628 788066 42656 790191
rect 42182 786542 42288 786570
rect 42352 788038 42656 788066
rect 42352 785958 42380 788038
rect 42522 787944 42578 787953
rect 42522 787879 42578 787888
rect 42168 785890 42196 785944
rect 42260 785930 42380 785958
rect 42260 785890 42288 785930
rect 42168 785862 42288 785890
rect 42536 785278 42564 787879
rect 42182 785250 42564 785278
rect 8588 775132 8616 775268
rect 9048 775132 9076 775268
rect 9508 775132 9536 775268
rect 9968 775132 9996 775268
rect 10428 775132 10456 775268
rect 10888 775132 10916 775268
rect 11348 775132 11376 775268
rect 11808 775132 11836 775268
rect 12268 775132 12296 775268
rect 12728 775132 12756 775268
rect 13188 775132 13216 775268
rect 13648 775132 13676 775268
rect 14108 775132 14136 775268
rect 40038 775024 40094 775033
rect 40038 774959 40094 774968
rect 40052 774382 40080 774959
rect 35808 774376 35860 774382
rect 35806 774344 35808 774353
rect 40040 774376 40092 774382
rect 35860 774344 35862 774353
rect 40040 774318 40092 774324
rect 35806 774279 35862 774288
rect 35806 773936 35862 773945
rect 35806 773871 35862 773880
rect 35346 773528 35402 773537
rect 35346 773463 35402 773472
rect 35360 772886 35388 773463
rect 35532 773424 35584 773430
rect 35532 773366 35584 773372
rect 35544 773129 35572 773366
rect 35820 773294 35848 773871
rect 40868 773424 40920 773430
rect 40868 773366 40920 773372
rect 35808 773288 35860 773294
rect 35808 773230 35860 773236
rect 35808 773152 35860 773158
rect 35530 773120 35586 773129
rect 35530 773055 35586 773064
rect 35806 773120 35808 773129
rect 40880 773129 40908 773366
rect 41696 773152 41748 773158
rect 35860 773120 35862 773129
rect 35806 773055 35862 773064
rect 40866 773120 40922 773129
rect 42064 773152 42116 773158
rect 41748 773100 42064 773106
rect 41696 773094 42116 773100
rect 41708 773078 42104 773094
rect 40866 773055 40922 773064
rect 41696 773016 41748 773022
rect 42064 773016 42116 773022
rect 41748 772964 42064 772970
rect 41696 772958 42116 772964
rect 41708 772942 42104 772958
rect 35348 772880 35400 772886
rect 35348 772822 35400 772828
rect 41696 772744 41748 772750
rect 42064 772744 42116 772750
rect 41748 772692 42064 772698
rect 41696 772686 42116 772692
rect 41708 772670 42104 772686
rect 42812 772313 42840 794866
rect 42996 790673 43024 794866
rect 42982 790664 43038 790673
rect 42982 790599 43038 790608
rect 43074 773120 43130 773129
rect 43074 773055 43130 773064
rect 35346 772304 35402 772313
rect 35346 772239 35402 772248
rect 39762 772304 39818 772313
rect 39762 772239 39818 772248
rect 42798 772304 42854 772313
rect 42798 772239 42854 772248
rect 35360 771458 35388 772239
rect 39776 772070 39804 772239
rect 35900 772064 35952 772070
rect 35900 772006 35952 772012
rect 39764 772064 39816 772070
rect 39764 772006 39816 772012
rect 35532 771928 35584 771934
rect 35530 771896 35532 771905
rect 35584 771896 35586 771905
rect 35530 771831 35586 771840
rect 35716 771656 35768 771662
rect 35716 771598 35768 771604
rect 35728 771497 35756 771598
rect 35912 771594 35940 772006
rect 39856 771928 39908 771934
rect 39856 771870 39908 771876
rect 35900 771588 35952 771594
rect 35900 771530 35952 771536
rect 35714 771488 35770 771497
rect 35348 771452 35400 771458
rect 35714 771423 35770 771432
rect 39118 771488 39174 771497
rect 39118 771423 39120 771432
rect 35348 771394 35400 771400
rect 39172 771423 39174 771432
rect 39120 771394 39172 771400
rect 39868 771089 39896 771870
rect 35438 771080 35494 771089
rect 35438 771015 35494 771024
rect 39854 771080 39910 771089
rect 39854 771015 39910 771024
rect 42890 771080 42946 771089
rect 42890 771015 42946 771024
rect 35452 770098 35480 771015
rect 35622 770672 35678 770681
rect 35622 770607 35678 770616
rect 35636 770234 35664 770607
rect 35808 770500 35860 770506
rect 35808 770442 35860 770448
rect 41420 770500 41472 770506
rect 41420 770442 41472 770448
rect 35820 770273 35848 770442
rect 41432 770273 41460 770442
rect 41696 770296 41748 770302
rect 35806 770264 35862 770273
rect 35624 770228 35676 770234
rect 35806 770199 35862 770208
rect 41418 770264 41474 770273
rect 42064 770296 42116 770302
rect 41748 770244 42064 770250
rect 41696 770238 42116 770244
rect 41708 770222 42104 770238
rect 41418 770199 41474 770208
rect 35624 770170 35676 770176
rect 41708 770098 42104 770114
rect 35440 770092 35492 770098
rect 35440 770034 35492 770040
rect 41696 770092 42116 770098
rect 41748 770086 42064 770092
rect 41696 770034 41748 770040
rect 42064 770034 42116 770040
rect 35346 769448 35402 769457
rect 35346 769383 35402 769392
rect 35360 768738 35388 769383
rect 35530 769040 35586 769049
rect 35530 768975 35586 768984
rect 35806 769040 35862 769049
rect 35806 768975 35808 768984
rect 35544 768874 35572 768975
rect 35860 768975 35862 768984
rect 39856 769004 39908 769010
rect 35808 768946 35860 768952
rect 39856 768946 39908 768952
rect 35532 768868 35584 768874
rect 35532 768810 35584 768816
rect 39304 768868 39356 768874
rect 39304 768810 39356 768816
rect 35348 768732 35400 768738
rect 35348 768674 35400 768680
rect 35806 767816 35862 767825
rect 35806 767751 35862 767760
rect 32402 767408 32458 767417
rect 35820 767378 35848 767751
rect 32402 767343 32458 767352
rect 35808 767372 35860 767378
rect 32416 759665 32444 767343
rect 35808 767314 35860 767320
rect 36544 767372 36596 767378
rect 36544 767314 36596 767320
rect 35162 767000 35218 767009
rect 35162 766935 35218 766944
rect 32402 759656 32458 759665
rect 32402 759591 32458 759600
rect 35176 758334 35204 766935
rect 35806 766592 35862 766601
rect 35806 766527 35862 766536
rect 35820 766358 35848 766527
rect 35808 766352 35860 766358
rect 35808 766294 35860 766300
rect 35806 766184 35862 766193
rect 35806 766119 35862 766128
rect 35820 765950 35848 766119
rect 35808 765944 35860 765950
rect 35808 765886 35860 765892
rect 35808 764720 35860 764726
rect 35808 764662 35860 764668
rect 35820 764561 35848 764662
rect 35806 764552 35862 764561
rect 35806 764487 35862 764496
rect 35622 764144 35678 764153
rect 35622 764079 35678 764088
rect 35636 763298 35664 764079
rect 35806 763736 35862 763745
rect 35806 763671 35808 763680
rect 35860 763671 35862 763680
rect 35808 763642 35860 763648
rect 35624 763292 35676 763298
rect 35624 763234 35676 763240
rect 35806 762920 35862 762929
rect 35806 762855 35862 762864
rect 35820 761938 35848 762855
rect 35808 761932 35860 761938
rect 35808 761874 35860 761880
rect 36556 759082 36584 767314
rect 37924 763700 37976 763706
rect 37924 763642 37976 763648
rect 36544 759076 36596 759082
rect 36544 759018 36596 759024
rect 35164 758328 35216 758334
rect 35164 758270 35216 758276
rect 37936 757790 37964 763642
rect 37924 757784 37976 757790
rect 39316 757761 39344 768810
rect 39868 768641 39896 768946
rect 40040 768732 40092 768738
rect 40040 768674 40092 768680
rect 39854 768632 39910 768641
rect 39854 768567 39910 768576
rect 40052 765406 40080 768674
rect 42706 768632 42762 768641
rect 42706 768567 42762 768576
rect 42246 768360 42302 768369
rect 42246 768295 42302 768304
rect 40408 766216 40460 766222
rect 40406 766184 40408 766193
rect 40460 766184 40462 766193
rect 40406 766119 40462 766128
rect 41696 766012 41748 766018
rect 41696 765954 41748 765960
rect 41708 765898 41736 765954
rect 42076 765950 42104 765981
rect 42064 765944 42116 765950
rect 41892 765898 42064 765914
rect 41708 765892 42064 765898
rect 41708 765886 42116 765892
rect 41708 765870 41920 765886
rect 40040 765400 40092 765406
rect 40040 765342 40092 765348
rect 41696 765400 41748 765406
rect 41696 765342 41748 765348
rect 40408 764720 40460 764726
rect 40408 764662 40460 764668
rect 40420 764561 40448 764662
rect 40406 764552 40462 764561
rect 40406 764487 40462 764496
rect 41510 763328 41566 763337
rect 41510 763263 41512 763272
rect 41564 763263 41566 763272
rect 41512 763234 41564 763240
rect 40500 761932 40552 761938
rect 40500 761874 40552 761880
rect 40512 760345 40540 761874
rect 40498 760336 40554 760345
rect 40498 760271 40554 760280
rect 41420 759076 41472 759082
rect 41420 759018 41472 759024
rect 40408 758328 40460 758334
rect 40406 758296 40408 758305
rect 40460 758296 40462 758305
rect 40406 758231 40462 758240
rect 37924 757726 37976 757732
rect 39302 757752 39358 757761
rect 39302 757687 39358 757696
rect 41432 757353 41460 759018
rect 41708 758010 41736 765342
rect 42260 763154 42288 768295
rect 42260 763126 42380 763154
rect 42352 761138 42380 763126
rect 42352 761110 42656 761138
rect 42430 758296 42486 758305
rect 42430 758231 42486 758240
rect 41708 757982 42380 758010
rect 41696 757784 41748 757790
rect 41748 757732 41828 757738
rect 41696 757726 41828 757732
rect 41708 757710 41828 757726
rect 41418 757344 41474 757353
rect 41418 757279 41474 757288
rect 41800 757058 41828 757710
rect 41800 757030 42288 757058
rect 41786 756664 41842 756673
rect 41786 756599 41842 756608
rect 41800 756226 41828 756599
rect 42168 755018 42196 755072
rect 42260 755018 42288 757030
rect 42168 754990 42288 755018
rect 42352 754882 42380 757982
rect 42168 754854 42380 754882
rect 42168 754392 42196 754854
rect 42444 754746 42472 758231
rect 42260 754718 42472 754746
rect 42062 754080 42118 754089
rect 42062 754015 42118 754024
rect 42076 753780 42104 754015
rect 42062 752992 42118 753001
rect 42062 752927 42118 752936
rect 42076 752556 42104 752927
rect 42260 751641 42288 754718
rect 42432 754520 42484 754526
rect 42432 754462 42484 754468
rect 42246 751632 42302 751641
rect 42246 751567 42302 751576
rect 42444 751482 42472 754462
rect 42168 751454 42472 751482
rect 42168 751369 42196 751454
rect 41786 751088 41842 751097
rect 42628 751074 42656 761110
rect 41786 751023 41842 751032
rect 42352 751046 42656 751074
rect 41800 750720 41828 751023
rect 41786 750408 41842 750417
rect 41786 750343 41842 750352
rect 41800 750108 41828 750343
rect 42352 749543 42380 751046
rect 42720 750802 42748 768567
rect 42628 750774 42748 750802
rect 42628 750666 42656 750774
rect 42628 750638 42840 750666
rect 42614 750544 42670 750553
rect 42614 750479 42670 750488
rect 42182 749515 42380 749543
rect 42430 749456 42486 749465
rect 42430 749391 42486 749400
rect 42248 748604 42300 748610
rect 42248 748546 42300 748552
rect 42260 747182 42288 748546
rect 42248 747176 42300 747182
rect 42248 747118 42300 747124
rect 42444 747062 42472 749391
rect 42182 747034 42472 747062
rect 42248 746904 42300 746910
rect 42248 746846 42300 746852
rect 42260 746415 42288 746846
rect 42628 746450 42656 750479
rect 42812 750394 42840 750638
rect 42182 746387 42288 746415
rect 42444 746422 42656 746450
rect 42720 750366 42840 750394
rect 42444 745770 42472 746422
rect 42182 745742 42472 745770
rect 42246 745648 42302 745657
rect 42246 745583 42302 745592
rect 42260 745346 42288 745583
rect 42248 745340 42300 745346
rect 42248 745282 42300 745288
rect 42720 745226 42748 750366
rect 42182 745198 42748 745226
rect 42248 745136 42300 745142
rect 42248 745078 42300 745084
rect 42430 745104 42486 745113
rect 41786 743744 41842 743753
rect 41786 743679 41842 743688
rect 41800 743376 41828 743679
rect 42260 743050 42288 745078
rect 42430 745039 42486 745048
rect 42168 743022 42288 743050
rect 42168 742696 42196 743022
rect 42444 742098 42472 745039
rect 42182 742070 42472 742098
rect 8588 731884 8616 732020
rect 9048 731884 9076 732020
rect 9508 731884 9536 732020
rect 9968 731884 9996 732020
rect 10428 731884 10456 732020
rect 10888 731884 10916 732020
rect 11348 731884 11376 732020
rect 11808 731884 11836 732020
rect 12268 731884 12296 732020
rect 12728 731884 12756 732020
rect 13188 731884 13216 732020
rect 13648 731884 13676 732020
rect 14108 731884 14136 732020
rect 42432 731196 42484 731202
rect 42432 731138 42484 731144
rect 42444 730969 42472 731138
rect 42430 730960 42486 730969
rect 42430 730895 42486 730904
rect 41142 730552 41198 730561
rect 41142 730487 41198 730496
rect 41156 730114 41184 730487
rect 41144 730108 41196 730114
rect 41144 730050 41196 730056
rect 41696 730108 41748 730114
rect 42064 730108 42116 730114
rect 41748 730068 42064 730096
rect 41696 730050 41748 730056
rect 42064 730050 42116 730056
rect 42904 729337 42932 771015
rect 43088 730153 43116 773055
rect 43272 770302 43300 813583
rect 43260 770296 43312 770302
rect 43260 770238 43312 770244
rect 43258 766184 43314 766193
rect 43258 766119 43314 766128
rect 43272 748610 43300 766119
rect 43456 754089 43484 870810
rect 44824 844620 44876 844626
rect 44824 844562 44876 844568
rect 44180 814292 44232 814298
rect 44180 814234 44232 814240
rect 43628 799060 43680 799066
rect 43628 799002 43680 799008
rect 43640 797337 43668 799002
rect 43626 797328 43682 797337
rect 43626 797263 43682 797272
rect 44192 771497 44220 814234
rect 44454 814056 44510 814065
rect 44454 813991 44510 814000
rect 44468 773158 44496 813991
rect 44638 807936 44694 807945
rect 44638 807871 44694 807880
rect 44652 796346 44680 807871
rect 44640 796340 44692 796346
rect 44640 796282 44692 796288
rect 44836 775033 44864 844562
rect 46216 819097 46244 896990
rect 46202 819088 46258 819097
rect 46202 819023 46258 819032
rect 46202 806304 46258 806313
rect 46202 806239 46258 806248
rect 44822 775024 44878 775033
rect 44822 774959 44878 774968
rect 44456 773152 44508 773158
rect 44456 773094 44508 773100
rect 44178 771488 44234 771497
rect 44178 771423 44234 771432
rect 44270 770264 44326 770273
rect 44270 770199 44326 770208
rect 43628 767372 43680 767378
rect 43628 767314 43680 767320
rect 43442 754080 43498 754089
rect 43442 754015 43498 754024
rect 43260 748604 43312 748610
rect 43260 748546 43312 748552
rect 43074 730144 43130 730153
rect 43074 730079 43130 730088
rect 42890 729328 42946 729337
rect 42890 729263 42946 729272
rect 40866 728682 40922 728691
rect 40866 728617 40922 728626
rect 40880 727326 40908 728617
rect 43074 728104 43130 728113
rect 43074 728039 43130 728048
rect 41708 727666 42104 727682
rect 41696 727660 42116 727666
rect 41748 727654 42064 727660
rect 41696 727602 41748 727608
rect 42064 727602 42116 727608
rect 42892 727660 42944 727666
rect 42892 727602 42944 727608
rect 41052 727592 41104 727598
rect 41052 727534 41104 727540
rect 41064 727467 41092 727534
rect 41708 727530 42104 727546
rect 41696 727524 42116 727530
rect 41748 727518 42064 727524
rect 41050 727458 41106 727467
rect 41050 727393 41106 727402
rect 41326 727458 41382 727467
rect 41696 727466 41748 727472
rect 42064 727466 42116 727472
rect 41326 727393 41382 727402
rect 40868 727320 40920 727326
rect 40868 727262 40920 727268
rect 41696 727320 41748 727326
rect 42064 727320 42116 727326
rect 41748 727268 42064 727274
rect 41696 727262 42116 727268
rect 41708 727246 42104 727262
rect 41142 726880 41198 726889
rect 41142 726815 41198 726824
rect 40958 726234 41014 726243
rect 40958 726169 41014 726178
rect 37922 725248 37978 725257
rect 37922 725183 37978 725192
rect 35162 724840 35218 724849
rect 35162 724775 35218 724784
rect 33046 724432 33102 724441
rect 33046 724367 33102 724376
rect 31758 720352 31814 720361
rect 31758 720287 31760 720296
rect 31812 720287 31814 720296
rect 31760 720258 31812 720264
rect 33060 716825 33088 724367
rect 33782 723786 33838 723795
rect 33782 723721 33838 723730
rect 33046 716816 33102 716825
rect 33046 716751 33102 716760
rect 33796 715290 33824 723721
rect 35176 715698 35204 724775
rect 35164 715692 35216 715698
rect 35164 715634 35216 715640
rect 37936 715426 37964 725183
rect 40682 723208 40738 723217
rect 40682 723143 40738 723152
rect 40040 720316 40092 720322
rect 40040 720258 40092 720264
rect 39212 715692 39264 715698
rect 39212 715634 39264 715640
rect 37924 715420 37976 715426
rect 37924 715362 37976 715368
rect 33784 715284 33836 715290
rect 33784 715226 33836 715232
rect 39224 715193 39252 715634
rect 39210 715184 39266 715193
rect 39210 715119 39266 715128
rect 40052 714241 40080 720258
rect 40696 714270 40724 723143
rect 40972 721754 41000 726169
rect 41156 726102 41184 726815
rect 41326 726234 41382 726243
rect 41326 726169 41382 726178
rect 41696 726232 41748 726238
rect 42064 726232 42116 726238
rect 41748 726192 42064 726220
rect 41696 726174 41748 726180
rect 42064 726174 42116 726180
rect 42524 726232 42576 726238
rect 42524 726174 42576 726180
rect 41144 726096 41196 726102
rect 41144 726038 41196 726044
rect 41604 726096 41656 726102
rect 41604 726038 41656 726044
rect 41616 725778 41644 726038
rect 41786 725792 41842 725801
rect 41616 725750 41786 725778
rect 41786 725727 41842 725736
rect 41326 725656 41382 725665
rect 41326 725591 41382 725600
rect 41142 721768 41198 721777
rect 40972 721726 41142 721754
rect 41142 721703 41198 721712
rect 41340 714513 41368 725591
rect 41786 722392 41842 722401
rect 41786 722327 41842 722336
rect 41800 718593 41828 722327
rect 41786 718584 41842 718593
rect 41786 718519 41842 718528
rect 41512 715420 41564 715426
rect 41512 715362 41564 715368
rect 41326 714504 41382 714513
rect 41326 714439 41382 714448
rect 40684 714264 40736 714270
rect 40038 714232 40094 714241
rect 41524 714241 41552 715362
rect 41696 715284 41748 715290
rect 41748 715244 41920 715272
rect 41696 715226 41748 715232
rect 41696 714264 41748 714270
rect 40684 714206 40736 714212
rect 41510 714232 41566 714241
rect 40038 714167 40094 714176
rect 41892 714252 41920 715244
rect 42536 715193 42564 726174
rect 42338 715184 42394 715193
rect 42338 715119 42394 715128
rect 42522 715184 42578 715193
rect 42522 715119 42578 715128
rect 42064 714264 42116 714270
rect 41892 714224 42064 714252
rect 41748 714212 41828 714218
rect 41696 714206 41828 714212
rect 42064 714206 42116 714212
rect 41708 714190 41828 714206
rect 41510 714167 41566 714176
rect 41800 713969 41828 714190
rect 41786 713960 41842 713969
rect 41786 713895 41842 713904
rect 42352 713810 42380 715119
rect 42522 714504 42578 714513
rect 42522 714439 42578 714448
rect 42352 713782 42472 713810
rect 42444 713062 42472 713782
rect 42536 713474 42564 714439
rect 42708 714264 42760 714270
rect 42708 714206 42760 714212
rect 42536 713446 42656 713474
rect 42182 713034 42472 713062
rect 41786 712192 41842 712201
rect 41786 712127 41842 712136
rect 41800 711824 41828 712127
rect 42154 711648 42210 711657
rect 42154 711583 42210 711592
rect 42168 711212 42196 711583
rect 42248 711136 42300 711142
rect 42248 711078 42300 711084
rect 42260 710575 42288 711078
rect 42182 710547 42288 710575
rect 42246 710424 42302 710433
rect 42246 710359 42302 710368
rect 42260 709390 42288 710359
rect 42182 709362 42288 709390
rect 42246 709200 42302 709209
rect 42246 709135 42302 709144
rect 41786 708520 41842 708529
rect 41786 708455 41842 708464
rect 41800 708152 41828 708455
rect 42062 707840 42118 707849
rect 42062 707775 42118 707784
rect 42076 707540 42104 707775
rect 42260 707146 42288 709135
rect 42430 707296 42486 707305
rect 42430 707231 42486 707240
rect 42168 707118 42288 707146
rect 42168 706860 42196 707118
rect 42062 706616 42118 706625
rect 42062 706551 42118 706560
rect 42248 706580 42300 706586
rect 42076 706316 42104 706551
rect 42248 706522 42300 706528
rect 42260 704274 42288 706522
rect 42248 704268 42300 704274
rect 42248 704210 42300 704216
rect 42444 704154 42472 707231
rect 42076 704126 42472 704154
rect 42076 703868 42104 704126
rect 42248 704064 42300 704070
rect 42248 704006 42300 704012
rect 42260 703338 42288 704006
rect 42168 703310 42288 703338
rect 42168 703188 42196 703310
rect 42628 703202 42656 713446
rect 42444 703174 42656 703202
rect 42156 702908 42208 702914
rect 42156 702850 42208 702856
rect 42168 702794 42196 702850
rect 41984 702766 42196 702794
rect 41984 702576 42012 702766
rect 42444 702434 42472 703174
rect 42720 702914 42748 714206
rect 42708 702908 42760 702914
rect 42708 702850 42760 702856
rect 42614 702536 42670 702545
rect 42614 702471 42670 702480
rect 42260 702406 42472 702434
rect 42168 701978 42196 702032
rect 42260 701978 42288 702406
rect 42168 701950 42288 701978
rect 42430 701448 42486 701457
rect 42430 701383 42486 701392
rect 42246 701176 42302 701185
rect 42246 701111 42302 701120
rect 42064 700596 42116 700602
rect 42064 700538 42116 700544
rect 42076 700165 42104 700538
rect 42260 699530 42288 701111
rect 42182 699502 42288 699530
rect 42444 698918 42472 701383
rect 42628 700602 42656 702471
rect 42904 702434 42932 727602
rect 42812 702406 42932 702434
rect 42616 700596 42668 700602
rect 42616 700538 42668 700544
rect 42168 698850 42196 698904
rect 42260 698890 42472 698918
rect 42260 698850 42288 698890
rect 42168 698822 42288 698850
rect 8588 688772 8616 688908
rect 9048 688772 9076 688908
rect 9508 688772 9536 688908
rect 9968 688772 9996 688908
rect 10428 688772 10456 688908
rect 10888 688772 10916 688908
rect 11348 688772 11376 688908
rect 11808 688772 11836 688908
rect 12268 688772 12296 688908
rect 12728 688772 12756 688908
rect 13188 688772 13216 688908
rect 13648 688772 13676 688908
rect 14108 688772 14136 688908
rect 40958 688392 41014 688401
rect 40958 688327 41014 688336
rect 40972 687274 41000 688327
rect 42524 687744 42576 687750
rect 42524 687686 42576 687692
rect 42536 687313 42564 687686
rect 42522 687304 42578 687313
rect 40960 687268 41012 687274
rect 40960 687210 41012 687216
rect 41696 687268 41748 687274
rect 42064 687268 42116 687274
rect 41748 687228 42064 687256
rect 41696 687210 41748 687216
rect 42522 687239 42578 687248
rect 42064 687210 42116 687216
rect 41142 686896 41198 686905
rect 41142 686831 41198 686840
rect 40866 685910 40922 685919
rect 41156 685914 41184 686831
rect 41696 686112 41748 686118
rect 42064 686112 42116 686118
rect 41748 686060 42064 686066
rect 41696 686054 42116 686060
rect 41328 686044 41380 686050
rect 41708 686038 42104 686054
rect 41328 685986 41380 685992
rect 41340 685919 41368 685986
rect 40866 685845 40922 685854
rect 41144 685908 41196 685914
rect 41144 685850 41196 685856
rect 41326 685910 41382 685919
rect 41326 685845 41382 685854
rect 41696 685908 41748 685914
rect 42064 685908 42116 685914
rect 41748 685868 42064 685896
rect 41696 685850 41748 685856
rect 42064 685850 42116 685856
rect 40880 684826 40908 685845
rect 41142 685264 41198 685273
rect 41142 685199 41198 685208
rect 40868 684820 40920 684826
rect 40868 684762 40920 684768
rect 40774 684686 40830 684695
rect 41156 684690 41184 685199
rect 41696 684752 41748 684758
rect 42064 684752 42116 684758
rect 41748 684700 42064 684706
rect 41696 684694 42116 684700
rect 40774 684621 40830 684630
rect 41144 684684 41196 684690
rect 41708 684678 42104 684694
rect 41144 684626 41196 684632
rect 40788 683330 40816 684621
rect 41708 684554 42104 684570
rect 41696 684548 42116 684554
rect 41748 684542 42064 684548
rect 41696 684490 41748 684496
rect 42064 684490 42116 684496
rect 41142 684040 41198 684049
rect 41142 683975 41198 683984
rect 40958 683632 41014 683641
rect 40958 683567 41014 683576
rect 40776 683324 40828 683330
rect 40776 683266 40828 683272
rect 34426 682408 34482 682417
rect 40972 682394 41000 683567
rect 41156 683194 41184 683975
rect 41708 683602 42104 683618
rect 41328 683596 41380 683602
rect 41328 683538 41380 683544
rect 41696 683596 42104 683602
rect 41748 683590 42104 683596
rect 41696 683538 41748 683544
rect 41340 683233 41368 683538
rect 42076 683534 42104 683590
rect 42064 683528 42116 683534
rect 42064 683470 42116 683476
rect 42524 683528 42576 683534
rect 42524 683470 42576 683476
rect 42064 683392 42116 683398
rect 41708 683340 42064 683346
rect 41708 683334 42116 683340
rect 41708 683330 42104 683334
rect 41696 683324 42104 683330
rect 41748 683318 42104 683324
rect 41696 683266 41748 683272
rect 41326 683224 41382 683233
rect 41144 683188 41196 683194
rect 41326 683159 41382 683168
rect 41696 683188 41748 683194
rect 41144 683130 41196 683136
rect 42064 683188 42116 683194
rect 41748 683148 42064 683176
rect 41696 683130 41748 683136
rect 42064 683130 42116 683136
rect 41326 682816 41382 682825
rect 41326 682751 41382 682760
rect 41340 682514 41368 682751
rect 41328 682508 41380 682514
rect 41328 682450 41380 682456
rect 41786 682408 41842 682417
rect 40972 682366 41786 682394
rect 34426 682343 34482 682352
rect 41786 682343 41842 682352
rect 32402 681184 32458 681193
rect 32402 681119 32458 681128
rect 31022 680776 31078 680785
rect 31022 680711 31078 680720
rect 31036 672722 31064 680711
rect 32416 672761 32444 681119
rect 34440 675510 34468 682343
rect 41328 682304 41380 682310
rect 41328 682246 41380 682252
rect 40682 682000 40738 682009
rect 40682 681935 40738 681944
rect 36542 681592 36598 681601
rect 36542 681527 36598 681536
rect 34428 675504 34480 675510
rect 34428 675446 34480 675452
rect 32402 672752 32458 672761
rect 31024 672716 31076 672722
rect 32402 672687 32458 672696
rect 31024 672658 31076 672664
rect 36556 672110 36584 681527
rect 40696 675617 40724 681935
rect 41340 680762 41368 682246
rect 41340 680734 41552 680762
rect 41524 680354 41552 680734
rect 41786 680368 41842 680377
rect 41524 680326 41786 680354
rect 41786 680303 41842 680312
rect 41142 677104 41198 677113
rect 41142 677039 41198 677048
rect 40682 675608 40738 675617
rect 40682 675543 40738 675552
rect 39764 675504 39816 675510
rect 39764 675446 39816 675452
rect 36544 672104 36596 672110
rect 36544 672046 36596 672052
rect 39776 670993 39804 675446
rect 40408 672716 40460 672722
rect 40408 672658 40460 672664
rect 40420 671265 40448 672658
rect 41156 672489 41184 677039
rect 42062 676696 42118 676705
rect 42062 676631 42118 676640
rect 42076 676394 42104 676631
rect 42064 676388 42116 676394
rect 42064 676330 42116 676336
rect 42064 675640 42116 675646
rect 42062 675608 42064 675617
rect 42116 675608 42118 675617
rect 42062 675543 42118 675552
rect 41142 672480 41198 672489
rect 41142 672415 41198 672424
rect 42338 672480 42394 672489
rect 42338 672415 42394 672424
rect 41696 672104 41748 672110
rect 41748 672052 42288 672058
rect 41696 672046 42288 672052
rect 41708 672030 42288 672046
rect 40406 671256 40462 671265
rect 40406 671191 40462 671200
rect 39762 670984 39818 670993
rect 39762 670919 39818 670928
rect 42260 670290 42288 672030
rect 42076 670262 42288 670290
rect 42076 669868 42104 670262
rect 42352 668658 42380 672415
rect 42182 668630 42380 668658
rect 42536 668250 42564 683470
rect 42812 683398 42840 702406
rect 43088 684758 43116 728039
rect 43258 723616 43314 723625
rect 43258 723551 43314 723560
rect 43272 706586 43300 723551
rect 43442 719944 43498 719953
rect 43442 719879 43498 719888
rect 43456 719166 43484 719879
rect 43444 719160 43496 719166
rect 43444 719102 43496 719108
rect 43260 706580 43312 706586
rect 43260 706522 43312 706528
rect 43442 687712 43498 687721
rect 43442 687647 43498 687656
rect 43456 687410 43484 687647
rect 43444 687404 43496 687410
rect 43444 687346 43496 687352
rect 43076 684752 43128 684758
rect 43076 684694 43128 684700
rect 43074 684584 43130 684593
rect 43074 684519 43130 684528
rect 42800 683392 42852 683398
rect 42800 683334 42852 683340
rect 42892 683188 42944 683194
rect 42892 683130 42944 683136
rect 42708 675640 42760 675646
rect 42760 675588 42840 675594
rect 42708 675582 42840 675588
rect 42720 675566 42840 675582
rect 42352 668222 42564 668250
rect 42352 668046 42380 668222
rect 42168 667978 42196 668032
rect 42260 668018 42380 668046
rect 42260 667978 42288 668018
rect 42168 667950 42288 667978
rect 42614 667992 42670 668001
rect 42614 667927 42670 667936
rect 42154 667720 42210 667729
rect 42154 667655 42210 667664
rect 42168 667352 42196 667655
rect 42430 667448 42486 667457
rect 42430 667383 42486 667392
rect 42248 667140 42300 667146
rect 42248 667082 42300 667088
rect 42260 666482 42288 667082
rect 42260 666454 42380 666482
rect 42154 666360 42210 666369
rect 42154 666295 42210 666304
rect 42168 666165 42196 666295
rect 42352 664986 42380 666454
rect 42182 664958 42380 664986
rect 42248 664896 42300 664902
rect 42248 664838 42300 664844
rect 42260 664339 42288 664838
rect 42182 664311 42288 664339
rect 41970 664048 42026 664057
rect 41970 663983 42026 663992
rect 41984 663680 42012 663983
rect 42248 663536 42300 663542
rect 42248 663478 42300 663484
rect 42260 663150 42288 663478
rect 42182 663122 42288 663150
rect 42248 662856 42300 662862
rect 42062 662824 42118 662833
rect 42300 662804 42380 662810
rect 42248 662798 42380 662804
rect 42260 662782 42380 662798
rect 42062 662759 42118 662768
rect 42076 662674 42104 662759
rect 42076 662646 42288 662674
rect 42260 661042 42288 662646
rect 42168 661014 42288 661042
rect 42168 660620 42196 661014
rect 42352 660022 42380 662782
rect 42182 659994 42380 660022
rect 42444 659818 42472 667383
rect 42628 663626 42656 667927
rect 42812 666554 42840 675566
rect 42536 663598 42656 663626
rect 42720 666526 42840 666554
rect 42536 663354 42564 663598
rect 42720 663542 42748 666526
rect 42708 663536 42760 663542
rect 42708 663478 42760 663484
rect 42536 663326 42656 663354
rect 42628 659818 42656 663326
rect 42260 659790 42472 659818
rect 42536 659790 42656 659818
rect 42260 659654 42288 659790
rect 42536 659654 42564 659790
rect 42706 659696 42762 659705
rect 41984 659626 42288 659654
rect 42444 659626 42564 659654
rect 42628 659640 42706 659654
rect 42628 659631 42762 659640
rect 42628 659626 42748 659631
rect 41984 659357 42012 659626
rect 42168 658838 42380 658866
rect 42168 658784 42196 658838
rect 42352 658798 42380 658838
rect 42444 658798 42472 659626
rect 42352 658770 42472 658798
rect 42430 658608 42486 658617
rect 42430 658543 42486 658552
rect 42154 658336 42210 658345
rect 42210 658294 42380 658322
rect 42154 658271 42210 658280
rect 42156 657416 42208 657422
rect 42156 657358 42208 657364
rect 42168 656948 42196 657358
rect 42352 656350 42380 658294
rect 42182 656322 42380 656350
rect 42168 655710 42288 655738
rect 42168 655656 42196 655710
rect 42260 655670 42288 655710
rect 42444 655670 42472 658543
rect 42628 657422 42656 659626
rect 42616 657416 42668 657422
rect 42616 657358 42668 657364
rect 42260 655642 42472 655670
rect 38842 646096 38898 646105
rect 38842 646031 38898 646040
rect 8588 645524 8616 645660
rect 9048 645524 9076 645660
rect 9508 645524 9536 645660
rect 9968 645524 9996 645660
rect 10428 645524 10456 645660
rect 10888 645524 10916 645660
rect 11348 645524 11376 645660
rect 11808 645524 11836 645660
rect 12268 645524 12296 645660
rect 12728 645524 12756 645660
rect 13188 645524 13216 645660
rect 13648 645524 13676 645660
rect 14108 645524 14136 645660
rect 38856 644774 38884 646031
rect 41234 645688 41290 645697
rect 41234 645623 41290 645632
rect 35808 644768 35860 644774
rect 35530 644736 35586 644745
rect 35530 644671 35586 644680
rect 35806 644736 35808 644745
rect 38844 644768 38896 644774
rect 35860 644736 35862 644745
rect 38844 644710 38896 644716
rect 39670 644736 39726 644745
rect 35806 644671 35862 644680
rect 39670 644671 39726 644680
rect 35544 644502 35572 644671
rect 35532 644496 35584 644502
rect 35532 644438 35584 644444
rect 35346 643920 35402 643929
rect 35346 643855 35402 643864
rect 35360 643142 35388 643855
rect 35808 643544 35860 643550
rect 35530 643512 35586 643521
rect 35530 643447 35586 643456
rect 35806 643512 35808 643521
rect 35860 643512 35862 643521
rect 35806 643447 35862 643456
rect 35544 643278 35572 643447
rect 35532 643272 35584 643278
rect 35532 643214 35584 643220
rect 35348 643136 35400 643142
rect 35348 643078 35400 643084
rect 35438 642696 35494 642705
rect 35438 642631 35494 642640
rect 35452 641918 35480 642631
rect 35622 642288 35678 642297
rect 35622 642223 35678 642232
rect 39026 642288 39082 642297
rect 39026 642223 39028 642232
rect 35440 641912 35492 641918
rect 35440 641854 35492 641860
rect 35636 641782 35664 642223
rect 39080 642223 39082 642232
rect 39028 642194 39080 642200
rect 35808 642184 35860 642190
rect 35808 642126 35860 642132
rect 35820 641889 35848 642126
rect 39684 641986 39712 644671
rect 41248 644502 41276 645623
rect 41236 644496 41288 644502
rect 41236 644438 41288 644444
rect 40316 643544 40368 643550
rect 40316 643486 40368 643492
rect 39672 641980 39724 641986
rect 39672 641922 39724 641928
rect 35806 641880 35862 641889
rect 35806 641815 35862 641824
rect 35624 641776 35676 641782
rect 35624 641718 35676 641724
rect 39764 641776 39816 641782
rect 39764 641718 39816 641724
rect 39776 641481 39804 641718
rect 35346 641472 35402 641481
rect 35346 641407 35402 641416
rect 39762 641472 39818 641481
rect 39762 641407 39818 641416
rect 35360 640354 35388 641407
rect 40328 641073 40356 643486
rect 41708 643346 42104 643362
rect 41696 643340 42116 643346
rect 41748 643334 42064 643340
rect 41696 643282 41748 643288
rect 42064 643282 42116 643288
rect 41696 643136 41748 643142
rect 42064 643136 42116 643142
rect 41748 643084 42064 643090
rect 41696 643078 42116 643084
rect 41708 643062 42104 643078
rect 35530 641064 35586 641073
rect 35530 640999 35586 641008
rect 35806 641064 35862 641073
rect 35806 640999 35862 641008
rect 40314 641064 40370 641073
rect 40314 640999 40370 641008
rect 35544 640490 35572 640999
rect 35820 640762 35848 640999
rect 42904 640966 42932 683130
rect 43088 642297 43116 684519
rect 43258 680640 43314 680649
rect 43258 680575 43314 680584
rect 43272 662862 43300 680575
rect 43442 678328 43498 678337
rect 43442 678263 43498 678272
rect 43456 667146 43484 678263
rect 43640 667729 43668 767314
rect 43812 754928 43864 754934
rect 43812 754870 43864 754876
rect 43824 753001 43852 754870
rect 43810 752992 43866 753001
rect 43810 752927 43866 752936
rect 44284 727530 44312 770199
rect 44548 770092 44600 770098
rect 44548 770034 44600 770040
rect 44272 727524 44324 727530
rect 44272 727466 44324 727472
rect 44560 727326 44588 770034
rect 45008 765944 45060 765950
rect 45008 765886 45060 765892
rect 44822 760336 44878 760345
rect 44822 760271 44878 760280
rect 44548 727320 44600 727326
rect 44548 727262 44600 727268
rect 44362 722800 44418 722809
rect 44362 722735 44418 722744
rect 44376 707849 44404 722735
rect 44362 707840 44418 707849
rect 44362 707775 44418 707784
rect 43812 688696 43864 688702
rect 43812 688638 43864 688644
rect 43626 667720 43682 667729
rect 43626 667655 43682 667664
rect 43444 667140 43496 667146
rect 43444 667082 43496 667088
rect 43444 666596 43496 666602
rect 43444 666538 43496 666544
rect 43456 664902 43484 666538
rect 43444 664896 43496 664902
rect 43444 664838 43496 664844
rect 43260 662856 43312 662862
rect 43260 662798 43312 662804
rect 43444 662448 43496 662454
rect 43444 662390 43496 662396
rect 43074 642288 43130 642297
rect 43074 642223 43130 642232
rect 42064 640960 42116 640966
rect 42064 640902 42116 640908
rect 42892 640960 42944 640966
rect 42892 640902 42944 640908
rect 35808 640756 35860 640762
rect 35808 640698 35860 640704
rect 39856 640756 39908 640762
rect 39856 640698 39908 640704
rect 35532 640484 35584 640490
rect 35532 640426 35584 640432
rect 35348 640348 35400 640354
rect 35348 640290 35400 640296
rect 39868 640257 39896 640698
rect 42076 640642 42104 640902
rect 41708 640614 42104 640642
rect 41708 640490 41736 640614
rect 41696 640484 41748 640490
rect 41696 640426 41748 640432
rect 41696 640348 41748 640354
rect 42064 640348 42116 640354
rect 41748 640306 42064 640334
rect 41696 640290 41748 640296
rect 42064 640290 42116 640296
rect 43168 640348 43220 640354
rect 43168 640290 43220 640296
rect 39854 640248 39910 640257
rect 39854 640183 39910 640192
rect 42890 640248 42946 640257
rect 42890 640183 42946 640192
rect 34426 639840 34482 639849
rect 34426 639775 34482 639784
rect 33782 638616 33838 638625
rect 33782 638551 33838 638560
rect 32402 638208 32458 638217
rect 32402 638143 32458 638152
rect 32416 629950 32444 638143
rect 33796 630086 33824 638551
rect 34440 638246 34468 639775
rect 35530 639432 35586 639441
rect 35530 639367 35586 639376
rect 35806 639432 35862 639441
rect 35806 639367 35862 639376
rect 35544 638994 35572 639367
rect 35820 639130 35848 639367
rect 35808 639124 35860 639130
rect 35808 639066 35860 639072
rect 40224 639124 40276 639130
rect 40224 639066 40276 639072
rect 35532 638988 35584 638994
rect 35532 638930 35584 638936
rect 40040 638988 40092 638994
rect 40040 638930 40092 638936
rect 34428 638240 34480 638246
rect 34428 638182 34480 638188
rect 35532 637968 35584 637974
rect 35532 637910 35584 637916
rect 35544 637809 35572 637910
rect 35530 637800 35586 637809
rect 35530 637735 35586 637744
rect 35806 637800 35862 637809
rect 35806 637735 35808 637744
rect 35860 637735 35862 637744
rect 35808 637706 35860 637712
rect 40052 637401 40080 638930
rect 40038 637392 40094 637401
rect 40038 637327 40094 637336
rect 35806 636576 35862 636585
rect 35806 636511 35862 636520
rect 35820 636410 35848 636511
rect 35808 636404 35860 636410
rect 35808 636346 35860 636352
rect 40236 635361 40264 639066
rect 41696 638240 41748 638246
rect 41748 638188 42104 638194
rect 41696 638182 42104 638188
rect 41708 638178 42104 638182
rect 41708 638172 42116 638178
rect 41708 638166 42064 638172
rect 42064 638114 42116 638120
rect 42708 638172 42760 638178
rect 42708 638114 42760 638120
rect 41696 637968 41748 637974
rect 41748 637916 42104 637922
rect 41696 637910 42104 637916
rect 41708 637906 42104 637910
rect 41708 637900 42116 637906
rect 41708 637894 42064 637900
rect 42064 637842 42116 637848
rect 41510 637800 41566 637809
rect 41510 637735 41512 637744
rect 41564 637735 41566 637744
rect 41512 637706 41564 637712
rect 41328 636404 41380 636410
rect 41328 636346 41380 636352
rect 41340 636177 41368 636346
rect 41326 636168 41382 636177
rect 41326 636103 41382 636112
rect 35622 635352 35678 635361
rect 35622 635287 35678 635296
rect 40222 635352 40278 635361
rect 40222 635287 40278 635296
rect 35636 634846 35664 635287
rect 35808 635112 35860 635118
rect 35808 635054 35860 635060
rect 39764 635112 39816 635118
rect 39764 635054 39816 635060
rect 35820 634953 35848 635054
rect 39776 634953 39804 635054
rect 35806 634944 35862 634953
rect 35806 634879 35862 634888
rect 39762 634944 39818 634953
rect 39762 634879 39818 634888
rect 35624 634840 35676 634846
rect 35624 634782 35676 634788
rect 39304 634840 39356 634846
rect 39304 634782 39356 634788
rect 35622 634536 35678 634545
rect 35622 634471 35678 634480
rect 35636 633486 35664 634471
rect 35806 633720 35862 633729
rect 35806 633655 35808 633664
rect 35860 633655 35862 633664
rect 35808 633626 35860 633632
rect 35624 633480 35676 633486
rect 35624 633422 35676 633428
rect 39316 631417 39344 634782
rect 42338 633856 42394 633865
rect 42338 633791 42394 633800
rect 41708 633690 42104 633706
rect 41696 633684 42116 633690
rect 41748 633678 42064 633684
rect 41696 633626 41748 633632
rect 42064 633626 42116 633632
rect 41696 633480 41748 633486
rect 42064 633480 42116 633486
rect 41748 633428 42064 633434
rect 41696 633422 42116 633428
rect 41708 633406 42104 633422
rect 39302 631408 39358 631417
rect 39302 631343 39358 631352
rect 33784 630080 33836 630086
rect 33784 630022 33836 630028
rect 41696 630080 41748 630086
rect 41748 630028 42104 630034
rect 41696 630022 42104 630028
rect 41708 630018 42104 630022
rect 41708 630012 42116 630018
rect 41708 630006 42064 630012
rect 42064 629954 42116 629960
rect 32404 629944 32456 629950
rect 32404 629886 32456 629892
rect 41696 629944 41748 629950
rect 41748 629892 42288 629898
rect 41696 629886 42288 629892
rect 41708 629870 42288 629886
rect 42260 627178 42288 629870
rect 42168 627150 42288 627178
rect 42168 626620 42196 627150
rect 42352 627042 42380 633791
rect 42720 630674 42748 638114
rect 42260 627014 42380 627042
rect 42444 630646 42748 630674
rect 42904 630674 42932 640183
rect 42904 630646 43024 630674
rect 42260 625954 42288 627014
rect 42444 626770 42472 630646
rect 42708 630012 42760 630018
rect 42708 629954 42760 629960
rect 42720 626793 42748 629954
rect 42352 626742 42472 626770
rect 42706 626784 42762 626793
rect 42352 626090 42380 626742
rect 42706 626719 42762 626728
rect 42616 626544 42668 626550
rect 42616 626486 42668 626492
rect 42352 626062 42472 626090
rect 42260 625926 42380 625954
rect 42352 625682 42380 625926
rect 42168 625654 42380 625682
rect 42168 625464 42196 625654
rect 42168 624838 42288 624866
rect 42168 624784 42196 624838
rect 42260 624798 42288 624838
rect 42444 624798 42472 626062
rect 42260 624770 42472 624798
rect 42628 624186 42656 626486
rect 42182 624158 42656 624186
rect 42340 623416 42392 623422
rect 42154 623384 42210 623393
rect 42340 623358 42392 623364
rect 42154 623319 42210 623328
rect 42168 622948 42196 623319
rect 42352 622146 42380 623358
rect 42076 622118 42380 622146
rect 42076 621792 42104 622118
rect 42432 622056 42484 622062
rect 42432 621998 42484 622004
rect 41970 621480 42026 621489
rect 41970 621415 42026 621424
rect 41984 621112 42012 621415
rect 42444 620514 42472 621998
rect 42168 620378 42196 620500
rect 42260 620486 42472 620514
rect 42260 620378 42288 620486
rect 42168 620350 42288 620378
rect 41970 620256 42026 620265
rect 41970 620191 42026 620200
rect 41984 619956 42012 620191
rect 42246 619848 42302 619857
rect 42246 619783 42302 619792
rect 42260 617454 42288 619783
rect 42430 619032 42486 619041
rect 42430 618967 42486 618976
rect 42182 617426 42288 617454
rect 42444 616842 42472 618967
rect 42616 618928 42668 618934
rect 42168 616706 42196 616828
rect 42260 616814 42472 616842
rect 42536 618876 42616 618882
rect 42536 618870 42668 618876
rect 42536 618854 42656 618870
rect 42260 616706 42288 616814
rect 42168 616678 42288 616706
rect 42536 616434 42564 618854
rect 42706 618760 42762 618769
rect 42706 618695 42762 618704
rect 42168 616406 42564 616434
rect 42168 616148 42196 616406
rect 42246 616040 42302 616049
rect 42246 615975 42302 615984
rect 42260 615738 42288 615975
rect 42248 615732 42300 615738
rect 42248 615674 42300 615680
rect 42720 615618 42748 618695
rect 42182 615590 42748 615618
rect 42248 615528 42300 615534
rect 42248 615470 42300 615476
rect 42260 613782 42288 615470
rect 42182 613754 42288 613782
rect 42156 613624 42208 613630
rect 42156 613566 42208 613572
rect 42168 613121 42196 613566
rect 41786 612776 41842 612785
rect 41786 612711 41842 612720
rect 41800 612476 41828 612711
rect 8588 602276 8616 602412
rect 9048 602276 9076 602412
rect 9508 602276 9536 602412
rect 9968 602276 9996 602412
rect 10428 602276 10456 602412
rect 10888 602276 10916 602412
rect 11348 602276 11376 602412
rect 11808 602276 11836 602412
rect 12268 602276 12296 602412
rect 12728 602276 12756 602412
rect 13188 602276 13216 602412
rect 13648 602276 13676 602412
rect 14108 602276 14136 602412
rect 35806 601760 35862 601769
rect 41708 601730 42104 601746
rect 35806 601695 35808 601704
rect 35860 601695 35862 601704
rect 41696 601724 42116 601730
rect 35808 601666 35860 601672
rect 41748 601718 42064 601724
rect 41696 601666 41748 601672
rect 42064 601666 42116 601672
rect 42614 600944 42670 600953
rect 42614 600879 42670 600888
rect 42628 600438 42656 600879
rect 42616 600432 42668 600438
rect 42616 600374 42668 600380
rect 41326 599312 41382 599321
rect 41326 599247 41382 599256
rect 41340 599010 41368 599247
rect 41328 599004 41380 599010
rect 41328 598946 41380 598952
rect 41696 599004 41748 599010
rect 42064 599004 42116 599010
rect 41748 598964 42064 598992
rect 41696 598946 41748 598952
rect 42064 598946 42116 598952
rect 40866 598496 40922 598505
rect 40866 598431 40922 598440
rect 40880 597582 40908 598431
rect 41050 597850 41106 597859
rect 41050 597785 41106 597794
rect 41326 597850 41382 597859
rect 41326 597785 41382 597794
rect 41696 597848 41748 597854
rect 42064 597848 42116 597854
rect 41748 597808 42064 597836
rect 41696 597790 41748 597796
rect 42064 597790 42116 597796
rect 42800 597848 42852 597854
rect 42800 597790 42852 597796
rect 41064 597718 41092 597785
rect 41052 597712 41104 597718
rect 41052 597654 41104 597660
rect 41696 597712 41748 597718
rect 42064 597712 42116 597718
rect 41748 597672 42064 597700
rect 41696 597654 41748 597660
rect 42064 597654 42116 597660
rect 40868 597576 40920 597582
rect 40868 597518 40920 597524
rect 41696 597576 41748 597582
rect 42064 597576 42116 597582
rect 41748 597524 42064 597530
rect 41696 597518 42116 597524
rect 41708 597502 42104 597518
rect 41142 597272 41198 597281
rect 41142 597207 41198 597216
rect 41156 596086 41184 597207
rect 41326 596864 41382 596873
rect 41326 596799 41382 596808
rect 41340 596494 41368 596799
rect 41328 596488 41380 596494
rect 41328 596430 41380 596436
rect 41696 596488 41748 596494
rect 41748 596436 42104 596442
rect 41696 596430 42104 596436
rect 41708 596414 42104 596430
rect 41144 596080 41196 596086
rect 41604 596080 41656 596086
rect 41144 596022 41196 596028
rect 41326 596048 41382 596057
rect 41786 596048 41842 596057
rect 41656 596028 41786 596034
rect 41604 596022 41786 596028
rect 41616 596006 41786 596022
rect 41326 595983 41382 595992
rect 41786 595983 41842 595992
rect 33046 595640 33102 595649
rect 33046 595575 33102 595584
rect 31022 594416 31078 594425
rect 31022 594351 31078 594360
rect 31036 585750 31064 594351
rect 33060 587042 33088 595575
rect 35162 595232 35218 595241
rect 35162 595167 35218 595176
rect 34426 594824 34482 594833
rect 34426 594759 34482 594768
rect 34440 587217 34468 594759
rect 34426 587208 34482 587217
rect 34426 587143 34482 587152
rect 33048 587036 33100 587042
rect 33048 586978 33100 586984
rect 35176 585954 35204 595167
rect 41340 594794 41368 595983
rect 41328 594788 41380 594794
rect 41328 594730 41380 594736
rect 41696 594788 41748 594794
rect 41748 594748 42012 594776
rect 41696 594730 41748 594736
rect 41786 594008 41842 594017
rect 41616 593966 41786 593994
rect 36542 593600 36598 593609
rect 36542 593535 36598 593544
rect 35164 585948 35216 585954
rect 35164 585890 35216 585896
rect 31024 585744 31076 585750
rect 31024 585686 31076 585692
rect 36556 585206 36584 593535
rect 41616 593094 41644 593966
rect 41786 593943 41842 593952
rect 40592 593088 40644 593094
rect 40592 593030 40644 593036
rect 41604 593088 41656 593094
rect 41604 593030 41656 593036
rect 39946 590744 40002 590753
rect 39946 590679 40002 590688
rect 39960 585410 39988 590679
rect 40604 589393 40632 593030
rect 41786 592920 41842 592929
rect 41616 592878 41786 592906
rect 41616 592754 41644 592878
rect 41786 592855 41842 592864
rect 40776 592748 40828 592754
rect 40776 592690 40828 592696
rect 41604 592748 41656 592754
rect 41604 592690 41656 592696
rect 40788 589665 40816 592690
rect 41786 592376 41842 592385
rect 41786 592311 41842 592320
rect 40774 589656 40830 589665
rect 40774 589591 40830 589600
rect 41800 589529 41828 592311
rect 41786 589520 41842 589529
rect 41786 589455 41842 589464
rect 40590 589384 40646 589393
rect 40590 589319 40646 589328
rect 41984 589274 42012 594748
rect 42076 592034 42104 596414
rect 42812 592034 42840 597790
rect 42996 597718 43024 630646
rect 43180 598913 43208 640290
rect 43166 598904 43222 598913
rect 43166 598839 43222 598848
rect 42984 597712 43036 597718
rect 42984 597654 43036 597660
rect 43076 597576 43128 597582
rect 43076 597518 43128 597524
rect 42076 592006 42472 592034
rect 42812 592006 42932 592034
rect 41984 589246 42104 589274
rect 40132 587036 40184 587042
rect 40132 586978 40184 586984
rect 39948 585404 40000 585410
rect 39948 585346 40000 585352
rect 36544 585200 36596 585206
rect 36544 585142 36596 585148
rect 39396 585200 39448 585206
rect 39396 585142 39448 585148
rect 39408 584633 39436 585142
rect 40144 584905 40172 586978
rect 41604 585948 41656 585954
rect 41604 585890 41656 585896
rect 41616 585834 41644 585890
rect 41616 585806 41828 585834
rect 41604 585744 41656 585750
rect 41604 585686 41656 585692
rect 41420 585404 41472 585410
rect 41420 585346 41472 585352
rect 41432 584905 41460 585346
rect 40130 584896 40186 584905
rect 40130 584831 40186 584840
rect 41418 584896 41474 584905
rect 41418 584831 41474 584840
rect 41616 584633 41644 585686
rect 39394 584624 39450 584633
rect 39394 584559 39450 584568
rect 41602 584624 41658 584633
rect 41602 584559 41658 584568
rect 41800 584361 41828 585806
rect 42076 584458 42104 589246
rect 42064 584452 42116 584458
rect 42064 584394 42116 584400
rect 41786 584352 41842 584361
rect 41786 584287 41842 584296
rect 41786 583944 41842 583953
rect 41786 583879 41842 583888
rect 41800 583440 41828 583879
rect 41970 582584 42026 582593
rect 41970 582519 42026 582528
rect 41984 582249 42012 582519
rect 42444 581618 42472 592006
rect 42708 584452 42760 584458
rect 42708 584394 42760 584400
rect 42720 584338 42748 584394
rect 42720 584310 42840 584338
rect 42182 581590 42472 581618
rect 42154 581224 42210 581233
rect 42154 581159 42210 581168
rect 42168 580961 42196 581159
rect 42432 580644 42484 580650
rect 42432 580586 42484 580592
rect 41786 580272 41842 580281
rect 41786 580207 41842 580216
rect 41800 579768 41828 580207
rect 42246 580000 42302 580009
rect 42246 579935 42302 579944
rect 42260 578746 42288 579935
rect 42248 578740 42300 578746
rect 42248 578682 42300 578688
rect 42168 578598 42288 578626
rect 42168 578544 42196 578598
rect 42260 578558 42288 578598
rect 42444 578558 42472 580586
rect 42614 580544 42670 580553
rect 42614 580479 42670 580488
rect 42628 579614 42656 580479
rect 42812 579614 42840 584310
rect 42260 578530 42472 578558
rect 42536 579586 42656 579614
rect 42720 579586 42840 579614
rect 42248 578468 42300 578474
rect 42248 578410 42300 578416
rect 42062 578232 42118 578241
rect 42062 578167 42118 578176
rect 42076 577932 42104 578167
rect 42260 577295 42288 578410
rect 42182 577267 42288 577295
rect 42536 576994 42564 579586
rect 42168 576966 42564 576994
rect 42168 576708 42196 576966
rect 42338 576600 42394 576609
rect 42338 576535 42394 576544
rect 42062 575648 42118 575657
rect 42118 575606 42288 575634
rect 42062 575583 42118 575592
rect 41786 574696 41842 574705
rect 41786 574631 41842 574640
rect 41800 574260 41828 574631
rect 42260 573866 42288 575606
rect 42168 573838 42288 573866
rect 42168 573580 42196 573838
rect 42352 573458 42380 576535
rect 42720 574138 42748 579586
rect 42168 573430 42380 573458
rect 42444 574110 42748 574138
rect 42168 572968 42196 573430
rect 42444 572714 42472 574110
rect 42706 574016 42762 574025
rect 42706 573951 42762 573960
rect 42720 572714 42748 573951
rect 42260 572686 42472 572714
rect 42628 572686 42748 572714
rect 42168 572370 42196 572424
rect 42260 572370 42288 572686
rect 42168 572342 42288 572370
rect 42246 572248 42302 572257
rect 42246 572183 42302 572192
rect 42064 570988 42116 570994
rect 42064 570930 42116 570936
rect 42076 570588 42104 570930
rect 42260 569922 42288 572183
rect 42430 571976 42486 571985
rect 42430 571911 42486 571920
rect 42182 569894 42288 569922
rect 42444 569310 42472 571911
rect 42628 570994 42656 572686
rect 42616 570988 42668 570994
rect 42616 570930 42668 570936
rect 42168 569242 42196 569296
rect 42260 569282 42472 569310
rect 42260 569242 42288 569282
rect 42168 569214 42288 569242
rect 42904 563054 42932 592006
rect 43088 563054 43116 597518
rect 43258 593192 43314 593201
rect 43258 593127 43314 593136
rect 43272 578241 43300 593127
rect 43456 581233 43484 662390
rect 43824 645697 43852 688638
rect 44270 686488 44326 686497
rect 44270 686423 44326 686432
rect 43810 645688 43866 645697
rect 43810 645623 43866 645632
rect 44284 643346 44312 686423
rect 44456 684548 44508 684554
rect 44456 684490 44508 684496
rect 44468 644745 44496 684490
rect 44638 679960 44694 679969
rect 44638 679895 44694 679904
rect 44652 666369 44680 679895
rect 44638 666360 44694 666369
rect 44638 666295 44694 666304
rect 44454 644736 44510 644745
rect 44454 644671 44510 644680
rect 44272 643340 44324 643346
rect 44272 643282 44324 643288
rect 44270 641472 44326 641481
rect 44270 641407 44326 641416
rect 43628 637900 43680 637906
rect 43628 637842 43680 637848
rect 43640 618934 43668 637842
rect 43994 636168 44050 636177
rect 43994 636103 44050 636112
rect 43810 634944 43866 634953
rect 43810 634879 43866 634888
rect 43824 623830 43852 634879
rect 43812 623824 43864 623830
rect 43812 623766 43864 623772
rect 44008 623393 44036 636103
rect 43994 623384 44050 623393
rect 43994 623319 44050 623328
rect 43628 618928 43680 618934
rect 43628 618870 43680 618876
rect 43628 609272 43680 609278
rect 43628 609214 43680 609220
rect 43442 581224 43498 581233
rect 43442 581159 43498 581168
rect 43258 578232 43314 578241
rect 43258 578167 43314 578176
rect 43444 571396 43496 571402
rect 43444 571338 43496 571344
rect 42904 563026 43024 563054
rect 43088 563026 43208 563054
rect 8588 559164 8616 559300
rect 9048 559164 9076 559300
rect 9508 559164 9536 559300
rect 9968 559164 9996 559300
rect 10428 559164 10456 559300
rect 10888 559164 10916 559300
rect 11348 559164 11376 559300
rect 11808 559164 11836 559300
rect 12268 559164 12296 559300
rect 12728 559164 12756 559300
rect 13188 559164 13216 559300
rect 13648 559164 13676 559300
rect 14108 559164 14136 559300
rect 41708 557802 42104 557818
rect 41696 557796 42116 557802
rect 41748 557790 42064 557796
rect 41696 557738 41748 557744
rect 42064 557738 42116 557744
rect 41328 557728 41380 557734
rect 41326 557696 41328 557705
rect 41380 557696 41382 557705
rect 41326 557631 41382 557640
rect 40590 556064 40646 556073
rect 40590 555999 40646 556008
rect 40604 554810 40632 555999
rect 41142 555656 41198 555665
rect 41142 555591 41198 555600
rect 41156 555354 41184 555591
rect 42064 555416 42116 555422
rect 41708 555364 42064 555370
rect 41708 555358 42116 555364
rect 41144 555348 41196 555354
rect 41144 555290 41196 555296
rect 41708 555342 42104 555358
rect 41708 555150 41736 555342
rect 42798 555248 42854 555257
rect 42798 555183 42854 555192
rect 41696 555144 41748 555150
rect 41050 555078 41106 555087
rect 41696 555086 41748 555092
rect 41050 555013 41106 555022
rect 41064 554946 41092 555013
rect 41052 554940 41104 554946
rect 41052 554882 41104 554888
rect 41696 554940 41748 554946
rect 42064 554940 42116 554946
rect 41748 554900 42064 554928
rect 41696 554882 41748 554888
rect 42064 554882 42116 554888
rect 41708 554810 42104 554826
rect 40592 554804 40644 554810
rect 40592 554746 40644 554752
rect 41696 554804 42116 554810
rect 41748 554798 42064 554804
rect 41696 554746 41748 554752
rect 42064 554746 42116 554752
rect 40038 553408 40094 553417
rect 40038 553343 40094 553352
rect 40958 553408 41014 553417
rect 40958 553343 41014 553352
rect 29642 551984 29698 551993
rect 29642 551919 29698 551928
rect 29656 544406 29684 551919
rect 40052 550458 40080 553343
rect 40040 550452 40092 550458
rect 40040 550394 40092 550400
rect 40972 548026 41000 553343
rect 42812 550634 42840 555183
rect 42996 554946 43024 563026
rect 43180 555422 43208 563026
rect 43456 558113 43484 571338
rect 43442 558104 43498 558113
rect 43442 558039 43498 558048
rect 43168 555416 43220 555422
rect 43168 555358 43220 555364
rect 42984 554940 43036 554946
rect 42984 554882 43036 554888
rect 43166 554432 43222 554441
rect 43166 554367 43222 554376
rect 42812 550606 42932 550634
rect 41708 550458 42104 550474
rect 41696 550452 42116 550458
rect 41748 550446 42064 550452
rect 41696 550394 41748 550400
rect 42064 550394 42116 550400
rect 42524 550452 42576 550458
rect 42524 550394 42576 550400
rect 41878 549944 41934 549953
rect 41878 549879 41934 549888
rect 40972 547998 41184 548026
rect 31758 547496 31814 547505
rect 31758 547431 31760 547440
rect 31812 547431 31814 547440
rect 38568 547460 38620 547466
rect 31760 547402 31812 547408
rect 38568 547402 38620 547408
rect 29644 544400 29696 544406
rect 29644 544342 29696 544348
rect 38580 542366 38608 547402
rect 41156 547346 41184 547998
rect 41156 547318 41368 547346
rect 41340 546417 41368 547318
rect 41326 546408 41382 546417
rect 41326 546343 41382 546352
rect 41892 545601 41920 549879
rect 42062 549536 42118 549545
rect 42062 549471 42118 549480
rect 41878 545592 41934 545601
rect 41878 545527 41934 545536
rect 42076 545329 42104 549471
rect 42338 548312 42394 548321
rect 42338 548247 42394 548256
rect 42352 547942 42380 548247
rect 42340 547936 42392 547942
rect 42340 547878 42392 547884
rect 42062 545320 42118 545329
rect 42062 545255 42118 545264
rect 41512 544400 41564 544406
rect 41512 544342 41564 544348
rect 38568 542360 38620 542366
rect 38568 542302 38620 542308
rect 41524 542042 41552 544342
rect 41696 542360 41748 542366
rect 41696 542302 41748 542308
rect 41708 542178 41736 542302
rect 41708 542150 42380 542178
rect 41524 542014 42288 542042
rect 42260 540682 42288 542014
rect 42168 540654 42288 540682
rect 42168 540260 42196 540654
rect 42352 539050 42380 542150
rect 42182 539022 42380 539050
rect 42536 538438 42564 550394
rect 42706 549128 42762 549137
rect 42706 549063 42762 549072
rect 42720 540974 42748 549063
rect 42720 540946 42840 540974
rect 42168 538370 42196 538424
rect 42260 538410 42564 538438
rect 42260 538370 42288 538410
rect 42168 538342 42288 538370
rect 42246 538248 42302 538257
rect 42246 538183 42302 538192
rect 42260 538098 42288 538183
rect 42260 538070 42380 538098
rect 42062 537976 42118 537985
rect 42062 537911 42118 537920
rect 42076 537744 42104 537911
rect 42352 537758 42380 538070
rect 42260 537730 42380 537758
rect 42168 536466 42196 536588
rect 42260 536466 42288 537730
rect 42430 537024 42486 537033
rect 42430 536959 42486 536968
rect 42168 536438 42288 536466
rect 42248 536308 42300 536314
rect 42248 536250 42300 536256
rect 42260 535378 42288 536250
rect 42182 535350 42288 535378
rect 42444 534766 42472 536959
rect 42812 536874 42840 540946
rect 42168 534698 42196 534752
rect 42260 534738 42472 534766
rect 42536 536846 42840 536874
rect 42260 534698 42288 534738
rect 42168 534670 42288 534698
rect 42536 534290 42564 536846
rect 42260 534262 42564 534290
rect 42260 534086 42288 534262
rect 42432 534200 42484 534206
rect 42432 534142 42484 534148
rect 42182 534058 42288 534086
rect 42444 533542 42472 534142
rect 42616 533996 42668 534002
rect 42616 533938 42668 533944
rect 42182 533514 42472 533542
rect 42246 533352 42302 533361
rect 42246 533287 42302 533296
rect 42260 531059 42288 533287
rect 42430 532672 42486 532681
rect 42430 532607 42486 532616
rect 42182 531031 42288 531059
rect 42248 530936 42300 530942
rect 42248 530878 42300 530884
rect 42260 530414 42288 530878
rect 42182 530386 42288 530414
rect 42248 530324 42300 530330
rect 42248 530266 42300 530272
rect 42260 529771 42288 530266
rect 42182 529743 42288 529771
rect 42444 529219 42472 532607
rect 42628 530942 42656 533938
rect 42616 530936 42668 530942
rect 42616 530878 42668 530884
rect 42616 530800 42668 530806
rect 42616 530742 42668 530748
rect 42628 530330 42656 530742
rect 42616 530324 42668 530330
rect 42616 530266 42668 530272
rect 42614 529816 42670 529825
rect 42614 529751 42670 529760
rect 42182 529191 42472 529219
rect 42432 529100 42484 529106
rect 42432 529042 42484 529048
rect 41786 527640 41842 527649
rect 41786 527575 41842 527584
rect 41800 527340 41828 527575
rect 42444 526742 42472 529042
rect 42628 528554 42656 529751
rect 42182 526714 42472 526742
rect 42536 528526 42656 528554
rect 42536 526091 42564 528526
rect 42182 526063 42564 526091
rect 42524 523728 42576 523734
rect 42524 523670 42576 523676
rect 42536 522753 42564 523670
rect 40682 522744 40738 522753
rect 40682 522679 40738 522688
rect 42522 522744 42578 522753
rect 42522 522679 42578 522688
rect 8588 431596 8616 431664
rect 9048 431596 9076 431664
rect 9508 431596 9536 431664
rect 9968 431596 9996 431664
rect 10428 431596 10456 431664
rect 10888 431596 10916 431664
rect 11348 431596 11376 431664
rect 11808 431596 11836 431664
rect 12268 431596 12296 431664
rect 12728 431596 12756 431664
rect 13188 431596 13216 431664
rect 13648 431596 13676 431664
rect 14108 431596 14136 431664
rect 40696 431225 40724 522679
rect 42064 518968 42116 518974
rect 42064 518910 42116 518916
rect 42076 437474 42104 518910
rect 41708 437446 42104 437474
rect 40682 431216 40738 431225
rect 40682 431151 40738 431160
rect 41326 430536 41382 430545
rect 41326 430471 41382 430480
rect 41142 430128 41198 430137
rect 41142 430063 41198 430072
rect 40958 429482 41014 429491
rect 41156 429486 41184 430063
rect 41340 429622 41368 430471
rect 41708 429622 41736 437446
rect 42904 431225 42932 550606
rect 42890 431216 42946 431225
rect 42890 431151 42946 431160
rect 41328 429616 41380 429622
rect 41328 429558 41380 429564
rect 41696 429616 41748 429622
rect 41696 429558 41748 429564
rect 40958 429417 41014 429426
rect 41144 429480 41196 429486
rect 41144 429422 41196 429428
rect 41326 429482 41382 429491
rect 41326 429417 41382 429426
rect 41696 429480 41748 429486
rect 42064 429480 42116 429486
rect 41748 429440 42064 429468
rect 41696 429422 41748 429428
rect 42064 429422 42116 429428
rect 40972 429214 41000 429417
rect 41340 429350 41368 429417
rect 41328 429344 41380 429350
rect 41328 429286 41380 429292
rect 41696 429344 41748 429350
rect 42064 429344 42116 429350
rect 41748 429304 42064 429332
rect 41696 429286 41748 429292
rect 42064 429286 42116 429292
rect 40960 429208 41012 429214
rect 40960 429150 41012 429156
rect 41696 429208 41748 429214
rect 42064 429208 42116 429214
rect 41748 429168 42064 429196
rect 41696 429150 41748 429156
rect 42064 429150 42116 429156
rect 42982 428224 43038 428233
rect 42982 428159 43038 428168
rect 41142 427680 41198 427689
rect 41142 427615 41198 427624
rect 41156 426494 41184 427615
rect 41144 426488 41196 426494
rect 41144 426430 41196 426436
rect 41696 426488 41748 426494
rect 42064 426488 42116 426494
rect 41748 426448 42064 426476
rect 41696 426430 41748 426436
rect 42064 426430 42116 426436
rect 41142 426048 41198 426057
rect 41142 425983 41198 425992
rect 40774 425232 40830 425241
rect 40774 425167 40830 425176
rect 40788 418441 40816 425167
rect 40774 418432 40830 418441
rect 40774 418367 40830 418376
rect 41156 418033 41184 425983
rect 41970 424416 42026 424425
rect 41970 424351 42026 424360
rect 41142 418024 41198 418033
rect 41142 417959 41198 417968
rect 41984 415394 42012 424351
rect 42798 423192 42854 423201
rect 42798 423127 42854 423136
rect 42246 419928 42302 419937
rect 42246 419863 42302 419872
rect 42260 417874 42288 419863
rect 42614 419520 42670 419529
rect 42614 419455 42670 419464
rect 42628 418198 42656 419455
rect 42616 418192 42668 418198
rect 42616 418134 42668 418140
rect 42430 418024 42486 418033
rect 42430 417959 42486 417968
rect 42260 417846 42380 417874
rect 42352 415394 42380 417846
rect 41984 415366 42104 415394
rect 42076 414338 42104 415366
rect 42260 415366 42380 415394
rect 42260 414610 42288 415366
rect 42260 414582 42380 414610
rect 42076 414310 42288 414338
rect 42260 413114 42288 414310
rect 42168 413086 42288 413114
rect 42168 412624 42196 413086
rect 42352 411618 42380 414582
rect 42260 411590 42380 411618
rect 42168 411346 42196 411468
rect 42260 411346 42288 411590
rect 42168 411318 42288 411346
rect 42168 410910 42288 410938
rect 42168 410788 42196 410910
rect 42260 410802 42288 410910
rect 42444 410802 42472 417959
rect 42260 410774 42472 410802
rect 42182 410162 42472 410190
rect 42248 409828 42300 409834
rect 42248 409770 42300 409776
rect 42260 408966 42288 409770
rect 42182 408938 42288 408966
rect 42444 408474 42472 410162
rect 42432 408468 42484 408474
rect 42432 408410 42484 408416
rect 42432 408332 42484 408338
rect 42432 408274 42484 408280
rect 42444 407810 42472 408274
rect 42168 407674 42196 407796
rect 42260 407782 42472 407810
rect 42260 407674 42288 407782
rect 42168 407646 42288 407674
rect 41786 407552 41842 407561
rect 41786 407487 41842 407496
rect 41800 407116 41828 407487
rect 42432 407108 42484 407114
rect 42432 407050 42484 407056
rect 42444 406518 42472 407050
rect 42168 406450 42196 406504
rect 42260 406490 42472 406518
rect 42260 406450 42288 406490
rect 42168 406422 42288 406450
rect 42182 405915 42472 405943
rect 42444 404190 42472 405915
rect 42432 404184 42484 404190
rect 42432 404126 42484 404132
rect 41786 403880 41842 403889
rect 41786 403815 41842 403824
rect 41800 403444 41828 403815
rect 42812 402974 42840 423127
rect 42996 408494 43024 428159
rect 43180 427281 43208 554367
rect 43442 547088 43498 547097
rect 43442 547023 43498 547032
rect 43456 546650 43484 547023
rect 43444 546644 43496 546650
rect 43444 546586 43496 546592
rect 43444 545148 43496 545154
rect 43444 545090 43496 545096
rect 43456 429486 43484 545090
rect 43640 537985 43668 609214
rect 44086 600128 44142 600137
rect 44086 600063 44142 600072
rect 44100 598934 44128 600063
rect 44284 599729 44312 641407
rect 44638 641064 44694 641073
rect 44638 640999 44694 641008
rect 44454 637800 44510 637809
rect 44454 637735 44510 637744
rect 44468 613630 44496 637735
rect 44456 613624 44508 613630
rect 44456 613566 44508 613572
rect 44652 600545 44680 640999
rect 44638 600536 44694 600545
rect 44638 600471 44694 600480
rect 44270 599720 44326 599729
rect 44270 599655 44326 599664
rect 44456 599004 44508 599010
rect 44456 598946 44508 598952
rect 44100 598906 44220 598934
rect 43810 591560 43866 591569
rect 43810 591495 43866 591504
rect 43824 590714 43852 591495
rect 43812 590708 43864 590714
rect 43812 590650 43864 590656
rect 43810 558512 43866 558521
rect 43810 558447 43866 558456
rect 43824 557598 43852 558447
rect 43812 557592 43864 557598
rect 43812 557534 43864 557540
rect 44192 557297 44220 598906
rect 44178 557288 44234 557297
rect 44178 557223 44234 557232
rect 44468 556481 44496 598946
rect 44638 591968 44694 591977
rect 44638 591903 44694 591912
rect 44652 580650 44680 591903
rect 44640 580644 44692 580650
rect 44640 580586 44692 580592
rect 44638 556880 44694 556889
rect 44638 556815 44694 556824
rect 44454 556472 44510 556481
rect 44454 556407 44510 556416
rect 44272 554804 44324 554810
rect 44272 554746 44324 554752
rect 43810 551576 43866 551585
rect 43810 551511 43866 551520
rect 43626 537976 43682 537985
rect 43626 537911 43682 537920
rect 43824 529106 43852 551511
rect 43994 550760 44050 550769
rect 43994 550695 44050 550704
rect 44008 534002 44036 550695
rect 43996 533996 44048 534002
rect 43996 533938 44048 533944
rect 43812 529100 43864 529106
rect 43812 529042 43864 529048
rect 43628 491972 43680 491978
rect 43628 491914 43680 491920
rect 43444 429480 43496 429486
rect 43444 429422 43496 429428
rect 43166 427272 43222 427281
rect 43166 427207 43222 427216
rect 43350 423600 43406 423609
rect 43350 423535 43406 423544
rect 43166 422784 43222 422793
rect 43166 422719 43222 422728
rect 43180 409834 43208 422719
rect 43168 409828 43220 409834
rect 43168 409770 43220 409776
rect 42536 402946 42840 402974
rect 42904 408466 43024 408494
rect 42536 402815 42564 402946
rect 42182 402787 42564 402815
rect 42432 402552 42484 402558
rect 42432 402494 42484 402500
rect 42444 402166 42472 402494
rect 42182 402138 42472 402166
rect 41786 401976 41842 401985
rect 41786 401911 41842 401920
rect 41800 401608 41828 401911
rect 41786 400072 41842 400081
rect 41786 400007 41842 400016
rect 41800 399772 41828 400007
rect 42182 399107 42472 399135
rect 41786 398848 41842 398857
rect 41786 398783 41842 398792
rect 41800 398480 41828 398783
rect 42444 397458 42472 399107
rect 42432 397452 42484 397458
rect 42432 397394 42484 397400
rect 8588 388348 8616 388484
rect 9048 388348 9076 388484
rect 9508 388348 9536 388484
rect 9968 388348 9996 388484
rect 10428 388348 10456 388484
rect 10888 388348 10916 388484
rect 11348 388348 11376 388484
rect 11808 388348 11836 388484
rect 12268 388348 12296 388484
rect 12728 388348 12756 388484
rect 13188 388348 13216 388484
rect 13648 388348 13676 388484
rect 14108 388348 14136 388484
rect 35346 387560 35402 387569
rect 39946 387560 40002 387569
rect 35346 387495 35402 387504
rect 35808 387524 35860 387530
rect 35360 386578 35388 387495
rect 39946 387495 39948 387504
rect 35808 387466 35860 387472
rect 40000 387495 40002 387504
rect 39948 387466 40000 387472
rect 35820 387161 35848 387466
rect 35530 387152 35586 387161
rect 35530 387087 35586 387096
rect 35806 387152 35862 387161
rect 35806 387087 35862 387096
rect 40130 387152 40186 387161
rect 40130 387087 40186 387096
rect 35348 386572 35400 386578
rect 35348 386514 35400 386520
rect 35544 386442 35572 387087
rect 40144 386850 40172 387087
rect 35808 386844 35860 386850
rect 35808 386786 35860 386792
rect 40132 386844 40184 386850
rect 40132 386786 40184 386792
rect 35532 386436 35584 386442
rect 35532 386378 35584 386384
rect 35820 386345 35848 386786
rect 40314 386744 40370 386753
rect 40314 386679 40370 386688
rect 40328 386578 40356 386679
rect 40316 386572 40368 386578
rect 40316 386514 40368 386520
rect 42064 386504 42116 386510
rect 41708 386452 42064 386458
rect 41708 386446 42116 386452
rect 41708 386442 42104 386446
rect 41696 386436 42104 386442
rect 41748 386430 42104 386436
rect 41696 386378 41748 386384
rect 35806 386336 35862 386345
rect 35806 386271 35862 386280
rect 35346 385928 35402 385937
rect 35346 385863 35402 385872
rect 35360 385082 35388 385863
rect 35530 385520 35586 385529
rect 35530 385455 35586 385464
rect 35806 385520 35862 385529
rect 35806 385455 35808 385464
rect 35544 385218 35572 385455
rect 35860 385455 35862 385464
rect 39580 385484 39632 385490
rect 35808 385426 35860 385432
rect 39580 385426 39632 385432
rect 35532 385212 35584 385218
rect 35532 385154 35584 385160
rect 39592 385121 39620 385426
rect 42904 385286 42932 408466
rect 43364 402558 43392 423535
rect 43352 402552 43404 402558
rect 43352 402494 43404 402500
rect 43640 387569 43668 491914
rect 43812 434036 43864 434042
rect 43812 433978 43864 433984
rect 43626 387560 43682 387569
rect 43626 387495 43682 387504
rect 41696 385280 41748 385286
rect 42064 385280 42116 385286
rect 41748 385228 42064 385234
rect 41696 385222 42116 385228
rect 42892 385280 42944 385286
rect 42892 385222 42944 385228
rect 41708 385206 42104 385222
rect 39578 385112 39634 385121
rect 35348 385076 35400 385082
rect 43074 385112 43130 385121
rect 41708 385082 42104 385098
rect 39578 385047 39634 385056
rect 41696 385076 42116 385082
rect 35348 385018 35400 385024
rect 41748 385070 42064 385076
rect 41696 385018 41748 385024
rect 43074 385047 43130 385056
rect 43260 385076 43312 385082
rect 42064 385018 42116 385024
rect 35622 384704 35678 384713
rect 35622 384639 35678 384648
rect 35636 383858 35664 384639
rect 35806 384296 35862 384305
rect 35806 384231 35862 384240
rect 35820 384130 35848 384231
rect 35808 384124 35860 384130
rect 35808 384066 35860 384072
rect 39672 384124 39724 384130
rect 39672 384066 39724 384072
rect 39684 383897 39712 384066
rect 42064 383920 42116 383926
rect 35806 383888 35862 383897
rect 35624 383852 35676 383858
rect 35806 383823 35862 383832
rect 39670 383888 39726 383897
rect 41708 383868 42064 383874
rect 41708 383862 42116 383868
rect 41708 383858 42104 383862
rect 39670 383823 39726 383832
rect 41696 383852 42104 383858
rect 35624 383794 35676 383800
rect 35820 383722 35848 383823
rect 41748 383846 42104 383852
rect 41696 383794 41748 383800
rect 41708 383722 42104 383738
rect 35808 383716 35860 383722
rect 35808 383658 35860 383664
rect 41696 383716 42116 383722
rect 41748 383710 42064 383716
rect 41696 383658 41748 383664
rect 42064 383658 42116 383664
rect 35346 383480 35402 383489
rect 35346 383415 35402 383424
rect 35360 382294 35388 383415
rect 35530 383072 35586 383081
rect 35530 383007 35586 383016
rect 35806 383072 35862 383081
rect 35806 383007 35862 383016
rect 35544 382702 35572 383007
rect 35532 382696 35584 382702
rect 35532 382638 35584 382644
rect 35820 382566 35848 383007
rect 40040 382696 40092 382702
rect 40040 382638 40092 382644
rect 35808 382560 35860 382566
rect 35808 382502 35860 382508
rect 35808 382424 35860 382430
rect 35808 382366 35860 382372
rect 35348 382288 35400 382294
rect 35820 382265 35848 382366
rect 40052 382265 40080 382638
rect 41696 382560 41748 382566
rect 41696 382502 41748 382508
rect 40224 382424 40276 382430
rect 40224 382366 40276 382372
rect 35348 382230 35400 382236
rect 35806 382256 35862 382265
rect 35806 382191 35862 382200
rect 40038 382256 40094 382265
rect 40038 382191 40094 382200
rect 35622 381848 35678 381857
rect 35622 381783 35678 381792
rect 32402 381440 32458 381449
rect 32402 381375 32458 381384
rect 28814 376544 28870 376553
rect 28814 376479 28870 376488
rect 28828 375902 28856 376479
rect 28816 375896 28868 375902
rect 28816 375838 28868 375844
rect 32416 371890 32444 381375
rect 35636 381070 35664 381783
rect 35806 381440 35862 381449
rect 35806 381375 35862 381384
rect 35624 381064 35676 381070
rect 35624 381006 35676 381012
rect 35820 380934 35848 381375
rect 40040 381064 40092 381070
rect 40040 381006 40092 381012
rect 35808 380928 35860 380934
rect 35808 380870 35860 380876
rect 39856 380928 39908 380934
rect 39856 380870 39908 380876
rect 39868 380633 39896 380870
rect 35622 380624 35678 380633
rect 35622 380559 35678 380568
rect 39854 380624 39910 380633
rect 39854 380559 39910 380568
rect 35438 380216 35494 380225
rect 35438 380151 35494 380160
rect 35452 379574 35480 380151
rect 35636 379982 35664 380559
rect 40052 380225 40080 381006
rect 35806 380216 35862 380225
rect 35806 380151 35862 380160
rect 40038 380216 40094 380225
rect 40038 380151 40094 380160
rect 35624 379976 35676 379982
rect 35624 379918 35676 379924
rect 35820 379710 35848 380151
rect 35808 379704 35860 379710
rect 35808 379646 35860 379652
rect 39764 379704 39816 379710
rect 39764 379646 39816 379652
rect 35440 379568 35492 379574
rect 35440 379510 35492 379516
rect 35806 378992 35862 379001
rect 35806 378927 35862 378936
rect 35820 378350 35848 378927
rect 35808 378344 35860 378350
rect 35808 378286 35860 378292
rect 39580 378344 39632 378350
rect 39580 378286 39632 378292
rect 35622 377768 35678 377777
rect 35622 377703 35678 377712
rect 35636 377058 35664 377703
rect 39592 377369 39620 378286
rect 39776 377777 39804 379646
rect 40236 379001 40264 382366
rect 41420 382288 41472 382294
rect 41420 382230 41472 382236
rect 41432 381857 41460 382230
rect 41418 381848 41474 381857
rect 41418 381783 41474 381792
rect 41052 379976 41104 379982
rect 41052 379918 41104 379924
rect 41064 379817 41092 379918
rect 41050 379808 41106 379817
rect 41050 379743 41106 379752
rect 41512 379568 41564 379574
rect 41512 379510 41564 379516
rect 41708 379514 41736 382502
rect 42798 380624 42854 380633
rect 42798 380559 42854 380568
rect 40222 378992 40278 379001
rect 40222 378927 40278 378936
rect 41524 378185 41552 379510
rect 41708 379486 42472 379514
rect 41510 378176 41566 378185
rect 41510 378111 41566 378120
rect 39762 377768 39818 377777
rect 39762 377703 39818 377712
rect 35806 377360 35862 377369
rect 35806 377295 35862 377304
rect 39578 377360 39634 377369
rect 39578 377295 39634 377304
rect 35624 377052 35676 377058
rect 35624 376994 35676 377000
rect 35820 376786 35848 377295
rect 41512 376984 41564 376990
rect 41510 376952 41512 376961
rect 41564 376952 41566 376961
rect 41510 376887 41566 376896
rect 42064 376848 42116 376854
rect 41708 376796 42064 376802
rect 41708 376790 42116 376796
rect 41708 376786 42104 376790
rect 35808 376780 35860 376786
rect 35808 376722 35860 376728
rect 41696 376780 42104 376786
rect 41748 376774 42104 376780
rect 41696 376722 41748 376728
rect 35806 376136 35862 376145
rect 35806 376071 35862 376080
rect 33784 375896 33836 375902
rect 33784 375838 33836 375844
rect 33796 373318 33824 375838
rect 35820 375630 35848 376071
rect 35808 375624 35860 375630
rect 35808 375566 35860 375572
rect 41696 375624 41748 375630
rect 41748 375572 42104 375578
rect 41696 375566 42104 375572
rect 41708 375562 42104 375566
rect 41708 375556 42116 375562
rect 41708 375550 42064 375556
rect 42064 375498 42116 375504
rect 33784 373312 33836 373318
rect 33784 373254 33836 373260
rect 41696 373312 41748 373318
rect 41696 373254 41748 373260
rect 41708 372858 41736 373254
rect 41708 372830 42288 372858
rect 32404 371884 32456 371890
rect 32404 371826 32456 371832
rect 41696 371884 41748 371890
rect 41696 371826 41748 371832
rect 41708 371770 41736 371826
rect 41708 371754 42104 371770
rect 41708 371748 42116 371754
rect 41708 371742 42064 371748
rect 42064 371690 42116 371696
rect 42062 369744 42118 369753
rect 42062 369679 42118 369688
rect 42076 369444 42104 369679
rect 42260 368263 42288 372830
rect 42182 368235 42288 368263
rect 42444 367622 42472 379486
rect 42616 371748 42668 371754
rect 42616 371690 42668 371696
rect 42628 369854 42656 371690
rect 42182 367594 42472 367622
rect 42536 369826 42656 369854
rect 42182 366947 42288 366975
rect 41800 365673 41828 365772
rect 41786 365664 41842 365673
rect 41786 365599 41842 365608
rect 42062 364984 42118 364993
rect 42062 364919 42118 364928
rect 42076 364548 42104 364919
rect 42260 364342 42288 366947
rect 42248 364336 42300 364342
rect 42248 364278 42300 364284
rect 42340 364132 42392 364138
rect 42340 364074 42392 364080
rect 42352 363950 42380 364074
rect 42182 363922 42380 363950
rect 41786 363760 41842 363769
rect 41786 363695 41842 363704
rect 41800 363256 41828 363695
rect 42168 362766 42288 362794
rect 42168 362712 42196 362766
rect 42260 362726 42288 362766
rect 42536 362726 42564 369826
rect 42812 369753 42840 380559
rect 43088 369854 43116 385047
rect 43260 385018 43312 385024
rect 42996 369826 43116 369854
rect 42798 369744 42854 369753
rect 42798 369679 42854 369688
rect 42260 362698 42564 362726
rect 41786 360632 41842 360641
rect 41786 360567 41842 360576
rect 41800 360264 41828 360567
rect 42432 360188 42484 360194
rect 42432 360130 42484 360136
rect 42156 359984 42208 359990
rect 42156 359926 42208 359932
rect 42168 359584 42196 359926
rect 42444 358986 42472 360130
rect 42182 358958 42472 358986
rect 41878 358728 41934 358737
rect 41878 358663 41934 358672
rect 41892 358428 41920 358663
rect 41786 356960 41842 356969
rect 41786 356895 41842 356904
rect 41800 356592 41828 356895
rect 42432 356040 42484 356046
rect 42432 355982 42484 355988
rect 42444 355926 42472 355982
rect 42182 355898 42472 355926
rect 41970 355736 42026 355745
rect 41970 355671 42026 355680
rect 41984 355300 42012 355671
rect 40406 345808 40462 345817
rect 40406 345743 40462 345752
rect 8588 345100 8616 345236
rect 9048 345100 9076 345236
rect 9508 345100 9536 345236
rect 9968 345100 9996 345236
rect 10428 345100 10456 345236
rect 10888 345100 10916 345236
rect 11348 345100 11376 345236
rect 11808 345100 11836 345236
rect 12268 345100 12296 345236
rect 12728 345100 12756 345236
rect 13188 345100 13216 345236
rect 13648 345100 13676 345236
rect 14108 345100 14136 345236
rect 39762 344992 39818 345001
rect 39762 344927 39818 344936
rect 39578 344720 39634 344729
rect 39578 344655 39634 344664
rect 35346 344312 35402 344321
rect 35346 344247 35402 344256
rect 35622 344312 35678 344321
rect 35622 344247 35678 344256
rect 35360 343670 35388 344247
rect 35636 343806 35664 344247
rect 39592 344078 39620 344655
rect 35808 344072 35860 344078
rect 35808 344014 35860 344020
rect 39580 344072 39632 344078
rect 39580 344014 39632 344020
rect 35820 343913 35848 344014
rect 35806 343904 35862 343913
rect 35806 343839 35862 343848
rect 35624 343800 35676 343806
rect 35624 343742 35676 343748
rect 35348 343664 35400 343670
rect 35348 343606 35400 343612
rect 39578 343496 39634 343505
rect 39578 343431 39634 343440
rect 35346 343088 35402 343097
rect 35346 343023 35402 343032
rect 35360 342446 35388 343023
rect 35808 342712 35860 342718
rect 35530 342680 35586 342689
rect 35530 342615 35586 342624
rect 35806 342680 35808 342689
rect 35860 342680 35862 342689
rect 35806 342615 35862 342624
rect 35348 342440 35400 342446
rect 35348 342382 35400 342388
rect 35544 342310 35572 342615
rect 39592 342514 39620 343431
rect 39580 342508 39632 342514
rect 39580 342450 39632 342456
rect 35532 342304 35584 342310
rect 35532 342246 35584 342252
rect 35622 341864 35678 341873
rect 35622 341799 35678 341808
rect 35636 341222 35664 341799
rect 39776 341494 39804 344927
rect 40420 343874 40448 345743
rect 40408 343868 40460 343874
rect 40408 343810 40460 343816
rect 41696 343664 41748 343670
rect 42064 343664 42116 343670
rect 41748 343612 42064 343618
rect 41696 343606 42116 343612
rect 41708 343590 42104 343606
rect 42996 343097 43024 369826
rect 43272 343505 43300 385018
rect 43442 377768 43498 377777
rect 43442 377703 43498 377712
rect 43456 359990 43484 377703
rect 43626 377360 43682 377369
rect 43626 377295 43682 377304
rect 43640 364138 43668 377295
rect 43628 364132 43680 364138
rect 43628 364074 43680 364080
rect 43444 359984 43496 359990
rect 43444 359926 43496 359932
rect 43824 344729 43852 433978
rect 43996 429344 44048 429350
rect 43996 429286 44048 429292
rect 44008 387161 44036 429286
rect 44284 428913 44312 554746
rect 44652 550634 44680 556815
rect 44560 550606 44680 550634
rect 44560 429214 44588 550606
rect 44548 429208 44600 429214
rect 44548 429150 44600 429156
rect 44270 428904 44326 428913
rect 44270 428839 44326 428848
rect 44178 426864 44234 426873
rect 44178 426799 44234 426808
rect 43994 387152 44050 387161
rect 43994 387087 44050 387096
rect 43994 383888 44050 383897
rect 43994 383823 44050 383832
rect 44008 345001 44036 383823
rect 44192 383722 44220 426799
rect 44548 426488 44600 426494
rect 44548 426430 44600 426436
rect 44362 421288 44418 421297
rect 44362 421223 44418 421232
rect 44376 408338 44404 421223
rect 44364 408332 44416 408338
rect 44364 408274 44416 408280
rect 44560 383926 44588 426430
rect 44548 383920 44600 383926
rect 44548 383862 44600 383868
rect 44180 383716 44232 383722
rect 44180 383658 44232 383664
rect 44178 381848 44234 381857
rect 44178 381783 44234 381792
rect 43994 344992 44050 345001
rect 43994 344927 44050 344936
rect 43810 344720 43866 344729
rect 43810 344655 43866 344664
rect 43258 343496 43314 343505
rect 43258 343431 43314 343440
rect 39946 343088 40002 343097
rect 39946 343023 40002 343032
rect 42982 343088 43038 343097
rect 42982 343023 43038 343032
rect 39960 342718 39988 343023
rect 39948 342712 40000 342718
rect 39948 342654 40000 342660
rect 40316 342304 40368 342310
rect 40314 342272 40316 342281
rect 40368 342272 40370 342281
rect 40314 342207 40370 342216
rect 43258 342272 43314 342281
rect 43258 342207 43314 342216
rect 35808 341488 35860 341494
rect 35806 341456 35808 341465
rect 39764 341488 39816 341494
rect 35860 341456 35862 341465
rect 39764 341430 39816 341436
rect 35806 341391 35862 341400
rect 40316 341284 40368 341290
rect 40316 341226 40368 341232
rect 35624 341216 35676 341222
rect 35624 341158 35676 341164
rect 35624 341080 35676 341086
rect 35622 341048 35624 341057
rect 40328 341057 40356 341226
rect 41696 341080 41748 341086
rect 35676 341048 35678 341057
rect 35622 340983 35678 340992
rect 40314 341048 40370 341057
rect 42064 341080 42116 341086
rect 41748 341028 42064 341034
rect 41696 341022 42116 341028
rect 42890 341048 42946 341057
rect 41708 341006 42104 341022
rect 40314 340983 40370 340992
rect 42890 340983 42946 340992
rect 35808 340944 35860 340950
rect 35808 340886 35860 340892
rect 41696 340944 41748 340950
rect 42064 340944 42116 340950
rect 41748 340892 42064 340898
rect 41696 340886 42116 340892
rect 35820 340649 35848 340886
rect 41708 340870 42104 340886
rect 35806 340640 35862 340649
rect 35806 340575 35862 340584
rect 35622 340232 35678 340241
rect 35622 340167 35678 340176
rect 35636 339658 35664 340167
rect 35624 339652 35676 339658
rect 35624 339594 35676 339600
rect 39580 339652 39632 339658
rect 39580 339594 39632 339600
rect 39592 339017 39620 339594
rect 35622 339008 35678 339017
rect 35622 338943 35678 338952
rect 39578 339008 39634 339017
rect 39578 338943 39634 338952
rect 35636 338162 35664 338943
rect 35806 338600 35862 338609
rect 35806 338535 35862 338544
rect 35820 338366 35848 338535
rect 35808 338360 35860 338366
rect 35808 338302 35860 338308
rect 41512 338360 41564 338366
rect 41512 338302 41564 338308
rect 41524 338201 41552 338302
rect 41510 338192 41566 338201
rect 35624 338156 35676 338162
rect 41708 338162 42104 338178
rect 41510 338127 41566 338136
rect 41696 338156 42116 338162
rect 35624 338098 35676 338104
rect 41748 338150 42064 338156
rect 41696 338098 41748 338104
rect 42064 338098 42116 338104
rect 35806 337784 35862 337793
rect 35806 337719 35862 337728
rect 35820 337210 35848 337719
rect 35808 337204 35860 337210
rect 35808 337146 35860 337152
rect 40040 337204 40092 337210
rect 40040 337146 40092 337152
rect 40052 336977 40080 337146
rect 41696 337000 41748 337006
rect 35530 336968 35586 336977
rect 35530 336903 35532 336912
rect 35584 336903 35586 336912
rect 35806 336968 35862 336977
rect 35806 336903 35862 336912
rect 40038 336968 40094 336977
rect 42064 337000 42116 337006
rect 41748 336948 42064 336954
rect 41696 336942 42116 336948
rect 41708 336926 42104 336942
rect 40038 336903 40094 336912
rect 35532 336874 35584 336880
rect 35820 336802 35848 336903
rect 41708 336802 42104 336818
rect 35808 336796 35860 336802
rect 35808 336738 35860 336744
rect 41696 336796 42116 336802
rect 41748 336790 42064 336796
rect 41696 336738 41748 336744
rect 42064 336738 42116 336744
rect 35622 336152 35678 336161
rect 35622 336087 35678 336096
rect 35636 335646 35664 336087
rect 35806 335744 35862 335753
rect 35806 335679 35862 335688
rect 35624 335640 35676 335646
rect 35624 335582 35676 335588
rect 35820 335374 35848 335679
rect 40316 335640 40368 335646
rect 40316 335582 40368 335588
rect 35808 335368 35860 335374
rect 39672 335368 39724 335374
rect 35808 335310 35860 335316
rect 39670 335336 39672 335345
rect 39724 335336 39726 335345
rect 39670 335271 39726 335280
rect 40328 334937 40356 335582
rect 35438 334928 35494 334937
rect 35438 334863 35494 334872
rect 35806 334928 35862 334937
rect 35806 334863 35862 334872
rect 40314 334928 40370 334937
rect 40314 334863 40370 334872
rect 35452 334150 35480 334863
rect 35622 334520 35678 334529
rect 35622 334455 35678 334464
rect 35440 334144 35492 334150
rect 35440 334086 35492 334092
rect 35636 334014 35664 334455
rect 35820 334422 35848 334863
rect 35808 334416 35860 334422
rect 35808 334358 35860 334364
rect 40316 334416 40368 334422
rect 40316 334358 40368 334364
rect 39580 334144 39632 334150
rect 39578 334112 39580 334121
rect 39632 334112 39634 334121
rect 39578 334047 39634 334056
rect 35624 334008 35676 334014
rect 35624 333950 35676 333956
rect 40328 333713 40356 334358
rect 42064 334144 42116 334150
rect 41708 334092 42064 334098
rect 41708 334086 42116 334092
rect 41708 334070 42104 334086
rect 41708 334014 41736 334070
rect 41696 334008 41748 334014
rect 41696 333950 41748 333956
rect 40314 333704 40370 333713
rect 40314 333639 40370 333648
rect 35622 333296 35678 333305
rect 35622 333231 35678 333240
rect 35636 332790 35664 333231
rect 35806 332888 35862 332897
rect 35806 332823 35862 332832
rect 35624 332784 35676 332790
rect 35624 332726 35676 332732
rect 35820 332654 35848 332823
rect 39580 332784 39632 332790
rect 39580 332726 39632 332732
rect 35808 332648 35860 332654
rect 35808 332590 35860 332596
rect 39592 330585 39620 332726
rect 41696 332648 41748 332654
rect 42064 332648 42116 332654
rect 41748 332596 42064 332602
rect 41696 332590 42116 332596
rect 41708 332574 42104 332590
rect 39578 330576 39634 330585
rect 39578 330511 39634 330520
rect 42432 327072 42484 327078
rect 42432 327014 42484 327020
rect 42444 326278 42472 327014
rect 42168 326210 42196 326264
rect 42260 326250 42472 326278
rect 42260 326210 42288 326250
rect 42168 326182 42288 326210
rect 42432 325644 42484 325650
rect 42432 325586 42484 325592
rect 42444 325054 42472 325586
rect 42182 325026 42472 325054
rect 41786 324864 41842 324873
rect 41786 324799 41842 324808
rect 41800 324428 41828 324799
rect 42432 324284 42484 324290
rect 42432 324226 42484 324232
rect 42444 323762 42472 324226
rect 42182 323734 42472 323762
rect 41786 322824 41842 322833
rect 41786 322759 41842 322768
rect 41800 322592 41828 322759
rect 42432 321564 42484 321570
rect 42432 321506 42484 321512
rect 42182 321354 42288 321382
rect 42260 321298 42288 321354
rect 42248 321292 42300 321298
rect 42248 321234 42300 321240
rect 42444 320739 42472 321506
rect 42182 320711 42472 320739
rect 42432 320136 42484 320142
rect 42182 320084 42432 320090
rect 42182 320078 42484 320084
rect 42182 320062 42472 320078
rect 42182 319518 42472 319546
rect 42444 318850 42472 319518
rect 42432 318844 42484 318850
rect 42432 318786 42484 318792
rect 42432 317416 42484 317422
rect 42432 317358 42484 317364
rect 42248 317280 42300 317286
rect 42248 317222 42300 317228
rect 42260 317059 42288 317222
rect 42182 317031 42288 317059
rect 42444 316418 42472 317358
rect 42182 316390 42472 316418
rect 42432 315920 42484 315926
rect 42432 315862 42484 315868
rect 42444 315771 42472 315862
rect 42182 315743 42472 315771
rect 41786 315616 41842 315625
rect 41786 315551 41842 315560
rect 41800 315180 41828 315551
rect 41786 313712 41842 313721
rect 41786 313647 41842 313656
rect 41800 313344 41828 313647
rect 41786 313032 41842 313041
rect 41786 312967 41842 312976
rect 41800 312732 41828 312967
rect 42168 312174 42288 312202
rect 42168 312052 42196 312174
rect 42260 312066 42288 312174
rect 42260 312038 42472 312066
rect 42444 310418 42472 312038
rect 42432 310412 42484 310418
rect 42432 310354 42484 310360
rect 8588 301988 8616 302124
rect 9048 301988 9076 302124
rect 9508 301988 9536 302124
rect 9968 301988 9996 302124
rect 10428 301988 10456 302124
rect 10888 301988 10916 302124
rect 11348 301988 11376 302124
rect 11808 301988 11836 302124
rect 12268 301988 12296 302124
rect 12728 301988 12756 302124
rect 13188 301988 13216 302124
rect 13648 301988 13676 302124
rect 14108 301988 14136 302124
rect 41142 299296 41198 299305
rect 41142 299231 41198 299240
rect 40958 298480 41014 298489
rect 40958 298415 41014 298424
rect 40972 298314 41000 298415
rect 41156 298314 41184 299231
rect 42706 298888 42762 298897
rect 42706 298823 42762 298832
rect 41696 298376 41748 298382
rect 42064 298376 42116 298382
rect 41748 298324 42064 298330
rect 41696 298318 42116 298324
rect 40960 298308 41012 298314
rect 40960 298250 41012 298256
rect 41144 298308 41196 298314
rect 41708 298302 42104 298318
rect 41144 298250 41196 298256
rect 42064 298240 42116 298246
rect 41708 298188 42064 298194
rect 41708 298182 42116 298188
rect 41708 298178 42104 298182
rect 41696 298172 42104 298178
rect 41748 298166 42104 298172
rect 41696 298114 41748 298120
rect 40958 298072 41014 298081
rect 40958 298007 41014 298016
rect 40972 296750 41000 298007
rect 40960 296744 41012 296750
rect 40960 296686 41012 296692
rect 41696 296744 41748 296750
rect 42064 296744 42116 296750
rect 41748 296704 42064 296732
rect 41696 296686 41748 296692
rect 42064 296686 42116 296692
rect 42062 295624 42118 295633
rect 42062 295559 42118 295568
rect 41786 295216 41842 295225
rect 41786 295151 41842 295160
rect 41800 294953 41828 295151
rect 41786 294944 41842 294953
rect 41786 294879 41842 294888
rect 35162 294808 35218 294817
rect 35162 294743 35218 294752
rect 35176 284986 35204 294743
rect 41786 293584 41842 293593
rect 41616 293542 41786 293570
rect 41616 292602 41644 293542
rect 41786 293519 41842 293528
rect 40500 292597 40552 292602
rect 40498 292596 40554 292597
rect 40498 292588 40500 292596
rect 40552 292588 40554 292596
rect 41604 292596 41656 292602
rect 41604 292538 41656 292544
rect 40498 292523 40554 292532
rect 42076 292369 42104 295559
rect 42062 292360 42118 292369
rect 42062 292295 42118 292304
rect 41142 290728 41198 290737
rect 41142 290663 41198 290672
rect 40958 290320 41014 290329
rect 40958 290255 41014 290264
rect 40972 289134 41000 290255
rect 41156 289882 41184 290663
rect 41786 290048 41842 290057
rect 41340 290006 41786 290034
rect 41144 289876 41196 289882
rect 41340 289837 41368 290006
rect 41786 289983 41842 289992
rect 41696 289876 41748 289882
rect 41144 289818 41196 289824
rect 41326 289828 41382 289837
rect 42064 289876 42116 289882
rect 41748 289836 42064 289864
rect 41696 289818 41748 289824
rect 42064 289818 42116 289824
rect 42720 289814 42748 298823
rect 42904 298382 42932 340983
rect 43076 337000 43128 337006
rect 43076 336942 43128 336948
rect 43088 315926 43116 336942
rect 43076 315920 43128 315926
rect 43076 315862 43128 315868
rect 43272 300121 43300 342207
rect 44192 340950 44220 381783
rect 44546 378176 44602 378185
rect 44546 378111 44602 378120
rect 44362 376952 44418 376961
rect 44362 376887 44418 376896
rect 44376 364993 44404 376887
rect 44362 364984 44418 364993
rect 44362 364919 44418 364928
rect 44560 360194 44588 378111
rect 44548 360188 44600 360194
rect 44548 360130 44600 360136
rect 44180 340944 44232 340950
rect 44180 340886 44232 340892
rect 44178 339008 44234 339017
rect 44178 338943 44234 338952
rect 43442 336968 43498 336977
rect 43442 336903 43498 336912
rect 43456 327078 43484 336903
rect 43812 336796 43864 336802
rect 43812 336738 43864 336744
rect 43626 334928 43682 334937
rect 43626 334863 43682 334872
rect 43444 327072 43496 327078
rect 43444 327014 43496 327020
rect 43640 321570 43668 334863
rect 43628 321564 43680 321570
rect 43628 321506 43680 321512
rect 43628 318096 43680 318102
rect 43628 318038 43680 318044
rect 43444 310548 43496 310554
rect 43444 310490 43496 310496
rect 43258 300112 43314 300121
rect 43258 300047 43314 300056
rect 42892 298376 42944 298382
rect 42892 298318 42944 298324
rect 43258 297256 43314 297265
rect 43258 297191 43314 297200
rect 43074 293992 43130 294001
rect 43074 293927 43130 293936
rect 42890 291136 42946 291145
rect 42890 291071 42946 291080
rect 42904 290018 42932 291071
rect 42892 290012 42944 290018
rect 42892 289954 42944 289960
rect 42720 289786 42932 289814
rect 41326 289763 41382 289772
rect 40960 289128 41012 289134
rect 40960 289070 41012 289076
rect 41696 289128 41748 289134
rect 41696 289070 41748 289076
rect 41708 288946 41736 289070
rect 41708 288918 42380 288946
rect 35164 284980 35216 284986
rect 35164 284922 35216 284928
rect 41696 284980 41748 284986
rect 41696 284922 41748 284928
rect 41708 284866 41736 284922
rect 41708 284838 42288 284866
rect 42260 283059 42288 284838
rect 42182 283031 42288 283059
rect 42352 281874 42380 288918
rect 42182 281846 42380 281874
rect 41970 281480 42026 281489
rect 41970 281415 42026 281424
rect 41984 281180 42012 281415
rect 42182 280554 42472 280582
rect 42248 280152 42300 280158
rect 42248 280094 42300 280100
rect 42260 279426 42288 280094
rect 42168 279398 42288 279426
rect 42168 279344 42196 279398
rect 42444 278594 42472 280554
rect 42432 278588 42484 278594
rect 42432 278530 42484 278536
rect 42432 278452 42484 278458
rect 42432 278394 42484 278400
rect 42444 278202 42472 278394
rect 42168 278066 42196 278188
rect 42260 278174 42472 278202
rect 42260 278066 42288 278174
rect 42168 278038 42288 278066
rect 42246 277944 42302 277953
rect 42246 277879 42302 277888
rect 41800 277409 41828 277508
rect 41786 277400 41842 277409
rect 41786 277335 41842 277344
rect 42062 277128 42118 277137
rect 42062 277063 42118 277072
rect 42076 276896 42104 277063
rect 42062 276584 42118 276593
rect 42062 276519 42118 276528
rect 42076 276352 42104 276519
rect 42260 273850 42288 277879
rect 42182 273822 42288 273850
rect 41786 273456 41842 273465
rect 41786 273391 41842 273400
rect 41800 273224 41828 273391
rect 42432 273216 42484 273222
rect 42432 273158 42484 273164
rect 42444 272558 42472 273158
rect 42182 272530 42472 272558
rect 41786 272368 41842 272377
rect 41786 272303 41842 272312
rect 41800 272000 41828 272303
rect 41786 270464 41842 270473
rect 41786 270399 41842 270408
rect 41800 270164 41828 270399
rect 42182 269507 42564 269535
rect 42340 269068 42392 269074
rect 42340 269010 42392 269016
rect 42352 268886 42380 269010
rect 42182 268858 42380 268886
rect 42536 267714 42564 269507
rect 42524 267708 42576 267714
rect 42524 267650 42576 267656
rect 40038 259448 40094 259457
rect 40038 259383 40094 259392
rect 8588 258740 8616 258876
rect 9048 258740 9076 258876
rect 9508 258740 9536 258876
rect 9968 258740 9996 258876
rect 10428 258740 10456 258876
rect 10888 258740 10916 258876
rect 11348 258740 11376 258876
rect 11808 258740 11836 258876
rect 12268 258740 12296 258876
rect 12728 258740 12756 258876
rect 13188 258740 13216 258876
rect 13648 258740 13676 258876
rect 14108 258740 14136 258876
rect 40052 258262 40080 259383
rect 40406 258904 40462 258913
rect 40406 258839 40462 258848
rect 35808 258256 35860 258262
rect 35808 258198 35860 258204
rect 40040 258256 40092 258262
rect 40040 258198 40092 258204
rect 35820 258097 35848 258198
rect 35806 258088 35862 258097
rect 35806 258023 35862 258032
rect 39578 257952 39634 257961
rect 39578 257887 39634 257896
rect 35622 257544 35678 257553
rect 35622 257479 35678 257488
rect 35636 256766 35664 257479
rect 39592 257174 39620 257887
rect 39946 257544 40002 257553
rect 39946 257479 40002 257488
rect 35808 257168 35860 257174
rect 35806 257136 35808 257145
rect 39580 257168 39632 257174
rect 35860 257136 35862 257145
rect 39580 257110 39632 257116
rect 35806 257071 35862 257080
rect 35808 256896 35860 256902
rect 35808 256838 35860 256844
rect 35624 256760 35676 256766
rect 35820 256737 35848 256838
rect 35624 256702 35676 256708
rect 35806 256728 35862 256737
rect 35806 256663 35862 256672
rect 35806 256320 35862 256329
rect 35806 256255 35862 256264
rect 35622 255912 35678 255921
rect 35622 255847 35678 255856
rect 35636 255474 35664 255847
rect 35820 255746 35848 256255
rect 35808 255740 35860 255746
rect 35808 255682 35860 255688
rect 35806 255504 35862 255513
rect 35624 255468 35676 255474
rect 35806 255439 35862 255448
rect 35624 255410 35676 255416
rect 35820 255338 35848 255439
rect 35808 255332 35860 255338
rect 35808 255274 35860 255280
rect 35346 255096 35402 255105
rect 35346 255031 35402 255040
rect 35162 254688 35218 254697
rect 35162 254623 35218 254632
rect 35176 253978 35204 254623
rect 35360 254114 35388 255031
rect 35532 254584 35584 254590
rect 35532 254526 35584 254532
rect 39304 254584 39356 254590
rect 39304 254526 39356 254532
rect 35544 254289 35572 254526
rect 35808 254312 35860 254318
rect 35530 254280 35586 254289
rect 35530 254215 35586 254224
rect 35806 254280 35808 254289
rect 35860 254280 35862 254289
rect 35806 254215 35862 254224
rect 35348 254108 35400 254114
rect 35348 254050 35400 254056
rect 35164 253972 35216 253978
rect 35164 253914 35216 253920
rect 35806 253464 35862 253473
rect 35806 253399 35862 253408
rect 35622 253056 35678 253065
rect 35622 252991 35678 253000
rect 35636 252754 35664 252991
rect 35820 252890 35848 253399
rect 39316 253065 39344 254526
rect 39960 254386 39988 257479
rect 40420 256970 40448 258839
rect 40408 256964 40460 256970
rect 40408 256906 40460 256912
rect 42064 256896 42116 256902
rect 41708 256844 42064 256850
rect 41708 256838 42116 256844
rect 41708 256834 42104 256838
rect 41696 256828 42104 256834
rect 41748 256822 42104 256828
rect 41696 256770 41748 256776
rect 40314 256728 40370 256737
rect 40314 256663 40370 256672
rect 39948 254380 40000 254386
rect 39948 254322 40000 254328
rect 40328 254182 40356 256663
rect 41420 255740 41472 255746
rect 41420 255682 41472 255688
rect 41432 255105 41460 255682
rect 42904 255542 42932 289786
rect 43088 273222 43116 293927
rect 43076 273216 43128 273222
rect 43076 273158 43128 273164
rect 43272 257553 43300 297191
rect 43258 257544 43314 257553
rect 43258 257479 43314 257488
rect 41696 255536 41748 255542
rect 42064 255536 42116 255542
rect 41748 255484 42064 255490
rect 41696 255478 42116 255484
rect 42892 255536 42944 255542
rect 42892 255478 42944 255484
rect 41708 255462 42104 255478
rect 41708 255338 42104 255354
rect 41696 255332 42116 255338
rect 41748 255326 42064 255332
rect 41696 255274 41748 255280
rect 42064 255274 42116 255280
rect 41418 255096 41474 255105
rect 41418 255031 41474 255040
rect 40316 254176 40368 254182
rect 40316 254118 40368 254124
rect 41696 253972 41748 253978
rect 42064 253972 42116 253978
rect 41748 253920 42064 253934
rect 41696 253914 42116 253920
rect 41708 253906 42104 253914
rect 39302 253056 39358 253065
rect 39302 252991 39358 253000
rect 42890 253056 42946 253065
rect 42890 252991 42946 253000
rect 41708 252890 42104 252906
rect 35808 252884 35860 252890
rect 35808 252826 35860 252832
rect 41696 252884 42116 252890
rect 41748 252878 42064 252884
rect 41696 252826 41748 252832
rect 42064 252826 42116 252832
rect 42708 252884 42760 252890
rect 42708 252826 42760 252832
rect 35624 252748 35676 252754
rect 35624 252690 35676 252696
rect 41696 252748 41748 252754
rect 41696 252690 41748 252696
rect 35806 252648 35862 252657
rect 35806 252583 35808 252592
rect 35860 252583 35862 252592
rect 41510 252648 41566 252657
rect 41510 252583 41512 252592
rect 35808 252554 35860 252560
rect 41564 252583 41566 252592
rect 41512 252554 41564 252560
rect 35806 252240 35862 252249
rect 35806 252175 35862 252184
rect 40590 252240 40646 252249
rect 40590 252175 40646 252184
rect 35622 251832 35678 251841
rect 35622 251767 35678 251776
rect 35636 251258 35664 251767
rect 35820 251666 35848 252175
rect 40604 251666 40632 252175
rect 41326 251832 41382 251841
rect 41326 251767 41382 251776
rect 35808 251660 35860 251666
rect 35808 251602 35860 251608
rect 40592 251660 40644 251666
rect 40592 251602 40644 251608
rect 35806 251424 35862 251433
rect 41340 251394 41368 251767
rect 41510 251424 41566 251433
rect 35806 251359 35808 251368
rect 35860 251359 35862 251368
rect 41328 251388 41380 251394
rect 35808 251330 35860 251336
rect 41510 251359 41566 251368
rect 41328 251330 41380 251336
rect 41524 251258 41552 251359
rect 35624 251252 35676 251258
rect 35624 251194 35676 251200
rect 41512 251252 41564 251258
rect 41512 251194 41564 251200
rect 35438 251016 35494 251025
rect 35438 250951 35494 250960
rect 35452 249830 35480 250951
rect 35622 250608 35678 250617
rect 35622 250543 35678 250552
rect 35636 249966 35664 250543
rect 35808 250232 35860 250238
rect 35806 250200 35808 250209
rect 39396 250232 39448 250238
rect 35860 250200 35862 250209
rect 35806 250135 35862 250144
rect 39394 250200 39396 250209
rect 39448 250200 39450 250209
rect 39394 250135 39450 250144
rect 40132 250028 40184 250034
rect 40132 249970 40184 249976
rect 35624 249960 35676 249966
rect 35624 249902 35676 249908
rect 35440 249824 35492 249830
rect 35440 249766 35492 249772
rect 39580 249824 39632 249830
rect 39580 249766 39632 249772
rect 35530 248976 35586 248985
rect 35530 248911 35586 248920
rect 35806 248976 35862 248985
rect 35806 248911 35862 248920
rect 35544 248742 35572 248911
rect 35532 248736 35584 248742
rect 35532 248678 35584 248684
rect 35820 248470 35848 248911
rect 35808 248464 35860 248470
rect 35808 248406 35860 248412
rect 35622 248160 35678 248169
rect 35622 248095 35678 248104
rect 35438 247752 35494 247761
rect 35438 247687 35494 247696
rect 35452 247110 35480 247687
rect 35636 247382 35664 248095
rect 35808 247580 35860 247586
rect 35808 247522 35860 247528
rect 35624 247376 35676 247382
rect 35820 247353 35848 247522
rect 35624 247318 35676 247324
rect 35806 247344 35862 247353
rect 35806 247279 35862 247288
rect 35624 247240 35676 247246
rect 35624 247182 35676 247188
rect 35440 247104 35492 247110
rect 35440 247046 35492 247052
rect 35636 246945 35664 247182
rect 35622 246936 35678 246945
rect 35622 246871 35678 246880
rect 39592 245585 39620 249766
rect 40144 248985 40172 249970
rect 40130 248976 40186 248985
rect 40130 248911 40186 248920
rect 39948 248736 40000 248742
rect 39948 248678 40000 248684
rect 39960 248577 39988 248678
rect 39946 248568 40002 248577
rect 39946 248503 40002 248512
rect 40132 248464 40184 248470
rect 40132 248406 40184 248412
rect 40144 248169 40172 248406
rect 40130 248160 40186 248169
rect 40130 248095 40186 248104
rect 41510 247752 41566 247761
rect 41510 247687 41566 247696
rect 41524 247586 41552 247687
rect 41512 247580 41564 247586
rect 41512 247522 41564 247528
rect 40132 247376 40184 247382
rect 40130 247344 40132 247353
rect 40184 247344 40186 247353
rect 40130 247279 40186 247288
rect 41052 247240 41104 247246
rect 41052 247182 41104 247188
rect 41064 246129 41092 247182
rect 41512 247104 41564 247110
rect 41512 247046 41564 247052
rect 41524 246945 41552 247046
rect 41510 246936 41566 246945
rect 41510 246871 41566 246880
rect 41050 246120 41106 246129
rect 41050 246055 41106 246064
rect 39578 245576 39634 245585
rect 39578 245511 39634 245520
rect 41708 244274 41736 252690
rect 42522 252240 42578 252249
rect 42522 252175 42578 252184
rect 42154 247752 42210 247761
rect 42154 247687 42210 247696
rect 42168 247518 42196 247687
rect 42156 247512 42208 247518
rect 42156 247454 42208 247460
rect 42064 247104 42116 247110
rect 42064 247046 42116 247052
rect 42076 246945 42104 247046
rect 42062 246936 42118 246945
rect 42062 246871 42118 246880
rect 41708 244246 42472 244274
rect 42248 240100 42300 240106
rect 42248 240042 42300 240048
rect 42260 239850 42288 240042
rect 42182 239822 42288 239850
rect 42182 238635 42288 238663
rect 42260 238513 42288 238635
rect 42246 238504 42302 238513
rect 42246 238439 42302 238448
rect 42444 238014 42472 244246
rect 42182 237986 42472 238014
rect 41786 236600 41842 236609
rect 41786 236535 41842 236544
rect 41800 236164 41828 236535
rect 42340 235952 42392 235958
rect 42340 235894 42392 235900
rect 42352 234983 42380 235894
rect 42182 234955 42380 234983
rect 42340 234592 42392 234598
rect 41786 234560 41842 234569
rect 42340 234534 42392 234540
rect 41786 234495 41842 234504
rect 41800 234328 41828 234495
rect 42352 233695 42380 234534
rect 42182 233667 42380 233695
rect 42168 233158 42380 233186
rect 42168 233104 42196 233158
rect 42352 232082 42380 233158
rect 42340 232076 42392 232082
rect 42340 232018 42392 232024
rect 42340 231804 42392 231810
rect 42340 231746 42392 231752
rect 42352 230670 42380 231746
rect 42182 230642 42380 230670
rect 42156 230444 42208 230450
rect 42156 230386 42208 230392
rect 42168 229976 42196 230386
rect 42340 230308 42392 230314
rect 42340 230250 42392 230256
rect 42352 229378 42380 230250
rect 42182 229350 42380 229378
rect 42536 228834 42564 252175
rect 42720 237425 42748 252826
rect 42706 237416 42762 237425
rect 42706 237351 42762 237360
rect 42182 228806 42564 228834
rect 42062 227352 42118 227361
rect 42062 227287 42118 227296
rect 42076 226984 42104 227287
rect 42168 226358 42288 226386
rect 42168 226304 42196 226358
rect 42260 226318 42288 226358
rect 42260 226290 42472 226318
rect 42182 225678 42288 225706
rect 41694 223680 41750 223689
rect 41694 223615 41750 223624
rect 40682 222592 40738 222601
rect 40682 222527 40738 222536
rect 28538 222320 28594 222329
rect 28538 222255 28594 222264
rect 8588 215492 8616 215628
rect 9048 215492 9076 215628
rect 9508 215492 9536 215628
rect 9968 215492 9996 215628
rect 10428 215492 10456 215628
rect 10888 215492 10916 215628
rect 11348 215492 11376 215628
rect 11808 215492 11836 215628
rect 12268 215492 12296 215628
rect 12728 215492 12756 215628
rect 13188 215492 13216 215628
rect 13648 215492 13676 215628
rect 14108 215492 14136 215628
rect 28552 212673 28580 222255
rect 39762 218376 39818 218385
rect 39762 218311 39818 218320
rect 39776 214742 39804 218311
rect 40222 218104 40278 218113
rect 40222 218039 40278 218048
rect 35532 214736 35584 214742
rect 35346 214704 35402 214713
rect 35532 214678 35584 214684
rect 39764 214736 39816 214742
rect 39764 214678 39816 214684
rect 35346 214639 35402 214648
rect 35360 213994 35388 214639
rect 35544 214305 35572 214678
rect 35808 214328 35860 214334
rect 35530 214296 35586 214305
rect 35530 214231 35586 214240
rect 35806 214296 35808 214305
rect 35860 214296 35862 214305
rect 35806 214231 35862 214240
rect 39762 214296 39818 214305
rect 39762 214231 39818 214240
rect 35348 213988 35400 213994
rect 35348 213930 35400 213936
rect 35806 213480 35862 213489
rect 35806 213415 35862 213424
rect 35622 213072 35678 213081
rect 35622 213007 35678 213016
rect 28538 212664 28594 212673
rect 28538 212599 28594 212608
rect 35636 212566 35664 213007
rect 35820 212974 35848 213415
rect 39302 213072 39358 213081
rect 39302 213007 39304 213016
rect 39356 213007 39358 213016
rect 39304 212978 39356 212984
rect 35808 212968 35860 212974
rect 35808 212910 35860 212916
rect 39776 212702 39804 214231
rect 40236 213994 40264 218039
rect 40696 214334 40724 222527
rect 40684 214328 40736 214334
rect 40684 214270 40736 214276
rect 40224 213988 40276 213994
rect 40224 213930 40276 213936
rect 35808 212696 35860 212702
rect 35806 212664 35808 212673
rect 39764 212696 39816 212702
rect 35860 212664 35862 212673
rect 39764 212638 39816 212644
rect 41234 212664 41290 212673
rect 35806 212599 35862 212608
rect 41234 212599 41236 212608
rect 41288 212599 41290 212608
rect 41236 212570 41288 212576
rect 35624 212560 35676 212566
rect 35624 212502 35676 212508
rect 41050 212256 41106 212265
rect 41050 212191 41106 212200
rect 35806 211848 35862 211857
rect 35806 211783 35862 211792
rect 35820 211614 35848 211783
rect 35808 211608 35860 211614
rect 35808 211550 35860 211556
rect 35622 211440 35678 211449
rect 35622 211375 35678 211384
rect 39670 211440 39726 211449
rect 39670 211375 39672 211384
rect 35636 211206 35664 211375
rect 39724 211375 39726 211384
rect 39672 211346 39724 211352
rect 35808 211336 35860 211342
rect 35808 211278 35860 211284
rect 35624 211200 35676 211206
rect 35624 211142 35676 211148
rect 35820 211041 35848 211278
rect 41064 211274 41092 212191
rect 41234 211848 41290 211857
rect 41234 211783 41290 211792
rect 41248 211614 41276 211783
rect 41236 211608 41288 211614
rect 41236 211550 41288 211556
rect 41052 211268 41104 211274
rect 41052 211210 41104 211216
rect 35806 211032 35862 211041
rect 35806 210967 35862 210976
rect 35622 210624 35678 210633
rect 35622 210559 35678 210568
rect 35636 209982 35664 210559
rect 35806 210216 35862 210225
rect 35806 210151 35862 210160
rect 35624 209976 35676 209982
rect 35624 209918 35676 209924
rect 35820 209846 35848 210151
rect 41708 209982 41736 223615
rect 42260 223582 42288 225678
rect 42444 224942 42472 226290
rect 42432 224936 42484 224942
rect 42432 224878 42484 224884
rect 42248 223576 42300 223582
rect 42248 223518 42300 223524
rect 42616 223032 42668 223038
rect 42616 222974 42668 222980
rect 42628 222601 42656 222974
rect 42614 222592 42670 222601
rect 42614 222527 42670 222536
rect 42156 212696 42208 212702
rect 42154 212664 42156 212673
rect 42208 212664 42210 212673
rect 42154 212599 42210 212608
rect 42904 211449 42932 252991
rect 43074 250200 43130 250209
rect 43074 250135 43130 250144
rect 43088 230450 43116 250135
rect 43258 248976 43314 248985
rect 43258 248911 43314 248920
rect 43076 230444 43128 230450
rect 43076 230386 43128 230392
rect 43272 230314 43300 248911
rect 43260 230308 43312 230314
rect 43260 230250 43312 230256
rect 43456 218385 43484 310490
rect 43640 257961 43668 318038
rect 43824 317422 43852 336738
rect 43994 335336 44050 335345
rect 43994 335271 44050 335280
rect 43812 317416 43864 317422
rect 43812 317358 43864 317364
rect 44008 317286 44036 335271
rect 43996 317280 44048 317286
rect 43996 317222 44048 317228
rect 43810 301608 43866 301617
rect 43810 301543 43866 301552
rect 43824 301238 43852 301543
rect 43812 301232 43864 301238
rect 43812 301174 43864 301180
rect 44192 297673 44220 338943
rect 44638 334112 44694 334121
rect 44638 334047 44694 334056
rect 44454 333704 44510 333713
rect 44454 333639 44510 333648
rect 44468 321298 44496 333639
rect 44456 321292 44508 321298
rect 44456 321234 44508 321240
rect 44652 320142 44680 334047
rect 44640 320136 44692 320142
rect 44640 320078 44692 320084
rect 44546 299704 44602 299713
rect 44546 299639 44602 299648
rect 44178 297664 44234 297673
rect 44178 297599 44234 297608
rect 43994 293176 44050 293185
rect 43994 293111 44050 293120
rect 43810 290048 43866 290057
rect 43810 289983 43866 289992
rect 43824 276690 43852 289983
rect 44008 280158 44036 293111
rect 44178 291816 44234 291825
rect 44178 291751 44234 291760
rect 43996 280152 44048 280158
rect 43996 280094 44048 280100
rect 44192 277137 44220 291751
rect 44362 291544 44418 291553
rect 44362 291479 44418 291488
rect 44376 278458 44404 291479
rect 44364 278452 44416 278458
rect 44364 278394 44416 278400
rect 44178 277128 44234 277137
rect 44178 277063 44234 277072
rect 43812 276684 43864 276690
rect 43812 276626 43864 276632
rect 44560 258913 44588 299639
rect 44546 258904 44602 258913
rect 44546 258839 44602 258848
rect 43626 257952 43682 257961
rect 43626 257887 43682 257896
rect 44178 255096 44234 255105
rect 44178 255031 44234 255040
rect 43812 253972 43864 253978
rect 43812 253914 43864 253920
rect 43626 248568 43682 248577
rect 43626 248503 43682 248512
rect 43640 231810 43668 248503
rect 43628 231804 43680 231810
rect 43628 231746 43680 231752
rect 43626 225040 43682 225049
rect 43626 224975 43682 224984
rect 43442 218376 43498 218385
rect 43442 218311 43498 218320
rect 43640 212265 43668 224975
rect 43626 212256 43682 212265
rect 43626 212191 43682 212200
rect 43824 211857 43852 253914
rect 44192 213081 44220 255031
rect 44546 248160 44602 248169
rect 44546 248095 44602 248104
rect 44362 247344 44418 247353
rect 44362 247279 44418 247288
rect 44376 235958 44404 247279
rect 44364 235952 44416 235958
rect 44364 235894 44416 235900
rect 44560 234598 44588 248095
rect 44548 234592 44600 234598
rect 44548 234534 44600 234540
rect 44836 231130 44864 760271
rect 45020 754934 45048 765886
rect 45190 764552 45246 764561
rect 45190 764487 45246 764496
rect 45008 754928 45060 754934
rect 45008 754870 45060 754876
rect 45204 754526 45232 764487
rect 45192 754520 45244 754526
rect 45192 754462 45244 754468
rect 45006 729736 45062 729745
rect 45006 729671 45062 729680
rect 45020 685914 45048 729671
rect 45190 728920 45246 728929
rect 45190 728855 45246 728864
rect 45204 686118 45232 728855
rect 45192 686112 45244 686118
rect 45192 686054 45244 686060
rect 45008 685908 45060 685914
rect 45008 685850 45060 685856
rect 45190 679552 45246 679561
rect 45190 679487 45246 679496
rect 45006 677920 45062 677929
rect 45006 677855 45062 677864
rect 44824 231124 44876 231130
rect 44824 231066 44876 231072
rect 45020 229809 45048 677855
rect 45204 666602 45232 679487
rect 45192 666596 45244 666602
rect 45192 666538 45244 666544
rect 45190 631408 45246 631417
rect 45190 631343 45246 631352
rect 45204 622470 45232 631343
rect 45192 622464 45244 622470
rect 45192 622406 45244 622412
rect 45558 552392 45614 552401
rect 45558 552327 45614 552336
rect 45190 551168 45246 551177
rect 45190 551103 45246 551112
rect 45204 531350 45232 551103
rect 45374 548720 45430 548729
rect 45572 548690 45600 552327
rect 45374 548655 45430 548664
rect 45560 548684 45612 548690
rect 45388 540974 45416 548655
rect 45560 548626 45612 548632
rect 45560 548548 45612 548554
rect 45560 548490 45612 548496
rect 45572 541090 45600 548490
rect 45296 540946 45416 540974
rect 45480 541062 45600 541090
rect 45296 536330 45324 540946
rect 45480 538642 45508 541062
rect 45480 538614 45784 538642
rect 45296 536314 45416 536330
rect 45296 536308 45428 536314
rect 45296 536302 45376 536308
rect 45376 536250 45428 536256
rect 45756 534206 45784 538614
rect 45744 534200 45796 534206
rect 45744 534142 45796 534148
rect 45192 531344 45244 531350
rect 45192 531286 45244 531292
rect 45558 424824 45614 424833
rect 45558 424759 45614 424768
rect 45374 421560 45430 421569
rect 45374 421495 45430 421504
rect 45190 420744 45246 420753
rect 45190 420679 45246 420688
rect 45204 419558 45232 420679
rect 45192 419552 45244 419558
rect 45192 419494 45244 419500
rect 45192 415472 45244 415478
rect 45192 415414 45244 415420
rect 45204 345817 45232 415414
rect 45388 407114 45416 421495
rect 45376 407108 45428 407114
rect 45376 407050 45428 407056
rect 45572 404190 45600 424759
rect 45560 404184 45612 404190
rect 45560 404126 45612 404132
rect 45374 379808 45430 379817
rect 45374 379743 45430 379752
rect 45388 356046 45416 379743
rect 45376 356040 45428 356046
rect 45376 355982 45428 355988
rect 45376 347064 45428 347070
rect 45376 347006 45428 347012
rect 45190 345808 45246 345817
rect 45190 345743 45246 345752
rect 45192 341080 45244 341086
rect 45192 341022 45244 341028
rect 45204 298246 45232 341022
rect 45388 300937 45416 347006
rect 45558 330576 45614 330585
rect 45558 330511 45614 330520
rect 45572 325650 45600 330511
rect 45560 325644 45612 325650
rect 45560 325586 45612 325592
rect 45374 300928 45430 300937
rect 45374 300863 45430 300872
rect 45192 298240 45244 298246
rect 45192 298182 45244 298188
rect 45192 296744 45244 296750
rect 45192 296686 45244 296692
rect 45204 256737 45232 296686
rect 45558 296032 45614 296041
rect 45558 295967 45614 295976
rect 45572 269074 45600 295967
rect 45742 294944 45798 294953
rect 45742 294879 45798 294888
rect 45756 276593 45784 294879
rect 45926 294400 45982 294409
rect 45926 294335 45982 294344
rect 45742 276584 45798 276593
rect 45742 276519 45798 276528
rect 45560 269068 45612 269074
rect 45560 269010 45612 269016
rect 45940 267714 45968 294335
rect 45928 267708 45980 267714
rect 45928 267650 45980 267656
rect 45190 256728 45246 256737
rect 45190 256663 45246 256672
rect 45560 255332 45612 255338
rect 45560 255274 45612 255280
rect 45190 251832 45246 251841
rect 45190 251767 45246 251776
rect 45204 240106 45232 251767
rect 45192 240100 45244 240106
rect 45192 240042 45244 240048
rect 45006 229800 45062 229809
rect 45006 229735 45062 229744
rect 45572 214305 45600 255274
rect 45834 251424 45890 251433
rect 45834 251359 45890 251368
rect 45848 232082 45876 251359
rect 46018 246120 46074 246129
rect 46018 246055 46074 246064
rect 46032 238513 46060 246055
rect 46018 238504 46074 238513
rect 46018 238439 46074 238448
rect 45836 232076 45888 232082
rect 45836 232018 45888 232024
rect 46216 231538 46244 806239
rect 47596 799066 47624 923238
rect 50344 909492 50396 909498
rect 50344 909434 50396 909440
rect 50356 815658 50384 909434
rect 51908 858424 51960 858430
rect 51908 858366 51960 858372
rect 51724 818372 51776 818378
rect 51724 818314 51776 818320
rect 50344 815652 50396 815658
rect 50344 815594 50396 815600
rect 48964 807356 49016 807362
rect 48964 807298 49016 807304
rect 47584 799060 47636 799066
rect 47584 799002 47636 799008
rect 47768 793620 47820 793626
rect 47768 793562 47820 793568
rect 47582 763328 47638 763337
rect 47582 763263 47638 763272
rect 46386 721168 46442 721177
rect 46386 721103 46442 721112
rect 46204 231532 46256 231538
rect 46204 231474 46256 231480
rect 46400 227497 46428 721103
rect 46572 446412 46624 446418
rect 46572 446354 46624 446360
rect 46584 324290 46612 446354
rect 46938 424008 46994 424017
rect 46938 423943 46994 423952
rect 46952 397458 46980 423943
rect 46940 397452 46992 397458
rect 46940 397394 46992 397400
rect 47030 338192 47086 338201
rect 47030 338127 47086 338136
rect 47216 338156 47268 338162
rect 46756 336796 46808 336802
rect 46756 336738 46808 336744
rect 46572 324284 46624 324290
rect 46572 324226 46624 324232
rect 46768 259457 46796 336738
rect 47044 318850 47072 338127
rect 47216 338098 47268 338104
rect 47032 318844 47084 318850
rect 47032 318786 47084 318792
rect 47228 310418 47256 338098
rect 47216 310412 47268 310418
rect 47216 310354 47268 310360
rect 46754 259448 46810 259457
rect 46754 259383 46810 259392
rect 46938 252648 46994 252657
rect 46938 252583 46994 252592
rect 46386 227488 46442 227497
rect 46386 227423 46442 227432
rect 46952 223582 46980 252583
rect 47122 245576 47178 245585
rect 47122 245511 47178 245520
rect 47136 224942 47164 245511
rect 47596 231402 47624 763263
rect 47780 731377 47808 793562
rect 47766 731368 47822 731377
rect 47766 731303 47822 731312
rect 47768 674892 47820 674898
rect 47768 674834 47820 674840
rect 47780 646105 47808 674834
rect 47766 646096 47822 646105
rect 47766 646031 47822 646040
rect 47768 623824 47820 623830
rect 47768 623766 47820 623772
rect 47780 601361 47808 623766
rect 47766 601352 47822 601361
rect 47766 601287 47822 601296
rect 47766 590336 47822 590345
rect 47766 590271 47822 590280
rect 47584 231396 47636 231402
rect 47584 231338 47636 231344
rect 47780 226953 47808 590271
rect 47952 480276 48004 480282
rect 47952 480218 48004 480224
rect 47964 386753 47992 480218
rect 48136 389292 48188 389298
rect 48136 389234 48188 389240
rect 47950 386744 48006 386753
rect 47950 386679 48006 386688
rect 48148 300529 48176 389234
rect 48134 300520 48190 300529
rect 48134 300455 48190 300464
rect 47952 298172 48004 298178
rect 47952 298114 48004 298120
rect 47766 226944 47822 226953
rect 47766 226879 47822 226888
rect 47124 224936 47176 224942
rect 47124 224878 47176 224884
rect 46940 223576 46992 223582
rect 46940 223518 46992 223524
rect 47582 221640 47638 221649
rect 47582 221575 47638 221584
rect 45558 214296 45614 214305
rect 45558 214231 45614 214240
rect 44178 213072 44234 213081
rect 44178 213007 44234 213016
rect 43810 211848 43866 211857
rect 43810 211783 43866 211792
rect 42890 211440 42946 211449
rect 42890 211375 42946 211384
rect 41696 209976 41748 209982
rect 41696 209918 41748 209924
rect 35808 209840 35860 209846
rect 35808 209782 35860 209788
rect 40040 209840 40092 209846
rect 40040 209782 40092 209788
rect 35622 209400 35678 209409
rect 35622 209335 35678 209344
rect 30286 208992 30342 209001
rect 30286 208927 30342 208936
rect 30300 200705 30328 208927
rect 35636 208418 35664 209335
rect 35806 208992 35862 209001
rect 35806 208927 35862 208936
rect 35820 208690 35848 208927
rect 35808 208684 35860 208690
rect 35808 208626 35860 208632
rect 39672 208616 39724 208622
rect 39670 208584 39672 208593
rect 39724 208584 39726 208593
rect 39670 208519 39726 208528
rect 35624 208412 35676 208418
rect 35624 208354 35676 208360
rect 39580 208412 39632 208418
rect 39580 208354 39632 208360
rect 35530 207360 35586 207369
rect 35530 207295 35586 207304
rect 35806 207360 35862 207369
rect 35806 207295 35808 207304
rect 35544 207058 35572 207295
rect 35860 207295 35862 207304
rect 35808 207266 35860 207272
rect 35532 207052 35584 207058
rect 35532 206994 35584 207000
rect 35622 206544 35678 206553
rect 35622 206479 35678 206488
rect 35636 205698 35664 206479
rect 35806 206136 35862 206145
rect 35806 206071 35862 206080
rect 35820 205970 35848 206071
rect 35808 205964 35860 205970
rect 35808 205906 35860 205912
rect 39396 205964 39448 205970
rect 39396 205906 39448 205912
rect 35624 205692 35676 205698
rect 35624 205634 35676 205640
rect 35622 205320 35678 205329
rect 35622 205255 35678 205264
rect 35636 204678 35664 205255
rect 35806 204912 35862 204921
rect 35806 204847 35808 204856
rect 35860 204847 35862 204856
rect 35808 204818 35860 204824
rect 35624 204672 35676 204678
rect 35624 204614 35676 204620
rect 39408 204513 39436 205906
rect 39592 205329 39620 208354
rect 39764 207324 39816 207330
rect 39764 207266 39816 207272
rect 39776 206961 39804 207266
rect 39762 206952 39818 206961
rect 39762 206887 39818 206896
rect 40052 205737 40080 209782
rect 43074 208584 43130 208593
rect 43074 208519 43130 208528
rect 40316 207052 40368 207058
rect 40316 206994 40368 207000
rect 40038 205728 40094 205737
rect 40038 205663 40094 205672
rect 39578 205320 39634 205329
rect 39578 205255 39634 205264
rect 40328 204921 40356 206994
rect 42890 206952 42946 206961
rect 42890 206887 42946 206896
rect 41144 205692 41196 205698
rect 41144 205634 41196 205640
rect 40314 204912 40370 204921
rect 39948 204876 40000 204882
rect 40314 204847 40370 204856
rect 39948 204818 40000 204824
rect 35530 204504 35586 204513
rect 35530 204439 35532 204448
rect 35584 204439 35586 204448
rect 35806 204504 35862 204513
rect 35806 204439 35862 204448
rect 39394 204504 39450 204513
rect 39394 204439 39450 204448
rect 35532 204410 35584 204416
rect 35820 204338 35848 204439
rect 35808 204332 35860 204338
rect 35808 204274 35860 204280
rect 39960 204105 39988 204818
rect 39946 204096 40002 204105
rect 39946 204031 40002 204040
rect 41156 203697 41184 205634
rect 41708 204610 42104 204626
rect 41696 204604 42116 204610
rect 41748 204598 42064 204604
rect 41696 204546 41748 204552
rect 42064 204546 42116 204552
rect 41708 204474 42104 204490
rect 41696 204468 42116 204474
rect 41748 204462 42064 204468
rect 41696 204410 41748 204416
rect 42064 204410 42116 204416
rect 41708 204338 42104 204354
rect 41696 204332 42116 204338
rect 41748 204326 42064 204332
rect 41696 204274 41748 204280
rect 42064 204274 42116 204280
rect 35622 203688 35678 203697
rect 35622 203623 35678 203632
rect 41142 203688 41198 203697
rect 41142 203623 41198 203632
rect 35636 203182 35664 203623
rect 35806 203280 35862 203289
rect 35806 203215 35862 203224
rect 41234 203280 41290 203289
rect 41234 203215 41236 203224
rect 35624 203176 35676 203182
rect 35624 203118 35676 203124
rect 35820 202910 35848 203215
rect 41288 203215 41290 203224
rect 41236 203186 41288 203192
rect 42064 203040 42116 203046
rect 41708 202988 42064 202994
rect 41708 202982 42116 202988
rect 41708 202966 42104 202982
rect 41708 202910 41736 202966
rect 35808 202904 35860 202910
rect 35808 202846 35860 202852
rect 41696 202904 41748 202910
rect 41696 202846 41748 202852
rect 30286 200696 30342 200705
rect 30286 200631 30342 200640
rect 41786 197160 41842 197169
rect 41786 197095 41842 197104
rect 41800 196656 41828 197095
rect 42904 195974 42932 206887
rect 43088 195974 43116 208519
rect 44178 205320 44234 205329
rect 44178 205255 44234 205264
rect 43258 204912 43314 204921
rect 43258 204847 43314 204856
rect 42812 195946 42932 195974
rect 42996 195946 43116 195974
rect 42432 195696 42484 195702
rect 42432 195638 42484 195644
rect 42168 195486 42288 195514
rect 42168 195432 42196 195486
rect 42260 195446 42288 195486
rect 42444 195446 42472 195638
rect 42260 195418 42472 195446
rect 41786 195256 41842 195265
rect 41786 195191 41842 195200
rect 41800 194820 41828 195191
rect 42432 193180 42484 193186
rect 42432 193122 42484 193128
rect 42444 192998 42472 193122
rect 42168 192930 42196 192984
rect 42260 192970 42472 192998
rect 42260 192930 42288 192970
rect 42168 192902 42288 192930
rect 42432 191820 42484 191826
rect 42182 191768 42432 191774
rect 42182 191762 42484 191768
rect 42182 191746 42472 191762
rect 42432 191684 42484 191690
rect 42432 191626 42484 191632
rect 41786 191584 41842 191593
rect 41786 191519 41842 191528
rect 41800 191148 41828 191519
rect 42444 190482 42472 191626
rect 42182 190454 42472 190482
rect 42432 190392 42484 190398
rect 42432 190334 42484 190340
rect 42444 189938 42472 190334
rect 42182 189910 42472 189938
rect 42432 187672 42484 187678
rect 42432 187614 42484 187620
rect 42444 187459 42472 187614
rect 42182 187431 42472 187459
rect 42812 186810 42840 195946
rect 42996 190398 43024 195946
rect 42984 190392 43036 190398
rect 42984 190334 43036 190340
rect 42182 186782 42840 186810
rect 43272 186314 43300 204847
rect 43442 204504 43498 204513
rect 43442 204439 43498 204448
rect 43456 187678 43484 204439
rect 43626 203688 43682 203697
rect 43626 203623 43682 203632
rect 43640 193186 43668 203623
rect 43810 203280 43866 203289
rect 43810 203215 43866 203224
rect 43824 195702 43852 203215
rect 43812 195696 43864 195702
rect 43812 195638 43864 195644
rect 43628 193180 43680 193186
rect 43628 193122 43680 193128
rect 43444 187672 43496 187678
rect 43444 187614 43496 187620
rect 43088 186286 43300 186314
rect 43088 186266 43116 186286
rect 42536 186238 43116 186266
rect 42536 186198 42564 186238
rect 42168 186130 42196 186184
rect 42260 186170 42564 186198
rect 42260 186130 42288 186170
rect 42168 186102 42288 186130
rect 41786 185872 41842 185881
rect 41786 185807 41842 185816
rect 41800 185605 41828 185807
rect 41786 184104 41842 184113
rect 41786 184039 41842 184048
rect 41800 183765 41828 184039
rect 44192 183530 44220 205255
rect 44364 204604 44416 204610
rect 44364 204546 44416 204552
rect 44376 191690 44404 204546
rect 47596 204474 47624 221575
rect 47964 218113 47992 298114
rect 48976 278089 49004 807298
rect 50344 805996 50396 806002
rect 50344 805938 50396 805944
rect 50356 730114 50384 805938
rect 50528 753568 50580 753574
rect 50528 753510 50580 753516
rect 50344 730108 50396 730114
rect 50344 730050 50396 730056
rect 50540 687750 50568 753510
rect 50712 714876 50764 714882
rect 50712 714818 50764 714824
rect 50528 687744 50580 687750
rect 50528 687686 50580 687692
rect 50344 676388 50396 676394
rect 50344 676330 50396 676336
rect 49148 636268 49200 636274
rect 49148 636210 49200 636216
rect 49160 601730 49188 636210
rect 49148 601724 49200 601730
rect 49148 601666 49200 601672
rect 49148 597576 49200 597582
rect 49148 597518 49200 597524
rect 49160 557802 49188 597518
rect 49148 557796 49200 557802
rect 49148 557738 49200 557744
rect 49148 546644 49200 546650
rect 49148 546586 49200 546592
rect 48962 278080 49018 278089
rect 48962 278015 49018 278024
rect 49160 228410 49188 546586
rect 49332 466472 49384 466478
rect 49332 466414 49384 466420
rect 49344 386510 49372 466414
rect 49332 386504 49384 386510
rect 49332 386446 49384 386452
rect 49332 375420 49384 375426
rect 49332 375362 49384 375368
rect 49344 301238 49372 375362
rect 49516 322992 49568 322998
rect 49516 322934 49568 322940
rect 49332 301232 49384 301238
rect 49332 301174 49384 301180
rect 49528 256902 49556 322934
rect 49516 256896 49568 256902
rect 49516 256838 49568 256844
rect 50356 228585 50384 676330
rect 50528 633480 50580 633486
rect 50528 633422 50580 633428
rect 50342 228576 50398 228585
rect 50342 228511 50398 228520
rect 49148 228404 49200 228410
rect 49148 228346 49200 228352
rect 50540 228313 50568 633422
rect 50724 626686 50752 714818
rect 51736 712298 51764 818314
rect 51920 772886 51948 858366
rect 51908 772880 51960 772886
rect 51908 772822 51960 772828
rect 51908 727320 51960 727326
rect 51908 727262 51960 727268
rect 51724 712292 51776 712298
rect 51724 712234 51776 712240
rect 51724 701072 51776 701078
rect 51724 701014 51776 701020
rect 51736 643142 51764 701014
rect 51920 687410 51948 727262
rect 51908 687404 51960 687410
rect 51908 687346 51960 687352
rect 51908 647896 51960 647902
rect 51908 647838 51960 647844
rect 51724 643136 51776 643142
rect 51724 643078 51776 643084
rect 51724 633684 51776 633690
rect 51724 633626 51776 633632
rect 50712 626680 50764 626686
rect 50712 626622 50764 626628
rect 50712 401668 50764 401674
rect 50712 401610 50764 401616
rect 50724 278594 50752 401610
rect 50712 278588 50764 278594
rect 50712 278530 50764 278536
rect 51736 231266 51764 633626
rect 51920 600370 51948 647838
rect 51908 600364 51960 600370
rect 51908 600306 51960 600312
rect 51908 583772 51960 583778
rect 51908 583714 51960 583720
rect 51920 557598 51948 583714
rect 51908 557592 51960 557598
rect 51908 557534 51960 557540
rect 52276 506524 52328 506530
rect 52276 506466 52328 506472
rect 51908 419552 51960 419558
rect 51908 419494 51960 419500
rect 51920 264246 51948 419494
rect 52092 375556 52144 375562
rect 52092 375498 52144 375504
rect 51908 264240 51960 264246
rect 51908 264182 51960 264188
rect 51724 231260 51776 231266
rect 51724 231202 51776 231208
rect 50526 228304 50582 228313
rect 50526 228239 50582 228248
rect 52104 227225 52132 375498
rect 52288 364342 52316 506466
rect 52276 364336 52328 364342
rect 52276 364278 52328 364284
rect 53116 231674 53144 931534
rect 53288 547936 53340 547942
rect 53288 547878 53340 547884
rect 53300 278186 53328 547878
rect 53472 376780 53524 376786
rect 53472 376722 53524 376728
rect 53288 278180 53340 278186
rect 53288 278122 53340 278128
rect 53484 276729 53512 376722
rect 53470 276720 53526 276729
rect 53470 276655 53526 276664
rect 54496 231810 54524 932894
rect 62118 923808 62174 923817
rect 62118 923743 62174 923752
rect 62132 923302 62160 923743
rect 62120 923296 62172 923302
rect 62120 923238 62172 923244
rect 62118 910752 62174 910761
rect 62118 910687 62174 910696
rect 62132 909498 62160 910687
rect 62120 909492 62172 909498
rect 62120 909434 62172 909440
rect 62118 897832 62174 897841
rect 62118 897767 62174 897776
rect 62132 897054 62160 897767
rect 62120 897048 62172 897054
rect 62120 896990 62172 896996
rect 62118 884776 62174 884785
rect 62118 884711 62120 884720
rect 62172 884711 62174 884720
rect 62120 884682 62172 884688
rect 62118 871720 62174 871729
rect 62118 871655 62174 871664
rect 62132 870874 62160 871655
rect 62120 870868 62172 870874
rect 62120 870810 62172 870816
rect 62118 858664 62174 858673
rect 62118 858599 62174 858608
rect 62132 858430 62160 858599
rect 62120 858424 62172 858430
rect 62120 858366 62172 858372
rect 62118 845608 62174 845617
rect 62118 845543 62174 845552
rect 62132 844626 62160 845543
rect 62120 844620 62172 844626
rect 62120 844562 62172 844568
rect 62118 832552 62174 832561
rect 62118 832487 62174 832496
rect 62132 832182 62160 832487
rect 55864 832176 55916 832182
rect 55864 832118 55916 832124
rect 62120 832176 62172 832182
rect 62120 832118 62172 832124
rect 55876 773022 55904 832118
rect 62118 819496 62174 819505
rect 62118 819431 62174 819440
rect 62132 818378 62160 819431
rect 62120 818372 62172 818378
rect 62120 818314 62172 818320
rect 62118 806576 62174 806585
rect 62118 806511 62174 806520
rect 62132 806002 62160 806511
rect 62120 805996 62172 806002
rect 62120 805938 62172 805944
rect 62118 793656 62174 793665
rect 62118 793591 62120 793600
rect 62172 793591 62174 793600
rect 62120 793562 62172 793568
rect 62118 780464 62174 780473
rect 62118 780399 62174 780408
rect 62132 780094 62160 780399
rect 56232 780088 56284 780094
rect 56232 780030 56284 780036
rect 62120 780088 62172 780094
rect 62120 780030 62172 780036
rect 55864 773016 55916 773022
rect 55864 772958 55916 772964
rect 56048 741124 56100 741130
rect 56048 741066 56100 741072
rect 55864 719160 55916 719166
rect 55864 719102 55916 719108
rect 54852 557592 54904 557598
rect 54852 557534 54904 557540
rect 54668 418192 54720 418198
rect 54668 418134 54720 418140
rect 54484 231804 54536 231810
rect 54484 231746 54536 231752
rect 53104 231668 53156 231674
rect 53104 231610 53156 231616
rect 54680 230081 54708 418134
rect 54864 408474 54892 557534
rect 54852 408468 54904 408474
rect 54852 408410 54904 408416
rect 54852 334008 54904 334014
rect 54852 333950 54904 333956
rect 54864 265577 54892 333950
rect 54850 265568 54906 265577
rect 54850 265503 54906 265512
rect 54666 230072 54722 230081
rect 54666 230007 54722 230016
rect 52090 227216 52146 227225
rect 52090 227151 52146 227160
rect 55876 226681 55904 719102
rect 56060 687274 56088 741066
rect 56244 731202 56272 780030
rect 62118 767408 62174 767417
rect 62118 767343 62120 767352
rect 62172 767343 62174 767352
rect 62120 767314 62172 767320
rect 62118 754352 62174 754361
rect 62118 754287 62174 754296
rect 62132 753574 62160 754287
rect 62120 753568 62172 753574
rect 62120 753510 62172 753516
rect 62118 741296 62174 741305
rect 62118 741231 62174 741240
rect 62132 741130 62160 741231
rect 62120 741124 62172 741130
rect 62120 741066 62172 741072
rect 56232 731196 56284 731202
rect 56232 731138 56284 731144
rect 62118 728240 62174 728249
rect 62118 728175 62174 728184
rect 62132 727326 62160 728175
rect 62120 727320 62172 727326
rect 62120 727262 62172 727268
rect 62118 715320 62174 715329
rect 62118 715255 62174 715264
rect 62132 714882 62160 715255
rect 62120 714876 62172 714882
rect 62120 714818 62172 714824
rect 62118 702264 62174 702273
rect 62118 702199 62174 702208
rect 62132 701078 62160 702199
rect 62120 701072 62172 701078
rect 62120 701014 62172 701020
rect 62118 689208 62174 689217
rect 62118 689143 62174 689152
rect 62132 688702 62160 689143
rect 62120 688696 62172 688702
rect 62120 688638 62172 688644
rect 56048 687268 56100 687274
rect 56048 687210 56100 687216
rect 62118 676152 62174 676161
rect 62118 676087 62174 676096
rect 62132 674898 62160 676087
rect 62120 674892 62172 674898
rect 62120 674834 62172 674840
rect 62118 663096 62174 663105
rect 62118 663031 62174 663040
rect 62132 662454 62160 663031
rect 62120 662448 62172 662454
rect 62120 662390 62172 662396
rect 62118 650040 62174 650049
rect 62118 649975 62174 649984
rect 62132 647902 62160 649975
rect 62120 647896 62172 647902
rect 62120 647838 62172 647844
rect 62118 637120 62174 637129
rect 62118 637055 62174 637064
rect 62132 636274 62160 637055
rect 62120 636268 62172 636274
rect 62120 636210 62172 636216
rect 62118 624064 62174 624073
rect 62118 623999 62174 624008
rect 62132 623830 62160 623999
rect 62120 623824 62172 623830
rect 62120 623766 62172 623772
rect 62118 611008 62174 611017
rect 62118 610943 62174 610952
rect 62132 609278 62160 610943
rect 62120 609272 62172 609278
rect 62120 609214 62172 609220
rect 62118 597952 62174 597961
rect 62118 597887 62174 597896
rect 62132 597582 62160 597887
rect 62120 597576 62172 597582
rect 62120 597518 62172 597524
rect 56048 590708 56100 590714
rect 56048 590650 56100 590656
rect 56060 277001 56088 590650
rect 62118 584896 62174 584905
rect 62118 584831 62174 584840
rect 62132 583778 62160 584831
rect 62120 583772 62172 583778
rect 62120 583714 62172 583720
rect 62118 571840 62174 571849
rect 62118 571775 62174 571784
rect 62132 571402 62160 571775
rect 62120 571396 62172 571402
rect 62120 571338 62172 571344
rect 62118 558784 62174 558793
rect 62118 558719 62174 558728
rect 62132 557598 62160 558719
rect 62120 557592 62172 557598
rect 62120 557534 62172 557540
rect 62118 545864 62174 545873
rect 62118 545799 62174 545808
rect 62132 545154 62160 545799
rect 62120 545148 62172 545154
rect 62120 545090 62172 545096
rect 62762 532808 62818 532817
rect 62762 532743 62818 532752
rect 62776 523734 62804 532743
rect 62764 523728 62816 523734
rect 62764 523670 62816 523676
rect 62118 519752 62174 519761
rect 62118 519687 62174 519696
rect 62132 518974 62160 519687
rect 62120 518968 62172 518974
rect 62120 518910 62172 518916
rect 62118 506696 62174 506705
rect 62118 506631 62174 506640
rect 62132 506530 62160 506631
rect 62120 506524 62172 506530
rect 62120 506466 62172 506472
rect 62118 493640 62174 493649
rect 62118 493575 62174 493584
rect 62132 491978 62160 493575
rect 62120 491972 62172 491978
rect 62120 491914 62172 491920
rect 62118 480584 62174 480593
rect 62118 480519 62174 480528
rect 62132 480282 62160 480519
rect 62120 480276 62172 480282
rect 62120 480218 62172 480224
rect 62118 467528 62174 467537
rect 62118 467463 62174 467472
rect 62132 466478 62160 467463
rect 62120 466472 62172 466478
rect 62120 466414 62172 466420
rect 62762 454608 62818 454617
rect 62762 454543 62818 454552
rect 62776 446418 62804 454543
rect 62764 446412 62816 446418
rect 62764 446354 62816 446360
rect 62118 441552 62174 441561
rect 62118 441487 62174 441496
rect 62132 434042 62160 441487
rect 62120 434036 62172 434042
rect 62120 433978 62172 433984
rect 62118 428496 62174 428505
rect 62118 428431 62174 428440
rect 62132 427854 62160 428431
rect 56232 427848 56284 427854
rect 56232 427790 56284 427796
rect 62120 427848 62172 427854
rect 62120 427790 62172 427796
rect 56244 343670 56272 427790
rect 62120 415472 62172 415478
rect 62118 415440 62120 415449
rect 62172 415440 62174 415449
rect 62118 415375 62174 415384
rect 62118 402384 62174 402393
rect 62118 402319 62174 402328
rect 62132 401674 62160 402319
rect 62120 401668 62172 401674
rect 62120 401610 62172 401616
rect 62118 389328 62174 389337
rect 62118 389263 62120 389272
rect 62172 389263 62174 389272
rect 62120 389234 62172 389240
rect 62118 376272 62174 376281
rect 62118 376207 62174 376216
rect 62132 375426 62160 376207
rect 62120 375420 62172 375426
rect 62120 375362 62172 375368
rect 62946 363352 63002 363361
rect 62946 363287 63002 363296
rect 62762 350296 62818 350305
rect 62762 350231 62818 350240
rect 56232 343664 56284 343670
rect 56232 343606 56284 343612
rect 62118 337240 62174 337249
rect 62118 337175 62174 337184
rect 62132 336802 62160 337175
rect 62120 336796 62172 336802
rect 62120 336738 62172 336744
rect 56232 332648 56284 332654
rect 56232 332590 56284 332596
rect 56244 278050 56272 332590
rect 62118 324184 62174 324193
rect 62118 324119 62174 324128
rect 62132 322998 62160 324119
rect 62120 322992 62172 322998
rect 62120 322934 62172 322940
rect 62776 318102 62804 350231
rect 62960 347070 62988 363287
rect 62948 347064 63000 347070
rect 62948 347006 63000 347012
rect 62764 318096 62816 318102
rect 62764 318038 62816 318044
rect 62118 311128 62174 311137
rect 62118 311063 62174 311072
rect 62132 310554 62160 311063
rect 62120 310548 62172 310554
rect 62120 310490 62172 310496
rect 62118 298208 62174 298217
rect 62118 298143 62120 298152
rect 62172 298143 62174 298152
rect 62120 298114 62172 298120
rect 64144 290012 64196 290018
rect 64144 289954 64196 289960
rect 61384 289876 61436 289882
rect 61384 289818 61436 289824
rect 61396 278322 61424 289818
rect 62762 285152 62818 285161
rect 62762 285087 62818 285096
rect 61384 278316 61436 278322
rect 61384 278258 61436 278264
rect 56232 278044 56284 278050
rect 56232 277986 56284 277992
rect 56046 276992 56102 277001
rect 56046 276927 56102 276936
rect 55862 226672 55918 226681
rect 55862 226607 55918 226616
rect 57888 225888 57940 225894
rect 57888 225830 57940 225836
rect 57244 224256 57296 224262
rect 57244 224198 57296 224204
rect 50342 223952 50398 223961
rect 50342 223887 50398 223896
rect 48964 219700 49016 219706
rect 48964 219642 49016 219648
rect 47950 218104 48006 218113
rect 47950 218039 48006 218048
rect 47584 204468 47636 204474
rect 47584 204410 47636 204416
rect 48976 204338 49004 219642
rect 48964 204332 49016 204338
rect 48964 204274 49016 204280
rect 44546 204096 44602 204105
rect 44546 204031 44602 204040
rect 44560 191826 44588 204031
rect 50356 203046 50384 223887
rect 50986 220008 51042 220017
rect 50986 219943 51042 219952
rect 51000 212702 51028 219943
rect 54206 219736 54262 219745
rect 54206 219671 54208 219680
rect 54260 219671 54262 219680
rect 54208 219642 54260 219648
rect 56508 218748 56560 218754
rect 56508 218690 56560 218696
rect 55680 218204 55732 218210
rect 55680 218146 55732 218152
rect 55692 217138 55720 218146
rect 56520 217138 56548 218690
rect 57256 218210 57284 224198
rect 57244 218204 57296 218210
rect 57244 218146 57296 218152
rect 57900 218074 57928 225830
rect 58990 225584 59046 225593
rect 58990 225519 59046 225528
rect 57336 218068 57388 218074
rect 57336 218010 57388 218016
rect 57888 218068 57940 218074
rect 57888 218010 57940 218016
rect 58164 218068 58216 218074
rect 58164 218010 58216 218016
rect 57348 217138 57376 218010
rect 58176 217138 58204 218010
rect 59004 217274 59032 225519
rect 62776 223038 62804 285087
rect 64156 278458 64184 289954
rect 499592 278730 499790 278746
rect 406936 278724 406988 278730
rect 406936 278666 406988 278672
rect 499580 278724 499790 278730
rect 499632 278718 499790 278724
rect 499580 278666 499632 278672
rect 64144 278452 64196 278458
rect 64144 278394 64196 278400
rect 65904 271182 65932 277780
rect 67022 277766 67588 277794
rect 65892 271176 65944 271182
rect 65892 271118 65944 271124
rect 67560 270094 67588 277766
rect 68204 275466 68232 277780
rect 68192 275460 68244 275466
rect 68192 275402 68244 275408
rect 67548 270088 67600 270094
rect 67548 270030 67600 270036
rect 69400 269822 69428 277780
rect 70596 275330 70624 277780
rect 70584 275324 70636 275330
rect 70584 275266 70636 275272
rect 71792 272950 71820 277780
rect 72988 273970 73016 277780
rect 72976 273964 73028 273970
rect 72976 273906 73028 273912
rect 71780 272944 71832 272950
rect 71780 272886 71832 272892
rect 74092 272542 74120 277780
rect 75302 277766 75868 277794
rect 76498 277766 77248 277794
rect 74080 272536 74132 272542
rect 74080 272478 74132 272484
rect 75840 269958 75868 277766
rect 75828 269952 75880 269958
rect 75828 269894 75880 269900
rect 69388 269816 69440 269822
rect 69388 269758 69440 269764
rect 77220 268802 77248 277766
rect 77680 274106 77708 277780
rect 77668 274100 77720 274106
rect 77668 274042 77720 274048
rect 78876 270366 78904 277780
rect 78864 270360 78916 270366
rect 78864 270302 78916 270308
rect 80072 270094 80100 277780
rect 81268 274990 81296 277780
rect 82386 277766 82768 277794
rect 83582 277766 84148 277794
rect 81256 274984 81308 274990
rect 81256 274926 81308 274932
rect 78220 270088 78272 270094
rect 78220 270030 78272 270036
rect 80060 270088 80112 270094
rect 80060 270030 80112 270036
rect 77208 268796 77260 268802
rect 77208 268738 77260 268744
rect 78232 267306 78260 270030
rect 82740 268394 82768 277766
rect 84120 269550 84148 277766
rect 84764 271318 84792 277780
rect 85960 275602 85988 277780
rect 85948 275596 86000 275602
rect 85948 275538 86000 275544
rect 86224 274984 86276 274990
rect 86224 274926 86276 274932
rect 84752 271312 84804 271318
rect 84752 271254 84804 271260
rect 84108 269544 84160 269550
rect 84108 269486 84160 269492
rect 82728 268388 82780 268394
rect 82728 268330 82780 268336
rect 78220 267300 78272 267306
rect 78220 267242 78272 267248
rect 86236 267170 86264 274926
rect 87156 268530 87184 277780
rect 88366 277766 88656 277794
rect 88628 271726 88656 277766
rect 89548 274718 89576 277780
rect 90666 277766 91048 277794
rect 89536 274712 89588 274718
rect 89536 274654 89588 274660
rect 88616 271720 88668 271726
rect 88616 271662 88668 271668
rect 87144 268524 87196 268530
rect 87144 268466 87196 268472
rect 86224 267164 86276 267170
rect 86224 267106 86276 267112
rect 91020 267034 91048 277766
rect 91848 272678 91876 277780
rect 92480 274712 92532 274718
rect 92480 274654 92532 274660
rect 91836 272672 91888 272678
rect 91836 272614 91888 272620
rect 92492 271454 92520 274654
rect 93044 274514 93072 277780
rect 93032 274508 93084 274514
rect 93032 274450 93084 274456
rect 92480 271448 92532 271454
rect 92480 271390 92532 271396
rect 94240 270230 94268 277780
rect 94228 270224 94280 270230
rect 94228 270166 94280 270172
rect 95436 268666 95464 277780
rect 96632 275738 96660 277780
rect 96620 275732 96672 275738
rect 96620 275674 96672 275680
rect 97736 272814 97764 277780
rect 97724 272808 97776 272814
rect 97724 272750 97776 272756
rect 98932 271590 98960 277780
rect 100142 277766 100708 277794
rect 98920 271584 98972 271590
rect 98920 271526 98972 271532
rect 95424 268660 95476 268666
rect 95424 268602 95476 268608
rect 100680 267442 100708 277766
rect 101324 271862 101352 277780
rect 102520 274242 102548 277780
rect 103716 275874 103744 277780
rect 103704 275868 103756 275874
rect 103704 275810 103756 275816
rect 102508 274236 102560 274242
rect 102508 274178 102560 274184
rect 101312 271856 101364 271862
rect 101312 271798 101364 271804
rect 104912 268938 104940 277780
rect 106016 274666 106044 277780
rect 107212 275194 107240 277780
rect 108422 277766 108988 277794
rect 109618 277766 110000 277794
rect 107200 275188 107252 275194
rect 107200 275130 107252 275136
rect 106016 274638 106320 274666
rect 104900 268932 104952 268938
rect 104900 268874 104952 268880
rect 106292 268802 106320 274638
rect 108960 270502 108988 277766
rect 109972 272950 110000 277766
rect 110800 276010 110828 277780
rect 110788 276004 110840 276010
rect 110788 275946 110840 275952
rect 111996 274378 112024 277780
rect 111984 274372 112036 274378
rect 111984 274314 112036 274320
rect 109684 272944 109736 272950
rect 109684 272886 109736 272892
rect 109960 272944 110012 272950
rect 109960 272886 110012 272892
rect 108948 270496 109000 270502
rect 108948 270438 109000 270444
rect 104900 268796 104952 268802
rect 104900 268738 104952 268744
rect 106280 268796 106332 268802
rect 106280 268738 106332 268744
rect 104912 267714 104940 268738
rect 104900 267708 104952 267714
rect 104900 267650 104952 267656
rect 100668 267436 100720 267442
rect 100668 267378 100720 267384
rect 91008 267028 91060 267034
rect 91008 266970 91060 266976
rect 109696 266762 109724 272886
rect 113192 272270 113220 277780
rect 113180 272264 113232 272270
rect 113180 272206 113232 272212
rect 114296 271046 114324 277780
rect 115506 277766 115796 277794
rect 114284 271040 114336 271046
rect 114284 270982 114336 270988
rect 115768 268258 115796 277766
rect 116688 274922 116716 277780
rect 117898 277766 118648 277794
rect 116676 274916 116728 274922
rect 116676 274858 116728 274864
rect 118620 269074 118648 277766
rect 119080 274514 119108 277780
rect 120276 274650 120304 277780
rect 119344 274644 119396 274650
rect 119344 274586 119396 274592
rect 120264 274644 120316 274650
rect 120264 274586 120316 274592
rect 119068 274508 119120 274514
rect 119068 274450 119120 274456
rect 118608 269068 118660 269074
rect 118608 269010 118660 269016
rect 115756 268252 115808 268258
rect 115756 268194 115808 268200
rect 119356 266898 119384 274586
rect 121380 273086 121408 277780
rect 122590 277766 122788 277794
rect 121368 273080 121420 273086
rect 121368 273022 121420 273028
rect 122760 269686 122788 277766
rect 123772 270910 123800 277780
rect 124968 273698 124996 277780
rect 126178 277766 126928 277794
rect 124956 273692 125008 273698
rect 124956 273634 125008 273640
rect 123760 270904 123812 270910
rect 123760 270846 123812 270852
rect 122748 269680 122800 269686
rect 122748 269622 122800 269628
rect 126900 269550 126928 277766
rect 127360 273222 127388 277780
rect 127348 273216 127400 273222
rect 127348 273158 127400 273164
rect 126704 269544 126756 269550
rect 126704 269486 126756 269492
rect 126888 269544 126940 269550
rect 126888 269486 126940 269492
rect 119344 266892 119396 266898
rect 119344 266834 119396 266840
rect 109684 266756 109736 266762
rect 109684 266698 109736 266704
rect 126716 266626 126744 269486
rect 128556 269278 128584 277780
rect 129384 277766 129674 277794
rect 129384 269414 129412 277766
rect 130856 273834 130884 277780
rect 132066 277766 132448 277794
rect 133262 277766 133828 277794
rect 130844 273828 130896 273834
rect 130844 273770 130896 273776
rect 129372 269408 129424 269414
rect 129372 269350 129424 269356
rect 128544 269272 128596 269278
rect 128544 269214 128596 269220
rect 132420 267578 132448 277766
rect 133800 270366 133828 277766
rect 134444 270774 134472 277780
rect 135260 275460 135312 275466
rect 135260 275402 135312 275408
rect 134432 270768 134484 270774
rect 134432 270710 134484 270716
rect 132592 270360 132644 270366
rect 132592 270302 132644 270308
rect 133788 270360 133840 270366
rect 133788 270302 133840 270308
rect 132408 267572 132460 267578
rect 132408 267514 132460 267520
rect 126704 266620 126756 266626
rect 126704 266562 126756 266568
rect 132604 266490 132632 270302
rect 135272 268122 135300 275402
rect 135640 274922 135668 277780
rect 135628 274916 135680 274922
rect 135628 274858 135680 274864
rect 136640 271176 136692 271182
rect 136640 271118 136692 271124
rect 135260 268116 135312 268122
rect 135260 268058 135312 268064
rect 132592 266484 132644 266490
rect 132592 266426 132644 266432
rect 136652 264316 136680 271118
rect 136836 270638 136864 277780
rect 137940 272406 137968 277780
rect 137928 272400 137980 272406
rect 137928 272342 137980 272348
rect 139136 271182 139164 277780
rect 139768 275324 139820 275330
rect 139768 275266 139820 275272
rect 139124 271176 139176 271182
rect 139124 271118 139176 271124
rect 136824 270632 136876 270638
rect 136824 270574 136876 270580
rect 138848 269816 138900 269822
rect 138848 269758 138900 269764
rect 138112 268116 138164 268122
rect 138112 268058 138164 268064
rect 137560 267776 137612 267782
rect 137560 267718 137612 267724
rect 137572 267306 137600 267718
rect 137376 267300 137428 267306
rect 137376 267242 137428 267248
rect 137560 267300 137612 267306
rect 137560 267242 137612 267248
rect 137388 264316 137416 267242
rect 138124 264316 138152 268058
rect 138860 264316 138888 269758
rect 139780 264330 139808 275266
rect 140332 274786 140360 277780
rect 141542 277766 141832 277794
rect 140320 274780 140372 274786
rect 140320 274722 140372 274728
rect 140780 274780 140832 274786
rect 140780 274722 140832 274728
rect 140044 271176 140096 271182
rect 140044 271118 140096 271124
rect 140056 267714 140084 271118
rect 140792 269822 140820 274722
rect 141804 273970 141832 277766
rect 142724 275058 142752 277780
rect 142712 275052 142764 275058
rect 142712 274994 142764 275000
rect 142988 274916 143040 274922
rect 142988 274858 143040 274864
rect 140964 273964 141016 273970
rect 140964 273906 141016 273912
rect 141792 273964 141844 273970
rect 141792 273906 141844 273912
rect 140780 269816 140832 269822
rect 140780 269758 140832 269764
rect 140044 267708 140096 267714
rect 140044 267650 140096 267656
rect 140320 266756 140372 266762
rect 140320 266698 140372 266704
rect 139610 264302 139808 264330
rect 140332 264316 140360 266698
rect 140976 264330 141004 273906
rect 142160 272536 142212 272542
rect 142160 272478 142212 272484
rect 141792 269952 141844 269958
rect 141792 269894 141844 269900
rect 140976 264302 141082 264330
rect 141804 264316 141832 269894
rect 142172 264330 142200 272478
rect 143000 272270 143028 274858
rect 143632 274100 143684 274106
rect 143632 274042 143684 274048
rect 142804 272264 142856 272270
rect 142804 272206 142856 272212
rect 142988 272264 143040 272270
rect 142988 272206 143040 272212
rect 142816 267714 142844 272206
rect 143448 267844 143500 267850
rect 143448 267786 143500 267792
rect 142804 267708 142856 267714
rect 142804 267650 142856 267656
rect 143460 267306 143488 267786
rect 143264 267300 143316 267306
rect 143264 267242 143316 267248
rect 143448 267300 143500 267306
rect 143448 267242 143500 267248
rect 142172 264302 142554 264330
rect 143276 264316 143304 267242
rect 143644 264330 143672 274042
rect 143920 269958 143948 277780
rect 145024 271182 145052 277780
rect 145564 271720 145616 271726
rect 145564 271662 145616 271668
rect 145012 271176 145064 271182
rect 145012 271118 145064 271124
rect 144460 270088 144512 270094
rect 144460 270030 144512 270036
rect 143908 269952 143960 269958
rect 143908 269894 143960 269900
rect 144472 264330 144500 270030
rect 145576 266898 145604 271662
rect 146220 267170 146248 277780
rect 147416 277394 147444 277780
rect 148626 277766 148916 277794
rect 147416 277366 147536 277394
rect 146944 268388 146996 268394
rect 146944 268330 146996 268336
rect 145932 267164 145984 267170
rect 145932 267106 145984 267112
rect 146208 267164 146260 267170
rect 146208 267106 146260 267112
rect 145564 266892 145616 266898
rect 145564 266834 145616 266840
rect 145472 266484 145524 266490
rect 145472 266426 145524 266432
rect 143644 264302 144026 264330
rect 144472 264302 144762 264330
rect 145484 264316 145512 266426
rect 145944 264330 145972 267106
rect 145944 264302 146234 264330
rect 146956 264316 146984 268330
rect 147508 268122 147536 277366
rect 147680 271312 147732 271318
rect 147680 271254 147732 271260
rect 147496 268116 147548 268122
rect 147496 268058 147548 268064
rect 147692 264316 147720 271254
rect 148888 268394 148916 277766
rect 149060 275596 149112 275602
rect 149060 275538 149112 275544
rect 148876 268388 148928 268394
rect 148876 268330 148928 268336
rect 148416 266620 148468 266626
rect 148416 266562 148468 266568
rect 148428 264316 148456 266562
rect 149072 264330 149100 275538
rect 149808 275330 149836 277780
rect 149796 275324 149848 275330
rect 149796 275266 149848 275272
rect 151004 274922 151032 277780
rect 152200 275194 152228 277780
rect 153304 275602 153332 277780
rect 153844 275732 153896 275738
rect 153844 275674 153896 275680
rect 153292 275596 153344 275602
rect 153292 275538 153344 275544
rect 151176 275188 151228 275194
rect 151176 275130 151228 275136
rect 152188 275188 152240 275194
rect 152188 275130 152240 275136
rect 150992 274916 151044 274922
rect 150992 274858 151044 274864
rect 150440 271448 150492 271454
rect 150440 271390 150492 271396
rect 149888 268524 149940 268530
rect 149888 268466 149940 268472
rect 149072 264302 149178 264330
rect 149900 264316 149928 268466
rect 150452 264330 150480 271390
rect 151188 266626 151216 275130
rect 152648 274916 152700 274922
rect 152648 274858 152700 274864
rect 152372 272672 152424 272678
rect 152372 272614 152424 272620
rect 152384 267734 152412 272614
rect 152660 270094 152688 274858
rect 153568 270224 153620 270230
rect 153568 270166 153620 270172
rect 152648 270088 152700 270094
rect 152648 270030 152700 270036
rect 152384 267706 152504 267734
rect 152096 267028 152148 267034
rect 152096 266970 152148 266976
rect 151360 266892 151412 266898
rect 151360 266834 151412 266840
rect 151176 266620 151228 266626
rect 151176 266562 151228 266568
rect 150452 264302 150650 264330
rect 151372 264316 151400 266834
rect 152108 264316 152136 266970
rect 152476 264330 152504 267706
rect 152476 264302 152858 264330
rect 153580 264316 153608 270166
rect 153856 266422 153884 275674
rect 154500 272542 154528 277780
rect 155408 272808 155460 272814
rect 155408 272750 155460 272756
rect 154488 272536 154540 272542
rect 154488 272478 154540 272484
rect 155040 268660 155092 268666
rect 155040 268602 155092 268608
rect 154304 266756 154356 266762
rect 154304 266698 154356 266704
rect 153844 266416 153896 266422
rect 153844 266358 153896 266364
rect 154316 264316 154344 266698
rect 155052 264316 155080 268602
rect 155420 264330 155448 272750
rect 155696 271318 155724 277780
rect 156420 276004 156472 276010
rect 156420 275946 156472 275952
rect 156236 271584 156288 271590
rect 156236 271526 156288 271532
rect 155684 271312 155736 271318
rect 155684 271254 155736 271260
rect 156248 267734 156276 271526
rect 156432 267734 156460 275946
rect 156892 275466 156920 277780
rect 156880 275460 156932 275466
rect 156880 275402 156932 275408
rect 156604 274780 156656 274786
rect 156604 274722 156656 274728
rect 156616 271454 156644 274722
rect 158088 274106 158116 277780
rect 159088 274236 159140 274242
rect 159088 274178 159140 274184
rect 158076 274100 158128 274106
rect 158076 274042 158128 274048
rect 157984 273692 158036 273698
rect 157984 273634 158036 273640
rect 157616 271856 157668 271862
rect 157616 271798 157668 271804
rect 156604 271448 156656 271454
rect 156604 271390 156656 271396
rect 156248 267706 156368 267734
rect 156432 267706 156552 267734
rect 156144 266416 156196 266422
rect 156144 266358 156196 266364
rect 156156 264330 156184 266358
rect 156340 264602 156368 267706
rect 156524 267034 156552 267706
rect 156512 267028 156564 267034
rect 156512 266970 156564 266976
rect 156340 264574 156920 264602
rect 156892 264330 156920 264574
rect 157628 264330 157656 271798
rect 157996 266898 158024 273634
rect 158720 267436 158772 267442
rect 158720 267378 158772 267384
rect 157984 266892 158036 266898
rect 157984 266834 158036 266840
rect 155420 264302 155802 264330
rect 156156 264302 156538 264330
rect 156892 264302 157274 264330
rect 157628 264302 158010 264330
rect 158732 264316 158760 267378
rect 159100 264330 159128 274178
rect 159284 272678 159312 277780
rect 160480 275738 160508 277780
rect 160652 275868 160704 275874
rect 160652 275810 160704 275816
rect 160468 275732 160520 275738
rect 160468 275674 160520 275680
rect 159272 272672 159324 272678
rect 159272 272614 159324 272620
rect 160192 268932 160244 268938
rect 160192 268874 160244 268880
rect 159100 264302 159482 264330
rect 160204 264316 160232 268874
rect 160664 264330 160692 275810
rect 161584 274718 161612 277780
rect 162584 275188 162636 275194
rect 162584 275130 162636 275136
rect 161572 274712 161624 274718
rect 161572 274654 161624 274660
rect 161434 274644 161486 274650
rect 161434 274586 161486 274592
rect 161446 274530 161474 274586
rect 161446 274502 161520 274530
rect 161492 273698 161520 274502
rect 161480 273692 161532 273698
rect 161480 273634 161532 273640
rect 162400 270496 162452 270502
rect 162400 270438 162452 270444
rect 161664 268796 161716 268802
rect 161664 268738 161716 268744
rect 160664 264302 160954 264330
rect 161676 264316 161704 268738
rect 162412 264316 162440 270438
rect 162596 268666 162624 275130
rect 162584 268660 162636 268666
rect 162584 268602 162636 268608
rect 162780 268530 162808 277780
rect 163976 274718 164004 277780
rect 163688 274712 163740 274718
rect 163688 274654 163740 274660
rect 163964 274712 164016 274718
rect 163964 274654 164016 274660
rect 163320 272944 163372 272950
rect 163320 272886 163372 272892
rect 162952 269272 163004 269278
rect 162952 269214 163004 269220
rect 162768 268524 162820 268530
rect 162768 268466 162820 268472
rect 162964 267442 162992 269214
rect 163332 267734 163360 272886
rect 163700 270230 163728 274654
rect 164240 274372 164292 274378
rect 164240 274314 164292 274320
rect 163688 270224 163740 270230
rect 163688 270166 163740 270172
rect 163332 267706 163544 267734
rect 162952 267436 163004 267442
rect 162952 267378 163004 267384
rect 163136 266620 163188 266626
rect 163136 266562 163188 266568
rect 163148 264316 163176 266562
rect 163516 264330 163544 267706
rect 164252 264330 164280 274314
rect 165172 271862 165200 277780
rect 166172 275460 166224 275466
rect 166172 275402 166224 275408
rect 165160 271856 165212 271862
rect 165160 271798 165212 271804
rect 164884 271040 164936 271046
rect 164884 270982 164936 270988
rect 164896 266422 164924 270982
rect 166184 268802 166212 275402
rect 166368 274242 166396 277780
rect 167564 275466 167592 277780
rect 167552 275460 167604 275466
rect 167552 275402 167604 275408
rect 167828 274712 167880 274718
rect 167828 274654 167880 274660
rect 166356 274236 166408 274242
rect 166356 274178 166408 274184
rect 167460 272264 167512 272270
rect 167460 272206 167512 272212
rect 166172 268796 166224 268802
rect 166172 268738 166224 268744
rect 166816 268252 166868 268258
rect 166816 268194 166868 268200
rect 166080 267708 166132 267714
rect 166080 267650 166132 267656
rect 165344 267028 165396 267034
rect 165344 266970 165396 266976
rect 164884 266416 164936 266422
rect 164884 266358 164936 266364
rect 163516 264302 163898 264330
rect 164252 264302 164634 264330
rect 165356 264316 165384 266970
rect 166092 264316 166120 267650
rect 166828 264316 166856 268194
rect 167472 267734 167500 272206
rect 167840 267734 167868 274654
rect 168472 274508 168524 274514
rect 168472 274450 168524 274456
rect 168484 267734 168512 274450
rect 168668 272814 168696 277780
rect 169878 277766 170168 277794
rect 169760 275052 169812 275058
rect 169760 274994 169812 275000
rect 169772 274514 169800 274994
rect 169760 274508 169812 274514
rect 169760 274450 169812 274456
rect 169944 273692 169996 273698
rect 169944 273634 169996 273640
rect 168656 272808 168708 272814
rect 168656 272750 168708 272756
rect 169760 269068 169812 269074
rect 169760 269010 169812 269016
rect 167472 267706 167776 267734
rect 167840 267706 167960 267734
rect 168484 267706 168696 267734
rect 167552 266416 167604 266422
rect 167552 266358 167604 266364
rect 167564 264316 167592 266358
rect 167748 264466 167776 267706
rect 167932 267034 167960 267706
rect 167920 267028 167972 267034
rect 167920 266970 167972 266976
rect 167748 264438 167960 264466
rect 167932 264330 167960 264438
rect 168668 264330 168696 267706
rect 167932 264302 168314 264330
rect 168668 264302 169050 264330
rect 169772 264316 169800 269010
rect 169956 267734 169984 273634
rect 170140 271590 170168 277766
rect 171060 276010 171088 277780
rect 172270 277766 172468 277794
rect 173466 277766 173848 277794
rect 171048 276004 171100 276010
rect 171048 275946 171100 275952
rect 171600 273080 171652 273086
rect 171600 273022 171652 273028
rect 170128 271584 170180 271590
rect 170128 271526 170180 271532
rect 171232 269680 171284 269686
rect 171232 269622 171284 269628
rect 169956 267706 170168 267734
rect 170140 264330 170168 267706
rect 170140 264302 170522 264330
rect 171244 264316 171272 269622
rect 171612 264330 171640 273022
rect 172440 269686 172468 277766
rect 172704 270904 172756 270910
rect 172704 270846 172756 270852
rect 172428 269680 172480 269686
rect 172428 269622 172480 269628
rect 171612 264302 171994 264330
rect 172716 264316 172744 270846
rect 173820 270502 173848 277766
rect 174648 275874 174676 277780
rect 175844 276010 175872 277780
rect 175648 276004 175700 276010
rect 175648 275946 175700 275952
rect 175832 276004 175884 276010
rect 175832 275946 175884 275952
rect 175660 275890 175688 275946
rect 174636 275868 174688 275874
rect 175660 275862 175964 275890
rect 174636 275810 174688 275816
rect 174452 275732 174504 275738
rect 174452 275674 174504 275680
rect 174268 273216 174320 273222
rect 174268 273158 174320 273164
rect 173808 270496 173860 270502
rect 173808 270438 173860 270444
rect 173440 269544 173492 269550
rect 173440 269486 173492 269492
rect 173452 264316 173480 269486
rect 174280 267734 174308 273158
rect 174464 273086 174492 275674
rect 174452 273080 174504 273086
rect 174452 273022 174504 273028
rect 174636 270632 174688 270638
rect 174636 270574 174688 270580
rect 174648 267734 174676 270574
rect 175648 269408 175700 269414
rect 175648 269350 175700 269356
rect 174280 267706 174584 267734
rect 174648 267706 174768 267734
rect 173900 267300 173952 267306
rect 173900 267242 173952 267248
rect 173912 266762 173940 267242
rect 174176 266892 174228 266898
rect 174176 266834 174228 266840
rect 173900 266756 173952 266762
rect 173900 266698 173952 266704
rect 174188 264316 174216 266834
rect 174556 264330 174584 267706
rect 174740 266422 174768 267706
rect 174728 266416 174780 266422
rect 174728 266358 174780 266364
rect 174556 264302 174938 264330
rect 175660 264316 175688 269350
rect 175936 267442 175964 275862
rect 176752 273828 176804 273834
rect 176752 273770 176804 273776
rect 175924 267436 175976 267442
rect 175924 267378 175976 267384
rect 176384 267300 176436 267306
rect 176384 267242 176436 267248
rect 176396 264316 176424 267242
rect 176764 264330 176792 273770
rect 176948 270502 176976 277780
rect 177396 276004 177448 276010
rect 177396 275946 177448 275952
rect 177408 274378 177436 275946
rect 178144 274990 178172 277780
rect 178132 274984 178184 274990
rect 178132 274926 178184 274932
rect 177396 274372 177448 274378
rect 177396 274314 177448 274320
rect 179340 271726 179368 277780
rect 180550 277766 180748 277794
rect 180064 274984 180116 274990
rect 180064 274926 180116 274932
rect 179328 271720 179380 271726
rect 179328 271662 179380 271668
rect 178960 270768 179012 270774
rect 178960 270710 179012 270716
rect 176936 270496 176988 270502
rect 176936 270438 176988 270444
rect 177580 270360 177632 270366
rect 177580 270302 177632 270308
rect 177592 264330 177620 270302
rect 178592 267572 178644 267578
rect 178592 267514 178644 267520
rect 176764 264302 177146 264330
rect 177592 264302 177882 264330
rect 178604 264316 178632 267514
rect 178972 264330 179000 270710
rect 180076 267578 180104 274926
rect 180720 274666 180748 277766
rect 181732 275738 181760 277780
rect 182942 277766 183508 277794
rect 184138 277766 184520 277794
rect 181720 275732 181772 275738
rect 181720 275674 181772 275680
rect 180720 274638 180840 274666
rect 180812 272950 180840 274638
rect 180800 272944 180852 272950
rect 180800 272886 180852 272892
rect 181168 272400 181220 272406
rect 181168 272342 181220 272348
rect 180800 271448 180852 271454
rect 180800 271390 180852 271396
rect 180064 267572 180116 267578
rect 180064 267514 180116 267520
rect 180064 266416 180116 266422
rect 180064 266358 180116 266364
rect 178972 264302 179354 264330
rect 180076 264316 180104 266358
rect 180812 264316 180840 271390
rect 181180 264330 181208 272342
rect 182272 269816 182324 269822
rect 182272 269758 182324 269764
rect 181180 264302 181562 264330
rect 182284 264316 182312 269758
rect 183480 269550 183508 277766
rect 184492 273970 184520 277766
rect 184756 275324 184808 275330
rect 184756 275266 184808 275272
rect 183744 273964 183796 273970
rect 183744 273906 183796 273912
rect 184480 273964 184532 273970
rect 184480 273906 184532 273912
rect 183468 269544 183520 269550
rect 183468 269486 183520 269492
rect 183008 266756 183060 266762
rect 183008 266698 183060 266704
rect 183020 264316 183048 266698
rect 183756 264316 183784 273906
rect 184768 269958 184796 275266
rect 185228 274718 185256 277780
rect 185768 275596 185820 275602
rect 185768 275538 185820 275544
rect 185216 274712 185268 274718
rect 185216 274654 185268 274660
rect 184940 274508 184992 274514
rect 184940 274450 184992 274456
rect 184480 269952 184532 269958
rect 184480 269894 184532 269900
rect 184756 269952 184808 269958
rect 184756 269894 184808 269900
rect 184492 264316 184520 269894
rect 184952 264330 184980 274450
rect 185584 271176 185636 271182
rect 185584 271118 185636 271124
rect 185596 264330 185624 271118
rect 185780 271046 185808 275538
rect 186424 274854 186452 277780
rect 187620 277394 187648 277780
rect 187528 277366 187648 277394
rect 186412 274848 186464 274854
rect 186412 274790 186464 274796
rect 186964 274712 187016 274718
rect 186964 274654 187016 274660
rect 185768 271040 185820 271046
rect 185768 270982 185820 270988
rect 186688 268116 186740 268122
rect 186688 268058 186740 268064
rect 184952 264302 185242 264330
rect 185596 264302 185978 264330
rect 186700 264316 186728 268058
rect 186976 267170 187004 274654
rect 187528 268938 187556 277366
rect 188816 275330 188844 277780
rect 190026 277766 190408 277794
rect 191222 277766 191788 277794
rect 188804 275324 188856 275330
rect 188804 275266 188856 275272
rect 188436 274848 188488 274854
rect 188436 274790 188488 274796
rect 187516 268932 187568 268938
rect 187516 268874 187568 268880
rect 188448 268394 188476 274790
rect 188896 270088 188948 270094
rect 188896 270030 188948 270036
rect 188160 268388 188212 268394
rect 188160 268330 188212 268336
rect 188436 268388 188488 268394
rect 188436 268330 188488 268336
rect 187424 267300 187476 267306
rect 187424 267242 187476 267248
rect 186964 267164 187016 267170
rect 186964 267106 187016 267112
rect 187436 264316 187464 267242
rect 188172 264316 188200 268330
rect 188908 264316 188936 270030
rect 189632 269952 189684 269958
rect 189632 269894 189684 269900
rect 189644 264316 189672 269894
rect 190380 268666 190408 277766
rect 190736 272536 190788 272542
rect 190736 272478 190788 272484
rect 190092 268660 190144 268666
rect 190092 268602 190144 268608
rect 190368 268660 190420 268666
rect 190368 268602 190420 268608
rect 190104 264330 190132 268602
rect 190748 264330 190776 272478
rect 191760 269822 191788 277766
rect 192312 277394 192340 277780
rect 192220 277366 192340 277394
rect 192220 271182 192248 277366
rect 193220 274100 193272 274106
rect 193220 274042 193272 274048
rect 192392 271312 192444 271318
rect 192392 271254 192444 271260
rect 192208 271176 192260 271182
rect 192208 271118 192260 271124
rect 192208 271040 192260 271046
rect 192208 270982 192260 270988
rect 191748 269816 191800 269822
rect 191748 269758 191800 269764
rect 192220 264330 192248 270982
rect 190104 264302 190394 264330
rect 190748 264302 191130 264330
rect 191866 264302 192248 264330
rect 192404 264330 192432 271254
rect 193232 264330 193260 274042
rect 193508 271318 193536 277780
rect 194704 277394 194732 277780
rect 194612 277366 194732 277394
rect 195716 277766 195914 277794
rect 193496 271312 193548 271318
rect 193496 271254 193548 271260
rect 194612 269958 194640 277366
rect 195716 272678 195744 277766
rect 196164 273080 196216 273086
rect 196164 273022 196216 273028
rect 194784 272672 194836 272678
rect 194784 272614 194836 272620
rect 195704 272672 195756 272678
rect 195704 272614 195756 272620
rect 194600 269952 194652 269958
rect 194600 269894 194652 269900
rect 194508 269544 194560 269550
rect 194508 269486 194560 269492
rect 194048 268796 194100 268802
rect 194048 268738 194100 268744
rect 192404 264302 192602 264330
rect 193232 264302 193338 264330
rect 194060 264316 194088 268738
rect 194520 267306 194548 269486
rect 194508 267300 194560 267306
rect 194508 267242 194560 267248
rect 194796 264316 194824 272614
rect 195520 270224 195572 270230
rect 195520 270166 195572 270172
rect 195532 264316 195560 270166
rect 196176 264330 196204 273022
rect 197096 272542 197124 277780
rect 197544 275868 197596 275874
rect 197544 275810 197596 275816
rect 197084 272536 197136 272542
rect 197084 272478 197136 272484
rect 197360 271856 197412 271862
rect 197360 271798 197412 271804
rect 196992 268524 197044 268530
rect 196992 268466 197044 268472
rect 196176 264302 196282 264330
rect 197004 264316 197032 268466
rect 197372 264330 197400 271798
rect 197556 270230 197584 275810
rect 198292 274106 198320 277780
rect 199488 275602 199516 277780
rect 199476 275596 199528 275602
rect 199476 275538 199528 275544
rect 200028 275460 200080 275466
rect 200028 275402 200080 275408
rect 200040 274530 200068 275402
rect 200040 274502 200252 274530
rect 198924 274236 198976 274242
rect 198924 274178 198976 274184
rect 198280 274100 198332 274106
rect 198280 274042 198332 274048
rect 198740 272808 198792 272814
rect 198740 272750 198792 272756
rect 197544 270224 197596 270230
rect 197544 270166 197596 270172
rect 198464 267028 198516 267034
rect 198464 266970 198516 266976
rect 197372 264302 197754 264330
rect 198476 264316 198504 266970
rect 198752 265946 198780 272750
rect 198740 265940 198792 265946
rect 198740 265882 198792 265888
rect 198936 264330 198964 274178
rect 200224 267734 200252 274502
rect 200592 274242 200620 277780
rect 200580 274236 200632 274242
rect 200580 274178 200632 274184
rect 201040 271584 201092 271590
rect 201040 271526 201092 271532
rect 200224 267706 200344 267734
rect 199660 265940 199712 265946
rect 199660 265882 199712 265888
rect 199672 264330 199700 265882
rect 200316 264330 200344 267706
rect 201052 264330 201080 271526
rect 201788 271454 201816 277780
rect 201776 271448 201828 271454
rect 201776 271390 201828 271396
rect 202984 270094 203012 277780
rect 203904 277766 204194 277794
rect 205390 277766 205588 277794
rect 203616 270496 203668 270502
rect 203616 270438 203668 270444
rect 202972 270088 203024 270094
rect 202972 270030 203024 270036
rect 202144 269680 202196 269686
rect 202144 269622 202196 269628
rect 198936 264302 199226 264330
rect 199672 264302 199962 264330
rect 200316 264302 200698 264330
rect 201052 264302 201434 264330
rect 202156 264316 202184 269622
rect 202880 267436 202932 267442
rect 202880 267378 202932 267384
rect 202892 264316 202920 267378
rect 203628 264316 203656 270438
rect 203904 268802 203932 277766
rect 204260 274372 204312 274378
rect 204260 274314 204312 274320
rect 203892 268796 203944 268802
rect 203892 268738 203944 268744
rect 204076 268660 204128 268666
rect 204076 268602 204128 268608
rect 204088 267442 204116 268602
rect 204076 267436 204128 267442
rect 204076 267378 204128 267384
rect 204272 264330 204300 274314
rect 204904 271720 204956 271726
rect 204904 271662 204956 271668
rect 204916 266422 204944 271662
rect 205560 270230 205588 277766
rect 206572 273970 206600 277780
rect 207020 275732 207072 275738
rect 207020 275674 207072 275680
rect 206284 273964 206336 273970
rect 206284 273906 206336 273912
rect 206560 273964 206612 273970
rect 206560 273906 206612 273912
rect 205824 270360 205876 270366
rect 205824 270302 205876 270308
rect 205088 270224 205140 270230
rect 205088 270166 205140 270172
rect 205548 270224 205600 270230
rect 205548 270166 205600 270172
rect 204904 266416 204956 266422
rect 204904 266358 204956 266364
rect 204272 264302 204378 264330
rect 205100 264316 205128 270166
rect 205836 264316 205864 270302
rect 206296 266762 206324 273906
rect 207032 270502 207060 275674
rect 207768 275466 207796 277780
rect 207756 275460 207808 275466
rect 207756 275402 207808 275408
rect 207480 272944 207532 272950
rect 207480 272886 207532 272892
rect 207020 270496 207072 270502
rect 207020 270438 207072 270444
rect 207492 267734 207520 272886
rect 208492 268932 208544 268938
rect 208492 268874 208544 268880
rect 207492 267706 207704 267734
rect 207296 267572 207348 267578
rect 207296 267514 207348 267520
rect 206284 266756 206336 266762
rect 206284 266698 206336 266704
rect 206560 266416 206612 266422
rect 206560 266358 206612 266364
rect 206572 264316 206600 266358
rect 207308 264316 207336 267514
rect 207676 264330 207704 267706
rect 208504 266490 208532 268874
rect 208872 268530 208900 277780
rect 210068 272678 210096 277780
rect 210976 275596 211028 275602
rect 210976 275538 211028 275544
rect 210608 272808 210660 272814
rect 210608 272750 210660 272756
rect 210056 272672 210108 272678
rect 210056 272614 210108 272620
rect 209504 270496 209556 270502
rect 209504 270438 209556 270444
rect 208860 268524 208912 268530
rect 208860 268466 208912 268472
rect 208768 267300 208820 267306
rect 208768 267242 208820 267248
rect 208492 266484 208544 266490
rect 208492 266426 208544 266432
rect 207676 264302 208058 264330
rect 208780 264316 208808 267242
rect 209516 264316 209544 270438
rect 210240 266756 210292 266762
rect 210240 266698 210292 266704
rect 210252 264316 210280 266698
rect 210620 266626 210648 272750
rect 210988 268394 211016 275538
rect 211264 275262 211292 277780
rect 212276 277766 212474 277794
rect 211252 275256 211304 275262
rect 211252 275198 211304 275204
rect 212276 270366 212304 277766
rect 212448 275256 212500 275262
rect 212448 275198 212500 275204
rect 212264 270360 212316 270366
rect 212264 270302 212316 270308
rect 211160 268796 211212 268802
rect 211160 268738 211212 268744
rect 210976 268388 211028 268394
rect 210976 268330 211028 268336
rect 210976 268252 211028 268258
rect 210976 268194 211028 268200
rect 210608 266620 210660 266626
rect 210608 266562 210660 266568
rect 210988 264316 211016 268194
rect 211172 267170 211200 268738
rect 211160 267164 211212 267170
rect 211160 267106 211212 267112
rect 212460 267034 212488 275198
rect 213184 274236 213236 274242
rect 213184 274178 213236 274184
rect 213196 267714 213224 274178
rect 213656 271590 213684 277780
rect 213920 275120 213972 275126
rect 213920 275062 213972 275068
rect 213644 271584 213696 271590
rect 213644 271526 213696 271532
rect 213184 267708 213236 267714
rect 213184 267650 213236 267656
rect 213184 267436 213236 267442
rect 213184 267378 213236 267384
rect 211712 267028 211764 267034
rect 211712 266970 211764 266976
rect 212448 267028 212500 267034
rect 212448 266970 212500 266976
rect 211724 264316 211752 266970
rect 212448 266484 212500 266490
rect 212448 266426 212500 266432
rect 212460 264316 212488 266426
rect 213196 264316 213224 267378
rect 213932 264316 213960 275062
rect 214852 274990 214880 277780
rect 214840 274984 214892 274990
rect 214840 274926 214892 274932
rect 215760 271312 215812 271318
rect 215760 271254 215812 271260
rect 215300 271176 215352 271182
rect 215300 271118 215352 271124
rect 214656 269816 214708 269822
rect 214656 269758 214708 269764
rect 214668 264316 214696 269758
rect 215312 264330 215340 271118
rect 215772 264330 215800 271254
rect 215956 271182 215984 277780
rect 217152 275942 217180 277780
rect 217140 275936 217192 275942
rect 217140 275878 217192 275884
rect 218348 275602 218376 277780
rect 219544 277394 219572 277780
rect 219544 277366 219664 277394
rect 218520 275936 218572 275942
rect 218520 275878 218572 275884
rect 218336 275596 218388 275602
rect 218336 275538 218388 275544
rect 216680 275460 216732 275466
rect 216680 275402 216732 275408
rect 215944 271176 215996 271182
rect 215944 271118 215996 271124
rect 216692 270502 216720 275402
rect 217968 274100 218020 274106
rect 217968 274042 218020 274048
rect 217980 273986 218008 274042
rect 217980 273958 218100 273986
rect 216680 270496 216732 270502
rect 216680 270438 216732 270444
rect 216864 269952 216916 269958
rect 216864 269894 216916 269900
rect 215312 264302 215418 264330
rect 215772 264302 216154 264330
rect 216876 264316 216904 269894
rect 217600 266620 217652 266626
rect 217600 266562 217652 266568
rect 217612 264316 217640 266562
rect 218072 265946 218100 273958
rect 218532 272542 218560 275878
rect 218520 272536 218572 272542
rect 218520 272478 218572 272484
rect 218244 272400 218296 272406
rect 218244 272342 218296 272348
rect 218060 265940 218112 265946
rect 218060 265882 218112 265888
rect 218256 264330 218284 272342
rect 219440 270360 219492 270366
rect 219440 270302 219492 270308
rect 219452 266422 219480 270302
rect 219636 269822 219664 277366
rect 219624 269816 219676 269822
rect 219624 269758 219676 269764
rect 220740 268394 220768 277780
rect 221936 275602 221964 277780
rect 221924 275596 221976 275602
rect 221924 275538 221976 275544
rect 222844 275460 222896 275466
rect 222844 275402 222896 275408
rect 221464 274984 221516 274990
rect 221464 274926 221516 274932
rect 221004 271448 221056 271454
rect 221004 271390 221056 271396
rect 219808 268388 219860 268394
rect 219808 268330 219860 268336
rect 220728 268388 220780 268394
rect 220728 268330 220780 268336
rect 219440 266416 219492 266422
rect 219440 266358 219492 266364
rect 218796 265940 218848 265946
rect 218796 265882 218848 265888
rect 218808 264330 218836 265882
rect 218256 264302 218362 264330
rect 218808 264302 219098 264330
rect 219820 264316 219848 268330
rect 220544 267708 220596 267714
rect 220544 267650 220596 267656
rect 220556 264316 220584 267650
rect 221016 264330 221044 271390
rect 221476 269958 221504 274926
rect 222016 270088 222068 270094
rect 222016 270030 222068 270036
rect 221464 269952 221516 269958
rect 221464 269894 221516 269900
rect 221016 264302 221306 264330
rect 222028 264316 222056 270030
rect 222856 267442 222884 275402
rect 223132 271318 223160 277780
rect 224236 273970 224264 277780
rect 223856 273964 223908 273970
rect 223856 273906 223908 273912
rect 224224 273964 224276 273970
rect 224224 273906 224276 273912
rect 223120 271312 223172 271318
rect 223120 271254 223172 271260
rect 223488 270224 223540 270230
rect 223488 270166 223540 270172
rect 222844 267436 222896 267442
rect 222844 267378 222896 267384
rect 222752 267164 222804 267170
rect 222752 267106 222804 267112
rect 222764 264316 222792 267106
rect 223500 264316 223528 270166
rect 223868 264330 223896 273906
rect 224960 270496 225012 270502
rect 224960 270438 225012 270444
rect 223868 264302 224250 264330
rect 224972 264316 225000 270438
rect 225432 269074 225460 277780
rect 226432 272672 226484 272678
rect 226432 272614 226484 272620
rect 225420 269068 225472 269074
rect 225420 269010 225472 269016
rect 225696 268524 225748 268530
rect 225696 268466 225748 268472
rect 225708 264316 225736 268466
rect 226444 264316 226472 272614
rect 226628 270094 226656 277780
rect 227824 275330 227852 277780
rect 228456 275596 228508 275602
rect 228456 275538 228508 275544
rect 227812 275324 227864 275330
rect 227812 275266 227864 275272
rect 228272 271584 228324 271590
rect 228272 271526 228324 271532
rect 226616 270088 226668 270094
rect 226616 270030 226668 270036
rect 227628 269068 227680 269074
rect 227628 269010 227680 269016
rect 227640 267034 227668 269010
rect 227168 267028 227220 267034
rect 227168 266970 227220 266976
rect 227628 267028 227680 267034
rect 227628 266970 227680 266976
rect 227180 264316 227208 266970
rect 227904 266416 227956 266422
rect 227904 266358 227956 266364
rect 227916 264316 227944 266358
rect 228284 264330 228312 271526
rect 228468 267306 228496 275538
rect 229020 271590 229048 277780
rect 230230 277766 230428 277794
rect 229008 271584 229060 271590
rect 229008 271526 229060 271532
rect 229744 271176 229796 271182
rect 229744 271118 229796 271124
rect 229376 269952 229428 269958
rect 229376 269894 229428 269900
rect 228456 267300 228508 267306
rect 228456 267242 228508 267248
rect 228284 264302 228666 264330
rect 229388 264316 229416 269894
rect 229756 264330 229784 271118
rect 230400 269958 230428 277766
rect 231412 272542 231440 277780
rect 232530 277766 233188 277794
rect 230572 272536 230624 272542
rect 230572 272478 230624 272484
rect 231400 272536 231452 272542
rect 231400 272478 231452 272484
rect 230388 269952 230440 269958
rect 230388 269894 230440 269900
rect 230584 264330 230612 272478
rect 233160 270494 233188 277766
rect 233712 271454 233740 277780
rect 234908 274174 234936 277780
rect 236104 275466 236132 277780
rect 237300 277394 237328 277780
rect 237208 277366 237328 277394
rect 236092 275460 236144 275466
rect 236092 275402 236144 275408
rect 234896 274168 234948 274174
rect 234896 274110 234948 274116
rect 234896 273964 234948 273970
rect 234896 273906 234948 273912
rect 233700 271448 233752 271454
rect 233700 271390 233752 271396
rect 234160 271312 234212 271318
rect 234160 271254 234212 271260
rect 233160 270466 233280 270494
rect 232320 269816 232372 269822
rect 232320 269758 232372 269764
rect 230756 268388 230808 268394
rect 230756 268330 230808 268336
rect 230768 266422 230796 268330
rect 231584 267436 231636 267442
rect 231584 267378 231636 267384
rect 230756 266416 230808 266422
rect 230756 266358 230808 266364
rect 229756 264302 230138 264330
rect 230584 264302 230874 264330
rect 231596 264316 231624 267378
rect 232332 264316 232360 269758
rect 233252 267170 233280 270466
rect 233792 267300 233844 267306
rect 233792 267242 233844 267248
rect 233240 267164 233292 267170
rect 233240 267106 233292 267112
rect 233056 266416 233108 266422
rect 233056 266358 233108 266364
rect 233068 264316 233096 266358
rect 233804 264316 233832 267242
rect 234172 264330 234200 271254
rect 234908 264330 234936 273906
rect 236736 270088 236788 270094
rect 236736 270030 236788 270036
rect 236000 267028 236052 267034
rect 236000 266970 236052 266976
rect 234172 264302 234554 264330
rect 234908 264302 235290 264330
rect 236012 264316 236040 266970
rect 236748 264316 236776 270030
rect 237208 269822 237236 277366
rect 238496 275330 238524 277780
rect 239600 277394 239628 277780
rect 240810 277766 241376 277794
rect 239600 277366 239720 277394
rect 237380 275324 237432 275330
rect 237380 275266 237432 275272
rect 238484 275324 238536 275330
rect 238484 275266 238536 275272
rect 237196 269816 237248 269822
rect 237196 269758 237248 269764
rect 237392 264330 237420 275266
rect 239496 274168 239548 274174
rect 239496 274110 239548 274116
rect 239312 272536 239364 272542
rect 239312 272478 239364 272484
rect 237840 271584 237892 271590
rect 237840 271526 237892 271532
rect 237852 264330 237880 271526
rect 238944 269952 238996 269958
rect 238944 269894 238996 269900
rect 237392 264302 237498 264330
rect 237852 264302 238234 264330
rect 238956 264316 238984 269894
rect 239324 264330 239352 272478
rect 239508 266422 239536 274110
rect 239692 272610 239720 277366
rect 239680 272604 239732 272610
rect 239680 272546 239732 272552
rect 240784 271448 240836 271454
rect 240784 271390 240836 271396
rect 240416 267164 240468 267170
rect 240416 267106 240468 267112
rect 239496 266416 239548 266422
rect 239496 266358 239548 266364
rect 239324 264302 239706 264330
rect 240428 264316 240456 267106
rect 240796 264330 240824 271390
rect 241348 266558 241376 277766
rect 241992 274718 242020 277780
rect 242256 275460 242308 275466
rect 242256 275402 242308 275408
rect 241980 274712 242032 274718
rect 241980 274654 242032 274660
rect 241336 266552 241388 266558
rect 241336 266494 241388 266500
rect 241888 266416 241940 266422
rect 241888 266358 241940 266364
rect 240796 264302 241178 264330
rect 241900 264316 241928 266358
rect 242268 264330 242296 275402
rect 243188 270366 243216 277780
rect 243728 275324 243780 275330
rect 243728 275266 243780 275272
rect 243176 270360 243228 270366
rect 243176 270302 243228 270308
rect 243360 269816 243412 269822
rect 243360 269758 243412 269764
rect 242268 264302 242650 264330
rect 243372 264316 243400 269758
rect 243740 264330 243768 275266
rect 244384 270502 244412 277780
rect 245580 275194 245608 277780
rect 245568 275188 245620 275194
rect 245568 275130 245620 275136
rect 246304 275188 246356 275194
rect 246304 275130 246356 275136
rect 246028 274712 246080 274718
rect 246028 274654 246080 274660
rect 244556 272604 244608 272610
rect 244556 272546 244608 272552
rect 244372 270496 244424 270502
rect 244372 270438 244424 270444
rect 244568 264330 244596 272546
rect 245568 266552 245620 266558
rect 245568 266494 245620 266500
rect 243740 264302 244122 264330
rect 244568 264302 244858 264330
rect 245580 264316 245608 266494
rect 246040 264330 246068 274654
rect 246316 266626 246344 275130
rect 246776 274718 246804 277780
rect 247894 277766 248368 277794
rect 246764 274712 246816 274718
rect 246764 274654 246816 274660
rect 247776 270496 247828 270502
rect 247776 270438 247828 270444
rect 247040 270360 247092 270366
rect 247040 270302 247092 270308
rect 246304 266620 246356 266626
rect 246304 266562 246356 266568
rect 246040 264302 246330 264330
rect 247052 264316 247080 270302
rect 247788 264316 247816 270438
rect 248340 269142 248368 277766
rect 249076 275058 249104 277780
rect 250272 277394 250300 277780
rect 250180 277366 250300 277394
rect 251192 277766 251482 277794
rect 249064 275052 249116 275058
rect 249064 274994 249116 275000
rect 248880 274712 248932 274718
rect 248880 274654 248932 274660
rect 248328 269136 248380 269142
rect 248328 269078 248380 269084
rect 248512 266620 248564 266626
rect 248512 266562 248564 266568
rect 248524 264316 248552 266562
rect 248892 264330 248920 274654
rect 250180 270502 250208 277366
rect 250352 275052 250404 275058
rect 250352 274994 250404 275000
rect 250168 270496 250220 270502
rect 250168 270438 250220 270444
rect 249984 269136 250036 269142
rect 249984 269078 250036 269084
rect 248892 264302 249274 264330
rect 249996 264316 250024 269078
rect 250364 264330 250392 274994
rect 251192 266422 251220 277766
rect 251456 270496 251508 270502
rect 251456 270438 251508 270444
rect 251180 266416 251232 266422
rect 251180 266358 251232 266364
rect 250364 264302 250746 264330
rect 251468 264316 251496 270438
rect 252192 266416 252244 266422
rect 252192 266358 252244 266364
rect 252204 264316 252232 266358
rect 252664 264330 252692 277780
rect 253032 277766 253874 277794
rect 254412 277766 255070 277794
rect 255332 277766 256174 277794
rect 256712 277766 257370 277794
rect 258092 277766 258566 277794
rect 259472 277766 259762 277794
rect 253032 267734 253060 277766
rect 253032 267706 253336 267734
rect 253308 264330 253336 267706
rect 252664 264302 252954 264330
rect 253308 264302 253690 264330
rect 254412 264316 254440 277766
rect 255332 267734 255360 277766
rect 255148 267706 255360 267734
rect 255148 264316 255176 267706
rect 256516 266892 256568 266898
rect 256516 266834 256568 266840
rect 255872 266416 255924 266422
rect 255872 266358 255924 266364
rect 255884 264316 255912 266358
rect 256528 264330 256556 266834
rect 256712 266422 256740 277766
rect 257344 267232 257396 267238
rect 257344 267174 257396 267180
rect 256700 266416 256752 266422
rect 256700 266358 256752 266364
rect 256528 264302 256634 264330
rect 257356 264316 257384 267174
rect 258092 266898 258120 277766
rect 258816 270496 258868 270502
rect 258816 270438 258868 270444
rect 258080 266892 258132 266898
rect 258080 266834 258132 266840
rect 258080 266416 258132 266422
rect 258080 266358 258132 266364
rect 258092 264316 258120 266358
rect 258828 264316 258856 270438
rect 259472 267238 259500 277766
rect 260944 277394 260972 277780
rect 260852 277366 260972 277394
rect 261312 277766 262154 277794
rect 262600 277766 263258 277794
rect 263612 277766 264454 277794
rect 264992 277766 265650 277794
rect 266372 277766 266846 277794
rect 260852 269550 260880 277366
rect 261312 270502 261340 277766
rect 261300 270496 261352 270502
rect 261300 270438 261352 270444
rect 261024 270360 261076 270366
rect 261024 270302 261076 270308
rect 259644 269544 259696 269550
rect 259644 269486 259696 269492
rect 260840 269544 260892 269550
rect 260840 269486 260892 269492
rect 259460 267232 259512 267238
rect 259460 267174 259512 267180
rect 259656 266422 259684 269486
rect 259920 266552 259972 266558
rect 259920 266494 259972 266500
rect 259644 266416 259696 266422
rect 259644 266358 259696 266364
rect 259932 264330 259960 266494
rect 260288 266416 260340 266422
rect 260288 266358 260340 266364
rect 259578 264302 259960 264330
rect 260300 264316 260328 266358
rect 261036 264316 261064 270302
rect 261760 269816 261812 269822
rect 261760 269758 261812 269764
rect 261772 266422 261800 269758
rect 262600 266558 262628 277766
rect 263416 271788 263468 271794
rect 263416 271730 263468 271736
rect 262864 267300 262916 267306
rect 262864 267242 262916 267248
rect 262588 266552 262640 266558
rect 262588 266494 262640 266500
rect 261760 266416 261812 266422
rect 261760 266358 261812 266364
rect 262128 266416 262180 266422
rect 262128 266358 262180 266364
rect 262140 264330 262168 266358
rect 262876 264330 262904 267242
rect 263428 264330 263456 271730
rect 263612 269822 263640 277766
rect 264992 270366 265020 277766
rect 265900 275324 265952 275330
rect 265900 275266 265952 275272
rect 264980 270360 265032 270366
rect 264980 270302 265032 270308
rect 263600 269816 263652 269822
rect 263600 269758 263652 269764
rect 265440 269816 265492 269822
rect 265440 269758 265492 269764
rect 264704 269340 264756 269346
rect 264704 269282 264756 269288
rect 263968 267776 264020 267782
rect 263968 267718 264020 267724
rect 261786 264302 262168 264330
rect 262522 264302 262904 264330
rect 263258 264302 263456 264330
rect 263980 264316 264008 267718
rect 264716 264316 264744 269282
rect 265452 264316 265480 269758
rect 265912 269346 265940 275266
rect 266176 270088 266228 270094
rect 266176 270030 266228 270036
rect 265900 269340 265952 269346
rect 265900 269282 265952 269288
rect 266188 264316 266216 270030
rect 266372 266422 266400 277766
rect 268028 277394 268056 277780
rect 267936 277366 268056 277394
rect 266912 269952 266964 269958
rect 266912 269894 266964 269900
rect 266360 266416 266412 266422
rect 266360 266358 266412 266364
rect 266924 264316 266952 269894
rect 267936 267306 267964 277366
rect 269224 271794 269252 277780
rect 269592 277766 270434 277794
rect 269212 271788 269264 271794
rect 269212 271730 269264 271736
rect 268844 271448 268896 271454
rect 268844 271390 268896 271396
rect 267924 267300 267976 267306
rect 267924 267242 267976 267248
rect 267648 267164 267700 267170
rect 267648 267106 267700 267112
rect 267660 264316 267688 267106
rect 268856 264330 268884 271390
rect 269120 269000 269172 269006
rect 269120 268942 269172 268948
rect 268410 264302 268884 264330
rect 269132 264316 269160 268942
rect 269592 267782 269620 277766
rect 271524 275330 271552 277780
rect 271892 277766 272734 277794
rect 273272 277766 273930 277794
rect 274652 277766 275126 277794
rect 271512 275324 271564 275330
rect 271512 275266 271564 275272
rect 271144 274712 271196 274718
rect 271144 274654 271196 274660
rect 269580 267776 269632 267782
rect 269580 267718 269632 267724
rect 271156 267170 271184 274654
rect 271696 272536 271748 272542
rect 271696 272478 271748 272484
rect 271708 267734 271736 272478
rect 271892 269822 271920 277766
rect 273076 271312 273128 271318
rect 273076 271254 273128 271260
rect 271880 269816 271932 269822
rect 271880 269758 271932 269764
rect 271880 269680 271932 269686
rect 271880 269622 271932 269628
rect 271892 267734 271920 269622
rect 271616 267706 271736 267734
rect 271800 267706 271920 267734
rect 271144 267164 271196 267170
rect 271144 267106 271196 267112
rect 269856 266552 269908 266558
rect 269856 266494 269908 266500
rect 269868 264316 269896 266494
rect 271616 266422 271644 267706
rect 270592 266416 270644 266422
rect 270592 266358 270644 266364
rect 271604 266416 271656 266422
rect 271604 266358 271656 266364
rect 270604 264316 270632 266358
rect 271800 264330 271828 267706
rect 272064 267164 272116 267170
rect 272064 267106 272116 267112
rect 271354 264302 271828 264330
rect 272076 264316 272104 267106
rect 273088 264330 273116 271254
rect 273272 270094 273300 277766
rect 274364 274236 274416 274242
rect 274364 274178 274416 274184
rect 273260 270088 273312 270094
rect 273260 270030 273312 270036
rect 273536 268388 273588 268394
rect 273536 268330 273588 268336
rect 272826 264302 273116 264330
rect 273548 264316 273576 268330
rect 274376 267734 274404 274178
rect 274652 269958 274680 277766
rect 276308 274718 276336 277780
rect 276296 274712 276348 274718
rect 276296 274654 276348 274660
rect 276664 274712 276716 274718
rect 276664 274654 276716 274660
rect 276480 270088 276532 270094
rect 276480 270030 276532 270036
rect 274640 269952 274692 269958
rect 274640 269894 274692 269900
rect 275008 269952 275060 269958
rect 275008 269894 275060 269900
rect 274640 269136 274692 269142
rect 274640 269078 274692 269084
rect 274284 267706 274404 267734
rect 274284 264316 274312 267706
rect 274652 266558 274680 269078
rect 274640 266552 274692 266558
rect 274640 266494 274692 266500
rect 275020 264316 275048 269894
rect 275744 267300 275796 267306
rect 275744 267242 275796 267248
rect 275756 264316 275784 267242
rect 276492 264316 276520 270030
rect 276676 269006 276704 274654
rect 277504 271454 277532 277780
rect 278412 275324 278464 275330
rect 278412 275266 278464 275272
rect 277492 271448 277544 271454
rect 277492 271390 277544 271396
rect 277308 271176 277360 271182
rect 277308 271118 277360 271124
rect 276664 269000 276716 269006
rect 276664 268942 276716 268948
rect 277320 267734 277348 271118
rect 277228 267706 277348 267734
rect 277228 264316 277256 267706
rect 278424 264330 278452 275266
rect 278700 274718 278728 277780
rect 278976 277766 279818 277794
rect 278688 274712 278740 274718
rect 278688 274654 278740 274660
rect 278976 269142 279004 277766
rect 280712 274712 280764 274718
rect 280712 274654 280764 274660
rect 279884 273964 279936 273970
rect 279884 273906 279936 273912
rect 278964 269136 279016 269142
rect 278964 269078 279016 269084
rect 278688 267028 278740 267034
rect 278688 266970 278740 266976
rect 277978 264302 278452 264330
rect 278700 264316 278728 266970
rect 279896 264330 279924 273906
rect 280724 267170 280752 274654
rect 281000 272542 281028 277780
rect 281552 277766 282210 277794
rect 280988 272536 281040 272542
rect 280988 272478 281040 272484
rect 280988 272400 281040 272406
rect 280988 272342 281040 272348
rect 281000 267306 281028 272342
rect 281552 269686 281580 277766
rect 282920 275596 282972 275602
rect 282920 275538 282972 275544
rect 282184 272536 282236 272542
rect 282184 272478 282236 272484
rect 281540 269680 281592 269686
rect 281540 269622 281592 269628
rect 281632 268524 281684 268530
rect 281632 268466 281684 268472
rect 280988 267300 281040 267306
rect 280988 267242 281040 267248
rect 280712 267164 280764 267170
rect 280712 267106 280764 267112
rect 280160 266552 280212 266558
rect 280160 266494 280212 266500
rect 279450 264302 279924 264330
rect 280172 264316 280200 266494
rect 280896 266416 280948 266422
rect 280896 266358 280948 266364
rect 280908 264316 280936 266358
rect 281644 264316 281672 268466
rect 282196 266422 282224 272478
rect 282932 268394 282960 275538
rect 283392 274718 283420 277780
rect 283380 274712 283432 274718
rect 283380 274654 283432 274660
rect 283932 274100 283984 274106
rect 283932 274042 283984 274048
rect 283104 269816 283156 269822
rect 283104 269758 283156 269764
rect 282920 268388 282972 268394
rect 282920 268330 282972 268336
rect 282368 267300 282420 267306
rect 282368 267242 282420 267248
rect 282184 266416 282236 266422
rect 282184 266358 282236 266364
rect 282380 264316 282408 267242
rect 283116 264316 283144 269758
rect 283944 267734 283972 274042
rect 284588 271318 284616 277780
rect 285784 275602 285812 277780
rect 285772 275596 285824 275602
rect 285772 275538 285824 275544
rect 285864 275460 285916 275466
rect 285864 275402 285916 275408
rect 285588 271448 285640 271454
rect 285588 271390 285640 271396
rect 284576 271312 284628 271318
rect 284576 271254 284628 271260
rect 284576 268796 284628 268802
rect 284576 268738 284628 268744
rect 283852 267706 283972 267734
rect 283852 264316 283880 267706
rect 284588 264316 284616 268738
rect 285600 264330 285628 271390
rect 285876 268802 285904 275402
rect 286888 274242 286916 277780
rect 287072 277766 288098 277794
rect 286876 274236 286928 274242
rect 286876 274178 286928 274184
rect 287072 269958 287100 277766
rect 289084 272672 289136 272678
rect 289084 272614 289136 272620
rect 287060 269952 287112 269958
rect 287060 269894 287112 269900
rect 287520 269952 287572 269958
rect 287520 269894 287572 269900
rect 285864 268796 285916 268802
rect 285864 268738 285916 268744
rect 285772 268660 285824 268666
rect 285772 268602 285824 268608
rect 285784 266558 285812 268602
rect 286784 268388 286836 268394
rect 286784 268330 286836 268336
rect 286048 267572 286100 267578
rect 286048 267514 286100 267520
rect 285772 266552 285824 266558
rect 285772 266494 285824 266500
rect 285338 264302 285628 264330
rect 286060 264316 286088 267514
rect 286796 264316 286824 268330
rect 287532 264316 287560 269894
rect 288256 267708 288308 267714
rect 288256 267650 288308 267656
rect 288268 264316 288296 267650
rect 289096 267306 289124 272614
rect 289280 272406 289308 277780
rect 289832 277766 290490 277794
rect 289268 272400 289320 272406
rect 289268 272342 289320 272348
rect 289636 271584 289688 271590
rect 289636 271526 289688 271532
rect 289084 267300 289136 267306
rect 289084 267242 289136 267248
rect 288992 266416 289044 266422
rect 288992 266358 289044 266364
rect 289004 264316 289032 266358
rect 289648 264330 289676 271526
rect 289832 270094 289860 277766
rect 290464 274236 290516 274242
rect 290464 274178 290516 274184
rect 289820 270088 289872 270094
rect 289820 270030 289872 270036
rect 290476 267578 290504 274178
rect 291672 271182 291700 277780
rect 292868 275330 292896 277780
rect 292856 275324 292908 275330
rect 292856 275266 292908 275272
rect 294064 274718 294092 277780
rect 293224 274712 293276 274718
rect 293224 274654 293276 274660
rect 294052 274712 294104 274718
rect 294052 274654 294104 274660
rect 291844 271312 291896 271318
rect 291844 271254 291896 271260
rect 291660 271176 291712 271182
rect 291660 271118 291712 271124
rect 290832 270224 290884 270230
rect 290832 270166 290884 270172
rect 290464 267572 290516 267578
rect 290464 267514 290516 267520
rect 290844 264330 290872 270166
rect 291200 266552 291252 266558
rect 291200 266494 291252 266500
rect 289648 264302 289754 264330
rect 290490 264302 290872 264330
rect 291212 264316 291240 266494
rect 291856 266422 291884 271254
rect 292396 271176 292448 271182
rect 292396 271118 292448 271124
rect 291844 266416 291896 266422
rect 291844 266358 291896 266364
rect 292408 264330 292436 271118
rect 292672 270496 292724 270502
rect 292672 270438 292724 270444
rect 291962 264302 292436 264330
rect 292684 264316 292712 270438
rect 293236 267034 293264 274654
rect 295168 273970 295196 277780
rect 295352 277766 296378 277794
rect 295156 273964 295208 273970
rect 295156 273906 295208 273912
rect 294604 273828 294656 273834
rect 294604 273770 294656 273776
rect 293408 267164 293460 267170
rect 293408 267106 293460 267112
rect 293224 267028 293276 267034
rect 293224 266970 293276 266976
rect 293420 264316 293448 267106
rect 294616 266558 294644 273770
rect 295156 273080 295208 273086
rect 295156 273022 295208 273028
rect 294880 267572 294932 267578
rect 294880 267514 294932 267520
rect 294604 266552 294656 266558
rect 294604 266494 294656 266500
rect 294144 266416 294196 266422
rect 294144 266358 294196 266364
rect 294156 264316 294184 266358
rect 294892 264316 294920 267514
rect 295168 266422 295196 273022
rect 295352 268666 295380 277766
rect 295524 274712 295576 274718
rect 295524 274654 295576 274660
rect 295340 268660 295392 268666
rect 295340 268602 295392 268608
rect 295536 268530 295564 274654
rect 297560 272542 297588 277780
rect 298008 275732 298060 275738
rect 298008 275674 298060 275680
rect 297548 272536 297600 272542
rect 297548 272478 297600 272484
rect 297364 271856 297416 271862
rect 297364 271798 297416 271804
rect 296628 271720 296680 271726
rect 296628 271662 296680 271668
rect 295524 268524 295576 268530
rect 295524 268466 295576 268472
rect 295616 267436 295668 267442
rect 295616 267378 295668 267384
rect 295156 266416 295208 266422
rect 295156 266358 295208 266364
rect 295628 264316 295656 267378
rect 296640 264330 296668 271662
rect 297088 268524 297140 268530
rect 297088 268466 297140 268472
rect 296378 264302 296668 264330
rect 297100 264316 297128 268466
rect 297376 267714 297404 271798
rect 298020 271590 298048 275674
rect 298756 274718 298784 277780
rect 299020 275596 299072 275602
rect 299020 275538 299072 275544
rect 298744 274712 298796 274718
rect 298744 274654 298796 274660
rect 299032 274106 299060 275538
rect 299204 274372 299256 274378
rect 299204 274314 299256 274320
rect 299020 274100 299072 274106
rect 299020 274042 299072 274048
rect 298008 271584 298060 271590
rect 298008 271526 298060 271532
rect 299216 269770 299244 274314
rect 299952 272678 299980 277780
rect 300872 277766 301162 277794
rect 300676 272808 300728 272814
rect 300676 272750 300728 272756
rect 299940 272672 299992 272678
rect 299940 272614 299992 272620
rect 300124 272672 300176 272678
rect 300124 272614 300176 272620
rect 299032 269742 299244 269770
rect 297364 267708 297416 267714
rect 297364 267650 297416 267656
rect 297824 266416 297876 266422
rect 297824 266358 297876 266364
rect 297836 264316 297864 266358
rect 299032 264330 299060 269742
rect 299296 268660 299348 268666
rect 299296 268602 299348 268608
rect 298586 264302 299060 264330
rect 299308 264316 299336 268602
rect 300136 267578 300164 272614
rect 300124 267572 300176 267578
rect 300124 267514 300176 267520
rect 300032 267028 300084 267034
rect 300032 266970 300084 266976
rect 300044 264316 300072 266970
rect 300688 264330 300716 272750
rect 300872 269822 300900 277766
rect 302344 275602 302372 277780
rect 302332 275596 302384 275602
rect 302332 275538 302384 275544
rect 303448 275466 303476 277780
rect 303436 275460 303488 275466
rect 303436 275402 303488 275408
rect 302240 275324 302292 275330
rect 302240 275266 302292 275272
rect 301504 275188 301556 275194
rect 301504 275130 301556 275136
rect 301516 271726 301544 275130
rect 302252 273086 302280 275266
rect 302240 273080 302292 273086
rect 302240 273022 302292 273028
rect 302884 272944 302936 272950
rect 302884 272886 302936 272892
rect 301504 271720 301556 271726
rect 301504 271662 301556 271668
rect 301964 270360 302016 270366
rect 301964 270302 302016 270308
rect 301228 270088 301280 270094
rect 301228 270030 301280 270036
rect 300860 269816 300912 269822
rect 300860 269758 300912 269764
rect 301240 266422 301268 270030
rect 301976 267442 302004 270302
rect 301964 267436 302016 267442
rect 301964 267378 302016 267384
rect 302896 267306 302924 272886
rect 303436 272536 303488 272542
rect 303436 272478 303488 272484
rect 302884 267300 302936 267306
rect 302884 267242 302936 267248
rect 302240 267164 302292 267170
rect 302240 267106 302292 267112
rect 301504 266552 301556 266558
rect 301504 266494 301556 266500
rect 301228 266416 301280 266422
rect 301228 266358 301280 266364
rect 300688 264302 300794 264330
rect 301516 264316 301544 266494
rect 302252 264316 302280 267106
rect 303448 264330 303476 272478
rect 304644 271454 304672 277780
rect 305092 275732 305144 275738
rect 305092 275674 305144 275680
rect 304908 271720 304960 271726
rect 304908 271662 304960 271668
rect 304632 271448 304684 271454
rect 304632 271390 304684 271396
rect 304172 268932 304224 268938
rect 304172 268874 304224 268880
rect 304184 266558 304212 268874
rect 304172 266552 304224 266558
rect 304172 266494 304224 266500
rect 304448 266552 304500 266558
rect 304448 266494 304500 266500
rect 303712 266416 303764 266422
rect 303712 266358 303764 266364
rect 303002 264302 303476 264330
rect 303724 264316 303752 266358
rect 304460 264316 304488 266494
rect 304920 266422 304948 271662
rect 305104 270502 305132 275674
rect 305840 274242 305868 277780
rect 306392 277766 307050 277794
rect 307772 277766 308246 277794
rect 306196 274508 306248 274514
rect 306196 274450 306248 274456
rect 305828 274236 305880 274242
rect 305828 274178 305880 274184
rect 305092 270496 305144 270502
rect 305092 270438 305144 270444
rect 305552 269816 305604 269822
rect 305552 269758 305604 269764
rect 305564 266558 305592 269758
rect 305920 267708 305972 267714
rect 305920 267650 305972 267656
rect 305552 266552 305604 266558
rect 305552 266494 305604 266500
rect 304908 266416 304960 266422
rect 304908 266358 304960 266364
rect 305184 266416 305236 266422
rect 305184 266358 305236 266364
rect 305196 264316 305224 266358
rect 305932 264316 305960 267650
rect 306208 266422 306236 274450
rect 306392 268394 306420 277766
rect 307576 274100 307628 274106
rect 307576 274042 307628 274048
rect 306380 268388 306432 268394
rect 306380 268330 306432 268336
rect 306656 267300 306708 267306
rect 306656 267242 306708 267248
rect 306196 266416 306248 266422
rect 306196 266358 306248 266364
rect 306668 264316 306696 267242
rect 307588 264330 307616 274042
rect 307772 269958 307800 277766
rect 309428 271862 309456 277780
rect 310060 274236 310112 274242
rect 310060 274178 310112 274184
rect 309416 271856 309468 271862
rect 309416 271798 309468 271804
rect 309048 271584 309100 271590
rect 309048 271526 309100 271532
rect 307760 269952 307812 269958
rect 307760 269894 307812 269900
rect 308128 267436 308180 267442
rect 308128 267378 308180 267384
rect 307418 264302 307616 264330
rect 308140 264316 308168 267378
rect 309060 264330 309088 271526
rect 310072 264330 310100 274178
rect 310532 271318 310560 277780
rect 311728 275602 311756 277780
rect 311912 277766 312938 277794
rect 311716 275596 311768 275602
rect 311716 275538 311768 275544
rect 311716 271448 311768 271454
rect 311716 271390 311768 271396
rect 310520 271312 310572 271318
rect 310520 271254 310572 271260
rect 310336 269952 310388 269958
rect 310336 269894 310388 269900
rect 308890 264302 309088 264330
rect 309626 264302 310100 264330
rect 310348 264316 310376 269894
rect 311532 269680 311584 269686
rect 311532 269622 311584 269628
rect 311544 267034 311572 269622
rect 311532 267028 311584 267034
rect 311532 266970 311584 266976
rect 311072 266892 311124 266898
rect 311072 266834 311124 266840
rect 311084 264316 311112 266834
rect 311728 264330 311756 271390
rect 311912 270230 311940 277766
rect 313280 275596 313332 275602
rect 313280 275538 313332 275544
rect 313292 274378 313320 275538
rect 313280 274372 313332 274378
rect 313280 274314 313332 274320
rect 314120 273970 314148 277780
rect 314108 273964 314160 273970
rect 314108 273906 314160 273912
rect 314476 273964 314528 273970
rect 314476 273906 314528 273912
rect 312544 271856 312596 271862
rect 312544 271798 312596 271804
rect 311900 270224 311952 270230
rect 311900 270166 311952 270172
rect 312556 267306 312584 271798
rect 312820 270224 312872 270230
rect 312820 270166 312872 270172
rect 312544 267300 312596 267306
rect 312544 267242 312596 267248
rect 312832 267170 312860 270166
rect 312820 267164 312872 267170
rect 312820 267106 312872 267112
rect 313280 267164 313332 267170
rect 313280 267106 313332 267112
rect 312544 267028 312596 267034
rect 312544 266970 312596 266976
rect 311728 264302 311834 264330
rect 312556 264316 312584 266970
rect 313292 264316 313320 267106
rect 314488 264330 314516 273906
rect 315316 271182 315344 277780
rect 316512 275738 316540 277780
rect 316776 275868 316828 275874
rect 316776 275810 316828 275816
rect 316500 275732 316552 275738
rect 316500 275674 316552 275680
rect 315948 271312 316000 271318
rect 315948 271254 316000 271260
rect 315304 271176 315356 271182
rect 315304 271118 315356 271124
rect 314752 268796 314804 268802
rect 314752 268738 314804 268744
rect 314042 264302 314516 264330
rect 314764 264316 314792 268738
rect 315960 264330 315988 271254
rect 316788 268666 316816 275810
rect 317328 275732 317380 275738
rect 317328 275674 317380 275680
rect 317144 273080 317196 273086
rect 317144 273022 317196 273028
rect 316776 268660 316828 268666
rect 316776 268602 316828 268608
rect 316960 268388 317012 268394
rect 316960 268330 317012 268336
rect 316224 266416 316276 266422
rect 316224 266358 316276 266364
rect 315514 264302 315988 264330
rect 316236 264316 316264 266358
rect 316972 264316 317000 268330
rect 317156 266422 317184 273022
rect 317340 272814 317368 275674
rect 317708 272950 317736 277780
rect 318812 275466 318840 277780
rect 319640 277766 320022 277794
rect 320284 277766 321218 277794
rect 318800 275460 318852 275466
rect 318800 275402 318852 275408
rect 318708 273828 318760 273834
rect 318708 273770 318760 273776
rect 317696 272944 317748 272950
rect 317696 272886 317748 272892
rect 317328 272808 317380 272814
rect 317328 272750 317380 272756
rect 317696 268660 317748 268666
rect 317696 268602 317748 268608
rect 317144 266416 317196 266422
rect 317144 266358 317196 266364
rect 317708 264316 317736 268602
rect 318720 264330 318748 273770
rect 319640 272678 319668 277766
rect 320088 275460 320140 275466
rect 320088 275402 320140 275408
rect 320100 274514 320128 275402
rect 320088 274508 320140 274514
rect 320088 274450 320140 274456
rect 319628 272672 319680 272678
rect 319628 272614 319680 272620
rect 319444 271040 319496 271046
rect 319444 270982 319496 270988
rect 319168 267572 319220 267578
rect 319168 267514 319220 267520
rect 318458 264302 318748 264330
rect 319180 264316 319208 267514
rect 319456 266898 319484 270982
rect 320284 270366 320312 277766
rect 322400 275330 322428 277780
rect 322952 277766 323610 277794
rect 324332 277766 324806 277794
rect 322388 275324 322440 275330
rect 322388 275266 322440 275272
rect 322572 275324 322624 275330
rect 322572 275266 322624 275272
rect 321468 272808 321520 272814
rect 321468 272750 321520 272756
rect 320272 270360 320324 270366
rect 320272 270302 320324 270308
rect 319444 266892 319496 266898
rect 319444 266834 319496 266840
rect 321284 266892 321336 266898
rect 321284 266834 321336 266840
rect 319904 266552 319956 266558
rect 319904 266494 319956 266500
rect 319916 264316 319944 266494
rect 320640 266416 320692 266422
rect 320640 266358 320692 266364
rect 320652 264316 320680 266358
rect 321296 264330 321324 266834
rect 321480 266422 321508 272750
rect 322584 272542 322612 275266
rect 322756 274372 322808 274378
rect 322756 274314 322808 274320
rect 322572 272536 322624 272542
rect 322572 272478 322624 272484
rect 322204 271176 322256 271182
rect 322204 271118 322256 271124
rect 322216 266558 322244 271118
rect 322204 266552 322256 266558
rect 322204 266494 322256 266500
rect 322480 266484 322532 266490
rect 322480 266426 322532 266432
rect 321468 266416 321520 266422
rect 321468 266358 321520 266364
rect 322492 264330 322520 266426
rect 321296 264302 321402 264330
rect 322138 264302 322520 264330
rect 322768 264330 322796 274314
rect 322952 268530 322980 277766
rect 323584 270496 323636 270502
rect 323584 270438 323636 270444
rect 322940 268524 322992 268530
rect 322940 268466 322992 268472
rect 322768 264302 322874 264330
rect 323596 264316 323624 270438
rect 324332 270094 324360 277766
rect 325988 275602 326016 277780
rect 327092 275874 327120 277780
rect 327276 277766 328302 277794
rect 327080 275868 327132 275874
rect 327080 275810 327132 275816
rect 325976 275596 326028 275602
rect 325976 275538 326028 275544
rect 326896 273216 326948 273222
rect 326896 273158 326948 273164
rect 325516 272944 325568 272950
rect 325516 272886 325568 272892
rect 324320 270088 324372 270094
rect 324320 270030 324372 270036
rect 324320 269068 324372 269074
rect 324320 269010 324372 269016
rect 324332 267714 324360 269010
rect 324688 268252 324740 268258
rect 324688 268194 324740 268200
rect 324320 267708 324372 267714
rect 324320 267650 324372 267656
rect 324700 264330 324728 268194
rect 325528 264330 325556 272886
rect 326712 272536 326764 272542
rect 326712 272478 326764 272484
rect 326724 266626 326752 272478
rect 325792 266620 325844 266626
rect 325792 266562 325844 266568
rect 326712 266620 326764 266626
rect 326712 266562 326764 266568
rect 324346 264302 324728 264330
rect 325082 264302 325556 264330
rect 325804 264316 325832 266562
rect 326908 264330 326936 273158
rect 327276 269686 327304 277766
rect 329484 275738 329512 277780
rect 329852 277766 330694 277794
rect 331416 277766 331890 277794
rect 329472 275732 329524 275738
rect 329472 275674 329524 275680
rect 329196 275596 329248 275602
rect 329196 275538 329248 275544
rect 327264 269680 327316 269686
rect 327264 269622 327316 269628
rect 328000 269408 328052 269414
rect 328000 269350 328052 269356
rect 327264 266756 327316 266762
rect 327264 266698 327316 266704
rect 326554 264302 326936 264330
rect 327276 264316 327304 266698
rect 328012 264316 328040 269350
rect 329208 264330 329236 275538
rect 329656 274508 329708 274514
rect 329656 274450 329708 274456
rect 329472 268524 329524 268530
rect 329472 268466 329524 268472
rect 329484 267442 329512 268466
rect 329472 267436 329524 267442
rect 329472 267378 329524 267384
rect 329668 264330 329696 274450
rect 329852 268938 329880 277766
rect 331220 275868 331272 275874
rect 331220 275810 331272 275816
rect 331232 274106 331260 275810
rect 331220 274100 331272 274106
rect 331220 274042 331272 274048
rect 331416 270230 331444 277766
rect 333072 275330 333100 277780
rect 333612 275596 333664 275602
rect 333612 275538 333664 275544
rect 333060 275324 333112 275330
rect 333060 275266 333112 275272
rect 332508 273556 332560 273562
rect 332508 273498 332560 273504
rect 331404 270224 331456 270230
rect 331404 270166 331456 270172
rect 332324 269680 332376 269686
rect 332324 269622 332376 269628
rect 330208 269544 330260 269550
rect 330208 269486 330260 269492
rect 329840 268932 329892 268938
rect 329840 268874 329892 268880
rect 328762 264302 329236 264330
rect 329498 264302 329696 264330
rect 330220 264316 330248 269486
rect 330484 267164 330536 267170
rect 330484 267106 330536 267112
rect 330496 266898 330524 267106
rect 330484 266892 330536 266898
rect 330484 266834 330536 266840
rect 330944 266756 330996 266762
rect 330944 266698 330996 266704
rect 330956 264316 330984 266698
rect 331680 266620 331732 266626
rect 331680 266562 331732 266568
rect 331692 264316 331720 266562
rect 332336 264330 332364 269622
rect 332520 266626 332548 273498
rect 333244 272672 333296 272678
rect 333244 272614 333296 272620
rect 333256 266762 333284 272614
rect 333244 266756 333296 266762
rect 333244 266698 333296 266704
rect 332508 266620 332560 266626
rect 332508 266562 332560 266568
rect 333624 264330 333652 275538
rect 334176 271726 334204 277780
rect 334164 271720 334216 271726
rect 334164 271662 334216 271668
rect 334624 270904 334676 270910
rect 334624 270846 334676 270852
rect 334636 267306 334664 270846
rect 334992 270360 335044 270366
rect 334992 270302 335044 270308
rect 334624 267300 334676 267306
rect 334624 267242 334676 267248
rect 333888 266892 333940 266898
rect 333888 266834 333940 266840
rect 332336 264302 332442 264330
rect 333178 264302 333652 264330
rect 333900 264316 333928 266834
rect 335004 264330 335032 270302
rect 335372 269822 335400 277780
rect 336568 275466 336596 277780
rect 336752 277766 337778 277794
rect 338592 277766 338974 277794
rect 336556 275460 336608 275466
rect 336556 275402 336608 275408
rect 336464 275188 336516 275194
rect 336464 275130 336516 275136
rect 336476 274242 336504 275130
rect 336464 274236 336516 274242
rect 336464 274178 336516 274184
rect 336556 274100 336608 274106
rect 336556 274042 336608 274048
rect 335360 269816 335412 269822
rect 335360 269758 335412 269764
rect 335728 267300 335780 267306
rect 335728 267242 335780 267248
rect 335740 264330 335768 267242
rect 336568 264330 336596 274042
rect 336752 269074 336780 277766
rect 338592 271862 338620 277766
rect 340156 275874 340184 277780
rect 340892 277766 341366 277794
rect 340144 275868 340196 275874
rect 340144 275810 340196 275816
rect 340236 275460 340288 275466
rect 340236 275402 340288 275408
rect 339224 274712 339276 274718
rect 339224 274654 339276 274660
rect 338580 271856 338632 271862
rect 338580 271798 338632 271804
rect 338948 271856 339000 271862
rect 338948 271798 339000 271804
rect 338028 271720 338080 271726
rect 338028 271662 338080 271668
rect 337200 270088 337252 270094
rect 337200 270030 337252 270036
rect 336740 269068 336792 269074
rect 336740 269010 336792 269016
rect 337212 264330 337240 270030
rect 338040 264330 338068 271662
rect 338488 269068 338540 269074
rect 338488 269010 338540 269016
rect 338500 267578 338528 269010
rect 338488 267572 338540 267578
rect 338488 267514 338540 267520
rect 338304 266756 338356 266762
rect 338304 266698 338356 266704
rect 334650 264302 335032 264330
rect 335386 264302 335768 264330
rect 336122 264302 336596 264330
rect 336858 264302 337240 264330
rect 337594 264302 338068 264330
rect 338316 264316 338344 266698
rect 338960 266490 338988 271798
rect 339236 269958 339264 274654
rect 339224 269952 339276 269958
rect 339224 269894 339276 269900
rect 339408 269952 339460 269958
rect 339408 269894 339460 269900
rect 338948 266484 339000 266490
rect 338948 266426 339000 266432
rect 339420 264330 339448 269894
rect 340248 264330 340276 275402
rect 340696 272128 340748 272134
rect 340696 272070 340748 272076
rect 340708 264330 340736 272070
rect 340892 268530 340920 277766
rect 342260 275324 342312 275330
rect 342260 275266 342312 275272
rect 342272 273970 342300 275266
rect 342260 273964 342312 273970
rect 342260 273906 342312 273912
rect 342456 271590 342484 277780
rect 343652 275194 343680 277780
rect 344008 276004 344060 276010
rect 344008 275946 344060 275952
rect 343824 275868 343876 275874
rect 343824 275810 343876 275816
rect 343640 275188 343692 275194
rect 343640 275130 343692 275136
rect 343548 273420 343600 273426
rect 343548 273362 343600 273368
rect 342444 271584 342496 271590
rect 342444 271526 342496 271532
rect 342536 270768 342588 270774
rect 342536 270710 342588 270716
rect 341248 269816 341300 269822
rect 341248 269758 341300 269764
rect 340880 268524 340932 268530
rect 340880 268466 340932 268472
rect 339066 264302 339448 264330
rect 339802 264302 340276 264330
rect 340538 264302 340736 264330
rect 341260 264316 341288 269758
rect 341984 267164 342036 267170
rect 341984 267106 342036 267112
rect 341996 264316 342024 267106
rect 342548 267034 342576 270710
rect 343364 267640 343416 267646
rect 343364 267582 343416 267588
rect 342536 267028 342588 267034
rect 342536 266970 342588 266976
rect 342720 266416 342772 266422
rect 342720 266358 342772 266364
rect 342732 264316 342760 266358
rect 343376 264330 343404 267582
rect 343560 266422 343588 273362
rect 343836 273222 343864 275810
rect 343824 273216 343876 273222
rect 343824 273158 343876 273164
rect 344020 273086 344048 275946
rect 344848 274718 344876 277780
rect 344836 274712 344888 274718
rect 344836 274654 344888 274660
rect 344008 273080 344060 273086
rect 344008 273022 344060 273028
rect 345664 272536 345716 272542
rect 345664 272478 345716 272484
rect 344192 267776 344244 267782
rect 344192 267718 344244 267724
rect 343548 266416 343600 266422
rect 343548 266358 343600 266364
rect 343376 264302 343482 264330
rect 344204 264316 344232 267718
rect 344928 267028 344980 267034
rect 344928 266970 344980 266976
rect 344940 264316 344968 266970
rect 345676 266626 345704 272478
rect 345848 271584 345900 271590
rect 345848 271526 345900 271532
rect 345860 267442 345888 271526
rect 346044 271046 346072 277780
rect 347044 275052 347096 275058
rect 347044 274994 347096 275000
rect 346032 271040 346084 271046
rect 346032 270982 346084 270988
rect 346400 270224 346452 270230
rect 346400 270166 346452 270172
rect 346412 267734 346440 270166
rect 347056 267782 347084 274994
rect 347240 271454 347268 277780
rect 348160 277766 348450 277794
rect 347228 271448 347280 271454
rect 347228 271390 347280 271396
rect 348160 270774 348188 277766
rect 348424 272264 348476 272270
rect 348424 272206 348476 272212
rect 348148 270768 348200 270774
rect 348148 270710 348200 270716
rect 347412 268932 347464 268938
rect 347412 268874 347464 268880
rect 346136 267706 346440 267734
rect 347044 267776 347096 267782
rect 347044 267718 347096 267724
rect 345848 267436 345900 267442
rect 345848 267378 345900 267384
rect 345664 266620 345716 266626
rect 345664 266562 345716 266568
rect 346136 264330 346164 267706
rect 346400 266416 346452 266422
rect 346400 266358 346452 266364
rect 345690 264302 346164 264330
rect 346412 264316 346440 266358
rect 347424 264330 347452 268874
rect 347688 267436 347740 267442
rect 347688 267378 347740 267384
rect 347700 266898 347728 267378
rect 348436 267306 348464 272206
rect 349632 270910 349660 277780
rect 350736 275330 350764 277780
rect 351946 277766 352144 277794
rect 350724 275324 350776 275330
rect 350724 275266 350776 275272
rect 350908 275324 350960 275330
rect 350908 275266 350960 275272
rect 350540 275188 350592 275194
rect 350540 275130 350592 275136
rect 350552 273834 350580 275130
rect 350920 275058 350948 275266
rect 350908 275052 350960 275058
rect 350908 274994 350960 275000
rect 351184 273964 351236 273970
rect 351184 273906 351236 273912
rect 350540 273828 350592 273834
rect 350540 273770 350592 273776
rect 350448 271040 350500 271046
rect 350448 270982 350500 270988
rect 349620 270904 349672 270910
rect 349620 270846 349672 270852
rect 349344 268524 349396 268530
rect 349344 268466 349396 268472
rect 348424 267300 348476 267306
rect 348424 267242 348476 267248
rect 347688 266892 347740 266898
rect 347688 266834 347740 266840
rect 347872 266892 347924 266898
rect 347872 266834 347924 266840
rect 347162 264302 347452 264330
rect 347884 264316 347912 266834
rect 348608 266552 348660 266558
rect 348608 266494 348660 266500
rect 348620 264316 348648 266494
rect 349356 264316 349384 268466
rect 350264 267572 350316 267578
rect 350264 267514 350316 267520
rect 350080 267300 350132 267306
rect 350080 267242 350132 267248
rect 350092 266422 350120 267242
rect 350276 267170 350304 267514
rect 350264 267164 350316 267170
rect 350264 267106 350316 267112
rect 350080 266416 350132 266422
rect 350080 266358 350132 266364
rect 350460 264330 350488 270982
rect 350816 267164 350868 267170
rect 350816 267106 350868 267112
rect 350106 264302 350488 264330
rect 350828 264316 350856 267106
rect 351196 267034 351224 273906
rect 351736 271992 351788 271998
rect 351736 271934 351788 271940
rect 351184 267028 351236 267034
rect 351184 266970 351236 266976
rect 351748 264330 351776 271934
rect 352116 268802 352144 277766
rect 353128 271318 353156 277780
rect 354324 276010 354352 277780
rect 354692 277766 355534 277794
rect 354312 276004 354364 276010
rect 354312 275946 354364 275952
rect 353944 274100 353996 274106
rect 353944 274042 353996 274048
rect 353116 271312 353168 271318
rect 353116 271254 353168 271260
rect 353208 270632 353260 270638
rect 353208 270574 353260 270580
rect 352104 268796 352156 268802
rect 352104 268738 352156 268744
rect 353024 267028 353076 267034
rect 353024 266970 353076 266976
rect 352288 266416 352340 266422
rect 352288 266358 352340 266364
rect 351578 264302 351776 264330
rect 352300 264316 352328 266358
rect 353036 264316 353064 266970
rect 353220 266422 353248 270574
rect 353956 267442 353984 274042
rect 354220 273828 354272 273834
rect 354220 273770 354272 273776
rect 353944 267436 353996 267442
rect 353944 267378 353996 267384
rect 353576 266892 353628 266898
rect 353576 266834 353628 266840
rect 353588 266626 353616 266834
rect 353576 266620 353628 266626
rect 353576 266562 353628 266568
rect 353208 266416 353260 266422
rect 353208 266358 353260 266364
rect 354232 264330 354260 273770
rect 354496 270768 354548 270774
rect 354496 270710 354548 270716
rect 353786 264302 354260 264330
rect 354508 264316 354536 270710
rect 354692 268394 354720 277766
rect 356716 274718 356744 277780
rect 356980 276004 357032 276010
rect 356980 275946 357032 275952
rect 355692 274712 355744 274718
rect 355692 274654 355744 274660
rect 356704 274712 356756 274718
rect 356704 274654 356756 274660
rect 355704 268666 355732 274654
rect 356992 271726 357020 275946
rect 357912 275194 357940 277780
rect 359016 277394 359044 277780
rect 359016 277366 359136 277394
rect 357900 275188 357952 275194
rect 357900 275130 357952 275136
rect 358728 274848 358780 274854
rect 358728 274790 358780 274796
rect 358740 274378 358768 274790
rect 358728 274372 358780 274378
rect 358728 274314 358780 274320
rect 358912 274372 358964 274378
rect 358912 274314 358964 274320
rect 358924 274258 358952 274314
rect 358740 274230 358952 274258
rect 358740 273290 358768 274230
rect 358176 273284 358228 273290
rect 358176 273226 358228 273232
rect 358728 273284 358780 273290
rect 358728 273226 358780 273232
rect 357992 273080 358044 273086
rect 357992 273022 358044 273028
rect 358004 272814 358032 273022
rect 357992 272808 358044 272814
rect 357992 272750 358044 272756
rect 356980 271720 357032 271726
rect 356980 271662 357032 271668
rect 357164 270904 357216 270910
rect 357164 270846 357216 270852
rect 355692 268660 355744 268666
rect 355692 268602 355744 268608
rect 354680 268388 354732 268394
rect 354680 268330 354732 268336
rect 354680 267980 354732 267986
rect 354680 267922 354732 267928
rect 354692 266626 354720 267922
rect 355968 267844 356020 267850
rect 355968 267786 356020 267792
rect 355232 267300 355284 267306
rect 355232 267242 355284 267248
rect 354680 266620 354732 266626
rect 354680 266562 354732 266568
rect 355244 264316 355272 267242
rect 355980 264316 356008 267786
rect 357176 264330 357204 270846
rect 358188 266762 358216 273226
rect 359108 269074 359136 277366
rect 359464 274644 359516 274650
rect 359464 274586 359516 274592
rect 359476 273970 359504 274586
rect 359464 273964 359516 273970
rect 359464 273906 359516 273912
rect 359464 272808 359516 272814
rect 359464 272750 359516 272756
rect 359476 272406 359504 272750
rect 359464 272400 359516 272406
rect 359464 272342 359516 272348
rect 360212 271318 360240 277780
rect 361212 273692 361264 273698
rect 361212 273634 361264 273640
rect 360200 271312 360252 271318
rect 360200 271254 360252 271260
rect 360108 271040 360160 271046
rect 360108 270982 360160 270988
rect 359096 269068 359148 269074
rect 359096 269010 359148 269016
rect 358544 268388 358596 268394
rect 358544 268330 358596 268336
rect 358176 266756 358228 266762
rect 358176 266698 358228 266704
rect 357440 266620 357492 266626
rect 357440 266562 357492 266568
rect 356730 264302 357204 264330
rect 357452 264316 357480 266562
rect 358556 264330 358584 268330
rect 359648 266892 359700 266898
rect 359648 266834 359700 266840
rect 358912 266620 358964 266626
rect 358912 266562 358964 266568
rect 358202 264302 358584 264330
rect 358924 264316 358952 266562
rect 359660 264316 359688 266834
rect 360120 266626 360148 270982
rect 361224 266626 361252 273634
rect 361408 273086 361436 277780
rect 361396 273080 361448 273086
rect 361396 273022 361448 273028
rect 361856 272400 361908 272406
rect 361856 272342 361908 272348
rect 361488 271448 361540 271454
rect 361488 271390 361540 271396
rect 360108 266620 360160 266626
rect 360108 266562 360160 266568
rect 360384 266620 360436 266626
rect 360384 266562 360436 266568
rect 361212 266620 361264 266626
rect 361212 266562 361264 266568
rect 360396 264316 360424 266562
rect 361500 264330 361528 271390
rect 361146 264302 361528 264330
rect 361868 264316 361896 272342
rect 362604 271590 362632 277780
rect 363800 271862 363828 277780
rect 364996 274854 365024 277780
rect 365824 277766 366114 277794
rect 367112 277766 367310 277794
rect 365628 275188 365680 275194
rect 365628 275130 365680 275136
rect 365260 274984 365312 274990
rect 365260 274926 365312 274932
rect 364984 274848 365036 274854
rect 364984 274790 365036 274796
rect 364340 273216 364392 273222
rect 364340 273158 364392 273164
rect 363788 271856 363840 271862
rect 363788 271798 363840 271804
rect 363696 271720 363748 271726
rect 363696 271662 363748 271668
rect 362592 271584 362644 271590
rect 362592 271526 362644 271532
rect 363236 267300 363288 267306
rect 363236 267242 363288 267248
rect 363248 266626 363276 267242
rect 363236 266620 363288 266626
rect 363236 266562 363288 266568
rect 362592 265804 362644 265810
rect 362592 265746 362644 265752
rect 362604 264316 362632 265746
rect 363708 264330 363736 271662
rect 364154 267744 364210 267753
rect 364154 267679 364210 267688
rect 364168 267578 364196 267679
rect 364156 267572 364208 267578
rect 364156 267514 364208 267520
rect 364352 266370 364380 273158
rect 365272 272814 365300 274926
rect 365640 274514 365668 275130
rect 365628 274508 365680 274514
rect 365628 274450 365680 274456
rect 365260 272808 365312 272814
rect 365260 272750 365312 272756
rect 365536 271584 365588 271590
rect 365536 271526 365588 271532
rect 365352 268116 365404 268122
rect 365352 268058 365404 268064
rect 364800 267708 364852 267714
rect 364800 267650 364852 267656
rect 364812 266490 364840 267650
rect 364984 267436 365036 267442
rect 364984 267378 365036 267384
rect 365168 267436 365220 267442
rect 365168 267378 365220 267384
rect 364996 267170 365024 267378
rect 364984 267164 365036 267170
rect 364984 267106 365036 267112
rect 365180 266762 365208 267378
rect 365168 266756 365220 266762
rect 365168 266698 365220 266704
rect 364800 266484 364852 266490
rect 364800 266426 364852 266432
rect 363354 264302 363736 264330
rect 364260 266342 364380 266370
rect 364260 264194 364288 266342
rect 365364 264330 365392 268058
rect 364826 264302 365392 264330
rect 365548 264316 365576 271526
rect 365824 270502 365852 277766
rect 366364 274508 366416 274514
rect 366364 274450 366416 274456
rect 365812 270496 365864 270502
rect 365812 270438 365864 270444
rect 365720 269408 365772 269414
rect 365720 269350 365772 269356
rect 365732 267578 365760 269350
rect 366376 267753 366404 274450
rect 367112 268258 367140 277766
rect 368020 274372 368072 274378
rect 368020 274314 368072 274320
rect 368032 273970 368060 274314
rect 368020 273964 368072 273970
rect 368020 273906 368072 273912
rect 368492 272950 368520 277780
rect 369688 274990 369716 277780
rect 370884 275874 370912 277780
rect 370872 275868 370924 275874
rect 370872 275810 370924 275816
rect 371056 275868 371108 275874
rect 371056 275810 371108 275816
rect 369676 274984 369728 274990
rect 369676 274926 369728 274932
rect 368848 273080 368900 273086
rect 368848 273022 368900 273028
rect 368480 272944 368532 272950
rect 368480 272886 368532 272892
rect 367744 270496 367796 270502
rect 367744 270438 367796 270444
rect 367100 268252 367152 268258
rect 367100 268194 367152 268200
rect 366362 267744 366418 267753
rect 366362 267679 366418 267688
rect 365720 267572 365772 267578
rect 365720 267514 365772 267520
rect 366272 267572 366324 267578
rect 366272 267514 366324 267520
rect 366284 264316 366312 267514
rect 367008 266756 367060 266762
rect 367008 266698 367060 266704
rect 367020 264316 367048 266698
rect 367756 264316 367784 270438
rect 368860 264330 368888 273022
rect 369952 271312 370004 271318
rect 369952 271254 370004 271260
rect 369216 268660 369268 268666
rect 369216 268602 369268 268608
rect 368506 264302 368888 264330
rect 369228 264316 369256 268602
rect 369964 264316 369992 271254
rect 371068 268530 371096 275810
rect 372080 272542 372108 277780
rect 372632 277766 373290 277794
rect 372632 273254 372660 277766
rect 374380 275738 374408 277780
rect 374368 275732 374420 275738
rect 374368 275674 374420 275680
rect 375576 275194 375604 277780
rect 376786 277766 376984 277794
rect 375564 275188 375616 275194
rect 375564 275130 375616 275136
rect 376024 275188 376076 275194
rect 376024 275130 376076 275136
rect 375288 275052 375340 275058
rect 375288 274994 375340 275000
rect 374552 274916 374604 274922
rect 374552 274858 374604 274864
rect 374564 273562 374592 274858
rect 374552 273556 374604 273562
rect 374552 273498 374604 273504
rect 372632 273226 372752 273254
rect 372068 272536 372120 272542
rect 372068 272478 372120 272484
rect 372528 269272 372580 269278
rect 372528 269214 372580 269220
rect 371056 268524 371108 268530
rect 371056 268466 371108 268472
rect 371424 268524 371476 268530
rect 371424 268466 371476 268472
rect 370504 267436 370556 267442
rect 370504 267378 370556 267384
rect 370688 267436 370740 267442
rect 370688 267378 370740 267384
rect 370516 266490 370544 267378
rect 370504 266484 370556 266490
rect 370504 266426 370556 266432
rect 370700 264316 370728 267378
rect 371436 264316 371464 268466
rect 372540 267714 372568 269214
rect 372724 269142 372752 273226
rect 374460 272536 374512 272542
rect 374460 272478 374512 272484
rect 374472 271998 374500 272478
rect 374644 272264 374696 272270
rect 374644 272206 374696 272212
rect 374828 272264 374880 272270
rect 374828 272206 374880 272212
rect 374656 271998 374684 272206
rect 374460 271992 374512 271998
rect 374460 271934 374512 271940
rect 374644 271992 374696 271998
rect 374644 271934 374696 271940
rect 374840 269770 374868 272206
rect 375300 272134 375328 274994
rect 375288 272128 375340 272134
rect 375288 272070 375340 272076
rect 374656 269742 374868 269770
rect 374460 269544 374512 269550
rect 374460 269486 374512 269492
rect 372712 269136 372764 269142
rect 372712 269078 372764 269084
rect 373908 269136 373960 269142
rect 373908 269078 373960 269084
rect 372528 267708 372580 267714
rect 372528 267650 372580 267656
rect 372896 267708 372948 267714
rect 372896 267650 372948 267656
rect 372160 266348 372212 266354
rect 372160 266290 372212 266296
rect 372172 264316 372200 266290
rect 372908 264316 372936 267650
rect 373920 267170 373948 269078
rect 374472 269006 374500 269486
rect 374460 269000 374512 269006
rect 374460 268942 374512 268948
rect 374460 267572 374512 267578
rect 374460 267514 374512 267520
rect 374472 267170 374500 267514
rect 373908 267164 373960 267170
rect 373908 267106 373960 267112
rect 374460 267164 374512 267170
rect 374460 267106 374512 267112
rect 373632 266212 373684 266218
rect 373632 266154 373684 266160
rect 373644 264316 373672 266154
rect 374656 264330 374684 269742
rect 374828 269680 374880 269686
rect 374828 269622 374880 269628
rect 374840 269414 374868 269622
rect 374828 269408 374880 269414
rect 374828 269350 374880 269356
rect 375012 269408 375064 269414
rect 375012 269350 375064 269356
rect 375024 269142 375052 269350
rect 375012 269136 375064 269142
rect 375012 269078 375064 269084
rect 375840 268932 375892 268938
rect 375840 268874 375892 268880
rect 375012 267708 375064 267714
rect 375012 267650 375064 267656
rect 375024 267458 375052 267650
rect 374840 267442 375052 267458
rect 374828 267436 375052 267442
rect 374880 267430 375052 267436
rect 374828 267378 374880 267384
rect 375472 267300 375524 267306
rect 375472 267242 375524 267248
rect 375484 264330 375512 267242
rect 374394 264302 374684 264330
rect 375130 264302 375512 264330
rect 375852 264316 375880 268874
rect 376036 268802 376064 275130
rect 376576 272808 376628 272814
rect 376576 272750 376628 272756
rect 376024 268796 376076 268802
rect 376024 268738 376076 268744
rect 376588 264316 376616 272750
rect 376760 272128 376812 272134
rect 376760 272070 376812 272076
rect 376772 267442 376800 272070
rect 376956 269142 376984 277766
rect 377968 272678 377996 277780
rect 379164 274922 379192 277780
rect 379532 277766 380374 277794
rect 379152 274916 379204 274922
rect 379152 274858 379204 274864
rect 378784 274780 378836 274786
rect 378784 274722 378836 274728
rect 378796 274242 378824 274722
rect 378784 274236 378836 274242
rect 378784 274178 378836 274184
rect 378784 273556 378836 273562
rect 378784 273498 378836 273504
rect 377956 272672 378008 272678
rect 377956 272614 378008 272620
rect 378140 272672 378192 272678
rect 378140 272614 378192 272620
rect 378152 272270 378180 272614
rect 378140 272264 378192 272270
rect 378140 272206 378192 272212
rect 376944 269136 376996 269142
rect 376944 269078 376996 269084
rect 378048 269068 378100 269074
rect 378048 269010 378100 269016
rect 377678 267472 377734 267481
rect 376760 267436 376812 267442
rect 377678 267407 377734 267416
rect 376760 267378 376812 267384
rect 377692 264330 377720 267407
rect 377338 264302 377720 264330
rect 378060 264316 378088 269010
rect 378796 266490 378824 273498
rect 379152 272264 379204 272270
rect 379152 272206 379204 272212
rect 378784 266484 378836 266490
rect 378784 266426 378836 266432
rect 379164 264330 379192 272206
rect 379532 269550 379560 277766
rect 380716 276956 380768 276962
rect 380716 276898 380768 276904
rect 379520 269544 379572 269550
rect 379520 269486 379572 269492
rect 379704 269544 379756 269550
rect 379704 269486 379756 269492
rect 379518 267472 379574 267481
rect 379518 267407 379574 267416
rect 379532 267306 379560 267407
rect 379520 267300 379572 267306
rect 379520 267242 379572 267248
rect 379716 267034 379744 269486
rect 379704 267028 379756 267034
rect 379704 266970 379756 266976
rect 379888 267028 379940 267034
rect 379888 266970 379940 266976
rect 379900 264330 379928 266970
rect 380728 264330 380756 276898
rect 380900 275732 380952 275738
rect 380900 275674 380952 275680
rect 380912 272542 380940 275674
rect 381556 275602 381584 277780
rect 381544 275596 381596 275602
rect 381544 275538 381596 275544
rect 382372 275052 382424 275058
rect 382372 274994 382424 275000
rect 381360 272944 381412 272950
rect 381360 272886 381412 272892
rect 380900 272536 380952 272542
rect 380900 272478 380952 272484
rect 381372 264330 381400 272886
rect 382384 271182 382412 274994
rect 382660 274106 382688 277780
rect 383672 277766 383870 277794
rect 382648 274100 382700 274106
rect 382648 274042 382700 274048
rect 383200 271448 383252 271454
rect 383200 271390 383252 271396
rect 382372 271176 382424 271182
rect 382372 271118 382424 271124
rect 382186 269648 382242 269657
rect 382186 269583 382242 269592
rect 382200 266626 382228 269583
rect 382464 268252 382516 268258
rect 382464 268194 382516 268200
rect 382188 266620 382240 266626
rect 382188 266562 382240 266568
rect 381728 266484 381780 266490
rect 381728 266426 381780 266432
rect 378810 264302 379192 264330
rect 379546 264302 379928 264330
rect 380282 264302 380756 264330
rect 381018 264302 381400 264330
rect 381740 264316 381768 266426
rect 382476 264316 382504 268194
rect 383212 264316 383240 271390
rect 383672 270366 383700 277766
rect 384488 272944 384540 272950
rect 384488 272886 384540 272892
rect 384500 272678 384528 272886
rect 384488 272672 384540 272678
rect 384488 272614 384540 272620
rect 385052 271998 385080 277780
rect 386248 274786 386276 277780
rect 386432 277766 387458 277794
rect 386236 274780 386288 274786
rect 386236 274722 386288 274728
rect 385040 271992 385092 271998
rect 385040 271934 385092 271940
rect 386432 270366 386460 277766
rect 387340 276820 387392 276826
rect 387340 276762 387392 276768
rect 383660 270360 383712 270366
rect 383660 270302 383712 270308
rect 383844 270360 383896 270366
rect 386420 270360 386472 270366
rect 383844 270302 383896 270308
rect 384946 270328 385002 270337
rect 383856 270094 383884 270302
rect 386604 270360 386656 270366
rect 386420 270302 386472 270308
rect 386602 270328 386604 270337
rect 386656 270328 386658 270337
rect 384946 270263 385002 270272
rect 386602 270263 386658 270272
rect 383844 270088 383896 270094
rect 383844 270030 383896 270036
rect 384120 270088 384172 270094
rect 384120 270030 384172 270036
rect 384132 269822 384160 270030
rect 384120 269816 384172 269822
rect 384120 269758 384172 269764
rect 384488 269680 384540 269686
rect 384486 269648 384488 269657
rect 384540 269648 384542 269657
rect 384486 269583 384542 269592
rect 384304 269068 384356 269074
rect 384304 269010 384356 269016
rect 384488 269068 384540 269074
rect 384488 269010 384540 269016
rect 384316 268802 384344 269010
rect 384304 268796 384356 268802
rect 384304 268738 384356 268744
rect 384500 268258 384528 269010
rect 384488 268252 384540 268258
rect 384488 268194 384540 268200
rect 384304 267436 384356 267442
rect 384304 267378 384356 267384
rect 384488 267436 384540 267442
rect 384488 267378 384540 267384
rect 383660 267300 383712 267306
rect 383660 267242 383712 267248
rect 383936 267300 383988 267306
rect 383936 267242 383988 267248
rect 383672 267073 383700 267242
rect 383658 267064 383714 267073
rect 383658 266999 383714 267008
rect 383948 264316 383976 267242
rect 384316 266490 384344 267378
rect 384500 267034 384528 267378
rect 384670 267064 384726 267073
rect 384488 267028 384540 267034
rect 384670 266999 384672 267008
rect 384488 266970 384540 266976
rect 384724 266999 384726 267008
rect 384672 266970 384724 266976
rect 384960 266626 384988 270263
rect 384948 266620 385000 266626
rect 384948 266562 385000 266568
rect 385408 266620 385460 266626
rect 385408 266562 385460 266568
rect 384304 266484 384356 266490
rect 384304 266426 384356 266432
rect 384672 265668 384724 265674
rect 384672 265610 384724 265616
rect 384684 264316 384712 265610
rect 385420 264316 385448 266562
rect 386144 264988 386196 264994
rect 386144 264930 386196 264936
rect 386156 264316 386184 264930
rect 387352 264330 387380 276762
rect 388640 276010 388668 277780
rect 388628 276004 388680 276010
rect 388628 275946 388680 275952
rect 388996 276004 389048 276010
rect 388996 275946 389048 275952
rect 387800 272944 387852 272950
rect 387800 272886 387852 272892
rect 387616 268252 387668 268258
rect 387616 268194 387668 268200
rect 386906 264302 387380 264330
rect 387628 264316 387656 268194
rect 387812 267034 387840 272886
rect 389008 267850 389036 275946
rect 389744 273970 389772 277780
rect 390572 277766 390954 277794
rect 390284 274508 390336 274514
rect 390284 274450 390336 274456
rect 389732 273964 389784 273970
rect 389732 273906 389784 273912
rect 389824 271176 389876 271182
rect 389824 271118 389876 271124
rect 388996 267844 389048 267850
rect 388996 267786 389048 267792
rect 388996 267300 389048 267306
rect 388996 267242 389048 267248
rect 389008 267073 389036 267242
rect 388994 267064 389050 267073
rect 387800 267028 387852 267034
rect 387800 266970 387852 266976
rect 388352 267028 388404 267034
rect 388994 266999 389050 267008
rect 388352 266970 388404 266976
rect 388364 264316 388392 266970
rect 389836 266626 389864 271118
rect 389824 266620 389876 266626
rect 389824 266562 389876 266568
rect 389088 265940 389140 265946
rect 389088 265882 389140 265888
rect 389100 264316 389128 265882
rect 390296 264330 390324 274450
rect 390572 269958 390600 277766
rect 392136 275466 392164 277780
rect 392124 275460 392176 275466
rect 392124 275402 392176 275408
rect 392308 275460 392360 275466
rect 392308 275402 392360 275408
rect 391848 273964 391900 273970
rect 391848 273906 391900 273912
rect 390560 269952 390612 269958
rect 390560 269894 390612 269900
rect 390744 269952 390796 269958
rect 390744 269894 390796 269900
rect 390756 266898 390784 269894
rect 390744 266892 390796 266898
rect 390744 266834 390796 266840
rect 391296 266892 391348 266898
rect 391296 266834 391348 266840
rect 390560 266620 390612 266626
rect 390560 266562 390612 266568
rect 389850 264302 390324 264330
rect 390572 264316 390600 266562
rect 391308 264316 391336 266834
rect 391860 266626 391888 273906
rect 392320 273426 392348 275402
rect 393332 274922 393360 277780
rect 393700 277766 394542 277794
rect 393320 274916 393372 274922
rect 393320 274858 393372 274864
rect 393228 274372 393280 274378
rect 393228 274314 393280 274320
rect 392308 273420 392360 273426
rect 392308 273362 392360 273368
rect 393240 267442 393268 274314
rect 393504 270224 393556 270230
rect 393504 270166 393556 270172
rect 393516 269906 393544 270166
rect 393700 270094 393728 277766
rect 394608 275596 394660 275602
rect 394608 275538 394660 275544
rect 394332 274236 394384 274242
rect 394332 274178 394384 274184
rect 393872 270224 393924 270230
rect 393872 270166 393924 270172
rect 393688 270088 393740 270094
rect 393688 270030 393740 270036
rect 393516 269878 393636 269906
rect 393608 269414 393636 269878
rect 393412 269408 393464 269414
rect 393412 269350 393464 269356
rect 393596 269408 393648 269414
rect 393596 269350 393648 269356
rect 393424 269249 393452 269350
rect 393410 269240 393466 269249
rect 393410 269175 393466 269184
rect 392032 267436 392084 267442
rect 392032 267378 392084 267384
rect 393228 267436 393280 267442
rect 393228 267378 393280 267384
rect 393412 267436 393464 267442
rect 393412 267378 393464 267384
rect 391848 266620 391900 266626
rect 391848 266562 391900 266568
rect 392044 264316 392072 267378
rect 393424 267322 393452 267378
rect 393148 267294 393452 267322
rect 393148 267034 393176 267294
rect 393318 267064 393374 267073
rect 393136 267028 393188 267034
rect 393318 266999 393320 267008
rect 393136 266970 393188 266976
rect 393372 266999 393374 267008
rect 393320 266970 393372 266976
rect 392216 266892 392268 266898
rect 392216 266834 392268 266840
rect 392768 266892 392820 266898
rect 392768 266834 392820 266840
rect 392228 266626 392256 266834
rect 392216 266620 392268 266626
rect 392216 266562 392268 266568
rect 392780 264316 392808 266834
rect 393884 264330 393912 270166
rect 394344 267734 394372 274178
rect 394620 273970 394648 275538
rect 395724 274106 395752 277780
rect 396920 275466 396948 277780
rect 397564 277766 398038 277794
rect 396908 275460 396960 275466
rect 396908 275402 396960 275408
rect 397092 275460 397144 275466
rect 397092 275402 397144 275408
rect 397104 274258 397132 275402
rect 397368 274916 397420 274922
rect 397368 274858 397420 274864
rect 396920 274230 397132 274258
rect 395712 274100 395764 274106
rect 395712 274042 395764 274048
rect 394608 273964 394660 273970
rect 394608 273906 394660 273912
rect 396724 273964 396776 273970
rect 396724 273906 396776 273912
rect 395436 273352 395488 273358
rect 395436 273294 395488 273300
rect 393530 264302 393912 264330
rect 394252 267706 394372 267734
rect 394252 264316 394280 267706
rect 395448 264330 395476 273294
rect 395988 270088 396040 270094
rect 395988 270030 396040 270036
rect 396000 264330 396028 270030
rect 396736 266762 396764 273906
rect 396920 273358 396948 274230
rect 397184 274100 397236 274106
rect 397184 274042 397236 274048
rect 396908 273352 396960 273358
rect 396908 273294 396960 273300
rect 397196 267734 397224 274042
rect 397380 273834 397408 274858
rect 397368 273828 397420 273834
rect 397368 273770 397420 273776
rect 397564 269822 397592 277766
rect 399220 275330 399248 277780
rect 399208 275324 399260 275330
rect 399208 275266 399260 275272
rect 399852 275324 399904 275330
rect 399852 275266 399904 275272
rect 398748 273828 398800 273834
rect 398748 273770 398800 273776
rect 398472 270224 398524 270230
rect 398472 270166 398524 270172
rect 397552 269816 397604 269822
rect 397552 269758 397604 269764
rect 398484 269498 398512 270166
rect 398300 269470 398512 269498
rect 398300 269414 398328 269470
rect 398288 269408 398340 269414
rect 398288 269350 398340 269356
rect 398472 269408 398524 269414
rect 398472 269350 398524 269356
rect 398104 269068 398156 269074
rect 398104 269010 398156 269016
rect 398288 269068 398340 269074
rect 398288 269010 398340 269016
rect 398116 268258 398144 269010
rect 397920 268252 397972 268258
rect 397920 268194 397972 268200
rect 398104 268252 398156 268258
rect 398104 268194 398156 268200
rect 397932 268138 397960 268194
rect 398300 268138 398328 269010
rect 397932 268110 398328 268138
rect 398484 267734 398512 269350
rect 398760 267734 398788 273770
rect 396920 267706 397224 267734
rect 398392 267706 398512 267734
rect 398668 267706 398788 267734
rect 396724 266756 396776 266762
rect 396724 266698 396776 266704
rect 396920 264330 396948 267706
rect 397184 266756 397236 266762
rect 397184 266698 397236 266704
rect 395002 264302 395476 264330
rect 395738 264302 396028 264330
rect 396474 264302 396948 264330
rect 397196 264316 397224 266698
rect 398392 264330 398420 267706
rect 397946 264302 398420 264330
rect 398668 264316 398696 267706
rect 399864 264330 399892 275266
rect 400416 274650 400444 277780
rect 401626 277766 401916 277794
rect 400404 274644 400456 274650
rect 400404 274586 400456 274592
rect 401324 274644 401376 274650
rect 401324 274586 401376 274592
rect 400126 269784 400182 269793
rect 400126 269719 400182 269728
rect 399418 264302 399892 264330
rect 400140 264316 400168 269719
rect 401138 267200 401194 267209
rect 401138 267135 401194 267144
rect 401152 266490 401180 267135
rect 401140 266484 401192 266490
rect 401140 266426 401192 266432
rect 401336 264330 401364 274586
rect 401888 270230 401916 277766
rect 402440 277766 402822 277794
rect 401876 270224 401928 270230
rect 401876 270166 401928 270172
rect 402244 270224 402296 270230
rect 402244 270166 402296 270172
rect 402256 267170 402284 270166
rect 402440 269249 402468 277766
rect 402796 276140 402848 276146
rect 402796 276082 402848 276088
rect 402426 269240 402482 269249
rect 402426 269175 402482 269184
rect 402612 267980 402664 267986
rect 402612 267922 402664 267928
rect 402624 267209 402652 267922
rect 402610 267200 402666 267209
rect 402244 267164 402296 267170
rect 402610 267135 402666 267144
rect 402244 267106 402296 267112
rect 402808 267016 402836 276082
rect 404004 275194 404032 277780
rect 404464 277766 405214 277794
rect 406120 277766 406318 277794
rect 403992 275188 404044 275194
rect 403992 275130 404044 275136
rect 404268 275188 404320 275194
rect 404268 275130 404320 275136
rect 404280 273698 404308 275130
rect 404268 273692 404320 273698
rect 404268 273634 404320 273640
rect 403992 270632 404044 270638
rect 403990 270600 403992 270609
rect 404176 270632 404228 270638
rect 404044 270600 404046 270609
rect 404176 270574 404228 270580
rect 403990 270535 404046 270544
rect 402980 267164 403032 267170
rect 402980 267106 403032 267112
rect 402348 266988 402836 267016
rect 401600 266484 401652 266490
rect 401600 266426 401652 266432
rect 400890 264302 401364 264330
rect 401612 264316 401640 266426
rect 402348 264316 402376 266988
rect 402992 266914 403020 267106
rect 402624 266886 403020 266914
rect 402624 266490 402652 266886
rect 404188 266762 404216 270574
rect 404464 267850 404492 277766
rect 405556 273692 405608 273698
rect 405556 273634 405608 273640
rect 404452 267844 404504 267850
rect 404452 267786 404504 267792
rect 402796 266756 402848 266762
rect 402796 266698 402848 266704
rect 403072 266756 403124 266762
rect 403072 266698 403124 266704
rect 404176 266756 404228 266762
rect 404176 266698 404228 266704
rect 402808 266490 402836 266698
rect 402612 266484 402664 266490
rect 402612 266426 402664 266432
rect 402796 266484 402848 266490
rect 402796 266426 402848 266432
rect 403084 264316 403112 266698
rect 404176 266076 404228 266082
rect 404176 266018 404228 266024
rect 404188 264330 404216 266018
rect 404544 265532 404596 265538
rect 404544 265474 404596 265480
rect 403834 264302 404216 264330
rect 404556 264316 404584 265474
rect 405568 264330 405596 273634
rect 406120 269278 406148 277766
rect 406108 269272 406160 269278
rect 406108 269214 406160 269220
rect 406016 266756 406068 266762
rect 406016 266698 406068 266704
rect 405306 264302 405596 264330
rect 406028 264316 406056 266698
rect 406948 264330 406976 278666
rect 590580 278594 590778 278610
rect 467564 278588 467616 278594
rect 467564 278530 467616 278536
rect 476488 278588 476540 278594
rect 476488 278530 476540 278536
rect 482284 278588 482336 278594
rect 482284 278530 482336 278536
rect 590568 278588 590778 278594
rect 590620 278582 590778 278588
rect 590568 278530 590620 278536
rect 437204 277840 437256 277846
rect 407500 275874 407528 277780
rect 407488 275868 407540 275874
rect 407488 275810 407540 275816
rect 408696 275058 408724 277780
rect 409328 277092 409380 277098
rect 409328 277034 409380 277040
rect 408684 275052 408736 275058
rect 408684 274994 408736 275000
rect 408868 275052 408920 275058
rect 408868 274994 408920 275000
rect 408880 274938 408908 274994
rect 408328 274910 408908 274938
rect 408328 270494 408356 274910
rect 408500 274780 408552 274786
rect 408500 274722 408552 274728
rect 408512 270609 408540 274722
rect 408498 270600 408554 270609
rect 408498 270535 408554 270544
rect 408328 270466 408448 270494
rect 407948 269816 408000 269822
rect 407948 269758 408000 269764
rect 408132 269816 408184 269822
rect 408132 269758 408184 269764
rect 407960 269550 407988 269758
rect 407948 269544 408000 269550
rect 407948 269486 408000 269492
rect 408144 269278 408172 269758
rect 408420 269362 408448 270466
rect 408420 269334 408540 269362
rect 408132 269272 408184 269278
rect 408132 269214 408184 269220
rect 408316 269272 408368 269278
rect 408316 269214 408368 269220
rect 407396 268388 407448 268394
rect 407396 268330 407448 268336
rect 407408 267850 407436 268330
rect 407948 268252 408000 268258
rect 407948 268194 408000 268200
rect 407960 267986 407988 268194
rect 407948 267980 408000 267986
rect 407948 267922 408000 267928
rect 407396 267844 407448 267850
rect 407396 267786 407448 267792
rect 408328 267734 408356 269214
rect 408512 269192 408540 269334
rect 407960 267706 408356 267734
rect 408420 269164 408540 269192
rect 407960 264330 407988 267706
rect 408420 264330 408448 269164
rect 409340 264330 409368 277034
rect 409892 272134 409920 277780
rect 410064 275868 410116 275874
rect 410064 275810 410116 275816
rect 409880 272128 409932 272134
rect 409880 272070 409932 272076
rect 409512 270632 409564 270638
rect 409512 270574 409564 270580
rect 409696 270632 409748 270638
rect 409696 270574 409748 270580
rect 409524 270473 409552 270574
rect 409510 270464 409566 270473
rect 409510 270399 409566 270408
rect 406778 264302 406976 264330
rect 407514 264302 407988 264330
rect 408250 264302 408448 264330
rect 408986 264302 409368 264330
rect 409708 264316 409736 270574
rect 410076 267850 410104 275810
rect 411088 275738 411116 277780
rect 411076 275732 411128 275738
rect 411076 275674 411128 275680
rect 412284 274786 412312 277780
rect 413388 277394 413416 277780
rect 413652 277568 413704 277574
rect 413652 277510 413704 277516
rect 413296 277366 413416 277394
rect 412456 275052 412508 275058
rect 412456 274994 412508 275000
rect 412468 274786 412496 274994
rect 412272 274780 412324 274786
rect 412272 274722 412324 274728
rect 412456 274780 412508 274786
rect 412456 274722 412508 274728
rect 412272 272128 412324 272134
rect 412272 272070 412324 272076
rect 410708 271992 410760 271998
rect 410708 271934 410760 271940
rect 410064 267844 410116 267850
rect 410064 267786 410116 267792
rect 410248 267844 410300 267850
rect 410248 267786 410300 267792
rect 410260 266762 410288 267786
rect 410720 267714 410748 271934
rect 412088 270768 412140 270774
rect 412086 270736 412088 270745
rect 412140 270736 412142 270745
rect 412086 270671 412142 270680
rect 411168 267980 411220 267986
rect 411168 267922 411220 267928
rect 410708 267708 410760 267714
rect 410708 267650 410760 267656
rect 410248 266756 410300 266762
rect 410248 266698 410300 266704
rect 410432 266756 410484 266762
rect 410432 266698 410484 266704
rect 410444 264316 410472 266698
rect 411180 264316 411208 267922
rect 412284 267734 412312 272070
rect 412638 271144 412694 271153
rect 412638 271079 412694 271088
rect 412652 270994 412680 271079
rect 412606 270966 412680 270994
rect 412606 270910 412634 270966
rect 412594 270904 412646 270910
rect 412594 270846 412646 270852
rect 412732 270904 412784 270910
rect 412732 270846 412784 270852
rect 412456 270768 412508 270774
rect 412744 270745 412772 270846
rect 412456 270710 412508 270716
rect 412730 270736 412786 270745
rect 412468 270473 412496 270710
rect 412730 270671 412786 270680
rect 412454 270464 412510 270473
rect 412454 270399 412510 270408
rect 412606 270286 412956 270314
rect 412606 270230 412634 270286
rect 412594 270224 412646 270230
rect 412594 270166 412646 270172
rect 412732 270224 412784 270230
rect 412732 270166 412784 270172
rect 412928 270178 412956 270286
rect 412744 270065 412772 270166
rect 412928 270150 413140 270178
rect 412454 270056 412510 270065
rect 412454 269991 412510 270000
rect 412730 270056 412786 270065
rect 412730 269991 412786 270000
rect 412468 269278 412496 269991
rect 413112 269686 413140 270150
rect 412732 269680 412784 269686
rect 412732 269622 412784 269628
rect 413100 269680 413152 269686
rect 413100 269622 413152 269628
rect 412744 269278 412772 269622
rect 413296 269498 413324 277366
rect 412928 269470 413324 269498
rect 412928 269414 412956 269470
rect 412916 269408 412968 269414
rect 412916 269350 412968 269356
rect 413100 269408 413152 269414
rect 413100 269350 413152 269356
rect 412456 269272 412508 269278
rect 412456 269214 412508 269220
rect 412732 269272 412784 269278
rect 412732 269214 412784 269220
rect 412284 267706 412404 267734
rect 411994 267608 412050 267617
rect 411994 267543 411996 267552
rect 412048 267543 412050 267552
rect 412180 267572 412232 267578
rect 411996 267514 412048 267520
rect 412180 267514 412232 267520
rect 412192 266778 412220 267514
rect 412376 266914 412404 267706
rect 412730 267608 412786 267617
rect 412594 267572 412646 267578
rect 412730 267543 412732 267552
rect 412594 267514 412646 267520
rect 412784 267543 412786 267552
rect 412732 267514 412784 267520
rect 412606 267458 412634 267514
rect 412606 267430 412680 267458
rect 412652 267345 412680 267430
rect 412638 267336 412694 267345
rect 412638 267271 412694 267280
rect 412100 266762 412220 266778
rect 412088 266756 412220 266762
rect 412140 266750 412220 266756
rect 412284 266886 412404 266914
rect 412088 266698 412140 266704
rect 412284 264330 412312 266886
rect 412456 266756 412508 266762
rect 412456 266698 412508 266704
rect 412468 266082 412496 266698
rect 412456 266076 412508 266082
rect 412456 266018 412508 266024
rect 413112 264330 413140 269350
rect 413664 264330 413692 277510
rect 414204 275732 414256 275738
rect 414204 275674 414256 275680
rect 414020 275052 414072 275058
rect 414020 274994 414072 275000
rect 414032 270910 414060 274994
rect 414020 270904 414072 270910
rect 414020 270846 414072 270852
rect 414216 269498 414244 275674
rect 414584 274922 414612 277780
rect 415780 275058 415808 277780
rect 416792 277766 416990 277794
rect 415768 275052 415820 275058
rect 415768 274994 415820 275000
rect 414572 274916 414624 274922
rect 414572 274858 414624 274864
rect 416136 273420 416188 273426
rect 416136 273362 416188 273368
rect 414664 270904 414716 270910
rect 414664 270846 414716 270852
rect 413940 269470 414244 269498
rect 413940 269414 413968 269470
rect 413928 269408 413980 269414
rect 413928 269350 413980 269356
rect 414112 269408 414164 269414
rect 414112 269350 414164 269356
rect 411930 264302 412312 264330
rect 412666 264302 413140 264330
rect 413402 264302 413692 264330
rect 414124 264316 414152 269350
rect 414676 267578 414704 270846
rect 415490 267880 415546 267889
rect 415308 267844 415360 267850
rect 415490 267815 415546 267824
rect 415308 267786 415360 267792
rect 415320 267714 415348 267786
rect 415308 267708 415360 267714
rect 415308 267650 415360 267656
rect 415122 267608 415178 267617
rect 414664 267572 414716 267578
rect 415122 267543 415178 267552
rect 415308 267572 415360 267578
rect 414664 267514 414716 267520
rect 415136 264330 415164 267543
rect 415308 267514 415360 267520
rect 415320 266762 415348 267514
rect 415504 267306 415532 267815
rect 415492 267300 415544 267306
rect 415492 267242 415544 267248
rect 415308 266756 415360 266762
rect 415308 266698 415360 266704
rect 415584 266756 415636 266762
rect 415584 266698 415636 266704
rect 414874 264302 415164 264330
rect 415596 264316 415624 266698
rect 416148 264330 416176 273362
rect 416792 269498 416820 277766
rect 418172 276010 418200 277780
rect 419000 277766 419382 277794
rect 418160 276004 418212 276010
rect 418160 275946 418212 275952
rect 418344 276004 418396 276010
rect 418344 275946 418396 275952
rect 418068 274916 418120 274922
rect 418068 274858 418120 274864
rect 417240 272400 417292 272406
rect 417240 272342 417292 272348
rect 417252 272116 417280 272342
rect 417700 272128 417752 272134
rect 417252 272088 417700 272116
rect 417700 272070 417752 272076
rect 417240 270904 417292 270910
rect 417240 270846 417292 270852
rect 417252 270609 417280 270846
rect 417238 270600 417294 270609
rect 417238 270535 417294 270544
rect 416424 269470 416820 269498
rect 416424 269278 416452 269470
rect 416412 269272 416464 269278
rect 416412 269214 416464 269220
rect 416688 269204 416740 269210
rect 416688 269146 416740 269152
rect 416318 267336 416374 267345
rect 416318 267271 416374 267280
rect 416332 267170 416360 267271
rect 416320 267164 416372 267170
rect 416320 267106 416372 267112
rect 416700 266762 416728 269146
rect 417424 268388 417476 268394
rect 417424 268330 417476 268336
rect 417608 268388 417660 268394
rect 417608 268330 417660 268336
rect 417054 268152 417110 268161
rect 417054 268087 417110 268096
rect 416688 266756 416740 266762
rect 416688 266698 416740 266704
rect 416148 264302 416346 264330
rect 417068 264316 417096 268087
rect 417436 267986 417464 268330
rect 417424 267980 417476 267986
rect 417424 267922 417476 267928
rect 417620 267850 417648 268330
rect 418080 268161 418108 274858
rect 418356 272134 418384 275946
rect 418344 272128 418396 272134
rect 418344 272070 418396 272076
rect 419000 271153 419028 277766
rect 420368 276412 420420 276418
rect 420368 276354 420420 276360
rect 418986 271144 419042 271153
rect 418986 271079 419042 271088
rect 418252 270768 418304 270774
rect 418252 270710 418304 270716
rect 418894 270736 418950 270745
rect 418264 270609 418292 270710
rect 418894 270671 418950 270680
rect 418250 270600 418306 270609
rect 418250 270535 418306 270544
rect 418066 268152 418122 268161
rect 418066 268087 418122 268096
rect 417790 267880 417846 267889
rect 417608 267844 417660 267850
rect 417790 267815 417792 267824
rect 417608 267786 417660 267792
rect 417844 267815 417846 267824
rect 417792 267786 417844 267792
rect 418342 267744 418398 267753
rect 417884 267708 417936 267714
rect 418342 267679 418344 267688
rect 417884 267650 417936 267656
rect 418396 267679 418398 267688
rect 418344 267650 418396 267656
rect 417896 266642 417924 267650
rect 418252 266756 418304 266762
rect 418252 266698 418304 266704
rect 418264 266642 418292 266698
rect 417896 266614 418292 266642
rect 417792 265260 417844 265266
rect 417792 265202 417844 265208
rect 417804 264316 417832 265202
rect 418908 264330 418936 270671
rect 419262 267336 419318 267345
rect 419262 267271 419318 267280
rect 418554 264302 418936 264330
rect 419276 264316 419304 267271
rect 420380 264330 420408 276354
rect 420564 273562 420592 277780
rect 421668 275874 421696 277780
rect 422496 277766 422878 277794
rect 423692 277766 424074 277794
rect 421932 277704 421984 277710
rect 421932 277646 421984 277652
rect 421656 275868 421708 275874
rect 421656 275810 421708 275816
rect 420552 273556 420604 273562
rect 420552 273498 420604 273504
rect 420734 269512 420790 269521
rect 420734 269447 420790 269456
rect 420026 264302 420408 264330
rect 420748 264316 420776 269447
rect 421102 267608 421158 267617
rect 421102 267543 421158 267552
rect 421472 267572 421524 267578
rect 421116 267442 421144 267543
rect 421472 267514 421524 267520
rect 421104 267436 421156 267442
rect 421104 267378 421156 267384
rect 421484 264316 421512 267514
rect 421944 264330 421972 277646
rect 422116 275052 422168 275058
rect 422116 274994 422168 275000
rect 422128 267578 422156 274994
rect 422496 271046 422524 277766
rect 423496 271992 423548 271998
rect 423496 271934 423548 271940
rect 422760 271720 422812 271726
rect 422812 271668 423352 271674
rect 422760 271662 423352 271668
rect 422772 271646 423352 271662
rect 423128 271584 423180 271590
rect 423128 271526 423180 271532
rect 422484 271040 422536 271046
rect 422484 270982 422536 270988
rect 423140 270774 423168 271526
rect 423324 270910 423352 271646
rect 423312 270904 423364 270910
rect 423312 270846 423364 270852
rect 423128 270768 423180 270774
rect 423312 270768 423364 270774
rect 423128 270710 423180 270716
rect 423310 270736 423312 270745
rect 423364 270736 423366 270745
rect 423310 270671 423366 270680
rect 422576 269544 422628 269550
rect 422628 269492 423168 269498
rect 422576 269486 423168 269492
rect 422588 269470 423168 269486
rect 423140 269414 423168 269470
rect 423128 269408 423180 269414
rect 423128 269350 423180 269356
rect 422300 267844 422352 267850
rect 422300 267786 422352 267792
rect 422944 267844 422996 267850
rect 422944 267786 422996 267792
rect 422312 267578 422340 267786
rect 422116 267572 422168 267578
rect 422116 267514 422168 267520
rect 422300 267572 422352 267578
rect 422300 267514 422352 267520
rect 421944 264302 422234 264330
rect 422956 264316 422984 267786
rect 423508 267578 423536 271934
rect 423692 269414 423720 277766
rect 425256 275194 425284 277780
rect 426072 275868 426124 275874
rect 426072 275810 426124 275816
rect 425244 275188 425296 275194
rect 425244 275130 425296 275136
rect 425428 275188 425480 275194
rect 425428 275130 425480 275136
rect 425440 275074 425468 275130
rect 424336 275046 425468 275074
rect 424336 273254 424364 275046
rect 424244 273226 424364 273254
rect 423680 269408 423732 269414
rect 423680 269350 423732 269356
rect 424244 267617 424272 273226
rect 424416 269408 424468 269414
rect 424416 269350 424468 269356
rect 424230 267608 424286 267617
rect 423496 267572 423548 267578
rect 423496 267514 423548 267520
rect 423680 267572 423732 267578
rect 424230 267543 424286 267552
rect 423680 267514 423732 267520
rect 423692 264316 423720 267514
rect 424428 264316 424456 269350
rect 424966 267608 425022 267617
rect 424966 267543 424968 267552
rect 425020 267543 425022 267552
rect 425152 267572 425204 267578
rect 424968 267514 425020 267520
rect 425152 267514 425204 267520
rect 425164 264316 425192 267514
rect 426084 264330 426112 275810
rect 426256 273556 426308 273562
rect 426256 273498 426308 273504
rect 426268 267578 426296 273498
rect 426452 270910 426480 277780
rect 427648 276010 427676 277780
rect 428200 277766 428858 277794
rect 429212 277766 429962 277794
rect 430776 277766 431158 277794
rect 432064 277766 432354 277794
rect 433352 277766 433550 277794
rect 427636 276004 427688 276010
rect 427636 275946 427688 275952
rect 428004 275868 428056 275874
rect 428004 275810 428056 275816
rect 428016 275194 428044 275810
rect 428004 275188 428056 275194
rect 428004 275130 428056 275136
rect 428200 273254 428228 277766
rect 428200 273226 428412 273254
rect 427818 272368 427874 272377
rect 427818 272303 427874 272312
rect 427832 272218 427860 272303
rect 427786 272190 427860 272218
rect 427786 272134 427814 272190
rect 427774 272128 427826 272134
rect 427774 272070 427826 272076
rect 427912 272128 427964 272134
rect 427912 272070 427964 272076
rect 427084 271992 427136 271998
rect 427082 271960 427084 271969
rect 427268 271992 427320 271998
rect 427136 271960 427138 271969
rect 427924 271969 427952 272070
rect 427268 271934 427320 271940
rect 427910 271960 427966 271969
rect 427082 271895 427138 271904
rect 426440 270904 426492 270910
rect 426440 270846 426492 270852
rect 426992 270768 427044 270774
rect 426992 270710 427044 270716
rect 426256 267572 426308 267578
rect 426256 267514 426308 267520
rect 426440 267572 426492 267578
rect 426440 267514 426492 267520
rect 426452 267170 426480 267514
rect 426440 267164 426492 267170
rect 426440 267106 426492 267112
rect 426624 267164 426676 267170
rect 426624 267106 426676 267112
rect 426636 266762 426664 267106
rect 426624 266756 426676 266762
rect 426624 266698 426676 266704
rect 427004 264330 427032 270710
rect 425914 264302 426112 264330
rect 426650 264302 427032 264330
rect 427280 264330 427308 271934
rect 427910 271895 427966 271904
rect 428188 271720 428240 271726
rect 428186 271688 428188 271697
rect 428240 271688 428242 271697
rect 428186 271623 428242 271632
rect 427818 270056 427874 270065
rect 427818 269991 427874 270000
rect 427832 269686 427860 269991
rect 427820 269680 427872 269686
rect 427820 269622 427872 269628
rect 428004 269680 428056 269686
rect 428004 269622 428056 269628
rect 427450 269512 427506 269521
rect 427506 269470 427860 269498
rect 427450 269447 427506 269456
rect 427832 269414 427860 269470
rect 427636 269408 427688 269414
rect 427636 269350 427688 269356
rect 427820 269408 427872 269414
rect 427820 269350 427872 269356
rect 427648 269249 427676 269350
rect 428016 269249 428044 269622
rect 427634 269240 427690 269249
rect 427634 269175 427690 269184
rect 428002 269240 428058 269249
rect 428002 269175 428058 269184
rect 427634 268152 427690 268161
rect 427634 268087 427690 268096
rect 427818 268152 427874 268161
rect 427818 268087 427874 268096
rect 427648 267986 427676 268087
rect 427832 267986 427860 268087
rect 427636 267980 427688 267986
rect 427636 267922 427688 267928
rect 427820 267980 427872 267986
rect 427820 267922 427872 267928
rect 427910 267608 427966 267617
rect 427774 267572 427826 267578
rect 427910 267543 427912 267552
rect 427774 267514 427826 267520
rect 427964 267543 427966 267552
rect 427912 267514 427964 267520
rect 427786 267458 427814 267514
rect 427786 267430 427952 267458
rect 427924 266626 427952 267430
rect 427912 266620 427964 266626
rect 427912 266562 427964 266568
rect 428384 265962 428412 273226
rect 428556 271856 428608 271862
rect 428556 271798 428608 271804
rect 428568 271318 428596 271798
rect 429212 271726 429240 277766
rect 430580 275188 430632 275194
rect 430580 275130 430632 275136
rect 429200 271720 429252 271726
rect 429384 271720 429436 271726
rect 429200 271662 429252 271668
rect 429382 271688 429384 271697
rect 429436 271688 429438 271697
rect 429382 271623 429438 271632
rect 429106 271416 429162 271425
rect 429106 271351 429162 271360
rect 428556 271312 428608 271318
rect 428556 271254 428608 271260
rect 428554 266928 428610 266937
rect 428554 266863 428610 266872
rect 428292 265934 428412 265962
rect 428292 265810 428320 265934
rect 428280 265804 428332 265810
rect 428280 265746 428332 265752
rect 428568 264330 428596 266863
rect 429120 264330 429148 271351
rect 430592 270586 430620 275130
rect 430776 273222 430804 277766
rect 430764 273216 430816 273222
rect 430764 273158 430816 273164
rect 430948 273216 431000 273222
rect 430948 273158 431000 273164
rect 430960 272377 430988 273158
rect 430946 272368 431002 272377
rect 430946 272303 431002 272312
rect 431774 271688 431830 271697
rect 431774 271623 431830 271632
rect 431406 271008 431462 271017
rect 431406 270943 431462 270952
rect 430500 270558 430620 270586
rect 429566 269512 429622 269521
rect 429566 269447 429622 269456
rect 427280 264302 427386 264330
rect 428122 264302 428596 264330
rect 428858 264302 429148 264330
rect 429580 264316 429608 269447
rect 430500 264330 430528 270558
rect 431224 267164 431276 267170
rect 431224 267106 431276 267112
rect 431236 267050 431264 267106
rect 430684 267034 431264 267050
rect 430672 267028 431264 267034
rect 430724 267022 431264 267028
rect 430672 266970 430724 266976
rect 431420 264330 431448 270943
rect 430330 264302 430528 264330
rect 431066 264302 431448 264330
rect 431788 264316 431816 271623
rect 432064 268122 432092 277766
rect 433154 272776 433210 272785
rect 433154 272711 433210 272720
rect 432604 271584 432656 271590
rect 432604 271526 432656 271532
rect 432788 271584 432840 271590
rect 432788 271526 432840 271532
rect 432616 271318 432644 271526
rect 432604 271312 432656 271318
rect 432604 271254 432656 271260
rect 432800 271046 432828 271526
rect 432788 271040 432840 271046
rect 432972 271040 433024 271046
rect 432788 270982 432840 270988
rect 432970 271008 432972 271017
rect 433024 271008 433026 271017
rect 432970 270943 433026 270952
rect 432604 268524 432656 268530
rect 432604 268466 432656 268472
rect 432616 268122 432644 268466
rect 432052 268116 432104 268122
rect 432052 268058 432104 268064
rect 432604 268116 432656 268122
rect 432604 268058 432656 268064
rect 433168 267866 433196 272711
rect 433352 271726 433380 277766
rect 434732 277394 434760 277780
rect 435192 277766 435942 277794
rect 436112 277766 437046 277794
rect 437204 277782 437256 277788
rect 434732 277366 434852 277394
rect 434442 274000 434498 274009
rect 434442 273935 434498 273944
rect 433340 271720 433392 271726
rect 433340 271662 433392 271668
rect 433524 271720 433576 271726
rect 433524 271662 433576 271668
rect 433536 271425 433564 271662
rect 433522 271416 433578 271425
rect 433522 271351 433578 271360
rect 432984 267838 433196 267866
rect 432604 266348 432656 266354
rect 432604 266290 432656 266296
rect 432616 266082 432644 266290
rect 432604 266076 432656 266082
rect 432604 266018 432656 266024
rect 432984 264330 433012 267838
rect 433246 267744 433302 267753
rect 433246 267679 433302 267688
rect 432538 264302 433012 264330
rect 433260 264316 433288 267679
rect 434456 264330 434484 273935
rect 434824 270065 434852 277366
rect 435192 273970 435220 277766
rect 435362 274000 435418 274009
rect 435180 273964 435232 273970
rect 435362 273935 435364 273944
rect 435180 273906 435232 273912
rect 435416 273935 435418 273944
rect 435364 273906 435416 273912
rect 436112 270502 436140 277766
rect 436744 276004 436796 276010
rect 436744 275946 436796 275952
rect 436928 276004 436980 276010
rect 436928 275946 436980 275952
rect 436756 275194 436784 275946
rect 436560 275188 436612 275194
rect 436560 275130 436612 275136
rect 436744 275188 436796 275194
rect 436744 275130 436796 275136
rect 436572 275074 436600 275130
rect 436940 275074 436968 275946
rect 436572 275046 436968 275074
rect 437216 273254 437244 277782
rect 437124 273226 437244 273254
rect 436928 273080 436980 273086
rect 436926 273048 436928 273057
rect 436980 273048 436982 273057
rect 436926 272983 436982 272992
rect 436100 270496 436152 270502
rect 436100 270438 436152 270444
rect 434810 270056 434866 270065
rect 434810 269991 434866 270000
rect 434720 268524 434772 268530
rect 434720 268466 434772 268472
rect 434732 267170 434760 268466
rect 436926 268424 436982 268433
rect 436926 268359 436982 268368
rect 436558 268016 436614 268025
rect 436558 267951 436614 267960
rect 434720 267164 434772 267170
rect 434720 267106 434772 267112
rect 436192 267164 436244 267170
rect 436192 267106 436244 267112
rect 435086 266248 435142 266257
rect 435086 266183 435142 266192
rect 435100 264330 435128 266183
rect 435456 264784 435508 264790
rect 435456 264726 435508 264732
rect 434010 264302 434484 264330
rect 434746 264302 435128 264330
rect 435468 264316 435496 264726
rect 436204 264316 436232 267106
rect 436572 266762 436600 267951
rect 436744 267028 436796 267034
rect 436744 266970 436796 266976
rect 436560 266756 436612 266762
rect 436560 266698 436612 266704
rect 436756 266529 436784 266970
rect 436742 266520 436798 266529
rect 436742 266455 436798 266464
rect 436940 264316 436968 268359
rect 437124 267170 437152 273226
rect 437434 273216 437486 273222
rect 437308 273164 437434 273170
rect 437308 273158 437486 273164
rect 437308 273142 437474 273158
rect 437308 272785 437336 273142
rect 438228 273057 438256 277780
rect 438872 277766 439438 277794
rect 438214 273048 438270 273057
rect 438214 272983 438270 272992
rect 437294 272776 437350 272785
rect 437294 272711 437350 272720
rect 438400 270496 438452 270502
rect 438400 270438 438452 270444
rect 437294 268696 437350 268705
rect 437294 268631 437296 268640
rect 437348 268631 437350 268640
rect 437434 268660 437486 268666
rect 437296 268602 437348 268608
rect 437434 268602 437486 268608
rect 437446 268546 437474 268602
rect 437308 268518 437474 268546
rect 437308 267986 437336 268518
rect 437296 267980 437348 267986
rect 437296 267922 437348 267928
rect 437434 267980 437486 267986
rect 437434 267922 437486 267928
rect 437446 267866 437474 267922
rect 437308 267838 437474 267866
rect 437308 267753 437336 267838
rect 437294 267744 437350 267753
rect 437294 267679 437350 267688
rect 437112 267164 437164 267170
rect 437112 267106 437164 267112
rect 437296 267164 437348 267170
rect 437296 267106 437348 267112
rect 437112 267028 437164 267034
rect 437112 266970 437164 266976
rect 437124 266626 437152 266970
rect 437308 266937 437336 267106
rect 437294 266928 437350 266937
rect 437294 266863 437350 266872
rect 437940 266756 437992 266762
rect 437940 266698 437992 266704
rect 437112 266620 437164 266626
rect 437112 266562 437164 266568
rect 437952 266529 437980 266698
rect 437938 266520 437994 266529
rect 437756 266484 437808 266490
rect 437938 266455 437994 266464
rect 437756 266426 437808 266432
rect 437768 266257 437796 266426
rect 437754 266248 437810 266257
rect 437754 266183 437810 266192
rect 437664 265804 437716 265810
rect 437664 265746 437716 265752
rect 437676 264316 437704 265746
rect 438412 264316 438440 270438
rect 438872 268705 438900 277766
rect 440620 271862 440648 277780
rect 441632 277766 441830 277794
rect 441632 273086 441660 277766
rect 442540 277228 442592 277234
rect 442540 277170 442592 277176
rect 441620 273080 441672 273086
rect 441620 273022 441672 273028
rect 442080 273080 442132 273086
rect 442080 273022 442132 273028
rect 442092 272542 442120 273022
rect 442080 272536 442132 272542
rect 442080 272478 442132 272484
rect 441526 272096 441582 272105
rect 441526 272031 441582 272040
rect 440608 271856 440660 271862
rect 440608 271798 440660 271804
rect 440976 271856 441028 271862
rect 440976 271798 441028 271804
rect 440988 271318 441016 271798
rect 441158 271416 441214 271425
rect 441158 271351 441214 271360
rect 440976 271312 441028 271318
rect 440976 271254 441028 271260
rect 439502 271144 439558 271153
rect 439502 271079 439558 271088
rect 438858 268696 438914 268705
rect 438858 268631 438914 268640
rect 439516 264330 439544 271079
rect 440424 268796 440476 268802
rect 440424 268738 440476 268744
rect 440436 268122 440464 268738
rect 440884 268524 440936 268530
rect 440620 268484 440884 268512
rect 440240 268116 440292 268122
rect 440240 268058 440292 268064
rect 440424 268116 440476 268122
rect 440424 268058 440476 268064
rect 440252 268002 440280 268058
rect 440620 268002 440648 268484
rect 440884 268466 440936 268472
rect 440252 267974 440648 268002
rect 439872 265124 439924 265130
rect 439872 265066 439924 265072
rect 439162 264302 439544 264330
rect 439884 264316 439912 265066
rect 441172 264330 441200 271351
rect 441540 264330 441568 272031
rect 442264 271584 442316 271590
rect 442264 271526 442316 271532
rect 442276 271318 442304 271526
rect 442264 271312 442316 271318
rect 442264 271254 442316 271260
rect 442264 267436 442316 267442
rect 442264 267378 442316 267384
rect 442276 267170 442304 267378
rect 442080 267164 442132 267170
rect 442080 267106 442132 267112
rect 442264 267164 442316 267170
rect 442264 267106 442316 267112
rect 442092 266490 442120 267106
rect 442080 266484 442132 266490
rect 442080 266426 442132 266432
rect 441710 266384 441766 266393
rect 441710 266319 441712 266328
rect 441764 266319 441766 266328
rect 441712 266290 441764 266296
rect 442264 266076 442316 266082
rect 442264 266018 442316 266024
rect 442276 265538 442304 266018
rect 442264 265532 442316 265538
rect 442264 265474 442316 265480
rect 442080 265396 442132 265402
rect 442080 265338 442132 265344
rect 440634 264302 441200 264330
rect 441370 264302 441568 264330
rect 442092 264316 442120 265338
rect 442552 264330 442580 277170
rect 442724 272400 442776 272406
rect 442724 272342 442776 272348
rect 442736 272134 442764 272342
rect 442724 272128 442776 272134
rect 442724 272070 442776 272076
rect 442724 271584 442776 271590
rect 442724 271526 442776 271532
rect 442736 271425 442764 271526
rect 442722 271416 442778 271425
rect 442722 271351 442778 271360
rect 443012 268682 443040 277780
rect 442828 268654 443040 268682
rect 443196 277766 444222 277794
rect 444576 277766 445326 277794
rect 446140 277766 446522 277794
rect 442828 268530 442856 268654
rect 442816 268524 442868 268530
rect 442816 268466 442868 268472
rect 443000 268524 443052 268530
rect 443000 268466 443052 268472
rect 443012 268025 443040 268466
rect 442998 268016 443054 268025
rect 442998 267951 443054 267960
rect 442724 267436 442776 267442
rect 442724 267378 442776 267384
rect 442736 266354 442764 267378
rect 442906 266384 442962 266393
rect 442724 266348 442776 266354
rect 442906 266319 442908 266328
rect 442724 266290 442776 266296
rect 442960 266319 442962 266328
rect 442908 266290 442960 266296
rect 443196 266218 443224 277766
rect 443368 272128 443420 272134
rect 443366 272096 443368 272105
rect 443420 272096 443422 272105
rect 443366 272031 443422 272040
rect 444576 271862 444604 277766
rect 445482 275496 445538 275505
rect 445482 275431 445538 275440
rect 445496 273222 445524 275431
rect 446140 273254 446168 277766
rect 446312 276548 446364 276554
rect 446312 276490 446364 276496
rect 445956 273226 446168 273254
rect 445484 273216 445536 273222
rect 445484 273158 445536 273164
rect 445390 273048 445446 273057
rect 445390 272983 445446 272992
rect 444564 271856 444616 271862
rect 444564 271798 444616 271804
rect 444748 271856 444800 271862
rect 444748 271798 444800 271804
rect 444760 271153 444788 271798
rect 444746 271144 444802 271153
rect 444746 271079 444802 271088
rect 443184 266212 443236 266218
rect 443184 266154 443236 266160
rect 443920 266212 443972 266218
rect 443920 266154 443972 266160
rect 443932 264330 443960 266154
rect 444288 265532 444340 265538
rect 444288 265474 444340 265480
rect 442552 264302 442842 264330
rect 443578 264302 443960 264330
rect 444300 264316 444328 265474
rect 445404 264330 445432 272983
rect 445956 266354 445984 273226
rect 446128 273080 446180 273086
rect 446128 273022 446180 273028
rect 446140 272134 446168 273022
rect 446324 272814 446352 276490
rect 446956 276276 447008 276282
rect 446956 276218 447008 276224
rect 446312 272808 446364 272814
rect 446312 272750 446364 272756
rect 446772 272400 446824 272406
rect 446770 272368 446772 272377
rect 446824 272368 446826 272377
rect 446770 272303 446826 272312
rect 446128 272128 446180 272134
rect 446128 272070 446180 272076
rect 446126 271144 446182 271153
rect 446126 271079 446182 271088
rect 445944 266348 445996 266354
rect 445944 266290 445996 266296
rect 446140 264330 446168 271079
rect 446770 268696 446826 268705
rect 446770 268631 446826 268640
rect 446784 268258 446812 268631
rect 446772 268252 446824 268258
rect 446772 268194 446824 268200
rect 446770 267608 446826 267617
rect 446770 267543 446826 267552
rect 446588 267436 446640 267442
rect 446588 267378 446640 267384
rect 446600 266801 446628 267378
rect 446784 267306 446812 267543
rect 446772 267300 446824 267306
rect 446772 267242 446824 267248
rect 446770 267064 446826 267073
rect 446770 266999 446772 267008
rect 446824 266999 446826 267008
rect 446772 266970 446824 266976
rect 446586 266792 446642 266801
rect 446586 266727 446642 266736
rect 446968 264330 446996 276218
rect 447704 273222 447732 277780
rect 448532 277766 448914 277794
rect 449912 277766 450110 277794
rect 448150 274000 448206 274009
rect 448150 273935 448206 273944
rect 447692 273216 447744 273222
rect 447692 273158 447744 273164
rect 447230 273048 447286 273057
rect 447286 273006 447456 273034
rect 447230 272983 447286 272992
rect 447428 272950 447456 273006
rect 447416 272944 447468 272950
rect 447416 272886 447468 272892
rect 447416 272536 447468 272542
rect 447416 272478 447468 272484
rect 447428 272377 447456 272478
rect 447414 272368 447470 272377
rect 447414 272303 447470 272312
rect 447598 272368 447654 272377
rect 447598 272303 447654 272312
rect 447414 267608 447470 267617
rect 447414 267543 447470 267552
rect 447232 267436 447284 267442
rect 447232 267378 447284 267384
rect 447244 267073 447272 267378
rect 447428 267306 447456 267543
rect 447416 267300 447468 267306
rect 447416 267242 447468 267248
rect 447230 267064 447286 267073
rect 447230 266999 447286 267008
rect 447612 264330 447640 272303
rect 448164 264330 448192 273935
rect 448532 268705 448560 277766
rect 449714 273184 449770 273193
rect 449714 273119 449770 273128
rect 448702 270192 448758 270201
rect 448702 270127 448758 270136
rect 448518 268696 448574 268705
rect 448518 268631 448574 268640
rect 448716 266506 448744 270127
rect 448532 266478 448744 266506
rect 448532 266218 448560 266478
rect 448520 266212 448572 266218
rect 448520 266154 448572 266160
rect 448704 266212 448756 266218
rect 448704 266154 448756 266160
rect 445050 264302 445432 264330
rect 445786 264302 446168 264330
rect 446522 264302 446996 264330
rect 447258 264302 447640 264330
rect 447994 264302 448192 264330
rect 448716 264316 448744 266154
rect 449728 264330 449756 273119
rect 449912 268938 449940 277766
rect 451292 276554 451320 277780
rect 452120 277766 452502 277794
rect 452672 277766 453606 277794
rect 454236 277766 454802 277794
rect 451280 276548 451332 276554
rect 451280 276490 451332 276496
rect 451370 274000 451426 274009
rect 451234 273964 451286 273970
rect 451370 273935 451372 273944
rect 451234 273906 451286 273912
rect 451424 273935 451426 273944
rect 451372 273906 451424 273912
rect 451246 273850 451274 273906
rect 451246 273822 451412 273850
rect 451384 273290 451412 273822
rect 451096 273284 451148 273290
rect 451096 273226 451148 273232
rect 451234 273284 451286 273290
rect 451234 273226 451286 273232
rect 451372 273284 451424 273290
rect 451372 273226 451424 273232
rect 451108 272950 451136 273226
rect 451246 273170 451274 273226
rect 451246 273142 451320 273170
rect 451096 272944 451148 272950
rect 451096 272886 451148 272892
rect 451292 272134 451320 273142
rect 451924 272944 451976 272950
rect 451924 272886 451976 272892
rect 451280 272128 451332 272134
rect 451280 272070 451332 272076
rect 449900 268932 449952 268938
rect 449900 268874 449952 268880
rect 451936 268410 451964 272886
rect 452120 272814 452148 277766
rect 452108 272808 452160 272814
rect 452108 272750 452160 272756
rect 451568 268382 451964 268410
rect 450910 267064 450966 267073
rect 450910 266999 450966 267008
rect 450544 266348 450596 266354
rect 450544 266290 450596 266296
rect 450556 264330 450584 266290
rect 449466 264302 449756 264330
rect 450202 264302 450584 264330
rect 450924 264316 450952 266999
rect 451568 264330 451596 268382
rect 452384 268252 452436 268258
rect 452384 268194 452436 268200
rect 451924 267164 451976 267170
rect 451924 267106 451976 267112
rect 451936 266762 451964 267106
rect 451924 266756 451976 266762
rect 451924 266698 451976 266704
rect 452108 266756 452160 266762
rect 452108 266698 452160 266704
rect 452120 266354 452148 266698
rect 452108 266348 452160 266354
rect 452108 266290 452160 266296
rect 451568 264302 451674 264330
rect 452396 264316 452424 268194
rect 452672 268122 452700 277766
rect 453856 272808 453908 272814
rect 453856 272750 453908 272756
rect 452660 268116 452712 268122
rect 452660 268058 452712 268064
rect 453120 264648 453172 264654
rect 453120 264590 453172 264596
rect 453132 264316 453160 264590
rect 453868 264316 453896 272750
rect 454236 272406 454264 277766
rect 455984 277394 456012 277780
rect 455892 277366 456012 277394
rect 454590 274136 454646 274145
rect 454590 274071 454646 274080
rect 454224 272400 454276 272406
rect 454408 272400 454460 272406
rect 454224 272342 454276 272348
rect 454406 272368 454408 272377
rect 454460 272368 454462 272377
rect 454406 272303 454462 272312
rect 454604 266762 454632 274071
rect 455892 272542 455920 277366
rect 457180 276962 457208 277780
rect 457168 276956 457220 276962
rect 457168 276898 457220 276904
rect 456984 276548 457036 276554
rect 456984 276490 457036 276496
rect 456996 273254 457024 276490
rect 456996 273226 457300 273254
rect 456616 272944 456668 272950
rect 456616 272886 456668 272892
rect 456628 272785 456656 272886
rect 456614 272776 456670 272785
rect 456614 272711 456670 272720
rect 455880 272536 455932 272542
rect 455880 272478 455932 272484
rect 456064 272536 456116 272542
rect 456064 272478 456116 272484
rect 455328 268932 455380 268938
rect 455328 268874 455380 268880
rect 454774 266792 454830 266801
rect 454592 266756 454644 266762
rect 454774 266727 454776 266736
rect 454592 266698 454644 266704
rect 454828 266727 454830 266736
rect 454776 266698 454828 266704
rect 454592 266212 454644 266218
rect 454592 266154 454644 266160
rect 454604 264316 454632 266154
rect 455340 264316 455368 268874
rect 456076 264316 456104 272478
rect 456800 271448 456852 271454
rect 456852 271396 457024 271402
rect 456800 271390 457024 271396
rect 456812 271374 457024 271390
rect 456614 271280 456670 271289
rect 456670 271238 456840 271266
rect 456614 271215 456670 271224
rect 456812 271182 456840 271238
rect 456996 271182 457024 271374
rect 456800 271176 456852 271182
rect 456800 271118 456852 271124
rect 456984 271176 457036 271182
rect 456984 271118 457036 271124
rect 456614 270600 456670 270609
rect 456614 270535 456670 270544
rect 456628 270366 456656 270535
rect 456616 270360 456668 270366
rect 456616 270302 456668 270308
rect 456754 270360 456806 270366
rect 456754 270302 456806 270308
rect 456614 270192 456670 270201
rect 456766 270178 456794 270302
rect 456670 270150 456794 270178
rect 456614 270127 456670 270136
rect 456430 268968 456486 268977
rect 456430 268903 456486 268912
rect 456444 268666 456472 268903
rect 456432 268660 456484 268666
rect 456432 268602 456484 268608
rect 456444 268530 457024 268546
rect 456432 268524 457036 268530
rect 456484 268518 456984 268524
rect 456432 268466 456484 268472
rect 456984 268466 457036 268472
rect 456628 268394 456840 268410
rect 456616 268388 456852 268394
rect 456668 268382 456800 268388
rect 456616 268330 456668 268336
rect 456800 268330 456852 268336
rect 456616 268252 456668 268258
rect 456616 268194 456668 268200
rect 456628 268025 456656 268194
rect 456614 268016 456670 268025
rect 456614 267951 456670 267960
rect 457272 267073 457300 273226
rect 457444 272808 457496 272814
rect 457442 272776 457444 272785
rect 457496 272776 457498 272785
rect 457442 272711 457498 272720
rect 458376 272678 458404 277780
rect 459586 277766 459968 277794
rect 458364 272672 458416 272678
rect 458364 272614 458416 272620
rect 458638 271960 458694 271969
rect 458638 271895 458694 271904
rect 457444 271448 457496 271454
rect 457444 271390 457496 271396
rect 457456 271017 457484 271390
rect 457442 271008 457498 271017
rect 457442 270943 457498 270952
rect 457536 268116 457588 268122
rect 457536 268058 457588 268064
rect 457258 267064 457314 267073
rect 457258 266999 457314 267008
rect 457166 266792 457222 266801
rect 457166 266727 457222 266736
rect 457180 264330 457208 266727
rect 456826 264302 457208 264330
rect 457548 264316 457576 268058
rect 458652 264330 458680 271895
rect 459940 270609 459968 277766
rect 460032 277766 460690 277794
rect 461412 277766 461886 277794
rect 462332 277766 463082 277794
rect 464080 277766 464278 277794
rect 465184 277766 465474 277794
rect 466670 277766 467328 277794
rect 460032 273254 460060 277766
rect 460754 273728 460810 273737
rect 460754 273663 460810 273672
rect 460768 273290 460796 273663
rect 460756 273284 460808 273290
rect 460032 273226 460152 273254
rect 460756 273226 460808 273232
rect 459926 270600 459982 270609
rect 459926 270535 459982 270544
rect 459006 270328 459062 270337
rect 459006 270263 459062 270272
rect 458298 264302 458680 264330
rect 459020 264316 459048 270263
rect 460124 268802 460152 273226
rect 460940 273216 460992 273222
rect 460938 273184 460940 273193
rect 460992 273184 460994 273193
rect 460938 273119 460994 273128
rect 460480 272672 460532 272678
rect 460480 272614 460532 272620
rect 460112 268796 460164 268802
rect 460112 268738 460164 268744
rect 460296 268660 460348 268666
rect 460296 268602 460348 268608
rect 460308 267734 460336 268602
rect 460124 267706 460336 267734
rect 460124 264330 460152 267706
rect 459770 264302 460152 264330
rect 460492 264316 460520 272614
rect 461412 271182 461440 277766
rect 461582 275224 461638 275233
rect 461582 275159 461638 275168
rect 461596 273254 461624 275159
rect 461596 273226 461716 273254
rect 461400 271176 461452 271182
rect 461400 271118 461452 271124
rect 461688 269090 461716 273226
rect 461860 271448 461912 271454
rect 461860 271390 461912 271396
rect 461872 271289 461900 271390
rect 461858 271280 461914 271289
rect 461858 271215 461914 271224
rect 461688 269062 461808 269090
rect 461400 268932 461452 268938
rect 461400 268874 461452 268880
rect 461030 268696 461086 268705
rect 461030 268631 461086 268640
rect 461044 268122 461072 268631
rect 461412 268122 461440 268874
rect 461584 268252 461636 268258
rect 461584 268194 461636 268200
rect 461032 268116 461084 268122
rect 461032 268058 461084 268064
rect 461400 268116 461452 268122
rect 461400 268058 461452 268064
rect 461596 268025 461624 268194
rect 461582 268016 461638 268025
rect 461582 267951 461638 267960
rect 461780 267594 461808 269062
rect 462332 268977 462360 277766
rect 464080 273254 464108 277766
rect 463988 273226 464108 273254
rect 462778 271416 462834 271425
rect 462778 271351 462834 271360
rect 462318 268968 462374 268977
rect 462318 268903 462374 268912
rect 462504 268932 462556 268938
rect 462504 268874 462556 268880
rect 462516 268705 462544 268874
rect 462502 268696 462558 268705
rect 461952 268660 462004 268666
rect 462502 268631 462558 268640
rect 461952 268602 462004 268608
rect 461412 267566 461808 267594
rect 461412 267034 461440 267566
rect 461584 267436 461636 267442
rect 461584 267378 461636 267384
rect 461768 267436 461820 267442
rect 461768 267378 461820 267384
rect 461596 267034 461624 267378
rect 461400 267028 461452 267034
rect 461400 266970 461452 266976
rect 461584 267028 461636 267034
rect 461584 266970 461636 266976
rect 461584 266076 461636 266082
rect 461584 266018 461636 266024
rect 461398 265840 461454 265849
rect 461398 265775 461454 265784
rect 461412 265674 461440 265775
rect 461596 265674 461624 266018
rect 461400 265668 461452 265674
rect 461400 265610 461452 265616
rect 461584 265668 461636 265674
rect 461584 265610 461636 265616
rect 461780 264330 461808 267378
rect 461242 264302 461808 264330
rect 461964 264316 461992 268602
rect 462792 266801 462820 271351
rect 462778 266792 462834 266801
rect 462778 266727 462834 266736
rect 463606 266792 463662 266801
rect 463606 266727 463662 266736
rect 462686 266112 462742 266121
rect 462136 266076 462188 266082
rect 462686 266047 462742 266056
rect 462136 266018 462188 266024
rect 462148 265849 462176 266018
rect 462134 265840 462190 265849
rect 462134 265775 462190 265784
rect 462700 264316 462728 266047
rect 463620 264330 463648 266727
rect 463988 266082 464016 273226
rect 464894 272232 464950 272241
rect 464894 272167 464950 272176
rect 463976 266076 464028 266082
rect 463976 266018 464028 266024
rect 464160 266076 464212 266082
rect 464160 266018 464212 266024
rect 463450 264302 463648 264330
rect 464172 264316 464200 266018
rect 464908 264316 464936 272167
rect 465184 271454 465212 277766
rect 466092 277364 466144 277370
rect 466092 277306 466144 277312
rect 465540 275868 465592 275874
rect 465540 275810 465592 275816
rect 465724 275868 465776 275874
rect 465724 275810 465776 275816
rect 465552 275074 465580 275810
rect 465736 275194 465764 275810
rect 465724 275188 465776 275194
rect 465724 275130 465776 275136
rect 465908 275188 465960 275194
rect 465908 275130 465960 275136
rect 465920 275074 465948 275130
rect 465552 275046 465948 275074
rect 465172 271448 465224 271454
rect 465172 271390 465224 271396
rect 465632 271448 465684 271454
rect 465632 271390 465684 271396
rect 465644 264316 465672 271390
rect 466104 267442 466132 277306
rect 466550 275224 466606 275233
rect 466414 275188 466466 275194
rect 466550 275159 466552 275168
rect 466414 275130 466466 275136
rect 466604 275159 466606 275168
rect 466552 275130 466604 275136
rect 466426 275074 466454 275130
rect 466426 275046 466500 275074
rect 466472 274961 466500 275046
rect 466458 274952 466514 274961
rect 466458 274887 466514 274896
rect 466412 274544 466468 274553
rect 466412 274479 466414 274488
rect 466466 274479 466468 274488
rect 466552 274508 466604 274514
rect 466414 274450 466466 274456
rect 466552 274450 466604 274456
rect 466564 273737 466592 274450
rect 466550 273728 466606 273737
rect 466550 273663 466606 273672
rect 466276 272672 466328 272678
rect 466276 272614 466328 272620
rect 466460 272672 466512 272678
rect 466460 272614 466512 272620
rect 466288 272513 466316 272614
rect 466274 272504 466330 272513
rect 466274 272439 466330 272448
rect 466472 272354 466500 272614
rect 466288 272326 466500 272354
rect 466288 271969 466316 272326
rect 466274 271960 466330 271969
rect 466274 271895 466330 271904
rect 466426 271510 466776 271538
rect 466426 271454 466454 271510
rect 466414 271448 466466 271454
rect 466552 271448 466604 271454
rect 466414 271390 466466 271396
rect 466550 271416 466552 271425
rect 466748 271425 466776 271510
rect 466604 271416 466606 271425
rect 466550 271351 466606 271360
rect 466734 271416 466790 271425
rect 466734 271351 466790 271360
rect 466274 269240 466330 269249
rect 466274 269175 466330 269184
rect 466458 269240 466514 269249
rect 466458 269175 466514 269184
rect 466288 269074 466316 269175
rect 466472 269074 466500 269175
rect 466276 269068 466328 269074
rect 466276 269010 466328 269016
rect 466460 269068 466512 269074
rect 466460 269010 466512 269016
rect 466288 268926 466592 268954
rect 466092 267436 466144 267442
rect 466092 267378 466144 267384
rect 466288 267186 466316 268926
rect 466564 268818 466592 268926
rect 466564 268790 467144 268818
rect 466734 268696 466790 268705
rect 467116 268666 467144 268790
rect 466734 268631 466790 268640
rect 467104 268660 467156 268666
rect 466748 268546 466776 268631
rect 467104 268602 467156 268608
rect 466426 268530 466776 268546
rect 466414 268524 466776 268530
rect 466466 268518 466776 268524
rect 466414 268466 466466 268472
rect 466104 267158 466316 267186
rect 466426 267294 466960 267322
rect 466426 267170 466454 267294
rect 466414 267164 466466 267170
rect 466104 264330 466132 267158
rect 466414 267106 466466 267112
rect 466552 267164 466604 267170
rect 466552 267106 466604 267112
rect 466274 267064 466330 267073
rect 466274 266999 466330 267008
rect 466288 266898 466316 266999
rect 466276 266892 466328 266898
rect 466276 266834 466328 266840
rect 466564 266801 466592 267106
rect 466734 267064 466790 267073
rect 466734 266999 466790 267008
rect 466550 266792 466606 266801
rect 466748 266762 466776 266999
rect 466550 266727 466606 266736
rect 466736 266756 466788 266762
rect 466736 266698 466788 266704
rect 466932 266626 466960 267294
rect 466552 266620 466604 266626
rect 466552 266562 466604 266568
rect 466920 266620 466972 266626
rect 466920 266562 466972 266568
rect 466564 266393 466592 266562
rect 466550 266384 466606 266393
rect 466550 266319 466606 266328
rect 467300 264994 467328 277766
rect 467288 264988 467340 264994
rect 467288 264930 467340 264936
rect 467576 264330 467604 278530
rect 467852 276826 467880 277780
rect 468128 277766 468970 277794
rect 469784 277766 470166 277794
rect 470704 277766 471362 277794
rect 472176 277766 472558 277794
rect 467840 276820 467892 276826
rect 467840 276762 467892 276768
rect 468128 269074 468156 277766
rect 469036 276820 469088 276826
rect 469036 276762 469088 276768
rect 468116 269068 468168 269074
rect 468116 269010 468168 269016
rect 467840 267572 467892 267578
rect 467840 267514 467892 267520
rect 466104 264302 466394 264330
rect 467130 264302 467604 264330
rect 467852 264316 467880 267514
rect 469048 264330 469076 276762
rect 469784 274961 469812 277766
rect 469954 276040 470010 276049
rect 469954 275975 470010 275984
rect 469770 274952 469826 274961
rect 469770 274887 469826 274896
rect 469678 269240 469734 269249
rect 469678 269175 469734 269184
rect 469692 264330 469720 269175
rect 469968 266880 469996 275975
rect 470506 275768 470562 275777
rect 470506 275703 470562 275712
rect 470520 275602 470548 275703
rect 470508 275596 470560 275602
rect 470508 275538 470560 275544
rect 469876 266852 469996 266880
rect 469876 266762 469904 266852
rect 469864 266756 469916 266762
rect 469864 266698 469916 266704
rect 470048 266756 470100 266762
rect 470048 266698 470100 266704
rect 468602 264302 469076 264330
rect 469338 264302 469720 264330
rect 470060 264316 470088 266698
rect 470704 266098 470732 277766
rect 471244 277364 471296 277370
rect 471244 277306 471296 277312
rect 471428 277364 471480 277370
rect 471428 277306 471480 277312
rect 471256 276962 471284 277306
rect 471244 276956 471296 276962
rect 471244 276898 471296 276904
rect 471440 276826 471468 277306
rect 471428 276820 471480 276826
rect 471428 276762 471480 276768
rect 471244 276004 471296 276010
rect 471244 275946 471296 275952
rect 471428 276004 471480 276010
rect 471428 275946 471480 275952
rect 470876 275868 470928 275874
rect 470876 275810 470928 275816
rect 471060 275868 471112 275874
rect 471060 275810 471112 275816
rect 470888 275346 470916 275810
rect 471072 275466 471100 275810
rect 471256 275602 471284 275946
rect 471440 275777 471468 275946
rect 471426 275768 471482 275777
rect 471426 275703 471482 275712
rect 471244 275596 471296 275602
rect 471244 275538 471296 275544
rect 471060 275460 471112 275466
rect 471060 275402 471112 275408
rect 471244 275460 471296 275466
rect 471244 275402 471296 275408
rect 471256 275346 471284 275402
rect 470888 275318 471284 275346
rect 472176 274553 472204 277766
rect 472900 276820 472952 276826
rect 472900 276762 472952 276768
rect 472162 274544 472218 274553
rect 471060 274508 471112 274514
rect 471060 274450 471112 274456
rect 471244 274508 471296 274514
rect 472162 274479 472218 274488
rect 471244 274450 471296 274456
rect 471072 274122 471100 274450
rect 471256 274242 471284 274450
rect 471244 274236 471296 274242
rect 471244 274178 471296 274184
rect 471428 274236 471480 274242
rect 471428 274178 471480 274184
rect 471440 274122 471468 274178
rect 471072 274094 471468 274122
rect 472254 270736 472310 270745
rect 472254 270671 472310 270680
rect 471244 269068 471296 269074
rect 471244 269010 471296 269016
rect 471256 268530 471284 269010
rect 471426 268696 471482 268705
rect 471426 268631 471482 268640
rect 471440 268530 471468 268631
rect 471244 268524 471296 268530
rect 471244 268466 471296 268472
rect 471428 268524 471480 268530
rect 471428 268466 471480 268472
rect 470612 266070 470732 266098
rect 470612 265946 470640 266070
rect 470600 265940 470652 265946
rect 470600 265882 470652 265888
rect 470784 265940 470836 265946
rect 470784 265882 470836 265888
rect 470796 264316 470824 265882
rect 471888 264512 471940 264518
rect 471888 264454 471940 264460
rect 471900 264330 471928 264454
rect 471546 264302 471928 264330
rect 472268 264316 472296 270671
rect 472912 264330 472940 276762
rect 473740 276010 473768 277780
rect 474752 277766 474950 277794
rect 473910 276040 473966 276049
rect 473728 276004 473780 276010
rect 473910 275975 473912 275984
rect 473728 275946 473780 275952
rect 473964 275975 473966 275984
rect 473912 275946 473964 275952
rect 473910 275768 473966 275777
rect 473910 275703 473966 275712
rect 473924 266393 473952 275703
rect 474752 268530 474780 277766
rect 475750 277536 475806 277545
rect 476132 277522 476160 277780
rect 476132 277494 476252 277522
rect 475750 277471 475806 277480
rect 475566 277264 475622 277273
rect 475566 277199 475622 277208
rect 475580 277098 475608 277199
rect 475568 277092 475620 277098
rect 475568 277034 475620 277040
rect 475764 276962 475792 277471
rect 475936 277432 475988 277438
rect 475936 277374 475988 277380
rect 475752 276956 475804 276962
rect 475752 276898 475804 276904
rect 475948 276826 475976 277374
rect 475752 276820 475804 276826
rect 475752 276762 475804 276768
rect 475936 276820 475988 276826
rect 475936 276762 475988 276768
rect 475764 276457 475792 276762
rect 475750 276448 475806 276457
rect 475750 276383 475806 276392
rect 475382 274544 475438 274553
rect 475382 274479 475438 274488
rect 474740 268524 474792 268530
rect 474740 268466 474792 268472
rect 475200 268524 475252 268530
rect 475200 268466 475252 268472
rect 474094 268152 474150 268161
rect 474094 268087 474150 268096
rect 473910 266384 473966 266393
rect 473910 266319 473966 266328
rect 474108 264330 474136 268087
rect 474646 267064 474702 267073
rect 474646 266999 474702 267008
rect 474660 264330 474688 266999
rect 472912 264302 473018 264330
rect 473754 264302 474136 264330
rect 474490 264302 474688 264330
rect 475212 264316 475240 268466
rect 475396 264466 475424 274479
rect 476224 274378 476252 277494
rect 476500 277438 476528 278530
rect 476670 277536 476726 277545
rect 476670 277471 476726 277480
rect 476488 277432 476540 277438
rect 476488 277374 476540 277380
rect 476394 277264 476450 277273
rect 476394 277199 476450 277208
rect 476408 277098 476436 277199
rect 476396 277092 476448 277098
rect 476396 277034 476448 277040
rect 476684 276962 476712 277471
rect 476672 276956 476724 276962
rect 476672 276898 476724 276904
rect 477236 276010 477264 277780
rect 477880 277766 478446 277794
rect 477224 276004 477276 276010
rect 477224 275946 477276 275952
rect 477408 276004 477460 276010
rect 477408 275946 477460 275952
rect 476212 274372 476264 274378
rect 476212 274314 476264 274320
rect 477420 273254 477448 275946
rect 476960 273226 477448 273254
rect 476762 272776 476818 272785
rect 476762 272711 476818 272720
rect 476776 272241 476804 272711
rect 476762 272232 476818 272241
rect 476762 272167 476818 272176
rect 475764 270422 476252 270450
rect 475764 270230 475792 270422
rect 475936 270360 475988 270366
rect 475936 270302 475988 270308
rect 475752 270224 475804 270230
rect 475752 270166 475804 270172
rect 475948 270094 475976 270302
rect 476224 270230 476252 270422
rect 476488 270360 476540 270366
rect 476488 270302 476540 270308
rect 476212 270224 476264 270230
rect 476212 270166 476264 270172
rect 475752 270088 475804 270094
rect 475750 270056 475752 270065
rect 475936 270088 475988 270094
rect 475804 270056 475806 270065
rect 475936 270030 475988 270036
rect 475750 269991 475806 270000
rect 476500 269249 476528 270302
rect 476486 269240 476542 269249
rect 476486 269175 476542 269184
rect 476670 269240 476726 269249
rect 476670 269175 476726 269184
rect 476210 268152 476266 268161
rect 476210 268087 476266 268096
rect 475750 267880 475806 267889
rect 476224 267850 476252 268087
rect 475750 267815 475752 267824
rect 475804 267815 475806 267824
rect 476212 267844 476264 267850
rect 475752 267786 475804 267792
rect 476212 267786 476264 267792
rect 475750 267608 475806 267617
rect 475750 267543 475752 267552
rect 475804 267543 475806 267552
rect 476118 267608 476174 267617
rect 476118 267543 476120 267552
rect 475752 267514 475804 267520
rect 476172 267543 476174 267552
rect 476302 267608 476358 267617
rect 476302 267543 476358 267552
rect 476120 267514 476172 267520
rect 476316 267186 476344 267543
rect 475764 267170 476344 267186
rect 475752 267164 476344 267170
rect 475804 267158 476344 267164
rect 475752 267106 475804 267112
rect 476210 267064 476266 267073
rect 476210 266999 476266 267008
rect 476396 267028 476448 267034
rect 476224 266626 476252 266999
rect 476396 266970 476448 266976
rect 476028 266620 476080 266626
rect 476028 266562 476080 266568
rect 476212 266620 476264 266626
rect 476212 266562 476264 266568
rect 476040 266506 476068 266562
rect 476408 266506 476436 266970
rect 476040 266478 476436 266506
rect 475396 264438 475608 264466
rect 475580 264330 475608 264438
rect 475580 264302 475962 264330
rect 476684 264316 476712 269175
rect 476960 267034 476988 273226
rect 477880 270065 477908 277766
rect 479628 274514 479656 277780
rect 480824 275874 480852 277780
rect 481652 277766 482034 277794
rect 480994 275904 481050 275913
rect 480812 275868 480864 275874
rect 480994 275839 480996 275848
rect 480812 275810 480864 275816
rect 481048 275839 481050 275848
rect 480996 275810 481048 275816
rect 481270 275224 481326 275233
rect 481270 275159 481326 275168
rect 480350 274544 480406 274553
rect 479616 274508 479668 274514
rect 480350 274479 480352 274488
rect 479616 274450 479668 274456
rect 480404 274479 480406 274488
rect 480352 274450 480404 274456
rect 478604 274372 478656 274378
rect 478604 274314 478656 274320
rect 477866 270056 477922 270065
rect 477866 269991 477922 270000
rect 477132 267300 477184 267306
rect 477132 267242 477184 267248
rect 477144 267034 477172 267242
rect 476948 267028 477000 267034
rect 476948 266970 477000 266976
rect 477132 267028 477184 267034
rect 477132 266970 477184 266976
rect 477408 264988 477460 264994
rect 477408 264930 477460 264936
rect 477420 264316 477448 264930
rect 478616 264330 478644 274314
rect 479982 270056 480038 270065
rect 479982 269991 480038 270000
rect 479246 265296 479302 265305
rect 479246 265231 479302 265240
rect 479260 264330 479288 265231
rect 479996 264330 480024 269991
rect 480904 268252 480956 268258
rect 480904 268194 480956 268200
rect 481088 268252 481140 268258
rect 481088 268194 481140 268200
rect 480916 267850 480944 268194
rect 480720 267844 480772 267850
rect 480720 267786 480772 267792
rect 480904 267844 480956 267850
rect 480904 267786 480956 267792
rect 480732 267730 480760 267786
rect 481100 267734 481128 268194
rect 481008 267730 481128 267734
rect 480732 267706 481128 267730
rect 480732 267702 481036 267706
rect 480352 267436 480404 267442
rect 480352 267378 480404 267384
rect 478170 264302 478644 264330
rect 478906 264302 479288 264330
rect 479642 264302 480024 264330
rect 480364 264316 480392 267378
rect 481284 264330 481312 275159
rect 481454 274408 481510 274417
rect 481454 274343 481510 274352
rect 481468 267442 481496 274343
rect 481652 269958 481680 277766
rect 481640 269952 481692 269958
rect 481640 269894 481692 269900
rect 482296 267617 482324 278530
rect 644662 278080 644718 278089
rect 644662 278015 644718 278024
rect 546684 277840 546736 277846
rect 483216 274106 483244 277780
rect 484122 275904 484178 275913
rect 484320 275874 484348 277780
rect 484688 277766 485530 277794
rect 484122 275839 484178 275848
rect 484308 275868 484360 275874
rect 483204 274100 483256 274106
rect 483204 274042 483256 274048
rect 484136 269249 484164 275839
rect 484308 275810 484360 275816
rect 484492 275868 484544 275874
rect 484492 275810 484544 275816
rect 484504 275330 484532 275810
rect 484492 275324 484544 275330
rect 484492 275266 484544 275272
rect 484306 274952 484362 274961
rect 484306 274887 484362 274896
rect 484320 273834 484348 274887
rect 484308 273828 484360 273834
rect 484308 273770 484360 273776
rect 484308 269952 484360 269958
rect 484308 269894 484360 269900
rect 484122 269240 484178 269249
rect 484122 269175 484178 269184
rect 482282 267608 482338 267617
rect 482282 267543 482338 267552
rect 481456 267436 481508 267442
rect 481456 267378 481508 267384
rect 481640 267436 481692 267442
rect 481640 267378 481692 267384
rect 481652 266626 481680 267378
rect 481640 266620 481692 266626
rect 481640 266562 481692 266568
rect 482560 266620 482612 266626
rect 482560 266562 482612 266568
rect 481822 265840 481878 265849
rect 481822 265775 481878 265784
rect 481114 264302 481312 264330
rect 481836 264316 481864 265775
rect 482572 264316 482600 266562
rect 483294 266520 483350 266529
rect 483294 266455 483350 266464
rect 483308 264316 483336 266455
rect 484320 264330 484348 269894
rect 484688 269822 484716 277766
rect 485870 276448 485926 276457
rect 485870 276383 485926 276392
rect 485884 276146 485912 276383
rect 485734 276140 485786 276146
rect 485734 276082 485786 276088
rect 485872 276140 485924 276146
rect 485872 276082 485924 276088
rect 485746 276026 485774 276082
rect 486054 276040 486110 276049
rect 485228 276004 485280 276010
rect 485746 275998 486054 276026
rect 486054 275975 486110 275984
rect 485228 275946 485280 275952
rect 485240 275602 485268 275946
rect 485870 275904 485926 275913
rect 485870 275839 485872 275848
rect 485924 275839 485926 275848
rect 485872 275810 485924 275816
rect 485228 275596 485280 275602
rect 485228 275538 485280 275544
rect 484860 275460 484912 275466
rect 484860 275402 484912 275408
rect 484872 275210 484900 275402
rect 484872 275194 485268 275210
rect 484872 275188 485280 275194
rect 484872 275182 485228 275188
rect 485228 275130 485280 275136
rect 486712 274961 486740 277780
rect 487908 276010 487936 277780
rect 488552 277766 489118 277794
rect 489932 277766 490314 277794
rect 487896 276004 487948 276010
rect 487896 275946 487948 275952
rect 487342 275768 487398 275777
rect 487342 275703 487398 275712
rect 487356 275330 487384 275703
rect 487344 275324 487396 275330
rect 487344 275266 487396 275272
rect 487528 275324 487580 275330
rect 487528 275266 487580 275272
rect 486698 274952 486754 274961
rect 486698 274887 486754 274896
rect 486698 274680 486754 274689
rect 486698 274615 486754 274624
rect 486422 274408 486478 274417
rect 486422 274343 486478 274352
rect 486436 274242 486464 274343
rect 484860 274236 484912 274242
rect 484860 274178 484912 274184
rect 485228 274236 485280 274242
rect 485228 274178 485280 274184
rect 486424 274236 486476 274242
rect 486424 274178 486476 274184
rect 484872 273834 484900 274178
rect 484860 273828 484912 273834
rect 484860 273770 484912 273776
rect 484858 270056 484914 270065
rect 484914 270014 485084 270042
rect 484858 269991 484914 270000
rect 485056 269958 485084 270014
rect 485044 269952 485096 269958
rect 485044 269894 485096 269900
rect 484676 269816 484728 269822
rect 484676 269758 484728 269764
rect 484674 268968 484730 268977
rect 484674 268903 484730 268912
rect 484688 268122 484716 268903
rect 484858 268696 484914 268705
rect 484858 268631 484914 268640
rect 484872 268258 484900 268631
rect 484860 268252 484912 268258
rect 484860 268194 484912 268200
rect 485042 268152 485098 268161
rect 484676 268116 484728 268122
rect 485042 268087 485098 268096
rect 484676 268058 484728 268064
rect 485056 267850 485084 268087
rect 485044 267844 485096 267850
rect 485044 267786 485096 267792
rect 485240 264330 485268 274178
rect 486712 273254 486740 274615
rect 486882 274408 486938 274417
rect 486882 274343 486938 274352
rect 486896 273698 486924 274343
rect 487066 273864 487122 273873
rect 487066 273799 487122 273808
rect 486884 273692 486936 273698
rect 486884 273634 486936 273640
rect 486712 273226 486924 273254
rect 485746 272326 486096 272354
rect 485746 272270 485774 272326
rect 485734 272264 485786 272270
rect 485872 272264 485924 272270
rect 485734 272206 485786 272212
rect 485870 272232 485872 272241
rect 486068 272241 486096 272326
rect 485924 272232 485926 272241
rect 485870 272167 485926 272176
rect 486054 272232 486110 272241
rect 486054 272167 486110 272176
rect 485778 271960 485834 271969
rect 485778 271895 485834 271904
rect 485792 271538 485820 271895
rect 485746 271510 485820 271538
rect 485746 271182 485774 271510
rect 485870 271416 485926 271425
rect 485870 271351 485926 271360
rect 485884 271182 485912 271351
rect 485734 271176 485786 271182
rect 485734 271118 485786 271124
rect 485872 271176 485924 271182
rect 485872 271118 485924 271124
rect 485502 271008 485558 271017
rect 485502 270943 485558 270952
rect 485516 268818 485544 270943
rect 486896 270745 486924 273226
rect 486882 270736 486938 270745
rect 486882 270671 486938 270680
rect 486606 269240 486662 269249
rect 486606 269175 486662 269184
rect 486422 268968 486478 268977
rect 486422 268903 486478 268912
rect 485424 268790 485544 268818
rect 485424 266642 485452 268790
rect 486238 268696 486294 268705
rect 486238 268631 486294 268640
rect 485688 268252 485740 268258
rect 485688 268194 485740 268200
rect 485872 268252 485924 268258
rect 485872 268194 485924 268200
rect 486056 268252 486108 268258
rect 486056 268194 486108 268200
rect 485700 267889 485728 268194
rect 485686 267880 485742 267889
rect 485686 267815 485742 267824
rect 485884 267753 485912 268194
rect 486068 268025 486096 268194
rect 486054 268016 486110 268025
rect 486054 267951 486110 267960
rect 486252 267850 486280 268631
rect 486436 268122 486464 268903
rect 486424 268116 486476 268122
rect 486424 268058 486476 268064
rect 486240 267844 486292 267850
rect 486240 267786 486292 267792
rect 485870 267744 485926 267753
rect 485870 267679 485926 267688
rect 485594 267064 485650 267073
rect 485594 266999 485650 267008
rect 484058 264302 484348 264330
rect 484794 264302 485268 264330
rect 485332 266614 485452 266642
rect 485608 266626 485636 266999
rect 485596 266620 485648 266626
rect 485332 264330 485360 266614
rect 485596 266562 485648 266568
rect 485780 266620 485832 266626
rect 485780 266562 485832 266568
rect 485792 266506 485820 266562
rect 485608 266478 485820 266506
rect 485608 265305 485636 266478
rect 485594 265296 485650 265305
rect 485594 265231 485650 265240
rect 486620 264330 486648 269175
rect 487080 268682 487108 273799
rect 485332 264302 485530 264330
rect 486266 264302 486648 264330
rect 486988 268654 487108 268682
rect 486988 264316 487016 268654
rect 487540 267034 487568 275266
rect 488354 270056 488410 270065
rect 488354 269991 488410 270000
rect 487528 267028 487580 267034
rect 487528 266970 487580 266976
rect 487712 267028 487764 267034
rect 487712 266970 487764 266976
rect 487724 264316 487752 266970
rect 488368 264330 488396 269991
rect 488552 269793 488580 277766
rect 489932 274802 489960 277766
rect 490564 276004 490616 276010
rect 490564 275946 490616 275952
rect 490576 275602 490604 275946
rect 490746 275768 490802 275777
rect 490746 275703 490802 275712
rect 490760 275602 490788 275703
rect 490564 275596 490616 275602
rect 490564 275538 490616 275544
rect 490748 275596 490800 275602
rect 490748 275538 490800 275544
rect 491496 275330 491524 277780
rect 492232 277766 492614 277794
rect 492968 277766 493810 277794
rect 492232 276049 492260 277766
rect 492218 276040 492274 276049
rect 492218 275975 492274 275984
rect 492586 275904 492642 275913
rect 492586 275839 492642 275848
rect 491484 275324 491536 275330
rect 491484 275266 491536 275272
rect 491668 275324 491720 275330
rect 491668 275266 491720 275272
rect 489840 274774 489960 274802
rect 491680 274786 491708 275266
rect 491668 274780 491720 274786
rect 489840 274650 489868 274774
rect 491668 274722 491720 274728
rect 491852 274780 491904 274786
rect 491852 274722 491904 274728
rect 489828 274644 489880 274650
rect 489828 274586 489880 274592
rect 490012 274644 490064 274650
rect 490012 274586 490064 274592
rect 488722 273864 488778 273873
rect 488722 273799 488724 273808
rect 488776 273799 488778 273808
rect 489366 273864 489422 273873
rect 489366 273799 489422 273808
rect 488724 273770 488776 273776
rect 488538 269784 488594 269793
rect 488538 269719 488594 269728
rect 489380 264330 489408 273799
rect 490024 267073 490052 274586
rect 491864 273254 491892 274722
rect 491404 273226 491892 273254
rect 491022 272776 491078 272785
rect 491022 272711 491078 272720
rect 490288 270224 490340 270230
rect 490288 270166 490340 270172
rect 490300 270042 490328 270166
rect 490300 270014 490880 270042
rect 490852 269958 490880 270014
rect 490196 269952 490248 269958
rect 490196 269894 490248 269900
rect 490840 269952 490892 269958
rect 490840 269894 490892 269900
rect 490208 269804 490236 269894
rect 490840 269816 490892 269822
rect 490208 269776 490840 269804
rect 490840 269758 490892 269764
rect 490194 268696 490250 268705
rect 490194 268631 490250 268640
rect 490208 267714 490236 268631
rect 491036 268138 491064 272711
rect 491404 269822 491432 273226
rect 491392 269816 491444 269822
rect 491392 269758 491444 269764
rect 491576 269816 491628 269822
rect 491576 269758 491628 269764
rect 491588 269249 491616 269758
rect 491574 269240 491630 269249
rect 491574 269175 491630 269184
rect 490392 268110 491064 268138
rect 490196 267708 490248 267714
rect 490196 267650 490248 267656
rect 490010 267064 490066 267073
rect 489828 267028 489880 267034
rect 490010 266999 490066 267008
rect 489828 266970 489880 266976
rect 489840 266914 489868 266970
rect 490194 266928 490250 266937
rect 489840 266886 490194 266914
rect 490194 266863 490250 266872
rect 490392 264330 490420 268110
rect 491574 268016 491630 268025
rect 491574 267951 491630 267960
rect 491392 267708 491444 267714
rect 491392 267650 491444 267656
rect 490576 267442 490880 267458
rect 490564 267436 490892 267442
rect 490616 267430 490840 267436
rect 490564 267378 490616 267384
rect 490840 267378 490892 267384
rect 490576 267306 490880 267322
rect 490564 267300 490892 267306
rect 490616 267294 490840 267300
rect 490564 267242 490616 267248
rect 490840 267242 490892 267248
rect 490576 267170 490880 267186
rect 490576 267164 490892 267170
rect 490576 267158 490840 267164
rect 490576 267102 490604 267158
rect 490840 267106 490892 267112
rect 490564 267096 490616 267102
rect 490564 267038 490616 267044
rect 491206 266928 491262 266937
rect 491206 266863 491208 266872
rect 491260 266863 491262 266872
rect 491208 266834 491260 266840
rect 491024 264376 491076 264382
rect 488368 264302 488474 264330
rect 489210 264302 489408 264330
rect 489946 264302 490420 264330
rect 490682 264324 491024 264330
rect 490682 264318 491076 264324
rect 490682 264302 491064 264318
rect 491404 264316 491432 267650
rect 491588 264382 491616 267951
rect 492600 267714 492628 275839
rect 492968 271969 492996 277766
rect 493138 276448 493194 276457
rect 493138 276383 493194 276392
rect 492954 271960 493010 271969
rect 492954 271895 493010 271904
rect 493152 269362 493180 276383
rect 494992 275602 495020 277780
rect 494980 275596 495032 275602
rect 494980 275538 495032 275544
rect 495164 275596 495216 275602
rect 495164 275538 495216 275544
rect 494150 274952 494206 274961
rect 494150 274887 494206 274896
rect 494164 274786 494192 274887
rect 495176 274802 495204 275538
rect 494152 274780 494204 274786
rect 494152 274722 494204 274728
rect 494336 274780 494388 274786
rect 494336 274722 494388 274728
rect 494992 274774 495204 274802
rect 493966 270872 494022 270881
rect 493966 270807 494022 270816
rect 493060 269334 493180 269362
rect 493060 268705 493088 269334
rect 493230 269240 493286 269249
rect 493230 269175 493286 269184
rect 493046 268696 493102 268705
rect 493046 268631 493102 268640
rect 492770 267744 492826 267753
rect 492588 267708 492640 267714
rect 492770 267679 492772 267688
rect 492588 267650 492640 267656
rect 492824 267679 492826 267688
rect 492772 267650 492824 267656
rect 492126 266792 492182 266801
rect 492126 266727 492182 266736
rect 491576 264376 491628 264382
rect 491576 264318 491628 264324
rect 492140 264316 492168 266727
rect 493244 264330 493272 269175
rect 493980 264330 494008 270807
rect 492890 264302 493272 264330
rect 493626 264302 494008 264330
rect 494348 264316 494376 274722
rect 494992 274689 495020 274774
rect 494978 274680 495034 274689
rect 494978 274615 495034 274624
rect 495254 274680 495310 274689
rect 495254 274615 495256 274624
rect 495308 274615 495310 274624
rect 495394 274644 495446 274650
rect 495256 274586 495308 274592
rect 495394 274586 495446 274592
rect 495406 274530 495434 274586
rect 495268 274502 495434 274530
rect 495268 274417 495296 274502
rect 495254 274408 495310 274417
rect 495254 274343 495310 274352
rect 494886 273320 494942 273329
rect 494886 273255 494942 273264
rect 494900 270494 494928 273255
rect 495898 273048 495954 273057
rect 495898 272983 495954 272992
rect 495912 272241 495940 272983
rect 495898 272232 495954 272241
rect 495898 272167 495954 272176
rect 496188 271538 496216 277780
rect 497016 277766 497398 277794
rect 497016 274650 497044 277766
rect 498580 276010 498608 277780
rect 499394 277264 499450 277273
rect 499394 277199 499450 277208
rect 499408 276146 499436 277199
rect 499396 276140 499448 276146
rect 499396 276082 499448 276088
rect 499534 276140 499586 276146
rect 499534 276082 499586 276088
rect 499546 276026 499574 276082
rect 498568 276004 498620 276010
rect 498568 275946 498620 275952
rect 498752 276004 498804 276010
rect 498752 275946 498804 275952
rect 499408 275998 499574 276026
rect 498764 275330 498792 275946
rect 499408 275913 499436 275998
rect 499394 275904 499450 275913
rect 499394 275839 499450 275848
rect 499408 275466 500172 275482
rect 499396 275460 500172 275466
rect 499448 275454 500172 275460
rect 499396 275402 499448 275408
rect 498752 275324 498804 275330
rect 498752 275266 498804 275272
rect 498936 275324 498988 275330
rect 498936 275266 498988 275272
rect 499672 275324 499724 275330
rect 499672 275266 499724 275272
rect 498948 274961 498976 275266
rect 499684 274961 499712 275266
rect 498934 274952 498990 274961
rect 498934 274887 498990 274896
rect 499394 274952 499450 274961
rect 499394 274887 499450 274896
rect 499670 274952 499726 274961
rect 499670 274887 499726 274896
rect 499408 274786 499436 274887
rect 500144 274786 500172 275454
rect 499396 274780 499448 274786
rect 499396 274722 499448 274728
rect 500132 274780 500184 274786
rect 500132 274722 500184 274728
rect 497186 274680 497242 274689
rect 497004 274644 497056 274650
rect 497186 274615 497188 274624
rect 497004 274586 497056 274592
rect 497240 274615 497242 274624
rect 497188 274586 497240 274592
rect 497462 273592 497518 273601
rect 497462 273527 497518 273536
rect 496004 271510 496216 271538
rect 495452 271374 495848 271402
rect 495452 271182 495480 271374
rect 495440 271176 495492 271182
rect 495440 271118 495492 271124
rect 495624 271176 495676 271182
rect 495820 271153 495848 271374
rect 495624 271118 495676 271124
rect 495806 271144 495862 271153
rect 495636 271046 495664 271118
rect 495806 271079 495862 271088
rect 495624 271040 495676 271046
rect 495624 270982 495676 270988
rect 495072 270904 495124 270910
rect 495808 270904 495860 270910
rect 495124 270852 495808 270858
rect 495072 270846 495860 270852
rect 495084 270830 495848 270846
rect 495072 270768 495124 270774
rect 496004 270722 496032 271510
rect 496544 271176 496596 271182
rect 496358 271144 496414 271153
rect 496544 271118 496596 271124
rect 496726 271144 496782 271153
rect 496358 271079 496414 271088
rect 495124 270716 495664 270722
rect 495072 270710 495664 270716
rect 495084 270694 495664 270710
rect 496004 270694 496124 270722
rect 495440 270632 495492 270638
rect 495438 270600 495440 270609
rect 495636 270620 495664 270694
rect 495900 270632 495952 270638
rect 495492 270600 495494 270609
rect 495636 270592 495900 270620
rect 495900 270574 495952 270580
rect 495438 270535 495494 270544
rect 496096 270494 496124 270694
rect 496372 270638 496400 271079
rect 496556 270881 496584 271118
rect 496726 271079 496782 271088
rect 496542 270872 496598 270881
rect 496542 270807 496598 270816
rect 496360 270632 496412 270638
rect 496360 270574 496412 270580
rect 496740 270494 496768 271079
rect 494900 270466 495296 270494
rect 495268 269958 495296 270466
rect 495912 270466 496124 270494
rect 496188 270466 496768 270494
rect 495256 269952 495308 269958
rect 495256 269894 495308 269900
rect 495532 269816 495584 269822
rect 494702 269784 494758 269793
rect 495532 269758 495584 269764
rect 494702 269719 494758 269728
rect 494518 268152 494574 268161
rect 494518 268087 494574 268096
rect 494532 267850 494560 268087
rect 494520 267844 494572 267850
rect 494520 267786 494572 267792
rect 494716 264330 494744 269719
rect 495544 269249 495572 269758
rect 495530 269240 495586 269249
rect 495530 269175 495586 269184
rect 495070 268696 495126 268705
rect 495070 268631 495126 268640
rect 495530 268696 495586 268705
rect 495530 268631 495586 268640
rect 495084 268394 495112 268631
rect 495544 268394 495572 268631
rect 495072 268388 495124 268394
rect 495072 268330 495124 268336
rect 495532 268388 495584 268394
rect 495532 268330 495584 268336
rect 494888 267708 494940 267714
rect 494888 267650 494940 267656
rect 494900 267306 494928 267650
rect 494888 267300 494940 267306
rect 494888 267242 494940 267248
rect 495912 265674 495940 270466
rect 495900 265668 495952 265674
rect 495900 265610 495952 265616
rect 496188 264330 496216 270466
rect 496544 267300 496596 267306
rect 496544 267242 496596 267248
rect 494716 264302 495098 264330
rect 495834 264302 496216 264330
rect 496556 264316 496584 267242
rect 497476 267170 497504 273527
rect 500880 273329 500908 277780
rect 501800 277766 502090 277794
rect 502352 277766 503286 277794
rect 504192 277766 504482 277794
rect 505296 277766 505678 277794
rect 506492 277766 506874 277794
rect 501800 276010 501828 277766
rect 502352 277098 502380 277766
rect 502522 277264 502578 277273
rect 502522 277199 502578 277208
rect 502536 277098 502564 277199
rect 502340 277092 502392 277098
rect 502340 277034 502392 277040
rect 502524 277092 502576 277098
rect 502524 277034 502576 277040
rect 501788 276004 501840 276010
rect 501788 275946 501840 275952
rect 501972 276004 502024 276010
rect 501972 275946 502024 275952
rect 500866 273320 500922 273329
rect 500866 273255 500922 273264
rect 500052 270286 500448 270314
rect 500052 269550 500080 270286
rect 500420 270230 500448 270286
rect 501984 270230 502012 275946
rect 504192 270609 504220 277766
rect 505296 273601 505324 277766
rect 505282 273592 505338 273601
rect 505282 273527 505338 273536
rect 504178 270600 504234 270609
rect 504178 270535 504234 270544
rect 500224 270224 500276 270230
rect 500224 270166 500276 270172
rect 500408 270224 500460 270230
rect 500408 270166 500460 270172
rect 501972 270224 502024 270230
rect 501972 270166 502024 270172
rect 502156 270224 502208 270230
rect 502156 270166 502208 270172
rect 500236 269550 500264 270166
rect 500040 269544 500092 269550
rect 500040 269486 500092 269492
rect 500224 269544 500276 269550
rect 500224 269486 500276 269492
rect 502168 267889 502196 270166
rect 506492 268705 506520 277766
rect 507964 277394 507992 277780
rect 507872 277366 507992 277394
rect 508700 277766 509174 277794
rect 507872 273057 507900 277366
rect 508700 275738 508728 277766
rect 510356 277574 510384 277780
rect 510344 277568 510396 277574
rect 510344 277510 510396 277516
rect 509422 277264 509478 277273
rect 508884 277222 509280 277250
rect 508884 276457 508912 277222
rect 509252 277098 509280 277222
rect 509422 277199 509478 277208
rect 509056 277092 509108 277098
rect 509056 277034 509108 277040
rect 509240 277092 509292 277098
rect 509240 277034 509292 277040
rect 509068 276842 509096 277034
rect 509436 276842 509464 277199
rect 509068 276814 509464 276842
rect 509056 276684 509108 276690
rect 509056 276626 509108 276632
rect 509240 276684 509292 276690
rect 509240 276626 509292 276632
rect 509068 276457 509096 276626
rect 509252 276457 509280 276626
rect 508870 276448 508926 276457
rect 508870 276383 508926 276392
rect 509054 276448 509110 276457
rect 509054 276383 509110 276392
rect 509238 276448 509294 276457
rect 509238 276383 509294 276392
rect 511552 276010 511580 277780
rect 512012 277766 512762 277794
rect 513392 277766 513958 277794
rect 512012 277098 512040 277766
rect 512182 277264 512238 277273
rect 512182 277199 512238 277208
rect 512196 277098 512224 277199
rect 512000 277092 512052 277098
rect 512000 277034 512052 277040
rect 512184 277092 512236 277098
rect 512184 277034 512236 277040
rect 511540 276004 511592 276010
rect 511540 275946 511592 275952
rect 508688 275732 508740 275738
rect 508688 275674 508740 275680
rect 511356 275732 511408 275738
rect 511356 275674 511408 275680
rect 507858 273048 507914 273057
rect 507858 272983 507914 272992
rect 511368 272785 511396 275674
rect 511354 272776 511410 272785
rect 511354 272711 511410 272720
rect 513392 269278 513420 277766
rect 515140 273426 515168 277780
rect 516244 274922 516272 277780
rect 516428 277766 517454 277794
rect 516232 274916 516284 274922
rect 516232 274858 516284 274864
rect 515128 273420 515180 273426
rect 515128 273362 515180 273368
rect 513852 270966 514248 270994
rect 513852 270910 513880 270966
rect 513840 270904 513892 270910
rect 513840 270846 513892 270852
rect 514024 270904 514076 270910
rect 514024 270846 514076 270852
rect 514036 270638 514064 270846
rect 514220 270638 514248 270966
rect 514024 270632 514076 270638
rect 514024 270574 514076 270580
rect 514208 270632 514260 270638
rect 514208 270574 514260 270580
rect 513380 269272 513432 269278
rect 513380 269214 513432 269220
rect 504914 268696 504970 268705
rect 504914 268631 504970 268640
rect 506478 268696 506534 268705
rect 506478 268631 506534 268640
rect 504928 268394 504956 268631
rect 504916 268388 504968 268394
rect 504916 268330 504968 268336
rect 505054 268388 505106 268394
rect 505054 268330 505106 268336
rect 505066 268274 505094 268330
rect 504928 268246 505094 268274
rect 504928 268161 504956 268246
rect 504914 268152 504970 268161
rect 504914 268087 504970 268096
rect 502154 267880 502210 267889
rect 502154 267815 502210 267824
rect 499946 267608 500002 267617
rect 499946 267543 500002 267552
rect 497464 267164 497516 267170
rect 497464 267106 497516 267112
rect 498752 267164 498804 267170
rect 498752 267106 498804 267112
rect 498014 267064 498070 267073
rect 498014 266999 498070 267008
rect 497648 264376 497700 264382
rect 497306 264324 497648 264330
rect 497306 264318 497700 264324
rect 497306 264302 497688 264318
rect 498028 264316 498056 266999
rect 498764 264316 498792 267106
rect 499960 266801 499988 267543
rect 504928 267430 505232 267458
rect 504928 267306 504956 267430
rect 504916 267300 504968 267306
rect 504916 267242 504968 267248
rect 505054 267300 505106 267306
rect 505054 267242 505106 267248
rect 505066 267186 505094 267242
rect 504836 267158 505094 267186
rect 504836 267073 504864 267158
rect 504822 267064 504878 267073
rect 504548 267028 504600 267034
rect 505204 267034 505232 267430
rect 504822 266999 504878 267008
rect 505192 267028 505244 267034
rect 504548 266970 504600 266976
rect 505192 266970 505244 266976
rect 504560 266914 504588 266970
rect 504560 266886 504956 266914
rect 499946 266792 500002 266801
rect 504928 266762 504956 266886
rect 499946 266727 500002 266736
rect 504732 266756 504784 266762
rect 504732 266698 504784 266704
rect 504916 266756 504968 266762
rect 504916 266698 504968 266704
rect 504744 266529 504772 266698
rect 504730 266520 504786 266529
rect 504730 266455 504786 266464
rect 507122 266520 507178 266529
rect 507122 266455 507178 266464
rect 499488 265668 499540 265674
rect 499488 265610 499540 265616
rect 499500 264316 499528 265610
rect 364090 264166 364288 264194
rect 507136 264110 507164 266455
rect 516428 265266 516456 277766
rect 518636 270638 518664 277780
rect 518912 277766 519846 277794
rect 518624 270632 518676 270638
rect 518624 270574 518676 270580
rect 518912 267345 518940 277766
rect 521028 276418 521056 277780
rect 521672 277766 522238 277794
rect 521016 276412 521068 276418
rect 521016 276354 521068 276360
rect 521672 269414 521700 277766
rect 523420 275058 523448 277780
rect 524340 277766 524538 277794
rect 524708 277766 525734 277794
rect 525996 277766 526930 277794
rect 527192 277766 528126 277794
rect 524340 277710 524368 277766
rect 524328 277704 524380 277710
rect 524328 277646 524380 277652
rect 523868 275188 523920 275194
rect 523868 275130 523920 275136
rect 523408 275052 523460 275058
rect 523408 274994 523460 275000
rect 523880 274922 523908 275130
rect 523868 274916 523920 274922
rect 523868 274858 523920 274864
rect 523684 274780 523736 274786
rect 523684 274722 523736 274728
rect 521660 269408 521712 269414
rect 521660 269350 521712 269356
rect 518898 267336 518954 267345
rect 518898 267271 518954 267280
rect 523696 265810 523724 274722
rect 524708 267850 524736 277766
rect 524696 267844 524748 267850
rect 524696 267786 524748 267792
rect 525996 267714 526024 277766
rect 527192 269686 527220 277766
rect 529308 273562 529336 277780
rect 530504 275058 530532 277780
rect 531228 276276 531280 276282
rect 531228 276218 531280 276224
rect 530492 275052 530544 275058
rect 530492 274994 530544 275000
rect 531240 274922 531268 276218
rect 531228 274916 531280 274922
rect 531228 274858 531280 274864
rect 529296 273556 529348 273562
rect 529296 273498 529348 273504
rect 531608 270774 531636 277780
rect 532804 271998 532832 277780
rect 532988 277766 534014 277794
rect 532792 271992 532844 271998
rect 532792 271934 532844 271940
rect 531596 270768 531648 270774
rect 531596 270710 531648 270716
rect 527180 269680 527232 269686
rect 527180 269622 527232 269628
rect 525984 267708 526036 267714
rect 525984 267650 526036 267656
rect 532988 266490 533016 277766
rect 535196 271726 535224 277780
rect 535472 277766 536406 277794
rect 535184 271720 535236 271726
rect 535184 271662 535236 271668
rect 535472 269521 535500 277766
rect 537588 275194 537616 277780
rect 538416 277766 538798 277794
rect 537576 275188 537628 275194
rect 537576 275130 537628 275136
rect 537760 275188 537812 275194
rect 537760 275130 537812 275136
rect 535458 269512 535514 269521
rect 535458 269447 535514 269456
rect 532976 266484 533028 266490
rect 532976 266426 533028 266432
rect 523684 265804 523736 265810
rect 523684 265746 523736 265752
rect 516416 265260 516468 265266
rect 516416 265202 516468 265208
rect 537772 265130 537800 275130
rect 538416 271046 538444 277766
rect 539888 271697 539916 277780
rect 541084 275505 541112 277780
rect 541360 277766 542294 277794
rect 541070 275496 541126 275505
rect 541070 275431 541126 275440
rect 539874 271688 539930 271697
rect 539874 271623 539930 271632
rect 538404 271040 538456 271046
rect 538404 270982 538456 270988
rect 538864 271040 538916 271046
rect 538864 270982 538916 270988
rect 538876 267578 538904 270982
rect 541360 267986 541388 277766
rect 543476 273698 543504 277780
rect 543752 277766 544686 277794
rect 545132 277766 545882 277794
rect 546736 277788 547078 277794
rect 546684 277782 547078 277788
rect 546696 277766 547078 277782
rect 547892 277766 548182 277794
rect 543464 273692 543516 273698
rect 543464 273634 543516 273640
rect 543004 271720 543056 271726
rect 543004 271662 543056 271668
rect 543016 270910 543044 271662
rect 543004 270904 543056 270910
rect 543004 270846 543056 270852
rect 543004 270496 543056 270502
rect 543004 270438 543056 270444
rect 543188 270496 543240 270502
rect 543188 270438 543240 270444
rect 543016 269686 543044 270438
rect 543004 269680 543056 269686
rect 543004 269622 543056 269628
rect 543200 269550 543228 270438
rect 543188 269544 543240 269550
rect 543188 269486 543240 269492
rect 541348 267980 541400 267986
rect 541348 267922 541400 267928
rect 538864 267572 538916 267578
rect 538864 267514 538916 267520
rect 543752 266762 543780 277766
rect 543740 266756 543792 266762
rect 543740 266698 543792 266704
rect 537760 265124 537812 265130
rect 537760 265066 537812 265072
rect 545132 264790 545160 277766
rect 547892 268433 547920 277766
rect 549364 275058 549392 277780
rect 549916 277766 550574 277794
rect 549352 275052 549404 275058
rect 549352 274994 549404 275000
rect 549916 269686 549944 277766
rect 551756 271862 551784 277780
rect 552952 275194 552980 277780
rect 553872 277766 554162 277794
rect 552940 275188 552992 275194
rect 552940 275130 552992 275136
rect 552664 274780 552716 274786
rect 552664 274722 552716 274728
rect 551744 271856 551796 271862
rect 551744 271798 551796 271804
rect 551928 271856 551980 271862
rect 551928 271798 551980 271804
rect 551940 271590 551968 271798
rect 551928 271584 551980 271590
rect 551928 271526 551980 271532
rect 549904 269680 549956 269686
rect 549904 269622 549956 269628
rect 547878 268424 547934 268433
rect 547878 268359 547934 268368
rect 550364 267300 550416 267306
rect 550364 267242 550416 267248
rect 550376 266762 550404 267242
rect 550364 266756 550416 266762
rect 550364 266698 550416 266704
rect 552676 265402 552704 274722
rect 553872 271862 553900 277766
rect 555252 273086 555280 277780
rect 556160 275188 556212 275194
rect 556160 275130 556212 275136
rect 555240 273080 555292 273086
rect 555240 273022 555292 273028
rect 556172 272134 556200 275130
rect 556448 274786 556476 277780
rect 557644 277234 557672 277780
rect 557828 277766 558854 277794
rect 559300 277766 560050 277794
rect 557632 277228 557684 277234
rect 557632 277170 557684 277176
rect 556436 274780 556488 274786
rect 556436 274722 556488 274728
rect 556160 272128 556212 272134
rect 556160 272070 556212 272076
rect 553860 271856 553912 271862
rect 553860 271798 553912 271804
rect 554044 271720 554096 271726
rect 554044 271662 554096 271668
rect 554056 266626 554084 271662
rect 557828 270502 557856 277766
rect 557816 270496 557868 270502
rect 557816 270438 557868 270444
rect 554044 266620 554096 266626
rect 554044 266562 554096 266568
rect 559300 265538 559328 277766
rect 561036 276004 561088 276010
rect 561036 275946 561088 275952
rect 561048 273970 561076 275946
rect 561232 275194 561260 277780
rect 562152 277766 562442 277794
rect 561220 275188 561272 275194
rect 561220 275130 561272 275136
rect 561036 273964 561088 273970
rect 561036 273906 561088 273912
rect 562152 271318 562180 277766
rect 563060 275052 563112 275058
rect 563060 274994 563112 275000
rect 562324 271584 562376 271590
rect 562324 271526 562376 271532
rect 562336 271318 562364 271526
rect 562140 271312 562192 271318
rect 562140 271254 562192 271260
rect 562324 271312 562376 271318
rect 562324 271254 562376 271260
rect 563072 268122 563100 274994
rect 563532 274922 563560 277780
rect 563520 274916 563572 274922
rect 563520 274858 563572 274864
rect 564728 272406 564756 277780
rect 565924 276010 565952 277780
rect 566292 277766 567134 277794
rect 565912 276004 565964 276010
rect 565912 275946 565964 275952
rect 564716 272400 564768 272406
rect 564716 272342 564768 272348
rect 563060 268116 563112 268122
rect 563060 268058 563112 268064
rect 566292 266354 566320 277766
rect 568316 273222 568344 277780
rect 569512 274145 569540 277780
rect 570708 276554 570736 277780
rect 570696 276548 570748 276554
rect 570696 276490 570748 276496
rect 569498 274136 569554 274145
rect 569498 274071 569554 274080
rect 568304 273216 568356 273222
rect 568304 273158 568356 273164
rect 571812 272814 571840 277780
rect 572732 277766 573022 277794
rect 571984 277092 572036 277098
rect 571984 277034 572036 277040
rect 571996 276554 572024 277034
rect 571984 276548 572036 276554
rect 571984 276490 572036 276496
rect 572168 273080 572220 273086
rect 572168 273022 572220 273028
rect 571800 272808 571852 272814
rect 571800 272750 571852 272756
rect 571984 272536 572036 272542
rect 571984 272478 572036 272484
rect 571996 272270 572024 272478
rect 571984 272264 572036 272270
rect 571984 272206 572036 272212
rect 572180 267442 572208 273022
rect 572732 268258 572760 277766
rect 574204 277394 574232 277780
rect 574112 277366 574232 277394
rect 572720 268252 572772 268258
rect 572720 268194 572772 268200
rect 572168 267436 572220 267442
rect 572168 267378 572220 267384
rect 566280 266348 566332 266354
rect 566280 266290 566332 266296
rect 559288 265532 559340 265538
rect 559288 265474 559340 265480
rect 552664 265396 552716 265402
rect 552664 265338 552716 265344
rect 545120 264784 545172 264790
rect 545120 264726 545172 264732
rect 574112 264654 574140 277366
rect 575400 272950 575428 277780
rect 575768 277766 576610 277794
rect 575388 272944 575440 272950
rect 575388 272886 575440 272892
rect 575768 266218 575796 277766
rect 577792 275058 577820 277780
rect 578528 277766 578910 277794
rect 577780 275052 577832 275058
rect 577780 274994 577832 275000
rect 578528 272406 578556 277766
rect 578884 272808 578936 272814
rect 578884 272750 578936 272756
rect 578516 272400 578568 272406
rect 578516 272342 578568 272348
rect 578896 267617 578924 272750
rect 580092 271454 580120 277780
rect 581012 277766 581302 277794
rect 580080 271448 580132 271454
rect 580080 271390 580132 271396
rect 581012 268938 581040 277766
rect 581644 276956 581696 276962
rect 581644 276898 581696 276904
rect 581656 276554 581684 276898
rect 581644 276548 581696 276554
rect 581644 276490 581696 276496
rect 582484 272678 582512 277780
rect 582760 277766 583694 277794
rect 583864 277766 584890 277794
rect 585612 277766 586086 277794
rect 582472 272672 582524 272678
rect 582472 272614 582524 272620
rect 582760 270337 582788 277766
rect 582746 270328 582802 270337
rect 582746 270263 582802 270272
rect 581000 268932 581052 268938
rect 581000 268874 581052 268880
rect 583864 268802 583892 277766
rect 585612 272542 585640 277766
rect 587176 277098 587204 277780
rect 587912 277766 588386 277794
rect 589292 277766 589582 277794
rect 591040 277766 591974 277794
rect 587164 277092 587216 277098
rect 587164 277034 587216 277040
rect 585600 272536 585652 272542
rect 585600 272478 585652 272484
rect 585784 272536 585836 272542
rect 585784 272478 585836 272484
rect 583852 268796 583904 268802
rect 583852 268738 583904 268744
rect 578882 267608 578938 267617
rect 578882 267543 578938 267552
rect 585796 267073 585824 272478
rect 587912 269074 587940 277766
rect 587900 269068 587952 269074
rect 587900 269010 587952 269016
rect 585782 267064 585838 267073
rect 585782 266999 585838 267008
rect 575756 266212 575808 266218
rect 575756 266154 575808 266160
rect 589292 266121 589320 277766
rect 589278 266112 589334 266121
rect 591040 266082 591068 277766
rect 593156 272513 593184 277780
rect 593142 272504 593198 272513
rect 593142 272439 593198 272448
rect 594352 271318 594380 277780
rect 594812 277766 595470 277794
rect 594340 271312 594392 271318
rect 594340 271254 594392 271260
rect 594812 268666 594840 277766
rect 596652 277438 596680 277780
rect 596640 277432 596692 277438
rect 596640 277374 596692 277380
rect 597848 271046 597876 277780
rect 599044 276826 599072 277780
rect 599412 277766 600254 277794
rect 600608 277766 601450 277794
rect 601712 277766 602554 277794
rect 603092 277766 603750 277794
rect 599032 276820 599084 276826
rect 599032 276762 599084 276768
rect 597836 271040 597888 271046
rect 597836 270982 597888 270988
rect 599412 270366 599440 277766
rect 599400 270360 599452 270366
rect 599400 270302 599452 270308
rect 594800 268660 594852 268666
rect 594800 268602 594852 268608
rect 594984 268660 595036 268666
rect 594984 268602 595036 268608
rect 594996 266762 595024 268602
rect 594984 266756 595036 266762
rect 594984 266698 595036 266704
rect 589278 266047 589334 266056
rect 591028 266076 591080 266082
rect 591028 266018 591080 266024
rect 574100 264648 574152 264654
rect 574100 264590 574152 264596
rect 600608 264110 600636 277766
rect 601712 265946 601740 277766
rect 601700 265940 601752 265946
rect 601700 265882 601752 265888
rect 603092 264518 603120 277766
rect 604932 275602 604960 277780
rect 606128 276962 606156 277780
rect 607324 277394 607352 277780
rect 607232 277366 607352 277394
rect 606116 276956 606168 276962
rect 606116 276898 606168 276904
rect 604920 275596 604972 275602
rect 604920 275538 604972 275544
rect 607232 268394 607260 277366
rect 608520 273086 608548 277780
rect 608704 277766 609730 277794
rect 608508 273080 608560 273086
rect 608508 273022 608560 273028
rect 608704 268530 608732 277766
rect 610820 274514 610848 277780
rect 612016 275874 612044 277780
rect 612752 277766 613226 277794
rect 612004 275868 612056 275874
rect 612004 275810 612056 275816
rect 610808 274508 610860 274514
rect 610808 274450 610860 274456
rect 608692 268524 608744 268530
rect 608692 268466 608744 268472
rect 607220 268388 607272 268394
rect 607220 268330 607272 268336
rect 612752 264994 612780 277766
rect 614408 274378 614436 277780
rect 614396 274372 614448 274378
rect 614396 274314 614448 274320
rect 615604 271726 615632 277780
rect 616800 275466 616828 277780
rect 616788 275460 616840 275466
rect 616788 275402 616840 275408
rect 617996 274242 618024 277780
rect 619100 275233 619128 277780
rect 619652 277766 620310 277794
rect 619086 275224 619142 275233
rect 619086 275159 619142 275168
rect 619456 274780 619508 274786
rect 619456 274722 619508 274728
rect 617984 274236 618036 274242
rect 617984 274178 618036 274184
rect 615592 271720 615644 271726
rect 615592 271662 615644 271668
rect 619468 270094 619496 274722
rect 619456 270088 619508 270094
rect 619456 270030 619508 270036
rect 619652 265849 619680 277766
rect 621492 274650 621520 277780
rect 621480 274644 621532 274650
rect 621480 274586 621532 274592
rect 622688 272542 622716 277780
rect 623884 274786 623912 277780
rect 623872 274780 623924 274786
rect 623872 274722 623924 274728
rect 625080 274106 625108 277780
rect 625068 274100 625120 274106
rect 625068 274042 625120 274048
rect 622676 272536 622728 272542
rect 622676 272478 622728 272484
rect 626184 271425 626212 277780
rect 626552 277766 627394 277794
rect 626170 271416 626226 271425
rect 626170 271351 626226 271360
rect 626552 269958 626580 277766
rect 628576 273834 628604 277780
rect 629312 277766 629786 277794
rect 630692 277766 630982 277794
rect 628564 273828 628616 273834
rect 628564 273770 628616 273776
rect 626540 269952 626592 269958
rect 626540 269894 626592 269900
rect 629312 266898 629340 277766
rect 630692 270065 630720 277766
rect 632164 273873 632192 277780
rect 633360 275738 633388 277780
rect 633636 277766 634478 277794
rect 633348 275732 633400 275738
rect 633348 275674 633400 275680
rect 632704 273964 632756 273970
rect 632704 273906 632756 273912
rect 632150 273864 632206 273873
rect 632150 273799 632206 273808
rect 630678 270056 630734 270065
rect 630678 269991 630734 270000
rect 632716 267034 632744 273906
rect 633636 270230 633664 277766
rect 635660 276010 635688 277780
rect 635648 276004 635700 276010
rect 635648 275946 635700 275952
rect 636856 272814 636884 277780
rect 637592 277766 638066 277794
rect 636844 272808 636896 272814
rect 636844 272750 636896 272756
rect 633624 270224 633676 270230
rect 633624 270166 633676 270172
rect 637592 269822 637620 277766
rect 639248 271182 639276 277780
rect 640444 275330 640472 277780
rect 640628 277766 641654 277794
rect 640432 275324 640484 275330
rect 640432 275266 640484 275272
rect 639236 271176 639288 271182
rect 639236 271118 639288 271124
rect 637580 269816 637632 269822
rect 637580 269758 637632 269764
rect 638316 269816 638368 269822
rect 640628 269793 640656 277766
rect 642744 271153 642772 277780
rect 643744 274712 643796 274718
rect 643744 274654 643796 274660
rect 642730 271144 642786 271153
rect 642730 271079 642786 271088
rect 638316 269758 638368 269764
rect 640614 269784 640670 269793
rect 638328 267170 638356 269758
rect 640614 269719 640670 269728
rect 638316 267164 638368 267170
rect 638316 267106 638368 267112
rect 632704 267028 632756 267034
rect 632704 266970 632756 266976
rect 629300 266892 629352 266898
rect 629300 266834 629352 266840
rect 619638 265840 619694 265849
rect 619638 265775 619694 265784
rect 612740 264988 612792 264994
rect 612740 264930 612792 264936
rect 603080 264512 603132 264518
rect 603080 264454 603132 264460
rect 643756 264382 643784 274654
rect 643940 273970 643968 277780
rect 643928 273964 643980 273970
rect 643928 273906 643980 273912
rect 643744 264376 643796 264382
rect 643744 264318 643796 264324
rect 507124 264104 507176 264110
rect 507124 264046 507176 264052
rect 600596 264104 600648 264110
rect 600596 264046 600648 264052
rect 511538 262712 511594 262721
rect 511538 262647 511594 262656
rect 511552 261526 511580 262647
rect 511540 261520 511592 261526
rect 511540 261462 511592 261468
rect 568580 261520 568632 261526
rect 568580 261462 568632 261468
rect 510986 260264 511042 260273
rect 510986 260199 511042 260208
rect 511000 259486 511028 260199
rect 510988 259480 511040 259486
rect 510988 259422 511040 259428
rect 514024 259480 514076 259486
rect 514024 259422 514076 259428
rect 510802 257816 510858 257825
rect 510802 257751 510858 257760
rect 510816 256766 510844 257751
rect 510804 256760 510856 256766
rect 510804 256702 510856 256708
rect 511538 255368 511594 255377
rect 511538 255303 511594 255312
rect 511552 250510 511580 255303
rect 511906 252920 511962 252929
rect 511906 252855 511962 252864
rect 511920 252618 511948 252855
rect 511908 252612 511960 252618
rect 511908 252554 511960 252560
rect 511540 250504 511592 250510
rect 510802 250472 510858 250481
rect 511540 250446 511592 250452
rect 510802 250407 510858 250416
rect 129096 247512 129148 247518
rect 129148 247460 129228 247466
rect 129096 247454 129228 247460
rect 129108 247438 129228 247454
rect 129004 247104 129056 247110
rect 129004 247046 129056 247052
rect 120724 230920 120776 230926
rect 120724 230862 120776 230868
rect 123300 230920 123352 230926
rect 123300 230862 123352 230868
rect 99288 230784 99340 230790
rect 99288 230726 99340 230732
rect 79322 230344 79378 230353
rect 79322 230279 79378 230288
rect 90364 230308 90416 230314
rect 77944 229900 77996 229906
rect 77944 229842 77996 229848
rect 67548 229764 67600 229770
rect 67548 229706 67600 229712
rect 66168 227180 66220 227186
rect 66168 227122 66220 227128
rect 63408 227044 63460 227050
rect 63408 226986 63460 226992
rect 62764 223032 62816 223038
rect 62764 222974 62816 222980
rect 62028 222896 62080 222902
rect 62028 222838 62080 222844
rect 60648 221604 60700 221610
rect 60648 221546 60700 221552
rect 59360 221468 59412 221474
rect 59360 221410 59412 221416
rect 59372 218074 59400 221410
rect 59820 219020 59872 219026
rect 59820 218962 59872 218968
rect 59360 218068 59412 218074
rect 59360 218010 59412 218016
rect 55646 217110 55720 217138
rect 56474 217110 56548 217138
rect 57302 217110 57376 217138
rect 58130 217110 58204 217138
rect 58958 217246 59032 217274
rect 55646 216988 55674 217110
rect 56474 216988 56502 217110
rect 57302 216988 57330 217110
rect 58130 216988 58158 217110
rect 58958 216988 58986 217246
rect 59832 217138 59860 218962
rect 60660 217274 60688 221546
rect 62040 218074 62068 222838
rect 63132 219428 63184 219434
rect 63132 219370 63184 219376
rect 61476 218068 61528 218074
rect 61476 218010 61528 218016
rect 62028 218068 62080 218074
rect 62028 218010 62080 218016
rect 62304 218068 62356 218074
rect 62304 218010 62356 218016
rect 59786 217110 59860 217138
rect 60614 217246 60688 217274
rect 59786 216988 59814 217110
rect 60614 216988 60642 217246
rect 61488 217138 61516 218010
rect 62316 217138 62344 218010
rect 63144 217138 63172 219370
rect 63420 218074 63448 226986
rect 64788 226296 64840 226302
rect 64788 226238 64840 226244
rect 64604 219156 64656 219162
rect 64604 219098 64656 219104
rect 63408 218068 63460 218074
rect 63408 218010 63460 218016
rect 63960 218068 64012 218074
rect 63960 218010 64012 218016
rect 63972 217138 64000 218010
rect 64616 217274 64644 219098
rect 64800 218074 64828 226238
rect 66180 218074 66208 227122
rect 67560 219434 67588 229706
rect 69572 228132 69624 228138
rect 69572 228074 69624 228080
rect 68928 227452 68980 227458
rect 68928 227394 68980 227400
rect 68742 222864 68798 222873
rect 68742 222799 68798 222808
rect 67284 219406 67588 219434
rect 66444 218204 66496 218210
rect 66444 218146 66496 218152
rect 64788 218068 64840 218074
rect 64788 218010 64840 218016
rect 65616 218068 65668 218074
rect 65616 218010 65668 218016
rect 66168 218068 66220 218074
rect 66168 218010 66220 218016
rect 64616 217246 64782 217274
rect 61442 217110 61516 217138
rect 62270 217110 62344 217138
rect 63098 217110 63172 217138
rect 63926 217110 64000 217138
rect 61442 216988 61470 217110
rect 62270 216988 62298 217110
rect 63098 216988 63126 217110
rect 63926 216988 63954 217110
rect 64754 216988 64782 217246
rect 65628 217138 65656 218010
rect 66456 217138 66484 218146
rect 67284 217274 67312 219406
rect 68756 218074 68784 222799
rect 68100 218068 68152 218074
rect 68100 218010 68152 218016
rect 68744 218068 68796 218074
rect 68744 218010 68796 218016
rect 65582 217110 65656 217138
rect 66410 217110 66484 217138
rect 67238 217246 67312 217274
rect 65582 216988 65610 217110
rect 66410 216988 66438 217110
rect 67238 216988 67266 217246
rect 68112 217138 68140 218010
rect 68940 217274 68968 227394
rect 69584 218210 69612 228074
rect 73712 227316 73764 227322
rect 73712 227258 73764 227264
rect 71410 223136 71466 223145
rect 71410 223071 71466 223080
rect 69756 220108 69808 220114
rect 69756 220050 69808 220056
rect 69572 218204 69624 218210
rect 69572 218146 69624 218152
rect 69768 217274 69796 220050
rect 70584 218884 70636 218890
rect 70584 218826 70636 218832
rect 68066 217110 68140 217138
rect 68894 217246 68968 217274
rect 69722 217246 69796 217274
rect 68066 216988 68094 217110
rect 68894 216988 68922 217246
rect 69722 216988 69750 217246
rect 70596 217138 70624 218826
rect 71424 217274 71452 223071
rect 73066 220144 73122 220153
rect 73066 220079 73122 220088
rect 72240 218068 72292 218074
rect 72240 218010 72292 218016
rect 70550 217110 70624 217138
rect 71378 217246 71452 217274
rect 70550 216988 70578 217110
rect 71378 216988 71406 217246
rect 72252 217138 72280 218010
rect 73080 217274 73108 220079
rect 73724 218074 73752 227258
rect 75736 225616 75788 225622
rect 75736 225558 75788 225564
rect 75552 223032 75604 223038
rect 75552 222974 75604 222980
rect 73896 221740 73948 221746
rect 73896 221682 73948 221688
rect 73712 218068 73764 218074
rect 73712 218010 73764 218016
rect 73908 217274 73936 221682
rect 75564 218074 75592 222974
rect 74724 218068 74776 218074
rect 74724 218010 74776 218016
rect 75552 218068 75604 218074
rect 75552 218010 75604 218016
rect 72206 217110 72280 217138
rect 73034 217246 73108 217274
rect 73862 217246 73936 217274
rect 72206 216988 72234 217110
rect 73034 216988 73062 217246
rect 73862 216988 73890 217246
rect 74736 217138 74764 218010
rect 75748 217274 75776 225558
rect 77956 221746 77984 229842
rect 79336 221746 79364 230279
rect 90364 230250 90416 230256
rect 83464 230036 83516 230042
rect 83464 229978 83516 229984
rect 82728 224392 82780 224398
rect 82728 224334 82780 224340
rect 81348 223168 81400 223174
rect 81348 223110 81400 223116
rect 79692 222080 79744 222086
rect 79692 222022 79744 222028
rect 77944 221740 77996 221746
rect 77944 221682 77996 221688
rect 79324 221740 79376 221746
rect 79324 221682 79376 221688
rect 78864 221604 78916 221610
rect 78864 221546 78916 221552
rect 76380 220244 76432 220250
rect 76380 220186 76432 220192
rect 76392 217274 76420 220186
rect 77206 218648 77262 218657
rect 77206 218583 77262 218592
rect 78036 218612 78088 218618
rect 74690 217110 74764 217138
rect 75518 217246 75776 217274
rect 76346 217246 76420 217274
rect 74690 216988 74718 217110
rect 75518 216988 75546 217246
rect 76346 216988 76374 217246
rect 77220 217138 77248 218583
rect 78036 218554 78088 218560
rect 78048 217138 78076 218554
rect 78876 217274 78904 221546
rect 79704 217274 79732 222022
rect 80520 221944 80572 221950
rect 80520 221886 80572 221892
rect 80532 217274 80560 221886
rect 81360 217274 81388 223110
rect 82740 218074 82768 224334
rect 83476 221950 83504 229978
rect 87604 229084 87656 229090
rect 87604 229026 87656 229032
rect 85488 228676 85540 228682
rect 85488 228618 85540 228624
rect 85304 224664 85356 224670
rect 85304 224606 85356 224612
rect 83464 221944 83516 221950
rect 83464 221886 83516 221892
rect 83004 221740 83056 221746
rect 83004 221682 83056 221688
rect 82176 218068 82228 218074
rect 82176 218010 82228 218016
rect 82728 218068 82780 218074
rect 82728 218010 82780 218016
rect 77174 217110 77248 217138
rect 78002 217110 78076 217138
rect 78830 217246 78904 217274
rect 79658 217246 79732 217274
rect 80486 217246 80560 217274
rect 81314 217246 81388 217274
rect 77174 216988 77202 217110
rect 78002 216988 78030 217110
rect 78830 216988 78858 217246
rect 79658 216988 79686 217246
rect 80486 216988 80514 217246
rect 81314 216988 81342 217246
rect 82188 217138 82216 218010
rect 83016 217274 83044 221682
rect 83188 220788 83240 220794
rect 83188 220730 83240 220736
rect 83200 219502 83228 220730
rect 83188 219496 83240 219502
rect 83188 219438 83240 219444
rect 83832 219020 83884 219026
rect 83832 218962 83884 218968
rect 82142 217110 82216 217138
rect 82970 217246 83044 217274
rect 82142 216988 82170 217110
rect 82970 216988 82998 217246
rect 83844 217138 83872 218962
rect 85316 218074 85344 224606
rect 84660 218068 84712 218074
rect 84660 218010 84712 218016
rect 85304 218068 85356 218074
rect 85304 218010 85356 218016
rect 84672 217138 84700 218010
rect 85500 217274 85528 228618
rect 87144 221332 87196 221338
rect 87144 221274 87196 221280
rect 86316 221196 86368 221202
rect 86316 221138 86368 221144
rect 86328 217274 86356 221138
rect 87156 217274 87184 221274
rect 87616 219162 87644 229026
rect 89628 224528 89680 224534
rect 89628 224470 89680 224476
rect 88984 222352 89036 222358
rect 88984 222294 89036 222300
rect 88800 222012 88852 222018
rect 88800 221954 88852 221960
rect 88812 221746 88840 221954
rect 88800 221740 88852 221746
rect 88800 221682 88852 221688
rect 88996 219298 89024 222294
rect 89260 221876 89312 221882
rect 89260 221818 89312 221824
rect 89272 221202 89300 221818
rect 89260 221196 89312 221202
rect 89260 221138 89312 221144
rect 88984 219292 89036 219298
rect 88984 219234 89036 219240
rect 87604 219156 87656 219162
rect 87604 219098 87656 219104
rect 87972 219156 88024 219162
rect 87972 219098 88024 219104
rect 83798 217110 83872 217138
rect 84626 217110 84700 217138
rect 85454 217246 85528 217274
rect 86282 217246 86356 217274
rect 87110 217246 87184 217274
rect 83798 216988 83826 217110
rect 84626 216988 84654 217110
rect 85454 216988 85482 217246
rect 86282 216988 86310 217246
rect 87110 216988 87138 217246
rect 87984 217138 88012 219098
rect 89444 218340 89496 218346
rect 89444 218282 89496 218288
rect 88800 218068 88852 218074
rect 88800 218010 88852 218016
rect 88812 217138 88840 218010
rect 89456 217274 89484 218282
rect 89640 218074 89668 224470
rect 90376 221338 90404 230250
rect 96436 228268 96488 228274
rect 96436 228210 96488 228216
rect 93768 227588 93820 227594
rect 93768 227530 93820 227536
rect 93584 225752 93636 225758
rect 93584 225694 93636 225700
rect 92112 223984 92164 223990
rect 92112 223926 92164 223932
rect 91284 222148 91336 222154
rect 91284 222090 91336 222096
rect 90364 221332 90416 221338
rect 90364 221274 90416 221280
rect 90456 218204 90508 218210
rect 90456 218146 90508 218152
rect 89628 218068 89680 218074
rect 89628 218010 89680 218016
rect 89456 217246 89622 217274
rect 87938 217110 88012 217138
rect 88766 217110 88840 217138
rect 87938 216988 87966 217110
rect 88766 216988 88794 217110
rect 89594 216988 89622 217246
rect 90468 217138 90496 218146
rect 91296 217274 91324 222090
rect 92124 217274 92152 223926
rect 93596 218074 93624 225694
rect 92940 218068 92992 218074
rect 92940 218010 92992 218016
rect 93584 218068 93636 218074
rect 93584 218010 93636 218016
rect 90422 217110 90496 217138
rect 91250 217246 91324 217274
rect 92078 217246 92152 217274
rect 90422 216988 90450 217110
rect 91250 216988 91278 217246
rect 92078 216988 92106 217246
rect 92952 217138 92980 218010
rect 93780 217274 93808 227530
rect 96252 224936 96304 224942
rect 96252 224878 96304 224884
rect 94596 220380 94648 220386
rect 94596 220322 94648 220328
rect 94608 217274 94636 220322
rect 96264 218346 96292 224878
rect 95424 218340 95476 218346
rect 95424 218282 95476 218288
rect 96252 218340 96304 218346
rect 96252 218282 96304 218288
rect 92906 217110 92980 217138
rect 93734 217246 93808 217274
rect 94562 217246 94636 217274
rect 92906 216988 92934 217110
rect 93734 216988 93762 217246
rect 94562 216988 94590 217246
rect 95436 217138 95464 218282
rect 96448 217274 96476 228210
rect 97908 223304 97960 223310
rect 97908 223246 97960 223252
rect 97724 221196 97776 221202
rect 97724 221138 97776 221144
rect 97736 219434 97764 221138
rect 97920 219434 97948 223246
rect 97080 219428 97132 219434
rect 97736 219406 97856 219434
rect 97920 219428 98052 219434
rect 97920 219406 98000 219428
rect 97080 219370 97132 219376
rect 95390 217110 95464 217138
rect 96218 217246 96476 217274
rect 95390 216988 95418 217110
rect 96218 216988 96246 217246
rect 97092 217138 97120 219370
rect 97828 217274 97856 219406
rect 98000 219370 98052 219376
rect 99300 218074 99328 230726
rect 113088 230648 113140 230654
rect 113088 230590 113140 230596
rect 107568 230444 107620 230450
rect 107568 230386 107620 230392
rect 100668 228540 100720 228546
rect 100668 228482 100720 228488
rect 100392 219292 100444 219298
rect 100392 219234 100444 219240
rect 98736 218068 98788 218074
rect 98736 218010 98788 218016
rect 99288 218068 99340 218074
rect 99288 218010 99340 218016
rect 99564 218068 99616 218074
rect 99564 218010 99616 218016
rect 97828 217246 97902 217274
rect 97046 217110 97120 217138
rect 97046 216988 97074 217110
rect 97874 216988 97902 217246
rect 98748 217138 98776 218010
rect 99576 217138 99604 218010
rect 100404 217138 100432 219234
rect 100680 218074 100708 228482
rect 107580 225894 107608 230386
rect 110328 228812 110380 228818
rect 110328 228754 110380 228760
rect 107568 225888 107620 225894
rect 107568 225830 107620 225836
rect 107568 225208 107620 225214
rect 107568 225150 107620 225156
rect 106188 224800 106240 224806
rect 106188 224742 106240 224748
rect 101404 224120 101456 224126
rect 101404 224062 101456 224068
rect 101416 219162 101444 224062
rect 102048 221332 102100 221338
rect 102048 221274 102100 221280
rect 101404 219156 101456 219162
rect 101404 219098 101456 219104
rect 100668 218068 100720 218074
rect 100668 218010 100720 218016
rect 101220 218068 101272 218074
rect 101220 218010 101272 218016
rect 101232 217138 101260 218010
rect 102060 217274 102088 221274
rect 104532 221060 104584 221066
rect 104532 221002 104584 221008
rect 103428 220516 103480 220522
rect 103428 220458 103480 220464
rect 103440 218074 103468 220458
rect 103704 218340 103756 218346
rect 103704 218282 103756 218288
rect 103428 218068 103480 218074
rect 103428 218010 103480 218016
rect 98702 217110 98776 217138
rect 99530 217110 99604 217138
rect 100358 217110 100432 217138
rect 101186 217110 101260 217138
rect 102014 217246 102088 217274
rect 102830 217252 102882 217258
rect 98702 216988 98730 217110
rect 99530 216988 99558 217110
rect 100358 216988 100386 217110
rect 101186 216988 101214 217110
rect 102014 216988 102042 217246
rect 102830 217194 102882 217200
rect 102842 216988 102870 217194
rect 103716 217138 103744 218282
rect 104544 217274 104572 221002
rect 106200 218074 106228 224742
rect 107580 218074 107608 225150
rect 108672 223440 108724 223446
rect 108672 223382 108724 223388
rect 107844 220652 107896 220658
rect 107844 220594 107896 220600
rect 105360 218068 105412 218074
rect 105360 218010 105412 218016
rect 106188 218068 106240 218074
rect 106188 218010 106240 218016
rect 107016 218068 107068 218074
rect 107016 218010 107068 218016
rect 107568 218068 107620 218074
rect 107568 218010 107620 218016
rect 103670 217110 103744 217138
rect 104498 217246 104572 217274
rect 103670 216988 103698 217110
rect 104498 216988 104526 217246
rect 105372 217138 105400 218010
rect 106188 217456 106240 217462
rect 106188 217398 106240 217404
rect 106200 217138 106228 217398
rect 107028 217138 107056 218010
rect 107856 217274 107884 220594
rect 108304 219428 108356 219434
rect 108304 219370 108356 219376
rect 108316 218618 108344 219370
rect 108304 218612 108356 218618
rect 108304 218554 108356 218560
rect 108684 217274 108712 223382
rect 110144 218476 110196 218482
rect 110144 218418 110196 218424
rect 109500 218068 109552 218074
rect 109500 218010 109552 218016
rect 105326 217110 105400 217138
rect 106154 217110 106228 217138
rect 106982 217110 107056 217138
rect 107810 217246 107884 217274
rect 108638 217246 108712 217274
rect 105326 216988 105354 217110
rect 106154 216988 106182 217110
rect 106982 216988 107010 217110
rect 107810 216988 107838 217246
rect 108638 216988 108666 217246
rect 109512 217138 109540 218010
rect 110156 217274 110184 218418
rect 110340 218074 110368 228754
rect 111708 227724 111760 227730
rect 111708 227666 111760 227672
rect 111720 218074 111748 227666
rect 113100 218618 113128 230590
rect 117872 230444 117924 230450
rect 117872 230386 117924 230392
rect 117228 226908 117280 226914
rect 117228 226850 117280 226856
rect 115296 225888 115348 225894
rect 115296 225830 115348 225836
rect 113824 223848 113876 223854
rect 113824 223790 113876 223796
rect 113836 219434 113864 223790
rect 113824 219428 113876 219434
rect 113824 219370 113876 219376
rect 114468 219428 114520 219434
rect 114468 219370 114520 219376
rect 113640 219156 113692 219162
rect 113640 219098 113692 219104
rect 111984 218612 112036 218618
rect 111984 218554 112036 218560
rect 113088 218612 113140 218618
rect 113088 218554 113140 218560
rect 110328 218068 110380 218074
rect 110328 218010 110380 218016
rect 111156 218068 111208 218074
rect 111156 218010 111208 218016
rect 111708 218068 111760 218074
rect 111708 218010 111760 218016
rect 110156 217246 110322 217274
rect 109466 217110 109540 217138
rect 109466 216988 109494 217110
rect 110294 216988 110322 217246
rect 111168 217138 111196 218010
rect 111996 217138 112024 218554
rect 112812 218068 112864 218074
rect 112812 218010 112864 218016
rect 112824 217138 112852 218010
rect 113652 217138 113680 219098
rect 114480 217138 114508 219370
rect 115308 217274 115336 225830
rect 116952 225072 117004 225078
rect 116952 225014 117004 225020
rect 116124 218476 116176 218482
rect 116124 218418 116176 218424
rect 111122 217110 111196 217138
rect 111950 217110 112024 217138
rect 112778 217110 112852 217138
rect 113606 217110 113680 217138
rect 114434 217110 114508 217138
rect 115262 217246 115336 217274
rect 111122 216988 111150 217110
rect 111950 216988 111978 217110
rect 112778 216988 112806 217110
rect 113606 216988 113634 217110
rect 114434 216988 114462 217110
rect 115262 216988 115290 217246
rect 116136 217138 116164 218418
rect 116964 217274 116992 225014
rect 117240 218482 117268 226850
rect 117884 225078 117912 230386
rect 119988 228948 120040 228954
rect 119988 228890 120040 228896
rect 118608 226160 118660 226166
rect 118608 226102 118660 226108
rect 117872 225072 117924 225078
rect 117872 225014 117924 225020
rect 117780 220924 117832 220930
rect 117780 220866 117832 220872
rect 117228 218476 117280 218482
rect 117228 218418 117280 218424
rect 117792 217274 117820 220866
rect 118620 217274 118648 226102
rect 120000 218482 120028 228890
rect 120356 218612 120408 218618
rect 120356 218554 120408 218560
rect 119436 218476 119488 218482
rect 119436 218418 119488 218424
rect 119988 218476 120040 218482
rect 119988 218418 120040 218424
rect 116090 217110 116164 217138
rect 116918 217246 116992 217274
rect 117746 217246 117820 217274
rect 118574 217246 118648 217274
rect 116090 216988 116118 217110
rect 116918 216988 116946 217246
rect 117746 216988 117774 217246
rect 118574 216988 118602 217246
rect 119448 217138 119476 218418
rect 120368 217274 120396 218554
rect 120736 218482 120764 230862
rect 123312 230518 123340 230862
rect 123300 230512 123352 230518
rect 123300 230454 123352 230460
rect 123116 230444 123168 230450
rect 123116 230386 123168 230392
rect 123128 230178 123156 230386
rect 122932 230172 122984 230178
rect 122932 230114 122984 230120
rect 123116 230172 123168 230178
rect 123116 230114 123168 230120
rect 122944 229634 122972 230114
rect 122932 229628 122984 229634
rect 122932 229570 122984 229576
rect 126888 229356 126940 229362
rect 126888 229298 126940 229304
rect 125692 226296 125744 226302
rect 125692 226238 125744 226244
rect 125876 226296 125928 226302
rect 125876 226238 125928 226244
rect 122748 226024 122800 226030
rect 122748 225966 122800 225972
rect 121092 223576 121144 223582
rect 121092 223518 121144 223524
rect 120908 219156 120960 219162
rect 120908 219098 120960 219104
rect 120920 218482 120948 219098
rect 120724 218476 120776 218482
rect 120724 218418 120776 218424
rect 120908 218476 120960 218482
rect 120908 218418 120960 218424
rect 121104 217274 121132 223518
rect 122760 219162 122788 225966
rect 125232 225480 125284 225486
rect 125232 225422 125284 225428
rect 124404 219972 124456 219978
rect 124404 219914 124456 219920
rect 121920 219156 121972 219162
rect 121920 219098 121972 219104
rect 122748 219156 122800 219162
rect 122748 219098 122800 219104
rect 123576 219156 123628 219162
rect 123576 219098 123628 219104
rect 119402 217110 119476 217138
rect 120230 217246 120396 217274
rect 121058 217246 121132 217274
rect 119402 216988 119430 217110
rect 120230 216988 120258 217246
rect 121058 216988 121086 217246
rect 121932 217138 121960 219098
rect 122748 217592 122800 217598
rect 122748 217534 122800 217540
rect 122760 217138 122788 217534
rect 123588 217138 123616 219098
rect 124416 217274 124444 219914
rect 125244 217274 125272 225422
rect 125704 225350 125732 226238
rect 125888 226030 125916 226238
rect 125876 226024 125928 226030
rect 125876 225966 125928 225972
rect 125692 225344 125744 225350
rect 125692 225286 125744 225292
rect 126060 219836 126112 219842
rect 126060 219778 126112 219784
rect 125520 219406 125732 219434
rect 125520 218618 125548 219406
rect 125704 218618 125732 219406
rect 125508 218612 125560 218618
rect 125508 218554 125560 218560
rect 125692 218612 125744 218618
rect 125692 218554 125744 218560
rect 126072 217274 126100 219778
rect 126426 219192 126482 219201
rect 126426 219127 126428 219136
rect 126480 219127 126482 219136
rect 126612 219156 126664 219162
rect 126428 219098 126480 219104
rect 126612 219098 126664 219104
rect 126624 218482 126652 219098
rect 126612 218476 126664 218482
rect 126612 218418 126664 218424
rect 126900 217274 126928 229298
rect 128268 222760 128320 222766
rect 128268 222702 128320 222708
rect 128280 218482 128308 222702
rect 129016 221785 129044 247046
rect 129200 230994 129228 247438
rect 510816 246362 510844 250407
rect 510986 248024 511042 248033
rect 510986 247959 511042 247968
rect 511000 247178 511028 247959
rect 510988 247172 511040 247178
rect 510988 247114 511040 247120
rect 512644 247172 512696 247178
rect 512644 247114 512696 247120
rect 510804 246356 510856 246362
rect 510804 246298 510856 246304
rect 131762 245712 131818 245721
rect 131762 245647 131818 245656
rect 129188 230988 129240 230994
rect 129188 230930 129240 230936
rect 130108 229492 130160 229498
rect 130108 229434 130160 229440
rect 129556 226636 129608 226642
rect 129556 226578 129608 226584
rect 129372 226296 129424 226302
rect 129372 226238 129424 226244
rect 129384 224954 129412 226238
rect 129568 224954 129596 226578
rect 130120 225214 130148 229434
rect 130108 225208 130160 225214
rect 130108 225150 130160 225156
rect 129292 224926 129412 224954
rect 129476 224926 129596 224954
rect 129002 221776 129058 221785
rect 129002 221711 129058 221720
rect 128452 219632 128504 219638
rect 128452 219574 128504 219580
rect 128464 219178 128492 219574
rect 128634 219192 128690 219201
rect 128464 219162 128538 219178
rect 128464 219156 128550 219162
rect 128464 219150 128498 219156
rect 128634 219127 128636 219136
rect 128498 219098 128550 219104
rect 128688 219127 128690 219136
rect 128636 219098 128688 219104
rect 129292 218482 129320 224926
rect 127716 218476 127768 218482
rect 127716 218418 127768 218424
rect 128268 218476 128320 218482
rect 128268 218418 128320 218424
rect 128544 218476 128596 218482
rect 128544 218418 128596 218424
rect 129280 218476 129332 218482
rect 129280 218418 129332 218424
rect 121886 217110 121960 217138
rect 122714 217110 122788 217138
rect 123542 217110 123616 217138
rect 124370 217246 124444 217274
rect 125198 217246 125272 217274
rect 126026 217246 126100 217274
rect 126854 217246 126928 217274
rect 121886 216988 121914 217110
rect 122714 216988 122742 217110
rect 123542 216988 123570 217110
rect 124370 216988 124398 217246
rect 125198 216988 125226 217246
rect 126026 216988 126054 217246
rect 126854 216988 126882 217246
rect 127728 217138 127756 218418
rect 128556 217138 128584 218418
rect 129476 217274 129504 224926
rect 129740 223712 129792 223718
rect 129740 223654 129792 223660
rect 129752 219638 129780 223654
rect 131028 222488 131080 222494
rect 131028 222430 131080 222436
rect 129740 219632 129792 219638
rect 129740 219574 129792 219580
rect 130198 218920 130254 218929
rect 130198 218855 130254 218864
rect 127682 217110 127756 217138
rect 128510 217110 128584 217138
rect 129338 217246 129504 217274
rect 127682 216988 127710 217110
rect 128510 216988 128538 217110
rect 129338 216988 129366 217246
rect 130212 217138 130240 218855
rect 131040 217138 131068 222430
rect 131776 222057 131804 245647
rect 511262 245576 511318 245585
rect 511262 245511 511318 245520
rect 511276 242214 511304 245511
rect 511906 243128 511962 243137
rect 511906 243063 511962 243072
rect 511264 242208 511316 242214
rect 511264 242150 511316 242156
rect 511920 240786 511948 243063
rect 511908 240780 511960 240786
rect 511908 240722 511960 240728
rect 511078 240680 511134 240689
rect 511078 240615 511134 240624
rect 510894 235784 510950 235793
rect 510894 235719 510950 235728
rect 510908 234054 510936 235719
rect 510896 234048 510948 234054
rect 510896 233990 510948 233996
rect 511092 233918 511120 240615
rect 511262 238232 511318 238241
rect 511262 238167 511318 238176
rect 511080 233912 511132 233918
rect 511080 233854 511132 233860
rect 507490 233064 507546 233073
rect 507490 232999 507546 233008
rect 164896 231946 165186 231962
rect 191392 231946 191682 231962
rect 157340 231940 157392 231946
rect 157340 231882 157392 231888
rect 164884 231940 165186 231946
rect 164936 231934 165186 231940
rect 190460 231940 190512 231946
rect 164884 231882 164936 231888
rect 190460 231882 190512 231888
rect 191380 231940 191682 231946
rect 191432 231934 191682 231940
rect 191380 231882 191432 231888
rect 147126 231296 147182 231305
rect 147126 231231 147182 231240
rect 144274 230888 144330 230897
rect 144274 230823 144330 230832
rect 132866 230616 132922 230625
rect 132866 230551 132922 230560
rect 132880 229634 132908 230551
rect 140778 230344 140834 230353
rect 140778 230279 140834 230288
rect 133052 229900 133104 229906
rect 133052 229842 133104 229848
rect 133236 229900 133288 229906
rect 133236 229842 133288 229848
rect 132868 229628 132920 229634
rect 132868 229570 132920 229576
rect 133064 229226 133092 229842
rect 133248 229498 133276 229842
rect 140792 229537 140820 230279
rect 140778 229528 140834 229537
rect 133236 229492 133288 229498
rect 140778 229463 140834 229472
rect 133236 229434 133288 229440
rect 133696 229356 133748 229362
rect 133696 229298 133748 229304
rect 133052 229220 133104 229226
rect 133052 229162 133104 229168
rect 133512 227996 133564 228002
rect 133512 227938 133564 227944
rect 132408 225208 132460 225214
rect 132408 225150 132460 225156
rect 131762 222048 131818 222057
rect 131762 221983 131818 221992
rect 132420 219434 132448 225150
rect 133524 224954 133552 227938
rect 133708 224954 133736 229298
rect 133880 229220 133932 229226
rect 133880 229162 133932 229168
rect 133892 225350 133920 229162
rect 136548 227860 136600 227866
rect 136548 227802 136600 227808
rect 133880 225344 133932 225350
rect 133880 225286 133932 225292
rect 135076 225072 135128 225078
rect 135076 225014 135128 225020
rect 133432 224926 133552 224954
rect 133616 224926 133736 224954
rect 133144 223440 133196 223446
rect 133144 223382 133196 223388
rect 133156 222630 133184 223382
rect 133144 222624 133196 222630
rect 133144 222566 133196 222572
rect 133432 219434 133460 224926
rect 131672 219428 131724 219434
rect 131672 219370 131724 219376
rect 131856 219428 131908 219434
rect 131856 219370 131908 219376
rect 132408 219428 132460 219434
rect 132408 219370 132460 219376
rect 132684 219428 132736 219434
rect 132684 219370 132736 219376
rect 133420 219428 133472 219434
rect 133420 219370 133472 219376
rect 131684 218482 131712 219370
rect 131672 218476 131724 218482
rect 131672 218418 131724 218424
rect 131868 217138 131896 219370
rect 132696 217138 132724 219370
rect 133616 217274 133644 224926
rect 133788 223440 133840 223446
rect 133788 223382 133840 223388
rect 133800 222494 133828 223382
rect 133788 222488 133840 222494
rect 133788 222430 133840 222436
rect 134340 217728 134392 217734
rect 134340 217670 134392 217676
rect 130166 217110 130240 217138
rect 130994 217110 131068 217138
rect 131822 217110 131896 217138
rect 132650 217110 132724 217138
rect 133478 217246 133644 217274
rect 130166 216988 130194 217110
rect 130994 216988 131022 217110
rect 131822 216988 131850 217110
rect 132650 216988 132678 217110
rect 133478 216988 133506 217246
rect 134352 217138 134380 217670
rect 135088 217274 135116 225014
rect 136560 219434 136588 227802
rect 139308 226500 139360 226506
rect 139308 226442 139360 226448
rect 137468 226296 137520 226302
rect 137468 226238 137520 226244
rect 137100 226160 137152 226166
rect 137100 226102 137152 226108
rect 137112 225350 137140 226102
rect 137100 225344 137152 225350
rect 137100 225286 137152 225292
rect 137480 225078 137508 226238
rect 137468 225072 137520 225078
rect 137468 225014 137520 225020
rect 139124 225072 139176 225078
rect 139124 225014 139176 225020
rect 137652 222488 137704 222494
rect 137652 222430 137704 222436
rect 135996 219428 136048 219434
rect 135996 219370 136048 219376
rect 136548 219428 136600 219434
rect 136548 219370 136600 219376
rect 136824 219428 136876 219434
rect 136824 219370 136876 219376
rect 135088 217246 135162 217274
rect 134306 217110 134380 217138
rect 134306 216988 134334 217110
rect 135134 216988 135162 217246
rect 136008 217138 136036 219370
rect 136836 217138 136864 219370
rect 137664 217138 137692 222430
rect 138296 219700 138348 219706
rect 138296 219642 138348 219648
rect 138308 219434 138336 219642
rect 138296 219428 138348 219434
rect 138296 219370 138348 219376
rect 138480 219428 138532 219434
rect 138480 219370 138532 219376
rect 138492 219201 138520 219370
rect 137926 219192 137982 219201
rect 137926 219127 137982 219136
rect 138478 219192 138534 219201
rect 138478 219127 138534 219136
rect 137940 218482 137968 219127
rect 139136 218482 139164 225014
rect 137928 218476 137980 218482
rect 137928 218418 137980 218424
rect 138480 218476 138532 218482
rect 138480 218418 138532 218424
rect 139124 218476 139176 218482
rect 139124 218418 139176 218424
rect 138492 217138 138520 218418
rect 139320 217274 139348 226442
rect 143446 226400 143502 226409
rect 143446 226335 143502 226344
rect 141606 225992 141662 226001
rect 141606 225927 141662 225936
rect 141620 225350 141648 225927
rect 141608 225344 141660 225350
rect 141608 225286 141660 225292
rect 141792 225344 141844 225350
rect 141792 225286 141844 225292
rect 140686 224224 140742 224233
rect 140686 224159 140742 224168
rect 140700 218482 140728 224159
rect 140964 219564 141016 219570
rect 140964 219506 141016 219512
rect 140136 218476 140188 218482
rect 140136 218418 140188 218424
rect 140688 218476 140740 218482
rect 140688 218418 140740 218424
rect 135962 217110 136036 217138
rect 136790 217110 136864 217138
rect 137618 217110 137692 217138
rect 138446 217110 138520 217138
rect 139274 217246 139348 217274
rect 135962 216988 135990 217110
rect 136790 216988 136818 217110
rect 137618 216988 137646 217110
rect 138446 216988 138474 217110
rect 139274 216988 139302 217246
rect 140148 217138 140176 218418
rect 140976 217274 141004 219506
rect 141148 219428 141200 219434
rect 141148 219370 141200 219376
rect 141160 218618 141188 219370
rect 141148 218612 141200 218618
rect 141148 218554 141200 218560
rect 141804 217274 141832 225286
rect 142158 224496 142214 224505
rect 142158 224431 142214 224440
rect 142172 224346 142200 224431
rect 142126 224318 142200 224346
rect 142126 224262 142154 224318
rect 142114 224256 142166 224262
rect 142252 224256 142304 224262
rect 142114 224198 142166 224204
rect 142250 224224 142252 224233
rect 142304 224224 142306 224233
rect 142250 224159 142306 224168
rect 142250 219192 142306 219201
rect 142250 219127 142306 219136
rect 142264 218618 142292 219127
rect 142252 218612 142304 218618
rect 142252 218554 142304 218560
rect 143460 218482 143488 226335
rect 143632 219700 143684 219706
rect 143632 219642 143684 219648
rect 143644 218482 143672 219642
rect 142620 218476 142672 218482
rect 142620 218418 142672 218424
rect 143448 218476 143500 218482
rect 143448 218418 143500 218424
rect 143632 218476 143684 218482
rect 143632 218418 143684 218424
rect 140102 217110 140176 217138
rect 140930 217246 141004 217274
rect 141758 217246 141832 217274
rect 140102 216988 140130 217110
rect 140930 216988 140958 217246
rect 141758 216988 141786 217246
rect 142632 217138 142660 218418
rect 143446 218104 143502 218113
rect 143446 218039 143502 218048
rect 143460 217138 143488 218039
rect 144288 217274 144316 230823
rect 147140 230518 147168 231231
rect 147310 230888 147366 230897
rect 148060 230874 148088 231676
rect 148520 231662 148626 231690
rect 149072 231662 149178 231690
rect 149440 231662 149730 231690
rect 149992 231662 150282 231690
rect 147366 230846 147536 230874
rect 148060 230846 148180 230874
rect 147310 230823 147366 230832
rect 147310 230616 147366 230625
rect 147310 230551 147366 230560
rect 147128 230512 147180 230518
rect 147128 230454 147180 230460
rect 147034 230344 147090 230353
rect 147034 230279 147036 230288
rect 147088 230279 147090 230288
rect 147324 230296 147352 230551
rect 147508 230382 147536 230846
rect 148152 230602 148180 230846
rect 148060 230574 148180 230602
rect 147496 230376 147548 230382
rect 147496 230318 147548 230324
rect 147324 230268 147444 230296
rect 147036 230250 147088 230256
rect 147416 230194 147444 230268
rect 147416 230166 147720 230194
rect 147692 229226 147720 230166
rect 147312 229220 147364 229226
rect 147312 229162 147364 229168
rect 147680 229220 147732 229226
rect 147680 229162 147732 229168
rect 147324 228857 147352 229162
rect 147494 229120 147550 229129
rect 147494 229055 147496 229064
rect 147548 229055 147550 229064
rect 147634 229084 147686 229090
rect 147496 229026 147548 229032
rect 147634 229026 147686 229032
rect 147646 228970 147674 229026
rect 147508 228942 147674 228970
rect 147310 228848 147366 228857
rect 147310 228783 147366 228792
rect 147508 228002 147536 228942
rect 148060 228256 148088 230574
rect 148520 228290 148548 231662
rect 148690 231296 148746 231305
rect 148690 231231 148746 231240
rect 148874 231296 148930 231305
rect 148874 231231 148930 231240
rect 148704 230625 148732 231231
rect 148690 230616 148746 230625
rect 148690 230551 148746 230560
rect 148336 228262 148548 228290
rect 148060 228228 148180 228256
rect 147956 228132 148008 228138
rect 147956 228074 148008 228080
rect 147496 227996 147548 228002
rect 147496 227938 147548 227944
rect 147680 227996 147732 228002
rect 147680 227938 147732 227944
rect 146116 226772 146168 226778
rect 146116 226714 146168 226720
rect 145930 222592 145986 222601
rect 145930 222527 145986 222536
rect 144734 220416 144790 220425
rect 144734 220351 144790 220360
rect 144460 219496 144512 219502
rect 144460 219438 144512 219444
rect 144472 218618 144500 219438
rect 144748 219201 144776 220351
rect 145012 219564 145064 219570
rect 145012 219506 145064 219512
rect 145024 219434 145052 219506
rect 144932 219406 145052 219434
rect 144734 219192 144790 219201
rect 144734 219127 144790 219136
rect 144932 218754 144960 219406
rect 144920 218748 144972 218754
rect 144920 218690 144972 218696
rect 144460 218612 144512 218618
rect 144460 218554 144512 218560
rect 145944 218482 145972 222527
rect 145104 218476 145156 218482
rect 145104 218418 145156 218424
rect 145932 218476 145984 218482
rect 145932 218418 145984 218424
rect 142586 217110 142660 217138
rect 143414 217110 143488 217138
rect 144242 217246 144316 217274
rect 142586 216988 142614 217110
rect 143414 216988 143442 217110
rect 144242 216988 144270 217246
rect 145116 217138 145144 218418
rect 146128 217274 146156 226714
rect 147692 226409 147720 227938
rect 147968 227905 147996 228074
rect 147954 227896 148010 227905
rect 147954 227831 148010 227840
rect 147678 226400 147734 226409
rect 147678 226335 147734 226344
rect 147956 226296 148008 226302
rect 147956 226238 148008 226244
rect 147968 225622 147996 226238
rect 147772 225616 147824 225622
rect 147772 225558 147824 225564
rect 147956 225616 148008 225622
rect 147956 225558 148008 225564
rect 147784 225457 147812 225558
rect 147770 225448 147826 225457
rect 147770 225383 147826 225392
rect 146666 224224 146722 224233
rect 146666 224159 146722 224168
rect 146680 222902 146708 224159
rect 146668 222896 146720 222902
rect 146668 222838 146720 222844
rect 146944 222896 146996 222902
rect 146944 222838 146996 222844
rect 146956 222630 146984 222838
rect 146944 222624 146996 222630
rect 147128 222624 147180 222630
rect 146944 222566 146996 222572
rect 147126 222592 147128 222601
rect 147180 222592 147182 222601
rect 147126 222527 147182 222536
rect 148152 222194 148180 228228
rect 147692 222166 148180 222194
rect 147036 221468 147088 221474
rect 147036 221410 147088 221416
rect 147220 221468 147272 221474
rect 147220 221410 147272 221416
rect 147048 221241 147076 221410
rect 147034 221232 147090 221241
rect 147034 221167 147090 221176
rect 147232 219298 147260 221410
rect 147692 219722 147720 222166
rect 148336 221241 148364 228262
rect 148508 226160 148560 226166
rect 148508 226102 148560 226108
rect 148520 226001 148548 226102
rect 148506 225992 148562 226001
rect 148506 225927 148562 225936
rect 148888 222358 148916 231231
rect 149072 224505 149100 231662
rect 149440 231033 149468 231662
rect 149426 231024 149482 231033
rect 149426 230959 149482 230968
rect 149336 230308 149388 230314
rect 149336 230250 149388 230256
rect 149348 229770 149376 230250
rect 149336 229764 149388 229770
rect 149336 229706 149388 229712
rect 149992 229129 150020 231662
rect 149978 229120 150034 229129
rect 149978 229055 150034 229064
rect 149244 228132 149296 228138
rect 149244 228074 149296 228080
rect 149058 224496 149114 224505
rect 149058 224431 149114 224440
rect 148876 222352 148928 222358
rect 148876 222294 148928 222300
rect 148322 221232 148378 221241
rect 148322 221167 148378 221176
rect 149256 220425 149284 228074
rect 149518 227760 149574 227769
rect 149518 227695 149574 227704
rect 149532 227186 149560 227695
rect 149520 227180 149572 227186
rect 149520 227122 149572 227128
rect 149888 227044 149940 227050
rect 149888 226986 149940 226992
rect 149242 220416 149298 220425
rect 149242 220351 149298 220360
rect 147416 219694 147720 219722
rect 147416 219570 147444 219694
rect 147404 219564 147456 219570
rect 147404 219506 147456 219512
rect 147588 219564 147640 219570
rect 147588 219506 147640 219512
rect 147220 219292 147272 219298
rect 147220 219234 147272 219240
rect 147404 219292 147456 219298
rect 147404 219234 147456 219240
rect 147416 218754 147444 219234
rect 147404 218748 147456 218754
rect 147404 218690 147456 218696
rect 146760 218612 146812 218618
rect 146760 218554 146812 218560
rect 145070 217110 145144 217138
rect 145898 217246 146156 217274
rect 145070 216988 145098 217110
rect 145898 216988 145926 217246
rect 146772 217138 146800 218554
rect 147600 217274 147628 219506
rect 149244 218748 149296 218754
rect 149244 218690 149296 218696
rect 148416 218476 148468 218482
rect 148416 218418 148468 218424
rect 146726 217110 146800 217138
rect 147554 217246 147628 217274
rect 146726 216988 146754 217110
rect 147554 216988 147582 217246
rect 148428 217138 148456 218418
rect 149256 217138 149284 218690
rect 149900 218482 149928 226986
rect 150820 224233 150848 231676
rect 151386 231662 151584 231690
rect 150992 229764 151044 229770
rect 150992 229706 151044 229712
rect 151004 228857 151032 229706
rect 150990 228848 151046 228857
rect 150990 228783 151046 228792
rect 151358 228848 151414 228857
rect 151358 228783 151414 228792
rect 151372 228138 151400 228783
rect 151360 228132 151412 228138
rect 151360 228074 151412 228080
rect 151082 226400 151138 226409
rect 151082 226335 151138 226344
rect 150806 224224 150862 224233
rect 150806 224159 150862 224168
rect 150716 221468 150768 221474
rect 150716 221410 150768 221416
rect 150900 221468 150952 221474
rect 150900 221410 150952 221416
rect 150728 221241 150756 221410
rect 150714 221232 150770 221241
rect 150714 221167 150770 221176
rect 149888 218476 149940 218482
rect 149888 218418 149940 218424
rect 150070 218376 150126 218385
rect 150070 218311 150126 218320
rect 150084 217138 150112 218311
rect 150912 217274 150940 221410
rect 151096 218618 151124 226335
rect 151556 225729 151584 231662
rect 151726 230344 151782 230353
rect 151726 230279 151782 230288
rect 151740 227186 151768 230279
rect 151924 229537 151952 231676
rect 152108 231662 152490 231690
rect 151910 229528 151966 229537
rect 151910 229463 151966 229472
rect 151728 227180 151780 227186
rect 151728 227122 151780 227128
rect 151542 225720 151598 225729
rect 151542 225655 151598 225664
rect 151280 222686 151768 222714
rect 151280 222630 151308 222686
rect 151268 222624 151320 222630
rect 151268 222566 151320 222572
rect 151452 222624 151504 222630
rect 151452 222566 151504 222572
rect 151464 219434 151492 222566
rect 151740 222442 151768 222686
rect 151910 222592 151966 222601
rect 151910 222527 151966 222536
rect 151740 222414 151814 222442
rect 151786 222358 151814 222414
rect 151774 222352 151826 222358
rect 151774 222294 151826 222300
rect 151924 221746 151952 222527
rect 151912 221740 151964 221746
rect 151912 221682 151964 221688
rect 152108 220794 152136 231662
rect 153028 231305 153056 231676
rect 153304 231662 153594 231690
rect 153014 231296 153070 231305
rect 153014 231231 153070 231240
rect 153304 230353 153332 231662
rect 153290 230344 153346 230353
rect 153290 230279 153346 230288
rect 154132 229770 154160 231676
rect 154684 229922 154712 231676
rect 154684 229894 154804 229922
rect 154120 229764 154172 229770
rect 154120 229706 154172 229712
rect 154580 229764 154632 229770
rect 154580 229706 154632 229712
rect 154118 229528 154174 229537
rect 153016 229492 153068 229498
rect 152568 229452 153016 229480
rect 152568 229362 152596 229452
rect 154118 229463 154174 229472
rect 153016 229434 153068 229440
rect 152556 229356 152608 229362
rect 152556 229298 152608 229304
rect 152464 229084 152516 229090
rect 152464 229026 152516 229032
rect 152924 229084 152976 229090
rect 152924 229026 152976 229032
rect 152476 228274 152504 229026
rect 152936 228857 152964 229026
rect 152922 228848 152978 228857
rect 152922 228783 152978 228792
rect 152464 228268 152516 228274
rect 152464 228210 152516 228216
rect 152278 224224 152334 224233
rect 152278 224159 152334 224168
rect 152292 223038 152320 224159
rect 152280 223032 152332 223038
rect 152280 222974 152332 222980
rect 152464 223032 152516 223038
rect 152464 222974 152516 222980
rect 152280 221740 152332 221746
rect 152280 221682 152332 221688
rect 152292 221241 152320 221682
rect 152278 221232 152334 221241
rect 152278 221167 152334 221176
rect 152096 220788 152148 220794
rect 152096 220730 152148 220736
rect 151464 219406 151768 219434
rect 151084 218612 151136 218618
rect 151084 218554 151136 218560
rect 151452 218612 151504 218618
rect 151452 218554 151504 218560
rect 151464 218113 151492 218554
rect 151450 218104 151506 218113
rect 151450 218039 151506 218048
rect 151740 217274 151768 219406
rect 151912 218748 151964 218754
rect 151912 218690 151964 218696
rect 151924 218385 151952 218690
rect 152476 218482 152504 222974
rect 153934 220416 153990 220425
rect 153934 220351 153990 220360
rect 153948 220250 153976 220351
rect 153936 220244 153988 220250
rect 153936 220186 153988 220192
rect 152464 218476 152516 218482
rect 152464 218418 152516 218424
rect 151910 218376 151966 218385
rect 154132 218346 154160 229463
rect 154592 227458 154620 229706
rect 154776 228041 154804 229894
rect 154762 228032 154818 228041
rect 154762 227967 154818 227976
rect 154580 227452 154632 227458
rect 154580 227394 154632 227400
rect 155236 222873 155264 231676
rect 155512 231662 155802 231690
rect 155512 227769 155540 231662
rect 156340 230314 156368 231676
rect 156524 231662 156906 231690
rect 156328 230308 156380 230314
rect 156328 230250 156380 230256
rect 156328 229356 156380 229362
rect 156328 229298 156380 229304
rect 156340 229129 156368 229298
rect 156326 229120 156382 229129
rect 156326 229055 156382 229064
rect 156524 228290 156552 231662
rect 157352 230058 157380 231882
rect 157458 231662 157932 231690
rect 157614 231160 157670 231169
rect 157614 231095 157670 231104
rect 157628 231010 157656 231095
rect 157306 230042 157380 230058
rect 157294 230036 157380 230042
rect 157346 230030 157380 230036
rect 157536 230982 157656 231010
rect 157294 229978 157346 229984
rect 157536 229786 157564 230982
rect 157904 229922 157932 231662
rect 157352 229758 157564 229786
rect 157812 229894 157932 229922
rect 156880 229356 156932 229362
rect 156880 229298 156932 229304
rect 156064 228262 156552 228290
rect 155498 227760 155554 227769
rect 155498 227695 155554 227704
rect 155684 227452 155736 227458
rect 155684 227394 155736 227400
rect 155222 222864 155278 222873
rect 155222 222799 155278 222808
rect 154304 220108 154356 220114
rect 154304 220050 154356 220056
rect 151910 218311 151966 218320
rect 153384 218340 153436 218346
rect 153384 218282 153436 218288
rect 154120 218340 154172 218346
rect 154120 218282 154172 218288
rect 152554 218240 152610 218249
rect 152554 218175 152610 218184
rect 148382 217110 148456 217138
rect 149210 217110 149284 217138
rect 150038 217110 150112 217138
rect 150866 217246 150940 217274
rect 151694 217246 151768 217274
rect 148382 216988 148410 217110
rect 149210 216988 149238 217110
rect 150038 216988 150066 217110
rect 150866 216988 150894 217246
rect 151694 216988 151722 217246
rect 152568 217138 152596 218175
rect 153396 217138 153424 218282
rect 154316 217274 154344 220050
rect 155696 219434 155724 227394
rect 155868 220788 155920 220794
rect 155868 220730 155920 220736
rect 155696 219406 155816 219434
rect 155040 218340 155092 218346
rect 155040 218282 155092 218288
rect 152522 217110 152596 217138
rect 153350 217110 153424 217138
rect 154178 217246 154344 217274
rect 152522 216988 152550 217110
rect 153350 216988 153378 217110
rect 154178 216988 154206 217246
rect 155052 217138 155080 218282
rect 155788 217274 155816 219406
rect 155880 218362 155908 220730
rect 156064 220250 156092 228262
rect 156696 227180 156748 227186
rect 156696 227122 156748 227128
rect 156512 226160 156564 226166
rect 156512 226102 156564 226108
rect 156524 226001 156552 226102
rect 156510 225992 156566 226001
rect 156510 225927 156566 225936
rect 156708 224262 156736 227122
rect 156892 226409 156920 229298
rect 157352 229242 157380 229758
rect 157614 229528 157670 229537
rect 157614 229463 157670 229472
rect 157306 229226 157380 229242
rect 157628 229226 157656 229463
rect 157294 229220 157380 229226
rect 157346 229214 157380 229220
rect 157616 229220 157668 229226
rect 157294 229162 157346 229168
rect 157616 229162 157668 229168
rect 156878 226400 156934 226409
rect 156878 226335 156934 226344
rect 157294 226296 157346 226302
rect 156984 226244 157294 226250
rect 156984 226238 157346 226244
rect 156984 226222 157334 226238
rect 156984 225622 157012 226222
rect 157430 225992 157486 226001
rect 157430 225927 157486 225936
rect 156972 225616 157024 225622
rect 156972 225558 157024 225564
rect 157156 225616 157208 225622
rect 157156 225558 157208 225564
rect 157292 225618 157348 225627
rect 157444 225622 157472 225927
rect 157168 225457 157196 225558
rect 157292 225553 157348 225562
rect 157432 225616 157484 225622
rect 157432 225558 157484 225564
rect 157154 225448 157210 225457
rect 157154 225383 157210 225392
rect 157812 224954 157840 229894
rect 157996 229770 158024 231676
rect 157984 229764 158036 229770
rect 157984 229706 158036 229712
rect 158168 229764 158220 229770
rect 158168 229706 158220 229712
rect 158180 229129 158208 229706
rect 158166 229120 158222 229129
rect 158166 229055 158222 229064
rect 157444 224926 157840 224954
rect 156696 224256 156748 224262
rect 156696 224198 156748 224204
rect 156972 224256 157024 224262
rect 156972 224198 157024 224204
rect 156420 223032 156472 223038
rect 156420 222974 156472 222980
rect 156432 222873 156460 222974
rect 156788 222896 156840 222902
rect 156418 222864 156474 222873
rect 156788 222838 156840 222844
rect 156418 222799 156474 222808
rect 156800 222714 156828 222838
rect 156432 222686 156828 222714
rect 156432 222630 156460 222686
rect 156420 222624 156472 222630
rect 156420 222566 156472 222572
rect 156604 222624 156656 222630
rect 156604 222566 156656 222572
rect 156616 222358 156644 222566
rect 156604 222352 156656 222358
rect 156604 222294 156656 222300
rect 156604 222012 156656 222018
rect 156604 221954 156656 221960
rect 156788 222012 156840 222018
rect 156788 221954 156840 221960
rect 156616 221746 156644 221954
rect 156420 221740 156472 221746
rect 156420 221682 156472 221688
rect 156604 221740 156656 221746
rect 156604 221682 156656 221688
rect 156432 221626 156460 221682
rect 156800 221626 156828 221954
rect 156432 221598 156828 221626
rect 156234 220416 156290 220425
rect 156234 220351 156290 220360
rect 156248 220250 156276 220351
rect 156052 220244 156104 220250
rect 156052 220186 156104 220192
rect 156236 220244 156288 220250
rect 156236 220186 156288 220192
rect 156984 219434 157012 224198
rect 157444 223281 157472 224926
rect 158548 224262 158576 231676
rect 158916 231662 159114 231690
rect 159284 231662 159666 231690
rect 158536 224256 158588 224262
rect 158536 224198 158588 224204
rect 158720 224256 158772 224262
rect 158720 224198 158772 224204
rect 158732 224074 158760 224198
rect 158364 224046 158760 224074
rect 157430 223272 157486 223281
rect 157430 223207 157486 223216
rect 156432 219406 157012 219434
rect 156432 218890 156460 219406
rect 156602 219192 156658 219201
rect 156602 219127 156658 219136
rect 156420 218884 156472 218890
rect 156420 218826 156472 218832
rect 156616 218657 156644 219127
rect 157524 218884 157576 218890
rect 157524 218826 157576 218832
rect 156602 218648 156658 218657
rect 156602 218583 156658 218592
rect 156696 218476 156748 218482
rect 156696 218418 156748 218424
rect 155880 218346 156000 218362
rect 155880 218340 156012 218346
rect 155880 218334 155960 218340
rect 155960 218282 156012 218288
rect 155788 217246 155862 217274
rect 155006 217110 155080 217138
rect 155006 216988 155034 217110
rect 155834 216988 155862 217246
rect 156708 217138 156736 218418
rect 157536 217138 157564 218826
rect 158364 217274 158392 224046
rect 158916 222442 158944 231662
rect 159284 224233 159312 231662
rect 159822 230752 159878 230761
rect 159822 230687 159878 230696
rect 159546 230616 159602 230625
rect 159546 230551 159602 230560
rect 159560 230382 159588 230551
rect 159548 230376 159600 230382
rect 159548 230318 159600 230324
rect 159836 228138 159864 230687
rect 159824 228132 159876 228138
rect 159824 228074 159876 228080
rect 160008 228132 160060 228138
rect 160008 228074 160060 228080
rect 159270 224224 159326 224233
rect 159270 224159 159326 224168
rect 158824 222414 158944 222442
rect 158824 220153 158852 222414
rect 158996 222352 159048 222358
rect 158996 222294 159048 222300
rect 158810 220144 158866 220153
rect 158810 220079 158866 220088
rect 159008 218346 159036 222294
rect 160020 218346 160048 228074
rect 160204 227322 160232 231676
rect 160756 229770 160784 231676
rect 160940 231662 161322 231690
rect 160744 229764 160796 229770
rect 160744 229706 160796 229712
rect 160940 228290 160968 231662
rect 161112 229764 161164 229770
rect 161112 229706 161164 229712
rect 160664 228262 160968 228290
rect 160192 227316 160244 227322
rect 160192 227258 160244 227264
rect 160466 223408 160522 223417
rect 160466 223343 160522 223352
rect 160480 223174 160508 223343
rect 160468 223168 160520 223174
rect 160468 223110 160520 223116
rect 160664 220250 160692 228262
rect 161124 224890 161152 229706
rect 160940 224862 161152 224890
rect 160940 222601 160968 224862
rect 161860 223854 161888 231676
rect 162320 231662 162426 231690
rect 162978 231662 163268 231690
rect 162124 230036 162176 230042
rect 162124 229978 162176 229984
rect 162136 229498 162164 229978
rect 162124 229492 162176 229498
rect 162124 229434 162176 229440
rect 162320 225593 162348 231662
rect 162306 225584 162362 225593
rect 162306 225519 162362 225528
rect 162674 225448 162730 225457
rect 162674 225383 162730 225392
rect 161848 223848 161900 223854
rect 161848 223790 161900 223796
rect 162492 223848 162544 223854
rect 162492 223790 162544 223796
rect 161480 223032 161532 223038
rect 161308 222980 161480 222986
rect 161308 222974 161532 222980
rect 161308 222958 161520 222974
rect 161110 222864 161166 222873
rect 161110 222799 161166 222808
rect 160926 222592 160982 222601
rect 160926 222527 160982 222536
rect 161124 222170 161152 222799
rect 161308 222358 161336 222958
rect 161570 222592 161626 222601
rect 161570 222527 161626 222536
rect 161296 222352 161348 222358
rect 161296 222294 161348 222300
rect 161434 222352 161486 222358
rect 161434 222294 161486 222300
rect 161446 222170 161474 222294
rect 161124 222142 161474 222170
rect 161584 222154 161612 222527
rect 161572 222148 161624 222154
rect 161572 222090 161624 222096
rect 161756 222148 161808 222154
rect 161756 222090 161808 222096
rect 161768 222034 161796 222090
rect 161446 222006 161796 222034
rect 161446 221882 161474 222006
rect 161434 221876 161486 221882
rect 161434 221818 161486 221824
rect 161572 221876 161624 221882
rect 161572 221818 161624 221824
rect 161584 221762 161612 221818
rect 161446 221734 161612 221762
rect 161446 221610 161474 221734
rect 161434 221604 161486 221610
rect 161434 221546 161486 221552
rect 161572 221604 161624 221610
rect 161572 221546 161624 221552
rect 161584 221241 161612 221546
rect 161386 221232 161442 221241
rect 161386 221167 161442 221176
rect 161570 221232 161626 221241
rect 161570 221167 161626 221176
rect 160652 220244 160704 220250
rect 160652 220186 160704 220192
rect 160836 220244 160888 220250
rect 160836 220186 160888 220192
rect 158996 218340 159048 218346
rect 158996 218282 159048 218288
rect 159180 218340 159232 218346
rect 159180 218282 159232 218288
rect 160008 218340 160060 218346
rect 160008 218282 160060 218288
rect 160192 218340 160244 218346
rect 160192 218282 160244 218288
rect 156662 217110 156736 217138
rect 157490 217110 157564 217138
rect 158318 217246 158392 217274
rect 156662 216988 156690 217110
rect 157490 216988 157518 217110
rect 158318 216988 158346 217246
rect 159192 217138 159220 218282
rect 160204 218226 160232 218282
rect 160020 218198 160232 218226
rect 160020 217274 160048 218198
rect 160848 217274 160876 220186
rect 161400 218890 161428 221167
rect 161756 219020 161808 219026
rect 161756 218962 161808 218968
rect 161388 218884 161440 218890
rect 161388 218826 161440 218832
rect 161768 218521 161796 218962
rect 161294 218512 161350 218521
rect 161754 218512 161810 218521
rect 161294 218447 161296 218456
rect 161348 218447 161350 218456
rect 161480 218476 161532 218482
rect 161296 218418 161348 218424
rect 161754 218447 161810 218456
rect 161480 218418 161532 218424
rect 161492 218362 161520 218418
rect 161308 218334 161520 218362
rect 161308 218249 161336 218334
rect 161294 218240 161350 218249
rect 161294 218175 161350 218184
rect 161478 218240 161534 218249
rect 161478 218175 161480 218184
rect 161532 218175 161534 218184
rect 161480 218146 161532 218152
rect 162504 218142 162532 223790
rect 161664 218136 161716 218142
rect 161664 218078 161716 218084
rect 162492 218136 162544 218142
rect 162492 218078 162544 218084
rect 159146 217110 159220 217138
rect 159974 217246 160048 217274
rect 160802 217246 160876 217274
rect 159146 216988 159174 217110
rect 159974 216988 160002 217246
rect 160802 216988 160830 217246
rect 161676 217138 161704 218078
rect 162688 217274 162716 225383
rect 163240 219201 163268 231662
rect 163516 229770 163544 231676
rect 163792 231662 164082 231690
rect 164436 231662 164634 231690
rect 163504 229764 163556 229770
rect 163504 229706 163556 229712
rect 163596 229492 163648 229498
rect 163596 229434 163648 229440
rect 163608 221746 163636 229434
rect 163792 223417 163820 231662
rect 163964 229764 164016 229770
rect 163964 229706 164016 229712
rect 163976 227186 164004 229706
rect 163964 227180 164016 227186
rect 163964 227122 164016 227128
rect 163778 223408 163834 223417
rect 163778 223343 163834 223352
rect 164436 221882 164464 231662
rect 165724 229498 165752 231676
rect 166000 231662 166290 231690
rect 166552 231662 166842 231690
rect 165712 229492 165764 229498
rect 165712 229434 165764 229440
rect 164790 228984 164846 228993
rect 164790 228919 164846 228928
rect 164606 222592 164662 222601
rect 164606 222527 164662 222536
rect 164620 221882 164648 222527
rect 164424 221876 164476 221882
rect 164424 221818 164476 221824
rect 164608 221876 164660 221882
rect 164608 221818 164660 221824
rect 163596 221740 163648 221746
rect 163596 221682 163648 221688
rect 164056 221740 164108 221746
rect 164056 221682 164108 221688
rect 163226 219192 163282 219201
rect 163226 219127 163282 219136
rect 163320 218204 163372 218210
rect 163320 218146 163372 218152
rect 161630 217110 161704 217138
rect 162458 217246 162716 217274
rect 161630 216988 161658 217110
rect 162458 216988 162486 217246
rect 163332 217138 163360 218146
rect 164068 217274 164096 221682
rect 164422 220008 164478 220017
rect 164422 219943 164478 219952
rect 164436 219162 164464 219943
rect 164424 219156 164476 219162
rect 164424 219098 164476 219104
rect 164608 219156 164660 219162
rect 164608 219098 164660 219104
rect 164620 218210 164648 219098
rect 164804 218346 164832 228919
rect 166000 224670 166028 231662
rect 166354 229256 166410 229265
rect 166354 229191 166410 229200
rect 166368 225758 166396 229191
rect 166356 225752 166408 225758
rect 166356 225694 166408 225700
rect 165988 224664 166040 224670
rect 165988 224606 166040 224612
rect 166264 224664 166316 224670
rect 166264 224606 166316 224612
rect 164792 218340 164844 218346
rect 164792 218282 164844 218288
rect 166276 218278 166304 224606
rect 166552 224398 166580 231662
rect 167184 230376 167236 230382
rect 167182 230344 167184 230353
rect 167236 230344 167238 230353
rect 167182 230279 167238 230288
rect 167000 229492 167052 229498
rect 167000 229434 167052 229440
rect 167012 228993 167040 229434
rect 166998 228984 167054 228993
rect 166998 228919 167054 228928
rect 167182 228848 167238 228857
rect 167012 228806 167182 228834
rect 167012 228562 167040 228806
rect 167182 228783 167238 228792
rect 166920 228546 167040 228562
rect 166908 228540 167040 228546
rect 166960 228534 167040 228540
rect 166908 228482 166960 228488
rect 166724 227452 166776 227458
rect 166724 227394 166776 227400
rect 166736 224954 166764 227394
rect 166736 224926 166856 224954
rect 166540 224392 166592 224398
rect 166540 224334 166592 224340
rect 166632 218340 166684 218346
rect 166632 218282 166684 218288
rect 164976 218272 165028 218278
rect 164976 218214 165028 218220
rect 166264 218272 166316 218278
rect 166264 218214 166316 218220
rect 164608 218204 164660 218210
rect 164608 218146 164660 218152
rect 164068 217246 164142 217274
rect 163286 217110 163360 217138
rect 163286 216988 163314 217110
rect 164114 216988 164142 217246
rect 164988 217138 165016 218214
rect 165804 218136 165856 218142
rect 165804 218078 165856 218084
rect 165816 217138 165844 218078
rect 166644 217138 166672 218282
rect 166828 218142 166856 224926
rect 167380 218890 167408 231676
rect 167656 231662 167946 231690
rect 168392 231662 168498 231690
rect 167656 222154 167684 231662
rect 167826 230752 167882 230761
rect 167826 230687 167882 230696
rect 167840 230382 167868 230687
rect 167828 230376 167880 230382
rect 167828 230318 167880 230324
rect 167828 228676 167880 228682
rect 167828 228618 167880 228624
rect 167840 227458 167868 228618
rect 167828 227452 167880 227458
rect 167828 227394 167880 227400
rect 168196 224392 168248 224398
rect 168196 224334 168248 224340
rect 167644 222148 167696 222154
rect 167644 222090 167696 222096
rect 167368 218884 167420 218890
rect 167368 218826 167420 218832
rect 167552 218884 167604 218890
rect 167552 218826 167604 218832
rect 167564 218249 167592 218826
rect 167550 218240 167606 218249
rect 167550 218175 167606 218184
rect 166816 218136 166868 218142
rect 166816 218078 166868 218084
rect 167276 217864 167328 217870
rect 167276 217806 167328 217812
rect 167460 217864 167512 217870
rect 167460 217806 167512 217812
rect 167288 217190 167316 217806
rect 164942 217110 165016 217138
rect 165770 217110 165844 217138
rect 166598 217110 166672 217138
rect 167276 217184 167328 217190
rect 167472 217138 167500 217806
rect 167276 217126 167328 217132
rect 167426 217110 167500 217138
rect 168208 217138 168236 224334
rect 168392 224126 168420 231662
rect 169036 228546 169064 231676
rect 169312 231662 169602 231690
rect 169312 231169 169340 231662
rect 169298 231160 169354 231169
rect 169298 231095 169354 231104
rect 169206 229528 169262 229537
rect 169206 229463 169262 229472
rect 169024 228540 169076 228546
rect 169024 228482 169076 228488
rect 169024 225616 169076 225622
rect 169024 225558 169076 225564
rect 169036 225457 169064 225558
rect 169022 225448 169078 225457
rect 169022 225383 169078 225392
rect 168380 224120 168432 224126
rect 168380 224062 168432 224068
rect 168564 224120 168616 224126
rect 168564 224062 168616 224068
rect 168576 220017 168604 224062
rect 168562 220008 168618 220017
rect 168562 219943 168618 219952
rect 169220 219434 169248 229463
rect 169208 219428 169260 219434
rect 169208 219370 169260 219376
rect 169944 219428 169996 219434
rect 169944 219370 169996 219376
rect 169116 218204 169168 218210
rect 169116 218146 169168 218152
rect 169128 217138 169156 218146
rect 169956 217138 169984 219370
rect 170140 218890 170168 231676
rect 170416 231662 170706 231690
rect 170416 221882 170444 231662
rect 171244 224534 171272 231676
rect 171428 231662 171810 231690
rect 171232 224528 171284 224534
rect 171232 224470 171284 224476
rect 171428 223530 171456 231662
rect 171612 230438 172008 230466
rect 171612 230382 171640 230438
rect 171600 230376 171652 230382
rect 171600 230318 171652 230324
rect 171784 230308 171836 230314
rect 171784 230250 171836 230256
rect 171796 230042 171824 230250
rect 171980 230042 172008 230438
rect 171784 230036 171836 230042
rect 171784 229978 171836 229984
rect 171968 230036 172020 230042
rect 171968 229978 172020 229984
rect 171784 229764 171836 229770
rect 171784 229706 171836 229712
rect 171968 229764 172020 229770
rect 171968 229706 172020 229712
rect 171796 229498 171824 229706
rect 171600 229492 171652 229498
rect 171600 229434 171652 229440
rect 171784 229492 171836 229498
rect 171784 229434 171836 229440
rect 171612 229378 171640 229434
rect 171980 229378 172008 229706
rect 171612 229350 172008 229378
rect 172348 229265 172376 231676
rect 172334 229256 172390 229265
rect 172334 229191 172390 229200
rect 171968 228676 172020 228682
rect 171968 228618 172020 228624
rect 172428 228676 172480 228682
rect 172428 228618 172480 228624
rect 171600 228540 171652 228546
rect 171600 228482 171652 228488
rect 171612 228274 171640 228482
rect 171600 228268 171652 228274
rect 171600 228210 171652 228216
rect 171980 228138 172008 228618
rect 171968 228132 172020 228138
rect 171968 228074 172020 228080
rect 171600 224936 171652 224942
rect 171600 224878 171652 224884
rect 171612 224534 171640 224878
rect 171968 224800 172020 224806
rect 171968 224742 172020 224748
rect 171600 224528 171652 224534
rect 171600 224470 171652 224476
rect 171980 224398 172008 224742
rect 171968 224392 172020 224398
rect 171968 224334 172020 224340
rect 172242 224360 172298 224369
rect 172242 224295 172298 224304
rect 172256 224126 172284 224295
rect 172244 224120 172296 224126
rect 172244 224062 172296 224068
rect 171244 223502 171456 223530
rect 170404 221876 170456 221882
rect 170404 221818 170456 221824
rect 170772 221876 170824 221882
rect 170772 221818 170824 221824
rect 170128 218884 170180 218890
rect 170128 218826 170180 218832
rect 170784 217138 170812 221818
rect 171244 217190 171272 223502
rect 171428 223366 171824 223394
rect 171428 223310 171456 223366
rect 171416 223304 171468 223310
rect 171416 223246 171468 223252
rect 171600 223304 171652 223310
rect 171600 223246 171652 223252
rect 171612 223038 171640 223246
rect 171796 223038 171824 223366
rect 171600 223032 171652 223038
rect 171600 222974 171652 222980
rect 171784 223032 171836 223038
rect 171784 222974 171836 222980
rect 171600 222148 171652 222154
rect 171600 222090 171652 222096
rect 171612 221338 171640 222090
rect 171784 221604 171836 221610
rect 171784 221546 171836 221552
rect 171968 221604 172020 221610
rect 171968 221546 172020 221552
rect 171796 221338 171824 221546
rect 171600 221332 171652 221338
rect 171600 221274 171652 221280
rect 171784 221332 171836 221338
rect 171784 221274 171836 221280
rect 171600 219156 171652 219162
rect 171600 219098 171652 219104
rect 171612 218890 171640 219098
rect 171600 218884 171652 218890
rect 171600 218826 171652 218832
rect 171980 217274 172008 221546
rect 172440 217274 172468 228618
rect 172612 224120 172664 224126
rect 172612 224062 172664 224068
rect 172624 217870 172652 224062
rect 172900 220386 172928 231676
rect 173084 231662 173466 231690
rect 173084 223990 173112 231662
rect 174004 227594 174032 231676
rect 174556 230042 174584 231676
rect 174740 231662 175122 231690
rect 174544 230036 174596 230042
rect 174544 229978 174596 229984
rect 173992 227588 174044 227594
rect 173992 227530 174044 227536
rect 173440 224800 173492 224806
rect 173440 224742 173492 224748
rect 173256 224392 173308 224398
rect 173256 224334 173308 224340
rect 173072 223984 173124 223990
rect 173072 223926 173124 223932
rect 172888 220380 172940 220386
rect 172888 220322 172940 220328
rect 172612 217864 172664 217870
rect 172612 217806 172664 217812
rect 171566 217246 172008 217274
rect 172394 217246 172468 217274
rect 168208 217110 168282 217138
rect 164942 216988 164970 217110
rect 165770 216988 165798 217110
rect 166598 216988 166626 217110
rect 167426 216988 167454 217110
rect 168254 216988 168282 217110
rect 169082 217110 169156 217138
rect 169910 217110 169984 217138
rect 170738 217110 170812 217138
rect 171232 217184 171284 217190
rect 171232 217126 171284 217132
rect 169082 216988 169110 217110
rect 169910 216988 169938 217110
rect 170738 216988 170766 217110
rect 171566 216988 171594 217246
rect 172394 216988 172422 217246
rect 173268 217138 173296 224334
rect 173452 224126 173480 224742
rect 173440 224120 173492 224126
rect 173440 224062 173492 224068
rect 173728 222006 174124 222034
rect 173728 221882 173756 222006
rect 173716 221876 173768 221882
rect 173716 221818 173768 221824
rect 173900 221876 173952 221882
rect 173900 221818 173952 221824
rect 173912 221354 173940 221818
rect 174096 221762 174124 222006
rect 174740 221882 174768 231662
rect 174912 230036 174964 230042
rect 174912 229978 174964 229984
rect 174924 228857 174952 229978
rect 174910 228848 174966 228857
rect 174910 228783 174966 228792
rect 175096 224800 175148 224806
rect 175096 224742 175148 224748
rect 174728 221876 174780 221882
rect 174728 221818 174780 221824
rect 174912 221876 174964 221882
rect 174912 221818 174964 221824
rect 174924 221762 174952 221818
rect 174096 221734 174952 221762
rect 173728 221326 173940 221354
rect 173728 221202 173756 221326
rect 173716 221196 173768 221202
rect 173716 221138 173768 221144
rect 173900 221196 173952 221202
rect 173900 221138 173952 221144
rect 173912 218210 173940 221138
rect 174084 220380 174136 220386
rect 174084 220322 174136 220328
rect 173900 218204 173952 218210
rect 173900 218146 173952 218152
rect 174096 217138 174124 220322
rect 175108 217274 175136 224742
rect 175660 224534 175688 231676
rect 176016 230784 176068 230790
rect 176014 230752 176016 230761
rect 176068 230752 176070 230761
rect 176014 230687 176070 230696
rect 175648 224528 175700 224534
rect 175648 224470 175700 224476
rect 176016 224392 176068 224398
rect 176016 224334 176068 224340
rect 176028 224126 176056 224334
rect 176016 224120 176068 224126
rect 176016 224062 176068 224068
rect 176212 223038 176240 231676
rect 176672 231662 176778 231690
rect 177040 231662 177330 231690
rect 177592 231662 177882 231690
rect 178144 231662 178434 231690
rect 178604 231662 178986 231690
rect 179432 231662 179538 231690
rect 179708 231662 180090 231690
rect 176672 231010 176700 231662
rect 176626 230982 176700 231010
rect 176842 231024 176898 231033
rect 176476 230784 176528 230790
rect 176626 230772 176654 230982
rect 176842 230959 176898 230968
rect 176856 230874 176884 230959
rect 176764 230858 176884 230874
rect 176752 230852 176884 230858
rect 176804 230846 176884 230852
rect 176752 230794 176804 230800
rect 176626 230744 176700 230772
rect 176476 230726 176528 230732
rect 176488 230466 176516 230726
rect 176396 230438 176516 230466
rect 176396 230353 176424 230438
rect 176382 230344 176438 230353
rect 176382 230279 176438 230288
rect 176672 230194 176700 230744
rect 176396 230166 176700 230194
rect 176396 230042 176424 230166
rect 176384 230036 176436 230042
rect 176384 229978 176436 229984
rect 176568 230036 176620 230042
rect 176568 229978 176620 229984
rect 176580 229537 176608 229978
rect 176566 229528 176622 229537
rect 176566 229463 176622 229472
rect 176568 227452 176620 227458
rect 176568 227394 176620 227400
rect 176382 224360 176438 224369
rect 176382 224295 176438 224304
rect 176396 224126 176424 224295
rect 176384 224120 176436 224126
rect 176384 224062 176436 224068
rect 176200 223032 176252 223038
rect 176200 222974 176252 222980
rect 176580 218210 176608 227394
rect 177040 220522 177068 231662
rect 177592 230761 177620 231662
rect 177578 230752 177634 230761
rect 177578 230687 177634 230696
rect 177948 223032 178000 223038
rect 177948 222974 178000 222980
rect 177028 220516 177080 220522
rect 177028 220458 177080 220464
rect 175740 218204 175792 218210
rect 175740 218146 175792 218152
rect 176568 218204 176620 218210
rect 176568 218146 176620 218152
rect 173222 217110 173296 217138
rect 174050 217110 174124 217138
rect 174878 217246 175136 217274
rect 173222 216988 173250 217110
rect 174050 216988 174078 217110
rect 174878 216988 174906 217246
rect 175752 217138 175780 218146
rect 177960 218142 177988 222974
rect 178144 222018 178172 231662
rect 178314 231024 178370 231033
rect 178314 230959 178370 230968
rect 178328 230858 178356 230959
rect 178316 230852 178368 230858
rect 178316 230794 178368 230800
rect 178604 224954 178632 231662
rect 179050 228848 179106 228857
rect 179050 228783 179106 228792
rect 178328 224926 178632 224954
rect 178132 222012 178184 222018
rect 178132 221954 178184 221960
rect 178328 219434 178356 224926
rect 178144 219406 178356 219434
rect 178592 219428 178644 219434
rect 177396 218136 177448 218142
rect 177396 218078 177448 218084
rect 177948 218136 178000 218142
rect 177948 218078 178000 218084
rect 176568 217864 176620 217870
rect 176568 217806 176620 217812
rect 176580 217138 176608 217806
rect 177408 217138 177436 218078
rect 178144 217410 178172 219406
rect 178592 219370 178644 219376
rect 178604 219162 178632 219370
rect 178408 219156 178460 219162
rect 178408 219098 178460 219104
rect 178592 219156 178644 219162
rect 178592 219098 178644 219104
rect 178420 218346 178448 219098
rect 178592 219020 178644 219026
rect 178592 218962 178644 218968
rect 178408 218340 178460 218346
rect 178408 218282 178460 218288
rect 178052 217382 178172 217410
rect 178052 217326 178080 217382
rect 178040 217320 178092 217326
rect 178604 217274 178632 218962
rect 179064 217274 179092 228783
rect 179432 221066 179460 231662
rect 179708 222154 179736 231662
rect 180628 223310 180656 231676
rect 181194 231662 181484 231690
rect 181258 225992 181314 226001
rect 181258 225927 181314 225936
rect 181272 225758 181300 225927
rect 181260 225752 181312 225758
rect 181260 225694 181312 225700
rect 181456 224210 181484 231662
rect 181180 224182 181484 224210
rect 181548 231662 181746 231690
rect 180616 223304 180668 223310
rect 180616 223246 180668 223252
rect 179696 222148 179748 222154
rect 179696 222090 179748 222096
rect 180064 222012 180116 222018
rect 180064 221954 180116 221960
rect 179420 221060 179472 221066
rect 179420 221002 179472 221008
rect 179880 221060 179932 221066
rect 179880 221002 179932 221008
rect 179892 217274 179920 221002
rect 180076 219026 180104 221954
rect 180708 220516 180760 220522
rect 180708 220458 180760 220464
rect 180064 219020 180116 219026
rect 180064 218962 180116 218968
rect 180248 219020 180300 219026
rect 180248 218962 180300 218968
rect 180260 217870 180288 218962
rect 180248 217864 180300 217870
rect 180248 217806 180300 217812
rect 180720 217274 180748 220458
rect 181180 217462 181208 224182
rect 181548 220658 181576 231662
rect 181996 226024 182048 226030
rect 181994 225992 181996 226001
rect 182048 225992 182050 226001
rect 181994 225927 182050 225936
rect 182284 224942 182312 231676
rect 182836 229906 182864 231676
rect 183112 231662 183402 231690
rect 182824 229900 182876 229906
rect 182824 229842 182876 229848
rect 183112 228818 183140 231662
rect 183468 229900 183520 229906
rect 183468 229842 183520 229848
rect 183282 228848 183338 228857
rect 183100 228812 183152 228818
rect 183282 228783 183284 228792
rect 183100 228754 183152 228760
rect 183336 228783 183338 228792
rect 183284 228754 183336 228760
rect 182824 227452 182876 227458
rect 182824 227394 182876 227400
rect 182272 224936 182324 224942
rect 182272 224878 182324 224884
rect 181536 220652 181588 220658
rect 181536 220594 181588 220600
rect 182836 218074 182864 227394
rect 183480 221066 183508 229842
rect 183940 227730 183968 231676
rect 183928 227724 183980 227730
rect 183928 227666 183980 227672
rect 184204 227588 184256 227594
rect 184204 227530 184256 227536
rect 183468 221060 183520 221066
rect 183468 221002 183520 221008
rect 184020 219428 184072 219434
rect 184020 219370 184072 219376
rect 183190 219192 183246 219201
rect 183190 219127 183246 219136
rect 181536 218068 181588 218074
rect 181536 218010 181588 218016
rect 182824 218068 182876 218074
rect 182824 218010 182876 218016
rect 183008 218068 183060 218074
rect 183008 218010 183060 218016
rect 181168 217456 181220 217462
rect 181168 217398 181220 217404
rect 178040 217262 178092 217268
rect 175706 217110 175780 217138
rect 176534 217110 176608 217138
rect 177362 217110 177436 217138
rect 178190 217246 178632 217274
rect 179018 217246 179092 217274
rect 179846 217246 179920 217274
rect 180674 217246 180748 217274
rect 175706 216988 175734 217110
rect 176534 216988 176562 217110
rect 177362 216988 177390 217110
rect 178190 216988 178218 217246
rect 179018 216988 179046 217246
rect 179846 216988 179874 217246
rect 180674 216988 180702 217246
rect 181548 217138 181576 218010
rect 183020 217274 183048 218010
rect 181502 217110 181576 217138
rect 182330 217246 183048 217274
rect 181502 216988 181530 217110
rect 182330 216988 182358 217246
rect 183204 217138 183232 219127
rect 183558 218512 183614 218521
rect 183558 218447 183560 218456
rect 183612 218447 183614 218456
rect 183560 218418 183612 218424
rect 184032 217138 184060 219370
rect 184216 218929 184244 227530
rect 184492 223174 184520 231676
rect 185044 230858 185072 231676
rect 185228 231662 185610 231690
rect 185872 231662 186162 231690
rect 185032 230852 185084 230858
rect 185032 230794 185084 230800
rect 184846 229528 184902 229537
rect 184846 229463 184902 229472
rect 184860 226914 184888 229463
rect 184848 226908 184900 226914
rect 184848 226850 184900 226856
rect 185228 224954 185256 231662
rect 185872 229090 185900 231662
rect 186700 230654 186728 231676
rect 186688 230648 186740 230654
rect 186688 230590 186740 230596
rect 186134 230344 186190 230353
rect 186134 230279 186190 230288
rect 186148 230178 186176 230279
rect 186136 230172 186188 230178
rect 186136 230114 186188 230120
rect 186274 230172 186326 230178
rect 186274 230114 186326 230120
rect 186286 230058 186314 230114
rect 186148 230030 186314 230058
rect 186148 229537 186176 230030
rect 186134 229528 186190 229537
rect 186134 229463 186190 229472
rect 185860 229084 185912 229090
rect 185860 229026 185912 229032
rect 186134 225448 186190 225457
rect 186134 225383 186190 225392
rect 185136 224926 185256 224954
rect 185400 224936 185452 224942
rect 184480 223168 184532 223174
rect 184480 223110 184532 223116
rect 184848 223168 184900 223174
rect 184848 223110 184900 223116
rect 184664 222148 184716 222154
rect 184664 222090 184716 222096
rect 184676 219434 184704 222090
rect 184860 219434 184888 223110
rect 184676 219406 184796 219434
rect 184860 219428 184992 219434
rect 184860 219406 184940 219428
rect 184202 218920 184258 218929
rect 184202 218855 184258 218864
rect 184768 217274 184796 219406
rect 184940 219370 184992 219376
rect 185136 217938 185164 224926
rect 185400 224878 185452 224884
rect 185412 224534 185440 224878
rect 185584 224800 185636 224806
rect 185584 224742 185636 224748
rect 185596 224534 185624 224742
rect 185400 224528 185452 224534
rect 185400 224470 185452 224476
rect 185584 224528 185636 224534
rect 185584 224470 185636 224476
rect 185308 219428 185360 219434
rect 185308 219370 185360 219376
rect 185320 218521 185348 219370
rect 185768 219020 185820 219026
rect 185768 218962 185820 218968
rect 185952 219020 186004 219026
rect 185952 218962 186004 218968
rect 185306 218512 185362 218521
rect 185306 218447 185362 218456
rect 185780 218210 185808 218962
rect 185768 218204 185820 218210
rect 185768 218146 185820 218152
rect 185676 218068 185728 218074
rect 185676 218010 185728 218016
rect 185124 217932 185176 217938
rect 185124 217874 185176 217880
rect 184768 217246 184842 217274
rect 183158 217110 183232 217138
rect 183986 217110 184060 217138
rect 183158 216988 183186 217110
rect 183986 216988 184014 217110
rect 184814 216988 184842 217246
rect 185688 217138 185716 218010
rect 185964 217938 185992 218962
rect 186148 218074 186176 225383
rect 187252 223718 187280 231676
rect 187804 230178 187832 231676
rect 187988 231662 188370 231690
rect 188632 231662 188922 231690
rect 189184 231662 189474 231690
rect 189736 231662 190026 231690
rect 187792 230172 187844 230178
rect 187792 230114 187844 230120
rect 187240 223712 187292 223718
rect 187240 223654 187292 223660
rect 187332 223304 187384 223310
rect 187332 223246 187384 223252
rect 186504 221060 186556 221066
rect 186504 221002 186556 221008
rect 186136 218068 186188 218074
rect 186136 218010 186188 218016
rect 185952 217932 186004 217938
rect 185952 217874 186004 217880
rect 186516 217274 186544 221002
rect 187344 217274 187372 223246
rect 187988 220930 188016 231662
rect 188632 225758 188660 231662
rect 189184 230353 189212 231662
rect 189170 230344 189226 230353
rect 189170 230279 189226 230288
rect 188988 229084 189040 229090
rect 188988 229026 189040 229032
rect 188620 225752 188672 225758
rect 188620 225694 188672 225700
rect 188804 223712 188856 223718
rect 188804 223654 188856 223660
rect 187976 220924 188028 220930
rect 187976 220866 188028 220872
rect 188816 218074 188844 223654
rect 188160 218068 188212 218074
rect 188160 218010 188212 218016
rect 188804 218068 188856 218074
rect 188804 218010 188856 218016
rect 185642 217110 185716 217138
rect 186470 217246 186544 217274
rect 187298 217246 187372 217274
rect 185642 216988 185670 217110
rect 186470 216988 186498 217246
rect 187298 216988 187326 217246
rect 188172 217138 188200 218010
rect 189000 217274 189028 229026
rect 189736 228954 189764 231662
rect 189908 230172 189960 230178
rect 189908 230114 189960 230120
rect 189724 228948 189776 228954
rect 189724 228890 189776 228896
rect 189920 226642 189948 230114
rect 190472 230058 190500 231882
rect 190380 230042 190500 230058
rect 190368 230036 190500 230042
rect 190420 230030 190500 230036
rect 190368 229978 190420 229984
rect 189908 226636 189960 226642
rect 189908 226578 189960 226584
rect 189736 225950 190408 225978
rect 189736 219434 189764 225950
rect 190380 225894 190408 225950
rect 190184 225888 190236 225894
rect 190184 225830 190236 225836
rect 190368 225888 190420 225894
rect 190368 225830 190420 225836
rect 190196 225729 190224 225830
rect 190414 225752 190466 225758
rect 190182 225720 190238 225729
rect 190414 225694 190466 225700
rect 190182 225655 190238 225664
rect 190426 225570 190454 225694
rect 190288 225542 190454 225570
rect 190288 225457 190316 225542
rect 190274 225448 190330 225457
rect 190274 225383 190330 225392
rect 190564 223582 190592 231676
rect 190748 231662 191130 231690
rect 190748 225729 190776 231662
rect 191380 230172 191432 230178
rect 191380 230114 191432 230120
rect 191392 229094 191420 230114
rect 191300 229066 191420 229094
rect 190734 225720 190790 225729
rect 190734 225655 190790 225664
rect 190552 223576 190604 223582
rect 190552 223518 190604 223524
rect 190644 220652 190696 220658
rect 190644 220594 190696 220600
rect 189724 219428 189776 219434
rect 189724 219370 189776 219376
rect 189908 219428 189960 219434
rect 189908 219370 189960 219376
rect 189920 219201 189948 219370
rect 189906 219192 189962 219201
rect 189906 219127 189962 219136
rect 189816 218068 189868 218074
rect 189816 218010 189868 218016
rect 188126 217110 188200 217138
rect 188954 217246 189028 217274
rect 188126 216988 188154 217110
rect 188954 216988 188982 217246
rect 189828 217138 189856 218010
rect 190656 217274 190684 220594
rect 191300 219842 191328 229066
rect 191472 224936 191524 224942
rect 191472 224878 191524 224884
rect 191288 219836 191340 219842
rect 191288 219778 191340 219784
rect 191484 217274 191512 224878
rect 192220 219434 192248 231676
rect 192496 231662 192786 231690
rect 192496 219978 192524 231662
rect 193034 230344 193090 230353
rect 193034 230279 193090 230288
rect 192666 228848 192722 228857
rect 192666 228783 192722 228792
rect 192484 219972 192536 219978
rect 192484 219914 192536 219920
rect 192680 219434 192708 228783
rect 193048 228546 193076 230279
rect 193036 228540 193088 228546
rect 193036 228482 193088 228488
rect 193324 226030 193352 231676
rect 193312 226024 193364 226030
rect 193312 225966 193364 225972
rect 193680 226024 193732 226030
rect 193680 225966 193732 225972
rect 193036 219836 193088 219842
rect 193036 219778 193088 219784
rect 192128 219406 192248 219434
rect 192496 219406 192708 219434
rect 191930 218648 191986 218657
rect 191930 218583 191932 218592
rect 191984 218583 191986 218592
rect 191932 218554 191984 218560
rect 192128 217598 192156 219406
rect 192496 219298 192524 219406
rect 192484 219292 192536 219298
rect 192484 219234 192536 219240
rect 192300 218612 192352 218618
rect 192300 218554 192352 218560
rect 192116 217592 192168 217598
rect 192116 217534 192168 217540
rect 189782 217110 189856 217138
rect 190610 217246 190684 217274
rect 191438 217246 191512 217274
rect 189782 216988 189810 217110
rect 190610 216988 190638 217246
rect 191438 216988 191466 217246
rect 192312 217138 192340 218554
rect 193048 217274 193076 219778
rect 193692 219434 193720 225966
rect 193876 224126 193904 231676
rect 194428 230178 194456 231676
rect 194784 230648 194836 230654
rect 194784 230590 194836 230596
rect 194598 230344 194654 230353
rect 194598 230279 194654 230288
rect 194612 230178 194640 230279
rect 194416 230172 194468 230178
rect 194416 230114 194468 230120
rect 194600 230172 194652 230178
rect 194600 230114 194652 230120
rect 194796 229634 194824 230590
rect 194784 229628 194836 229634
rect 194784 229570 194836 229576
rect 194232 228948 194284 228954
rect 194232 228890 194284 228896
rect 193864 224120 193916 224126
rect 193864 224062 193916 224068
rect 194244 221066 194272 228890
rect 194784 224800 194836 224806
rect 194784 224742 194836 224748
rect 194796 224126 194824 224742
rect 194784 224120 194836 224126
rect 194784 224062 194836 224068
rect 194416 223576 194468 223582
rect 194416 223518 194468 223524
rect 194232 221060 194284 221066
rect 194232 221002 194284 221008
rect 193692 219406 193812 219434
rect 193784 218618 193812 219406
rect 194428 218618 194456 223518
rect 194980 222766 195008 231676
rect 195244 229628 195296 229634
rect 195244 229570 195296 229576
rect 195256 229226 195284 229570
rect 195244 229220 195296 229226
rect 195244 229162 195296 229168
rect 195244 229084 195296 229090
rect 195244 229026 195296 229032
rect 195256 228546 195284 229026
rect 195244 228540 195296 228546
rect 195244 228482 195296 228488
rect 195532 225486 195560 231676
rect 195992 231662 196098 231690
rect 195992 230654 196020 231662
rect 195980 230648 196032 230654
rect 195980 230590 196032 230596
rect 196636 230042 196664 231676
rect 196624 230036 196676 230042
rect 196624 229978 196676 229984
rect 196808 230036 196860 230042
rect 196808 229978 196860 229984
rect 196532 229220 196584 229226
rect 196532 229162 196584 229168
rect 195704 229084 195756 229090
rect 195704 229026 195756 229032
rect 195716 228857 195744 229026
rect 195702 228848 195758 228857
rect 195702 228783 195758 228792
rect 196544 227866 196572 229162
rect 196820 228954 196848 229978
rect 196808 228948 196860 228954
rect 196808 228890 196860 228896
rect 196532 227860 196584 227866
rect 196532 227802 196584 227808
rect 196624 227724 196676 227730
rect 196624 227666 196676 227672
rect 195704 226024 195756 226030
rect 195704 225966 195756 225972
rect 195888 226024 195940 226030
rect 195888 225966 195940 225972
rect 195716 225486 195744 225966
rect 195520 225480 195572 225486
rect 195520 225422 195572 225428
rect 195704 225480 195756 225486
rect 195704 225422 195756 225428
rect 195244 224800 195296 224806
rect 195244 224742 195296 224748
rect 195256 223718 195284 224742
rect 195244 223712 195296 223718
rect 195244 223654 195296 223660
rect 194968 222760 195020 222766
rect 194968 222702 195020 222708
rect 195612 221332 195664 221338
rect 195612 221274 195664 221280
rect 195624 221066 195652 221274
rect 195612 221060 195664 221066
rect 195612 221002 195664 221008
rect 195612 219292 195664 219298
rect 195612 219234 195664 219240
rect 193772 218612 193824 218618
rect 193772 218554 193824 218560
rect 193956 218612 194008 218618
rect 193956 218554 194008 218560
rect 194416 218612 194468 218618
rect 194416 218554 194468 218560
rect 194784 218612 194836 218618
rect 194784 218554 194836 218560
rect 193048 217246 193122 217274
rect 192266 217110 192340 217138
rect 192266 216988 192294 217110
rect 193094 216988 193122 217246
rect 193968 217138 193996 218554
rect 194796 217138 194824 218554
rect 195624 217138 195652 219234
rect 195900 218618 195928 225966
rect 196636 218657 196664 227666
rect 197188 223446 197216 231676
rect 197740 226166 197768 231676
rect 198292 227594 198320 231676
rect 198844 230178 198872 231676
rect 199028 231662 199410 231690
rect 199672 231662 199962 231690
rect 198832 230172 198884 230178
rect 198832 230114 198884 230120
rect 199028 229094 199056 231662
rect 199200 230172 199252 230178
rect 199200 230114 199252 230120
rect 199212 229094 199240 230114
rect 198648 229084 198700 229090
rect 199028 229066 199148 229094
rect 199212 229066 199332 229094
rect 198648 229026 198700 229032
rect 198280 227588 198332 227594
rect 198280 227530 198332 227536
rect 197728 226160 197780 226166
rect 197728 226102 197780 226108
rect 197912 226160 197964 226166
rect 197912 226102 197964 226108
rect 197924 225570 197952 226102
rect 197740 225542 197952 225570
rect 197740 225486 197768 225542
rect 197728 225480 197780 225486
rect 197728 225422 197780 225428
rect 197912 225480 197964 225486
rect 197912 225422 197964 225428
rect 197176 223440 197228 223446
rect 197176 223382 197228 223388
rect 197268 222760 197320 222766
rect 197268 222702 197320 222708
rect 196622 218648 196678 218657
rect 195888 218612 195940 218618
rect 195888 218554 195940 218560
rect 196256 218612 196308 218618
rect 196622 218583 196678 218592
rect 196256 218554 196308 218560
rect 196268 218346 196296 218554
rect 196256 218340 196308 218346
rect 196256 218282 196308 218288
rect 196440 218340 196492 218346
rect 196440 218282 196492 218288
rect 196452 217138 196480 218282
rect 197280 217138 197308 222702
rect 197728 221468 197780 221474
rect 197728 221410 197780 221416
rect 197740 221066 197768 221410
rect 197728 221060 197780 221066
rect 197728 221002 197780 221008
rect 197924 219298 197952 225422
rect 198660 224126 198688 229026
rect 198648 224120 198700 224126
rect 198648 224062 198700 224068
rect 198096 223440 198148 223446
rect 198096 223382 198148 223388
rect 197912 219292 197964 219298
rect 197912 219234 197964 219240
rect 198108 217138 198136 223382
rect 198924 219292 198976 219298
rect 198924 219234 198976 219240
rect 198936 217138 198964 219234
rect 199120 217734 199148 229066
rect 199304 226506 199332 229066
rect 199476 227588 199528 227594
rect 199476 227530 199528 227536
rect 199292 226500 199344 226506
rect 199292 226442 199344 226448
rect 199292 226024 199344 226030
rect 199290 225992 199292 226001
rect 199344 225992 199346 226001
rect 199290 225927 199346 225936
rect 199488 224954 199516 227530
rect 199672 225214 199700 231662
rect 200500 230314 200528 231676
rect 200672 230376 200724 230382
rect 200672 230318 200724 230324
rect 200488 230308 200540 230314
rect 200488 230250 200540 230256
rect 200488 229628 200540 229634
rect 200488 229570 200540 229576
rect 200118 229392 200174 229401
rect 200086 229362 200118 229378
rect 200074 229356 200118 229362
rect 200500 229362 200528 229570
rect 200684 229498 200712 230318
rect 200672 229492 200724 229498
rect 200672 229434 200724 229440
rect 200856 229492 200908 229498
rect 200856 229434 200908 229440
rect 200126 229327 200174 229336
rect 200488 229356 200540 229362
rect 200074 229298 200126 229304
rect 200488 229298 200540 229304
rect 200120 226160 200172 226166
rect 200040 226108 200120 226114
rect 200040 226102 200172 226108
rect 200040 226086 200160 226102
rect 199842 225992 199898 226001
rect 199842 225927 199898 225936
rect 199856 225214 199884 225927
rect 199660 225208 199712 225214
rect 199660 225150 199712 225156
rect 199844 225208 199896 225214
rect 199844 225150 199896 225156
rect 199488 224926 199700 224954
rect 199108 217728 199160 217734
rect 199108 217670 199160 217676
rect 199672 217274 199700 224926
rect 200040 219298 200068 226086
rect 200580 219972 200632 219978
rect 200580 219914 200632 219920
rect 200028 219292 200080 219298
rect 200028 219234 200080 219240
rect 200212 219292 200264 219298
rect 200212 219234 200264 219240
rect 200224 218906 200252 219234
rect 199856 218878 200252 218906
rect 199856 218618 199884 218878
rect 200212 218748 200264 218754
rect 200212 218690 200264 218696
rect 199844 218612 199896 218618
rect 199844 218554 199896 218560
rect 200224 218346 200252 218690
rect 200212 218340 200264 218346
rect 200212 218282 200264 218288
rect 199672 217246 199746 217274
rect 193922 217110 193996 217138
rect 194750 217110 194824 217138
rect 195578 217110 195652 217138
rect 196406 217110 196480 217138
rect 197234 217110 197308 217138
rect 198062 217110 198136 217138
rect 198890 217110 198964 217138
rect 193922 216988 193950 217110
rect 194750 216988 194778 217110
rect 195578 216988 195606 217110
rect 196406 216988 196434 217110
rect 197234 216988 197262 217110
rect 198062 216988 198090 217110
rect 198890 216988 198918 217110
rect 199718 216988 199746 217246
rect 200592 217138 200620 219914
rect 200868 219842 200896 229434
rect 201052 229226 201080 231676
rect 201224 229628 201276 229634
rect 201224 229570 201276 229576
rect 201040 229220 201092 229226
rect 201040 229162 201092 229168
rect 201236 229090 201264 229570
rect 201406 229392 201462 229401
rect 201406 229327 201462 229336
rect 201420 229226 201448 229327
rect 201408 229220 201460 229226
rect 201408 229162 201460 229168
rect 201224 229084 201276 229090
rect 201224 229026 201276 229032
rect 201040 227860 201092 227866
rect 201040 227802 201092 227808
rect 200856 219836 200908 219842
rect 200856 219778 200908 219784
rect 201052 219298 201080 227802
rect 201604 222494 201632 231676
rect 202156 226302 202184 231676
rect 202432 231662 202722 231690
rect 202432 228954 202460 231662
rect 203260 230178 203288 231676
rect 203536 231662 203826 231690
rect 203248 230172 203300 230178
rect 203248 230114 203300 230120
rect 202420 228948 202472 228954
rect 202420 228890 202472 228896
rect 202604 228948 202656 228954
rect 202604 228890 202656 228896
rect 202144 226296 202196 226302
rect 202144 226238 202196 226244
rect 202616 224954 202644 228890
rect 202248 224926 202644 224954
rect 201592 222488 201644 222494
rect 201592 222430 201644 222436
rect 201040 219292 201092 219298
rect 201040 219234 201092 219240
rect 201408 218340 201460 218346
rect 201408 218282 201460 218288
rect 201420 217138 201448 218282
rect 202248 217274 202276 224926
rect 203536 219706 203564 231662
rect 204168 230376 204220 230382
rect 204168 230318 204220 230324
rect 204180 228002 204208 230318
rect 204168 227996 204220 228002
rect 204168 227938 204220 227944
rect 204364 225078 204392 231676
rect 204916 230246 204944 231676
rect 205468 230382 205496 231676
rect 206020 230518 206048 231676
rect 206008 230512 206060 230518
rect 206008 230454 206060 230460
rect 205456 230376 205508 230382
rect 205456 230318 205508 230324
rect 205732 230376 205784 230382
rect 205732 230318 205784 230324
rect 204904 230240 204956 230246
rect 204904 230182 204956 230188
rect 205548 230172 205600 230178
rect 205548 230114 205600 230120
rect 205272 227996 205324 228002
rect 205272 227938 205324 227944
rect 204536 225888 204588 225894
rect 204536 225830 204588 225836
rect 204720 225888 204772 225894
rect 204720 225830 204772 225836
rect 204548 225078 204576 225830
rect 204732 225486 204760 225830
rect 204720 225480 204772 225486
rect 204720 225422 204772 225428
rect 204904 225480 204956 225486
rect 204904 225422 204956 225428
rect 204916 225214 204944 225422
rect 204904 225208 204956 225214
rect 204904 225150 204956 225156
rect 205088 225208 205140 225214
rect 205088 225150 205140 225156
rect 204352 225072 204404 225078
rect 204352 225014 204404 225020
rect 204536 225072 204588 225078
rect 204536 225014 204588 225020
rect 205100 224954 205128 225150
rect 205284 224954 205312 227938
rect 205560 227594 205588 230114
rect 205548 227588 205600 227594
rect 205548 227530 205600 227536
rect 205456 227044 205508 227050
rect 205456 226986 205508 226992
rect 205468 224954 205496 226986
rect 205744 226778 205772 230318
rect 205916 227588 205968 227594
rect 205916 227530 205968 227536
rect 205928 227050 205956 227530
rect 205916 227044 205968 227050
rect 205916 226986 205968 226992
rect 205732 226772 205784 226778
rect 205732 226714 205784 226720
rect 206100 226364 206152 226370
rect 206100 226306 206152 226312
rect 205008 224926 205128 224954
rect 205192 224926 205312 224954
rect 205376 224926 205496 224954
rect 205008 224777 205036 224926
rect 203890 224768 203946 224777
rect 203890 224703 203946 224712
rect 204994 224768 205050 224777
rect 204994 224703 205050 224712
rect 203524 219700 203576 219706
rect 203524 219642 203576 219648
rect 202878 218784 202934 218793
rect 202878 218719 202880 218728
rect 202932 218719 202934 218728
rect 202880 218690 202932 218696
rect 200546 217110 200620 217138
rect 201374 217110 201448 217138
rect 202202 217246 202276 217274
rect 203018 217252 203070 217258
rect 200546 216988 200574 217110
rect 201374 216988 201402 217110
rect 202202 216988 202230 217246
rect 203018 217194 203070 217200
rect 203030 216988 203058 217194
rect 203904 217138 203932 224703
rect 205192 219178 205220 224926
rect 205376 219706 205404 224926
rect 205640 222488 205692 222494
rect 205640 222430 205692 222436
rect 205364 219700 205416 219706
rect 205364 219642 205416 219648
rect 204732 219150 205220 219178
rect 204732 217274 204760 219150
rect 205500 218784 205556 218793
rect 205500 218719 205502 218728
rect 205554 218719 205556 218728
rect 205502 218690 205554 218696
rect 205652 218521 205680 222430
rect 205824 219700 205876 219706
rect 205824 219642 205876 219648
rect 205454 218512 205510 218521
rect 205454 218447 205456 218456
rect 205508 218447 205510 218456
rect 205638 218512 205694 218521
rect 205638 218447 205694 218456
rect 205456 218418 205508 218424
rect 205456 218340 205508 218346
rect 205456 218282 205508 218288
rect 205640 218340 205692 218346
rect 205640 218282 205692 218288
rect 205468 217938 205496 218282
rect 205652 217938 205680 218282
rect 205456 217932 205508 217938
rect 205456 217874 205508 217880
rect 205640 217932 205692 217938
rect 205640 217874 205692 217880
rect 205836 217274 205864 219642
rect 206112 218550 206140 226306
rect 206572 225350 206600 231676
rect 207124 227730 207152 231676
rect 207676 230382 207704 231676
rect 207860 231662 208242 231690
rect 207664 230376 207716 230382
rect 207664 230318 207716 230324
rect 207112 227724 207164 227730
rect 207112 227666 207164 227672
rect 206560 225344 206612 225350
rect 206560 225286 206612 225292
rect 207204 219836 207256 219842
rect 207204 219778 207256 219784
rect 206100 218544 206152 218550
rect 206100 218486 206152 218492
rect 206376 218476 206428 218482
rect 206376 218418 206428 218424
rect 203858 217110 203932 217138
rect 204686 217246 204760 217274
rect 205514 217246 205864 217274
rect 203858 216988 203886 217110
rect 204686 216988 204714 217246
rect 205514 216988 205542 217246
rect 206388 217138 206416 218418
rect 207216 217138 207244 219778
rect 207860 219570 207888 231662
rect 208032 230308 208084 230314
rect 208032 230250 208084 230256
rect 208044 229498 208072 230250
rect 208032 229492 208084 229498
rect 208032 229434 208084 229440
rect 208216 229492 208268 229498
rect 208216 229434 208268 229440
rect 208228 229226 208256 229434
rect 208216 229220 208268 229226
rect 208216 229162 208268 229168
rect 208400 229220 208452 229226
rect 208400 229162 208452 229168
rect 208412 228274 208440 229162
rect 208400 228268 208452 228274
rect 208400 228210 208452 228216
rect 208032 225344 208084 225350
rect 208032 225286 208084 225292
rect 207848 219564 207900 219570
rect 207848 219506 207900 219512
rect 207848 218612 207900 218618
rect 207848 218554 207900 218560
rect 207860 217258 207888 218554
rect 208044 217274 208072 225286
rect 208780 222630 208808 231676
rect 209332 229498 209360 231676
rect 209320 229492 209372 229498
rect 209320 229434 209372 229440
rect 209596 227724 209648 227730
rect 209596 227666 209648 227672
rect 208768 222624 208820 222630
rect 208768 222566 208820 222572
rect 209608 219298 209636 227666
rect 209884 222358 209912 231676
rect 210068 231662 210450 231690
rect 210712 231662 211002 231690
rect 209872 222352 209924 222358
rect 209872 222294 209924 222300
rect 210068 221338 210096 231662
rect 210712 226914 210740 231662
rect 211160 229492 211212 229498
rect 211160 229434 211212 229440
rect 211172 228138 211200 229434
rect 211160 228132 211212 228138
rect 211160 228074 211212 228080
rect 210976 227044 211028 227050
rect 210976 226986 211028 226992
rect 210700 226908 210752 226914
rect 210700 226850 210752 226856
rect 210424 223984 210476 223990
rect 210424 223926 210476 223932
rect 210436 223718 210464 223926
rect 210424 223712 210476 223718
rect 210424 223654 210476 223660
rect 210332 222624 210384 222630
rect 210332 222566 210384 222572
rect 210056 221332 210108 221338
rect 210056 221274 210108 221280
rect 210344 219298 210372 222566
rect 210988 219298 211016 226986
rect 211540 226370 211568 231676
rect 211528 226364 211580 226370
rect 211528 226306 211580 226312
rect 212092 225078 212120 231676
rect 212264 229084 212316 229090
rect 212264 229026 212316 229032
rect 212080 225072 212132 225078
rect 212080 225014 212132 225020
rect 212276 224954 212304 229026
rect 212184 224926 212304 224954
rect 211344 221332 211396 221338
rect 211344 221274 211396 221280
rect 208860 219292 208912 219298
rect 208860 219234 208912 219240
rect 209596 219292 209648 219298
rect 209596 219234 209648 219240
rect 209780 219292 209832 219298
rect 209780 219234 209832 219240
rect 210332 219292 210384 219298
rect 210332 219234 210384 219240
rect 210516 219292 210568 219298
rect 210516 219234 210568 219240
rect 210976 219292 211028 219298
rect 210976 219234 211028 219240
rect 207848 217252 207900 217258
rect 207848 217194 207900 217200
rect 207998 217246 208072 217274
rect 206342 217110 206416 217138
rect 207170 217110 207244 217138
rect 206342 216988 206370 217110
rect 207170 216988 207198 217110
rect 207998 216988 208026 217246
rect 208872 217138 208900 219234
rect 209792 219042 209820 219234
rect 209148 219026 209820 219042
rect 209136 219020 209820 219026
rect 209188 219014 209820 219020
rect 209136 218962 209188 218968
rect 209688 218884 209740 218890
rect 209688 218826 209740 218832
rect 209700 217138 209728 218826
rect 210528 217138 210556 219234
rect 211356 217138 211384 221274
rect 212184 217274 212212 224926
rect 212644 220114 212672 231676
rect 213196 222902 213224 231676
rect 213552 230444 213604 230450
rect 213552 230386 213604 230392
rect 213184 222896 213236 222902
rect 213184 222838 213236 222844
rect 213368 221060 213420 221066
rect 213368 221002 213420 221008
rect 212632 220108 212684 220114
rect 212632 220050 212684 220056
rect 213000 219292 213052 219298
rect 213000 219234 213052 219240
rect 208826 217110 208900 217138
rect 209654 217110 209728 217138
rect 210482 217110 210556 217138
rect 211310 217110 211384 217138
rect 212138 217246 212212 217274
rect 208826 216988 208854 217110
rect 209654 216988 209682 217110
rect 210482 216988 210510 217110
rect 211310 216988 211338 217110
rect 212138 216988 212166 217246
rect 213012 217138 213040 219234
rect 213380 217274 213408 221002
rect 213564 219298 213592 230386
rect 213748 229362 213776 231676
rect 213736 229356 213788 229362
rect 213736 229298 213788 229304
rect 213828 228676 213880 228682
rect 213828 228618 213880 228624
rect 213840 228274 213868 228618
rect 213828 228268 213880 228274
rect 213828 228210 213880 228216
rect 214300 227186 214328 231676
rect 214484 231662 214866 231690
rect 214288 227180 214340 227186
rect 214288 227122 214340 227128
rect 214484 226386 214512 231662
rect 214748 228540 214800 228546
rect 214748 228482 214800 228488
rect 214760 228002 214788 228482
rect 214748 227996 214800 228002
rect 214748 227938 214800 227944
rect 215208 227180 215260 227186
rect 215208 227122 215260 227128
rect 214024 226358 214512 226386
rect 214024 221474 214052 226358
rect 214380 226296 214432 226302
rect 214380 226238 214432 226244
rect 214196 225616 214248 225622
rect 214196 225558 214248 225564
rect 214208 225078 214236 225558
rect 214392 225214 214420 226238
rect 214564 225888 214616 225894
rect 214564 225830 214616 225836
rect 214576 225622 214604 225830
rect 214564 225616 214616 225622
rect 214564 225558 214616 225564
rect 214380 225208 214432 225214
rect 214380 225150 214432 225156
rect 214196 225072 214248 225078
rect 214196 225014 214248 225020
rect 214012 221468 214064 221474
rect 214012 221410 214064 221416
rect 213920 219700 213972 219706
rect 213920 219642 213972 219648
rect 213552 219292 213604 219298
rect 213552 219234 213604 219240
rect 213736 219292 213788 219298
rect 213736 219234 213788 219240
rect 213748 218754 213776 219234
rect 213932 219162 213960 219642
rect 215220 219162 215248 227122
rect 215404 220794 215432 231676
rect 215680 231662 215970 231690
rect 215680 222494 215708 231662
rect 216508 229226 216536 231676
rect 216876 231662 217074 231690
rect 216496 229220 216548 229226
rect 216496 229162 216548 229168
rect 216496 224120 216548 224126
rect 216496 224062 216548 224068
rect 215944 222896 215996 222902
rect 215944 222838 215996 222844
rect 215668 222488 215720 222494
rect 215668 222430 215720 222436
rect 215392 220788 215444 220794
rect 215392 220730 215444 220736
rect 213920 219156 213972 219162
rect 213920 219098 213972 219104
rect 214656 219156 214708 219162
rect 214656 219098 214708 219104
rect 215208 219156 215260 219162
rect 215208 219098 215260 219104
rect 214104 218884 214156 218890
rect 214104 218826 214156 218832
rect 213736 218748 213788 218754
rect 213736 218690 213788 218696
rect 214116 218482 214144 218826
rect 214104 218476 214156 218482
rect 214104 218418 214156 218424
rect 213380 217246 213822 217274
rect 212966 217110 213040 217138
rect 212966 216988 212994 217110
rect 213794 216988 213822 217246
rect 214668 217138 214696 219098
rect 215956 219026 215984 222838
rect 215944 219020 215996 219026
rect 215944 218962 215996 218968
rect 216312 218476 216364 218482
rect 216312 218418 216364 218424
rect 215206 218240 215262 218249
rect 215206 218175 215208 218184
rect 215260 218175 215262 218184
rect 215484 218204 215536 218210
rect 215208 218146 215260 218152
rect 215484 218146 215536 218152
rect 215496 217138 215524 218146
rect 216324 217138 216352 218418
rect 216508 218210 216536 224062
rect 216876 220250 216904 231662
rect 217324 225208 217376 225214
rect 217324 225150 217376 225156
rect 216864 220244 216916 220250
rect 216864 220186 216916 220192
rect 217140 220108 217192 220114
rect 217140 220050 217192 220056
rect 216496 218204 216548 218210
rect 216496 218146 216548 218152
rect 217152 217274 217180 220050
rect 217336 218249 217364 225150
rect 217612 224262 217640 231676
rect 218164 229770 218192 231676
rect 218152 229764 218204 229770
rect 218152 229706 218204 229712
rect 218716 225078 218744 231676
rect 218900 231662 219282 231690
rect 219452 231662 219834 231690
rect 218704 225072 218756 225078
rect 218704 225014 218756 225020
rect 217600 224256 217652 224262
rect 217600 224198 217652 224204
rect 218900 221746 218928 231662
rect 219452 229106 219480 231662
rect 219360 229078 219480 229106
rect 220372 229094 220400 231676
rect 220544 229764 220596 229770
rect 220544 229706 220596 229712
rect 220556 229094 220584 229706
rect 220924 229498 220952 231676
rect 221108 231662 221490 231690
rect 221660 231662 222042 231690
rect 220912 229492 220964 229498
rect 220912 229434 220964 229440
rect 220820 229356 220872 229362
rect 220820 229298 220872 229304
rect 219360 223990 219388 229078
rect 220280 229066 220400 229094
rect 220464 229066 220584 229094
rect 219348 223984 219400 223990
rect 219348 223926 219400 223932
rect 219348 223848 219400 223854
rect 219348 223790 219400 223796
rect 218888 221740 218940 221746
rect 218888 221682 218940 221688
rect 217968 219020 218020 219026
rect 217968 218962 218020 218968
rect 217322 218240 217378 218249
rect 217322 218175 217378 218184
rect 214622 217110 214696 217138
rect 215450 217110 215524 217138
rect 216278 217110 216352 217138
rect 217106 217246 217180 217274
rect 214622 216988 214650 217110
rect 215450 216988 215478 217110
rect 216278 216988 216306 217110
rect 217106 216988 217134 217246
rect 217980 217138 218008 218962
rect 219360 218210 219388 223790
rect 220280 222902 220308 229066
rect 220268 222896 220320 222902
rect 220268 222838 220320 222844
rect 220464 219434 220492 229066
rect 220832 228274 220860 229298
rect 220820 228268 220872 228274
rect 220820 228210 220872 228216
rect 221108 223718 221136 231662
rect 221660 224670 221688 231662
rect 222016 228268 222068 228274
rect 222016 228210 222068 228216
rect 221648 224664 221700 224670
rect 221648 224606 221700 224612
rect 221280 224528 221332 224534
rect 221280 224470 221332 224476
rect 221464 224528 221516 224534
rect 221464 224470 221516 224476
rect 221292 223990 221320 224470
rect 221280 223984 221332 223990
rect 221280 223926 221332 223932
rect 221096 223712 221148 223718
rect 221096 223654 221148 223660
rect 221280 222896 221332 222902
rect 221280 222838 221332 222844
rect 220636 221468 220688 221474
rect 220636 221410 220688 221416
rect 220648 219434 220676 221410
rect 220372 219406 220492 219434
rect 220556 219406 220676 219434
rect 220372 218210 220400 219406
rect 218796 218204 218848 218210
rect 218796 218146 218848 218152
rect 219348 218204 219400 218210
rect 219348 218146 219400 218152
rect 219624 218204 219676 218210
rect 219624 218146 219676 218152
rect 220360 218204 220412 218210
rect 220360 218146 220412 218152
rect 218808 217138 218836 218146
rect 219636 217138 219664 218146
rect 220556 217274 220584 219406
rect 221292 217274 221320 222838
rect 221476 219026 221504 224470
rect 221464 219020 221516 219026
rect 221464 218962 221516 218968
rect 217934 217110 218008 217138
rect 218762 217110 218836 217138
rect 219590 217110 219664 217138
rect 220418 217246 220584 217274
rect 221246 217246 221320 217274
rect 222028 217274 222056 228210
rect 222580 227866 222608 231676
rect 222764 231662 223146 231690
rect 223698 231662 223988 231690
rect 222568 227860 222620 227866
rect 222568 227802 222620 227808
rect 222764 221202 222792 231662
rect 222936 229220 222988 229226
rect 222936 229162 222988 229168
rect 222752 221196 222804 221202
rect 222752 221138 222804 221144
rect 222948 219434 222976 229162
rect 223960 221882 223988 231662
rect 224236 224398 224264 231676
rect 224512 231662 224802 231690
rect 224512 229094 224540 231662
rect 225340 229362 225368 231676
rect 225524 231662 225906 231690
rect 225328 229356 225380 229362
rect 225328 229298 225380 229304
rect 224420 229066 224540 229094
rect 224224 224392 224276 224398
rect 224224 224334 224276 224340
rect 223948 221876 224000 221882
rect 223948 221818 224000 221824
rect 223764 221740 223816 221746
rect 223764 221682 223816 221688
rect 222856 219406 222976 219434
rect 222856 218890 222884 219406
rect 222844 218884 222896 218890
rect 222844 218826 222896 218832
rect 222936 218204 222988 218210
rect 222936 218146 222988 218152
rect 222028 217246 222102 217274
rect 217934 216988 217962 217110
rect 218762 216988 218790 217110
rect 219590 216988 219618 217110
rect 220418 216988 220446 217246
rect 221246 216988 221274 217246
rect 222074 216988 222102 217246
rect 222948 217138 222976 218146
rect 223776 217274 223804 221682
rect 224420 219706 224448 229066
rect 224592 224256 224644 224262
rect 224592 224198 224644 224204
rect 224408 219700 224460 219706
rect 224408 219642 224460 219648
rect 224224 219156 224276 219162
rect 224224 219098 224276 219104
rect 224236 218482 224264 219098
rect 224224 218476 224276 218482
rect 224224 218418 224276 218424
rect 224408 218476 224460 218482
rect 224408 218418 224460 218424
rect 224420 218210 224448 218418
rect 224408 218204 224460 218210
rect 224408 218146 224460 218152
rect 224604 217274 224632 224198
rect 225524 220386 225552 231662
rect 225972 229492 226024 229498
rect 225972 229434 226024 229440
rect 225984 228818 226012 229434
rect 225972 228812 226024 228818
rect 225972 228754 226024 228760
rect 226248 227860 226300 227866
rect 226248 227802 226300 227808
rect 226064 224392 226116 224398
rect 226064 224334 226116 224340
rect 225512 220380 225564 220386
rect 225512 220322 225564 220328
rect 226076 218210 226104 224334
rect 225420 218204 225472 218210
rect 225420 218146 225472 218152
rect 226064 218204 226116 218210
rect 226064 218146 226116 218152
rect 222902 217110 222976 217138
rect 223730 217246 223804 217274
rect 224558 217246 224632 217274
rect 222902 216988 222930 217110
rect 223730 216988 223758 217246
rect 224558 216988 224586 217246
rect 225432 217138 225460 218146
rect 226260 217274 226288 227802
rect 226444 221610 226472 231676
rect 226996 229634 227024 231676
rect 226984 229628 227036 229634
rect 226984 229570 227036 229576
rect 226984 229356 227036 229362
rect 226984 229298 227036 229304
rect 226996 228682 227024 229298
rect 226984 228676 227036 228682
rect 226984 228618 227036 228624
rect 227548 227322 227576 231676
rect 227536 227316 227588 227322
rect 227536 227258 227588 227264
rect 228100 223038 228128 231676
rect 228652 223990 228680 231676
rect 228824 227316 228876 227322
rect 228824 227258 228876 227264
rect 228640 223984 228692 223990
rect 228640 223926 228692 223932
rect 228088 223032 228140 223038
rect 228088 222974 228140 222980
rect 227076 221876 227128 221882
rect 227076 221818 227128 221824
rect 226432 221604 226484 221610
rect 226432 221546 226484 221552
rect 226892 220244 226944 220250
rect 226892 220186 226944 220192
rect 226904 219502 226932 220186
rect 226892 219496 226944 219502
rect 226892 219438 226944 219444
rect 227088 217274 227116 221818
rect 227904 221604 227956 221610
rect 227904 221546 227956 221552
rect 227916 217274 227944 221546
rect 228836 219434 228864 227258
rect 229204 225214 229232 231676
rect 229756 229498 229784 231676
rect 229940 231662 230322 231690
rect 230492 231662 230874 231690
rect 229744 229492 229796 229498
rect 229744 229434 229796 229440
rect 229192 225208 229244 225214
rect 229192 225150 229244 225156
rect 229940 220522 229968 231662
rect 230492 222018 230520 231662
rect 231412 229906 231440 231676
rect 231400 229900 231452 229906
rect 231400 229842 231452 229848
rect 230664 229628 230716 229634
rect 230664 229570 230716 229576
rect 230676 227866 230704 229570
rect 231676 228676 231728 228682
rect 231676 228618 231728 228624
rect 230664 227860 230716 227866
rect 230664 227802 230716 227808
rect 230480 222012 230532 222018
rect 230480 221954 230532 221960
rect 229928 220516 229980 220522
rect 229928 220458 229980 220464
rect 230388 220380 230440 220386
rect 230388 220322 230440 220328
rect 228744 219406 228864 219434
rect 228744 217274 228772 219406
rect 229560 218884 229612 218890
rect 229560 218826 229612 218832
rect 225386 217110 225460 217138
rect 226214 217246 226288 217274
rect 227042 217246 227116 217274
rect 227870 217246 227944 217274
rect 228698 217246 228772 217274
rect 225386 216988 225414 217110
rect 226214 216988 226242 217246
rect 227042 216988 227070 217246
rect 227870 216988 227898 217246
rect 228698 216988 228726 217246
rect 229572 217138 229600 218826
rect 230400 217274 230428 220322
rect 231688 218074 231716 228618
rect 231964 222630 231992 231676
rect 232516 223174 232544 231676
rect 233068 227458 233096 231676
rect 233436 231662 233634 231690
rect 233240 229900 233292 229906
rect 233240 229842 233292 229848
rect 233056 227452 233108 227458
rect 233056 227394 233108 227400
rect 233252 226386 233280 229842
rect 232884 226358 233280 226386
rect 232504 223168 232556 223174
rect 232504 223110 232556 223116
rect 231952 222624 232004 222630
rect 231952 222566 232004 222572
rect 231216 218068 231268 218074
rect 231216 218010 231268 218016
rect 231676 218068 231728 218074
rect 231676 218010 231728 218016
rect 232044 218068 232096 218074
rect 232044 218010 232096 218016
rect 229526 217110 229600 217138
rect 230354 217246 230428 217274
rect 229526 216988 229554 217110
rect 230354 216988 230382 217246
rect 231228 217138 231256 218010
rect 232056 217138 232084 218010
rect 232884 217274 232912 226358
rect 233056 223032 233108 223038
rect 233056 222974 233108 222980
rect 233068 218074 233096 222974
rect 233436 220250 233464 231662
rect 234172 225758 234200 231676
rect 234436 227452 234488 227458
rect 234436 227394 234488 227400
rect 234160 225752 234212 225758
rect 234160 225694 234212 225700
rect 233700 220516 233752 220522
rect 233700 220458 233752 220464
rect 233424 220244 233476 220250
rect 233424 220186 233476 220192
rect 233056 218068 233108 218074
rect 233056 218010 233108 218016
rect 233712 217274 233740 220458
rect 231182 217110 231256 217138
rect 232010 217110 232084 217138
rect 232838 217246 232912 217274
rect 233666 217246 233740 217274
rect 234448 217274 234476 227394
rect 234724 223310 234752 231676
rect 235000 231662 235290 231690
rect 234712 223304 234764 223310
rect 234712 223246 234764 223252
rect 235000 222154 235028 231662
rect 235828 230042 235856 231676
rect 235816 230036 235868 230042
rect 235816 229978 235868 229984
rect 236380 229362 236408 231676
rect 236564 231662 236946 231690
rect 236368 229356 236420 229362
rect 236368 229298 236420 229304
rect 236564 229094 236592 231662
rect 236472 229066 236592 229094
rect 235908 225752 235960 225758
rect 235908 225694 235960 225700
rect 234988 222148 235040 222154
rect 234988 222090 235040 222096
rect 235920 218074 235948 225694
rect 236472 220658 236500 229066
rect 236644 227860 236696 227866
rect 236644 227802 236696 227808
rect 236460 220652 236512 220658
rect 236460 220594 236512 220600
rect 236184 219428 236236 219434
rect 236184 219370 236236 219376
rect 235356 218068 235408 218074
rect 235356 218010 235408 218016
rect 235908 218068 235960 218074
rect 235908 218010 235960 218016
rect 234448 217246 234522 217274
rect 231182 216988 231210 217110
rect 232010 216988 232038 217110
rect 232838 216988 232866 217246
rect 233666 216988 233694 217246
rect 234494 216988 234522 217246
rect 235368 217138 235396 218010
rect 236196 217138 236224 219370
rect 236656 218210 236684 227802
rect 237484 224806 237512 231676
rect 238036 227866 238064 231676
rect 238312 231662 238602 231690
rect 238024 227860 238076 227866
rect 238024 227802 238076 227808
rect 238312 226030 238340 231662
rect 238576 228812 238628 228818
rect 238576 228754 238628 228760
rect 238300 226024 238352 226030
rect 238300 225966 238352 225972
rect 237472 224800 237524 224806
rect 237472 224742 237524 224748
rect 237012 223168 237064 223174
rect 237012 223110 237064 223116
rect 236644 218204 236696 218210
rect 236644 218146 236696 218152
rect 237024 217274 237052 223110
rect 237840 220244 237892 220250
rect 237840 220186 237892 220192
rect 237852 217274 237880 220186
rect 235322 217110 235396 217138
rect 236150 217110 236224 217138
rect 236978 217246 237052 217274
rect 237806 217246 237880 217274
rect 238588 217274 238616 228754
rect 239140 223582 239168 231676
rect 239692 224942 239720 231676
rect 240244 230314 240272 231676
rect 240232 230308 240284 230314
rect 240232 230250 240284 230256
rect 240048 227860 240100 227866
rect 240048 227802 240100 227808
rect 239680 224936 239732 224942
rect 239680 224878 239732 224884
rect 239128 223576 239180 223582
rect 239128 223518 239180 223524
rect 239312 222760 239364 222766
rect 239312 222702 239364 222708
rect 239324 219298 239352 222702
rect 239312 219292 239364 219298
rect 239312 219234 239364 219240
rect 240060 218074 240088 227802
rect 240796 225622 240824 231676
rect 241072 231662 241362 231690
rect 241072 229094 241100 231662
rect 241612 230036 241664 230042
rect 241612 229978 241664 229984
rect 240980 229066 241100 229094
rect 240784 225616 240836 225622
rect 240784 225558 240836 225564
rect 240980 222630 241008 229066
rect 241624 227866 241652 229978
rect 241612 227860 241664 227866
rect 241612 227802 241664 227808
rect 241152 225616 241204 225622
rect 241152 225558 241204 225564
rect 240968 222624 241020 222630
rect 240968 222566 241020 222572
rect 240324 220788 240376 220794
rect 240324 220730 240376 220736
rect 239496 218068 239548 218074
rect 239496 218010 239548 218016
rect 240048 218068 240100 218074
rect 240048 218010 240100 218016
rect 238588 217246 238662 217274
rect 235322 216988 235350 217110
rect 236150 216988 236178 217110
rect 236978 216988 237006 217246
rect 237806 216988 237834 217246
rect 238634 216988 238662 217246
rect 239508 217138 239536 218010
rect 240336 217274 240364 220730
rect 241164 217274 241192 225558
rect 241900 225486 241928 231676
rect 241888 225480 241940 225486
rect 241888 225422 241940 225428
rect 242164 223372 242216 223378
rect 242164 223314 242216 223320
rect 242176 218346 242204 223314
rect 242452 222766 242480 231676
rect 243004 226166 243032 231676
rect 243280 231662 243570 231690
rect 243832 231662 244122 231690
rect 242992 226160 243044 226166
rect 242992 226102 243044 226108
rect 242440 222760 242492 222766
rect 242440 222702 242492 222708
rect 242808 222760 242860 222766
rect 242808 222702 242860 222708
rect 242624 219020 242676 219026
rect 242624 218962 242676 218968
rect 242164 218340 242216 218346
rect 242164 218282 242216 218288
rect 241980 218068 242032 218074
rect 241980 218010 242032 218016
rect 239462 217110 239536 217138
rect 240290 217246 240364 217274
rect 241118 217246 241192 217274
rect 239462 216988 239490 217110
rect 240290 216988 240318 217246
rect 241118 216988 241146 217246
rect 241992 217138 242020 218010
rect 242636 217274 242664 218962
rect 242820 218074 242848 222702
rect 243280 219978 243308 231662
rect 243832 223514 243860 231662
rect 244660 230178 244688 231676
rect 244924 230308 244976 230314
rect 244924 230250 244976 230256
rect 244648 230172 244700 230178
rect 244648 230114 244700 230120
rect 244188 225888 244240 225894
rect 244188 225830 244240 225836
rect 243820 223508 243872 223514
rect 243820 223450 243872 223456
rect 243268 219972 243320 219978
rect 243268 219914 243320 219920
rect 243544 218748 243596 218754
rect 243544 218690 243596 218696
rect 243556 218346 243584 218690
rect 243544 218340 243596 218346
rect 243544 218282 243596 218288
rect 244200 218074 244228 225830
rect 244936 218618 244964 230250
rect 245212 228954 245240 231676
rect 245200 228948 245252 228954
rect 245200 228890 245252 228896
rect 245476 228948 245528 228954
rect 245476 228890 245528 228896
rect 245292 223508 245344 223514
rect 245292 223450 245344 223456
rect 244924 218612 244976 218618
rect 244924 218554 244976 218560
rect 245304 218074 245332 223450
rect 242808 218068 242860 218074
rect 242808 218010 242860 218016
rect 243636 218068 243688 218074
rect 243636 218010 243688 218016
rect 244188 218068 244240 218074
rect 244188 218010 244240 218016
rect 244464 218068 244516 218074
rect 244464 218010 244516 218016
rect 245292 218068 245344 218074
rect 245292 218010 245344 218016
rect 242636 217246 242802 217274
rect 241946 217110 242020 217138
rect 241946 216988 241974 217110
rect 242774 216988 242802 217246
rect 243648 217138 243676 218010
rect 244476 217138 244504 218010
rect 245488 217274 245516 228890
rect 245764 226302 245792 231676
rect 245752 226296 245804 226302
rect 245752 226238 245804 226244
rect 246316 223378 246344 231676
rect 246868 230314 246896 231676
rect 246856 230308 246908 230314
rect 246856 230250 246908 230256
rect 247420 227594 247448 231676
rect 247604 231662 247986 231690
rect 247408 227588 247460 227594
rect 247408 227530 247460 227536
rect 246856 226024 246908 226030
rect 246856 225966 246908 225972
rect 246672 223576 246724 223582
rect 246672 223518 246724 223524
rect 246304 223372 246356 223378
rect 246304 223314 246356 223320
rect 246684 222766 246712 223518
rect 246672 222760 246724 222766
rect 246672 222702 246724 222708
rect 246120 218068 246172 218074
rect 246120 218010 246172 218016
rect 243602 217110 243676 217138
rect 244430 217110 244504 217138
rect 245258 217246 245516 217274
rect 243602 216988 243630 217110
rect 244430 216988 244458 217110
rect 245258 216988 245286 217246
rect 246132 217138 246160 218010
rect 246868 217274 246896 225966
rect 247604 219858 247632 231662
rect 247776 230172 247828 230178
rect 247776 230114 247828 230120
rect 247788 229094 247816 230114
rect 247512 219842 247632 219858
rect 247500 219836 247632 219842
rect 247552 219830 247632 219836
rect 247696 229066 247816 229094
rect 247500 219778 247552 219784
rect 247696 219434 247724 229066
rect 248524 228546 248552 231676
rect 249076 229498 249104 231676
rect 249064 229492 249116 229498
rect 249064 229434 249116 229440
rect 248512 228540 248564 228546
rect 248512 228482 248564 228488
rect 249064 227792 249116 227798
rect 249064 227734 249116 227740
rect 247868 220652 247920 220658
rect 247868 220594 247920 220600
rect 247880 219434 247908 220594
rect 247604 219406 247724 219434
rect 247788 219406 247908 219434
rect 247604 218074 247632 219406
rect 247592 218068 247644 218074
rect 247592 218010 247644 218016
rect 247788 217274 247816 219406
rect 249076 218346 249104 227734
rect 249628 227662 249656 231676
rect 249616 227656 249668 227662
rect 249616 227598 249668 227604
rect 250180 227050 250208 231676
rect 250168 227044 250220 227050
rect 250168 226986 250220 226992
rect 249616 226908 249668 226914
rect 249616 226850 249668 226856
rect 249432 219292 249484 219298
rect 249432 219234 249484 219240
rect 249064 218340 249116 218346
rect 249064 218282 249116 218288
rect 248604 218068 248656 218074
rect 248604 218010 248656 218016
rect 246868 217246 246942 217274
rect 246086 217110 246160 217138
rect 246086 216988 246114 217110
rect 246914 216988 246942 217246
rect 247742 217246 247816 217274
rect 247742 216988 247770 217246
rect 248616 217138 248644 218010
rect 249444 217138 249472 219234
rect 249628 218074 249656 226850
rect 250732 225350 250760 231676
rect 251284 227798 251312 231676
rect 251836 229090 251864 231676
rect 252020 231662 252402 231690
rect 252664 231662 252954 231690
rect 252020 229094 252048 231662
rect 251824 229084 251876 229090
rect 252020 229066 252140 229094
rect 251824 229026 251876 229032
rect 251272 227792 251324 227798
rect 251272 227734 251324 227740
rect 251732 227792 251784 227798
rect 251732 227734 251784 227740
rect 251088 227656 251140 227662
rect 251088 227598 251140 227604
rect 250720 225344 250772 225350
rect 250720 225286 250772 225292
rect 250904 224528 250956 224534
rect 250904 224470 250956 224476
rect 250916 219434 250944 224470
rect 250916 219406 251036 219434
rect 249616 218068 249668 218074
rect 249616 218010 249668 218016
rect 250260 218068 250312 218074
rect 250260 218010 250312 218016
rect 250272 217138 250300 218010
rect 251008 217274 251036 219406
rect 251100 218090 251128 227598
rect 251744 219162 251772 227734
rect 251916 222012 251968 222018
rect 251916 221954 251968 221960
rect 251732 219156 251784 219162
rect 251732 219098 251784 219104
rect 251100 218074 251220 218090
rect 251100 218068 251232 218074
rect 251100 218062 251180 218068
rect 251180 218010 251232 218016
rect 251928 217274 251956 221954
rect 252112 221066 252140 229066
rect 252664 221338 252692 231662
rect 253492 230450 253520 231676
rect 253480 230444 253532 230450
rect 253480 230386 253532 230392
rect 253572 228540 253624 228546
rect 253572 228482 253624 228488
rect 252652 221332 252704 221338
rect 252652 221274 252704 221280
rect 252100 221060 252152 221066
rect 252100 221002 252152 221008
rect 252744 219156 252796 219162
rect 252744 219098 252796 219104
rect 251008 217246 251082 217274
rect 248570 217110 248644 217138
rect 249398 217110 249472 217138
rect 250226 217110 250300 217138
rect 248570 216988 248598 217110
rect 249398 216988 249426 217110
rect 250226 216988 250254 217110
rect 251054 216988 251082 217246
rect 251882 217246 251956 217274
rect 251882 216988 251910 217246
rect 252756 217138 252784 219098
rect 253584 217274 253612 228482
rect 254044 224126 254072 231676
rect 254320 231662 254610 231690
rect 254032 224120 254084 224126
rect 254032 224062 254084 224068
rect 253848 220924 253900 220930
rect 253848 220866 253900 220872
rect 253860 218482 253888 220866
rect 254320 220114 254348 231662
rect 255148 227186 255176 231676
rect 255700 227798 255728 231676
rect 255964 230308 256016 230314
rect 255964 230250 256016 230256
rect 255688 227792 255740 227798
rect 255688 227734 255740 227740
rect 255136 227180 255188 227186
rect 255136 227122 255188 227128
rect 255228 224800 255280 224806
rect 255228 224742 255280 224748
rect 254308 220108 254360 220114
rect 254308 220050 254360 220056
rect 254400 218680 254452 218686
rect 254400 218622 254452 218628
rect 253848 218476 253900 218482
rect 253848 218418 253900 218424
rect 252710 217110 252784 217138
rect 253538 217246 253612 217274
rect 252710 216988 252738 217110
rect 253538 216988 253566 217246
rect 254412 217138 254440 218622
rect 255240 217274 255268 224742
rect 255976 219162 256004 230250
rect 256252 229094 256280 231676
rect 256252 229066 256372 229094
rect 256148 227044 256200 227050
rect 256148 226986 256200 226992
rect 255964 219156 256016 219162
rect 255964 219098 256016 219104
rect 256160 218686 256188 226986
rect 256344 223854 256372 229066
rect 256516 227588 256568 227594
rect 256516 227530 256568 227536
rect 256528 226914 256556 227530
rect 256516 226908 256568 226914
rect 256516 226850 256568 226856
rect 256332 223848 256384 223854
rect 256332 223790 256384 223796
rect 256804 221474 256832 231676
rect 257356 224670 257384 231676
rect 257908 229770 257936 231676
rect 257896 229764 257948 229770
rect 257896 229706 257948 229712
rect 258460 228274 258488 231676
rect 258644 231662 259026 231690
rect 258448 228268 258500 228274
rect 258448 228210 258500 228216
rect 257344 224664 257396 224670
rect 257344 224606 257396 224612
rect 258172 222148 258224 222154
rect 258172 222090 258224 222096
rect 258184 221882 258212 222090
rect 258644 221882 258672 231662
rect 259276 227860 259328 227866
rect 259276 227802 259328 227808
rect 258172 221876 258224 221882
rect 258172 221818 258224 221824
rect 258632 221876 258684 221882
rect 258632 221818 258684 221824
rect 258540 221740 258592 221746
rect 258540 221682 258592 221688
rect 256792 221468 256844 221474
rect 256792 221410 256844 221416
rect 257712 221468 257764 221474
rect 257712 221410 257764 221416
rect 256884 220108 256936 220114
rect 256884 220050 256936 220056
rect 256148 218680 256200 218686
rect 256148 218622 256200 218628
rect 256056 218544 256108 218550
rect 256056 218486 256108 218492
rect 254366 217110 254440 217138
rect 255194 217246 255268 217274
rect 254366 216988 254394 217110
rect 255194 216988 255222 217246
rect 256068 217138 256096 218486
rect 256896 217274 256924 220050
rect 257724 217274 257752 221410
rect 258552 217274 258580 221682
rect 256022 217110 256096 217138
rect 256850 217246 256924 217274
rect 257678 217246 257752 217274
rect 258506 217246 258580 217274
rect 259288 217274 259316 227802
rect 259564 222902 259592 231676
rect 259840 231662 260130 231690
rect 260392 231662 260682 231690
rect 261036 231662 261234 231690
rect 259552 222896 259604 222902
rect 259552 222838 259604 222844
rect 259840 220930 259868 231662
rect 260392 224398 260420 231662
rect 260380 224392 260432 224398
rect 260380 224334 260432 224340
rect 260196 224120 260248 224126
rect 260196 224062 260248 224068
rect 259828 220924 259880 220930
rect 259828 220866 259880 220872
rect 260208 217274 260236 224062
rect 261036 222154 261064 231662
rect 261576 229764 261628 229770
rect 261576 229706 261628 229712
rect 261588 227866 261616 229706
rect 261576 227860 261628 227866
rect 261576 227802 261628 227808
rect 261772 224262 261800 231676
rect 262324 229634 262352 231676
rect 262312 229628 262364 229634
rect 262312 229570 262364 229576
rect 262036 229084 262088 229090
rect 262036 229026 262088 229032
rect 261760 224256 261812 224262
rect 261760 224198 261812 224204
rect 261852 222896 261904 222902
rect 261852 222838 261904 222844
rect 261024 222148 261076 222154
rect 261024 222090 261076 222096
rect 261864 218074 261892 222838
rect 261024 218068 261076 218074
rect 261024 218010 261076 218016
rect 261852 218068 261904 218074
rect 261852 218010 261904 218016
rect 259288 217246 259362 217274
rect 256022 216988 256050 217110
rect 256850 216988 256878 217246
rect 257678 216988 257706 217246
rect 258506 216988 258534 217246
rect 259334 216988 259362 217246
rect 260162 217246 260236 217274
rect 260162 216988 260190 217246
rect 261036 217138 261064 218010
rect 262048 217274 262076 229026
rect 262876 227322 262904 231676
rect 263060 231662 263442 231690
rect 263796 231662 263994 231690
rect 262864 227316 262916 227322
rect 262864 227258 262916 227264
rect 262680 224256 262732 224262
rect 262680 224198 262732 224204
rect 262692 218890 262720 224198
rect 263060 220386 263088 231662
rect 263508 221876 263560 221882
rect 263508 221818 263560 221824
rect 263048 220380 263100 220386
rect 263048 220322 263100 220328
rect 262864 219156 262916 219162
rect 262864 219098 262916 219104
rect 262680 218884 262732 218890
rect 262680 218826 262732 218832
rect 262680 218748 262732 218754
rect 262680 218690 262732 218696
rect 260990 217110 261064 217138
rect 261818 217246 262076 217274
rect 260990 216988 261018 217110
rect 261818 216988 261846 217246
rect 262692 217138 262720 218690
rect 262876 218550 262904 219098
rect 262864 218544 262916 218550
rect 262864 218486 262916 218492
rect 263520 217274 263548 221818
rect 263796 221610 263824 231662
rect 264532 224262 264560 231676
rect 264520 224256 264572 224262
rect 264520 224198 264572 224204
rect 265084 223038 265112 231676
rect 265360 231662 265650 231690
rect 265072 223032 265124 223038
rect 265072 222974 265124 222980
rect 263784 221604 263836 221610
rect 263784 221546 263836 221552
rect 265360 220522 265388 231662
rect 266188 228682 266216 231676
rect 266740 229906 266768 231676
rect 266728 229900 266780 229906
rect 266728 229842 266780 229848
rect 267004 229900 267056 229906
rect 267004 229842 267056 229848
rect 266176 228676 266228 228682
rect 266176 228618 266228 228624
rect 266360 228676 266412 228682
rect 266360 228618 266412 228624
rect 266372 228562 266400 228618
rect 266280 228534 266400 228562
rect 265992 222148 266044 222154
rect 265992 222090 266044 222096
rect 265348 220516 265400 220522
rect 265348 220458 265400 220464
rect 264336 220380 264388 220386
rect 264336 220322 264388 220328
rect 264348 217274 264376 220322
rect 265164 218068 265216 218074
rect 265164 218010 265216 218016
rect 262646 217110 262720 217138
rect 263474 217246 263548 217274
rect 264302 217246 264376 217274
rect 262646 216988 262674 217110
rect 263474 216988 263502 217246
rect 264302 216988 264330 217246
rect 265176 217138 265204 218010
rect 266004 217274 266032 222090
rect 266280 218074 266308 228534
rect 267016 222154 267044 229842
rect 267292 225758 267320 231676
rect 267844 229094 267872 231676
rect 268396 229094 268424 231676
rect 268672 231662 268962 231690
rect 268672 229094 268700 231662
rect 267844 229066 268148 229094
rect 267280 225752 267332 225758
rect 267280 225694 267332 225700
rect 267648 225752 267700 225758
rect 267648 225694 267700 225700
rect 267464 223440 267516 223446
rect 267464 223382 267516 223388
rect 267004 222148 267056 222154
rect 267004 222090 267056 222096
rect 267476 218074 267504 223382
rect 266268 218068 266320 218074
rect 266268 218010 266320 218016
rect 266820 218068 266872 218074
rect 266820 218010 266872 218016
rect 267464 218068 267516 218074
rect 267464 218010 267516 218016
rect 265130 217110 265204 217138
rect 265958 217246 266032 217274
rect 265130 216988 265158 217110
rect 265958 216988 265986 217246
rect 266832 217138 266860 218010
rect 267660 217274 267688 225694
rect 268120 223174 268148 229066
rect 268304 229066 268424 229094
rect 268488 229066 268700 229094
rect 268304 227458 268332 229066
rect 268292 227452 268344 227458
rect 268292 227394 268344 227400
rect 268108 223168 268160 223174
rect 268108 223110 268160 223116
rect 268488 222986 268516 229066
rect 269500 228818 269528 231676
rect 269776 231662 270066 231690
rect 269488 228812 269540 228818
rect 269488 228754 269540 228760
rect 267936 222958 268516 222986
rect 267936 219434 267964 222958
rect 269776 220794 269804 231662
rect 270132 226160 270184 226166
rect 270132 226102 270184 226108
rect 269764 220788 269816 220794
rect 269764 220730 269816 220736
rect 268476 220516 268528 220522
rect 268476 220458 268528 220464
rect 267924 219428 267976 219434
rect 267924 219370 267976 219376
rect 268488 217274 268516 220458
rect 269304 219428 269356 219434
rect 269304 219370 269356 219376
rect 266786 217110 266860 217138
rect 267614 217246 267688 217274
rect 268442 217246 268516 217274
rect 266786 216988 266814 217110
rect 267614 216988 267642 217246
rect 268442 216988 268470 217246
rect 269316 217138 269344 219370
rect 270144 217274 270172 226102
rect 270604 220250 270632 231676
rect 271156 230042 271184 231676
rect 271144 230036 271196 230042
rect 271144 229978 271196 229984
rect 271708 223582 271736 231676
rect 272260 225894 272288 231676
rect 272432 227316 272484 227322
rect 272432 227258 272484 227264
rect 272248 225888 272300 225894
rect 272248 225830 272300 225836
rect 271696 223576 271748 223582
rect 271696 223518 271748 223524
rect 271788 223032 271840 223038
rect 271788 222974 271840 222980
rect 270592 220244 270644 220250
rect 270592 220186 270644 220192
rect 271604 220244 271656 220250
rect 271604 220186 271656 220192
rect 271616 219434 271644 220186
rect 271616 219406 271736 219434
rect 270960 218068 271012 218074
rect 270960 218010 271012 218016
rect 269270 217110 269344 217138
rect 270098 217246 270172 217274
rect 269270 216988 269298 217110
rect 270098 216988 270126 217246
rect 270972 217138 271000 218010
rect 271708 217274 271736 219406
rect 271800 218090 271828 222974
rect 272444 219162 272472 227258
rect 272812 225622 272840 231676
rect 273364 229094 273392 231676
rect 273364 229066 273484 229094
rect 272800 225616 272852 225622
rect 272800 225558 272852 225564
rect 273168 225004 273220 225010
rect 273168 224946 273220 224952
rect 272432 219156 272484 219162
rect 272432 219098 272484 219104
rect 271800 218074 271920 218090
rect 273180 218074 273208 224946
rect 273456 219026 273484 229066
rect 273916 228954 273944 231676
rect 273904 228948 273956 228954
rect 273904 228890 273956 228896
rect 274468 226030 274496 231676
rect 274456 226024 274508 226030
rect 274456 225966 274508 225972
rect 274548 225616 274600 225622
rect 274548 225558 274600 225564
rect 273444 219020 273496 219026
rect 273444 218962 273496 218968
rect 274272 218204 274324 218210
rect 274272 218146 274324 218152
rect 271800 218068 271932 218074
rect 271800 218062 271880 218068
rect 271880 218010 271932 218016
rect 272616 218068 272668 218074
rect 272616 218010 272668 218016
rect 273168 218068 273220 218074
rect 273168 218010 273220 218016
rect 273444 218068 273496 218074
rect 273444 218010 273496 218016
rect 271708 217246 271782 217274
rect 270926 217110 271000 217138
rect 270926 216988 270954 217110
rect 271754 216988 271782 217246
rect 272628 217138 272656 218010
rect 273456 217138 273484 218010
rect 274284 217138 274312 218146
rect 274560 218074 274588 225558
rect 275020 223310 275048 231676
rect 275572 230178 275600 231676
rect 275560 230172 275612 230178
rect 275560 230114 275612 230120
rect 275652 230036 275704 230042
rect 275652 229978 275704 229984
rect 275664 225010 275692 229978
rect 275836 228812 275888 228818
rect 275836 228754 275888 228760
rect 275652 225004 275704 225010
rect 275652 224946 275704 224952
rect 275284 224256 275336 224262
rect 275284 224198 275336 224204
rect 275008 223304 275060 223310
rect 275008 223246 275060 223252
rect 275296 218210 275324 224198
rect 275652 219020 275704 219026
rect 275652 218962 275704 218968
rect 275284 218204 275336 218210
rect 275284 218146 275336 218152
rect 274548 218068 274600 218074
rect 274548 218010 274600 218016
rect 275100 218068 275152 218074
rect 275100 218010 275152 218016
rect 275112 217138 275140 218010
rect 275664 217274 275692 218962
rect 275848 218074 275876 228754
rect 276124 227594 276152 231676
rect 276676 227730 276704 231676
rect 276952 231662 277242 231690
rect 277596 231662 277794 231690
rect 278056 231662 278346 231690
rect 276664 227724 276716 227730
rect 276664 227666 276716 227672
rect 276112 227588 276164 227594
rect 276112 227530 276164 227536
rect 276952 220658 276980 231662
rect 277216 227180 277268 227186
rect 277216 227122 277268 227128
rect 276940 220652 276992 220658
rect 276940 220594 276992 220600
rect 277228 218074 277256 227122
rect 277596 218890 277624 231662
rect 278056 222018 278084 231662
rect 278884 228546 278912 231676
rect 278872 228540 278924 228546
rect 278872 228482 278924 228488
rect 279436 224534 279464 231676
rect 279988 230314 280016 231676
rect 279976 230308 280028 230314
rect 279976 230250 280028 230256
rect 279792 230172 279844 230178
rect 279792 230114 279844 230120
rect 279424 224528 279476 224534
rect 279424 224470 279476 224476
rect 278044 222012 278096 222018
rect 278044 221954 278096 221960
rect 278412 221604 278464 221610
rect 278412 221546 278464 221552
rect 277584 218884 277636 218890
rect 277584 218826 277636 218832
rect 277584 218204 277636 218210
rect 277584 218146 277636 218152
rect 275836 218068 275888 218074
rect 275836 218010 275888 218016
rect 276756 218068 276808 218074
rect 276756 218010 276808 218016
rect 277216 218068 277268 218074
rect 277216 218010 277268 218016
rect 275664 217246 275922 217274
rect 272582 217110 272656 217138
rect 273410 217110 273484 217138
rect 274238 217110 274312 217138
rect 275066 217110 275140 217138
rect 272582 216988 272610 217110
rect 273410 216988 273438 217110
rect 274238 216988 274266 217110
rect 275066 216988 275094 217110
rect 275894 216988 275922 217246
rect 276768 217138 276796 218010
rect 277596 217138 277624 218146
rect 278424 217274 278452 221546
rect 279804 218074 279832 230114
rect 280540 224806 280568 231676
rect 280724 231662 281106 231690
rect 280528 224800 280580 224806
rect 280528 224742 280580 224748
rect 279976 224528 280028 224534
rect 279976 224470 280028 224476
rect 279240 218068 279292 218074
rect 279240 218010 279292 218016
rect 279792 218068 279844 218074
rect 279792 218010 279844 218016
rect 276722 217110 276796 217138
rect 277550 217110 277624 217138
rect 278378 217246 278452 217274
rect 276722 216988 276750 217110
rect 277550 216988 277578 217110
rect 278378 216988 278406 217246
rect 279252 217138 279280 218010
rect 279988 217274 280016 224470
rect 280724 220114 280752 231662
rect 281644 227050 281672 231676
rect 282196 227322 282224 231676
rect 282472 231662 282762 231690
rect 282184 227316 282236 227322
rect 282184 227258 282236 227264
rect 281632 227044 281684 227050
rect 281632 226986 281684 226992
rect 280896 222012 280948 222018
rect 280896 221954 280948 221960
rect 280712 220108 280764 220114
rect 280712 220050 280764 220056
rect 280908 217274 280936 221954
rect 282472 221746 282500 231662
rect 282736 227044 282788 227050
rect 282736 226986 282788 226992
rect 282460 221740 282512 221746
rect 282460 221682 282512 221688
rect 281264 220108 281316 220114
rect 281264 220050 281316 220056
rect 281276 218210 281304 220050
rect 282552 218884 282604 218890
rect 282552 218826 282604 218832
rect 281264 218204 281316 218210
rect 281264 218146 281316 218152
rect 281724 218068 281776 218074
rect 281724 218010 281776 218016
rect 279988 217246 280062 217274
rect 279206 217110 279280 217138
rect 279206 216988 279234 217110
rect 280034 216988 280062 217246
rect 280862 217246 280936 217274
rect 280862 216988 280890 217246
rect 281736 217138 281764 218010
rect 282564 217138 282592 218826
rect 282748 218074 282776 226986
rect 283300 224398 283328 231676
rect 283484 231662 283866 231690
rect 283288 224392 283340 224398
rect 283288 224334 283340 224340
rect 283484 224210 283512 231662
rect 284404 229770 284432 231676
rect 284392 229764 284444 229770
rect 284392 229706 284444 229712
rect 284956 229090 284984 231676
rect 285140 231662 285522 231690
rect 284944 229084 284996 229090
rect 284944 229026 284996 229032
rect 283208 224182 283512 224210
rect 283208 221474 283236 224182
rect 284208 223168 284260 223174
rect 284208 223110 284260 223116
rect 283196 221468 283248 221474
rect 283196 221410 283248 221416
rect 283380 221468 283432 221474
rect 283380 221410 283432 221416
rect 282736 218068 282788 218074
rect 282736 218010 282788 218016
rect 283392 217274 283420 221410
rect 284220 217274 284248 223110
rect 285140 221882 285168 231662
rect 285312 230308 285364 230314
rect 285312 230250 285364 230256
rect 285128 221876 285180 221882
rect 285128 221818 285180 221824
rect 285324 219434 285352 230250
rect 285588 228540 285640 228546
rect 285588 228482 285640 228488
rect 284944 219428 285352 219434
rect 284996 219406 285352 219428
rect 284944 219370 284996 219376
rect 285600 218074 285628 228482
rect 286060 222902 286088 231676
rect 286244 231662 286626 231690
rect 286048 222896 286100 222902
rect 286048 222838 286100 222844
rect 286244 219434 286272 231662
rect 286692 228948 286744 228954
rect 286692 228890 286744 228896
rect 286060 219406 286272 219434
rect 285864 219156 285916 219162
rect 285864 219098 285916 219104
rect 285036 218068 285088 218074
rect 285036 218010 285088 218016
rect 285588 218068 285640 218074
rect 285588 218010 285640 218016
rect 281690 217110 281764 217138
rect 282518 217110 282592 217138
rect 283346 217246 283420 217274
rect 284174 217246 284248 217274
rect 281690 216988 281718 217110
rect 282518 216988 282546 217110
rect 283346 216988 283374 217246
rect 284174 216988 284202 217246
rect 285048 217138 285076 218010
rect 285876 217138 285904 219098
rect 286060 218754 286088 219406
rect 286048 218748 286100 218754
rect 286048 218690 286100 218696
rect 286704 217274 286732 228890
rect 287164 228682 287192 231676
rect 287152 228676 287204 228682
rect 287152 228618 287204 228624
rect 287716 223446 287744 231676
rect 287900 231662 288282 231690
rect 287704 223440 287756 223446
rect 287704 223382 287756 223388
rect 287900 220386 287928 231662
rect 288820 229906 288848 231676
rect 289004 231662 289386 231690
rect 288808 229900 288860 229906
rect 288808 229842 288860 229848
rect 288348 220652 288400 220658
rect 288348 220594 288400 220600
rect 287888 220380 287940 220386
rect 287888 220322 287940 220328
rect 287520 218068 287572 218074
rect 287520 218010 287572 218016
rect 285002 217110 285076 217138
rect 285830 217110 285904 217138
rect 286658 217246 286732 217274
rect 285002 216988 285030 217110
rect 285830 216988 285858 217110
rect 286658 216988 286686 217246
rect 287532 217138 287560 218010
rect 288360 217274 288388 220594
rect 289004 220522 289032 231662
rect 289728 229764 289780 229770
rect 289728 229706 289780 229712
rect 288992 220516 289044 220522
rect 288992 220458 289044 220464
rect 288532 220380 288584 220386
rect 288532 220322 288584 220328
rect 288544 218074 288572 220322
rect 289740 218074 289768 229706
rect 289924 226166 289952 231676
rect 290200 231662 290490 231690
rect 289912 226160 289964 226166
rect 289912 226102 289964 226108
rect 290200 225758 290228 231662
rect 291028 230314 291056 231676
rect 291396 231662 291594 231690
rect 291016 230308 291068 230314
rect 291016 230250 291068 230256
rect 290464 229424 290516 229430
rect 290464 229366 290516 229372
rect 290188 225752 290240 225758
rect 290188 225694 290240 225700
rect 290476 219026 290504 229366
rect 291016 225752 291068 225758
rect 291016 225694 291068 225700
rect 290464 219020 290516 219026
rect 290464 218962 290516 218968
rect 290832 218204 290884 218210
rect 290832 218146 290884 218152
rect 288532 218068 288584 218074
rect 288532 218010 288584 218016
rect 289176 218068 289228 218074
rect 289176 218010 289228 218016
rect 289728 218068 289780 218074
rect 289728 218010 289780 218016
rect 290004 218068 290056 218074
rect 290004 218010 290056 218016
rect 287486 217110 287560 217138
rect 288314 217246 288388 217274
rect 287486 216988 287514 217110
rect 288314 216988 288342 217246
rect 289188 217138 289216 218010
rect 290016 217138 290044 218010
rect 290844 217138 290872 218146
rect 291028 218074 291056 225694
rect 291396 220250 291424 231662
rect 292132 225622 292160 231676
rect 292488 228676 292540 228682
rect 292488 228618 292540 228624
rect 292120 225616 292172 225622
rect 292120 225558 292172 225564
rect 291384 220244 291436 220250
rect 291384 220186 291436 220192
rect 292304 218748 292356 218754
rect 292304 218690 292356 218696
rect 291016 218068 291068 218074
rect 291016 218010 291068 218016
rect 291660 218068 291712 218074
rect 291660 218010 291712 218016
rect 291672 217138 291700 218010
rect 292316 217274 292344 218690
rect 292500 218074 292528 228618
rect 292684 223038 292712 231676
rect 293236 230042 293264 231676
rect 293224 230036 293276 230042
rect 293224 229978 293276 229984
rect 293788 228818 293816 231676
rect 293776 228812 293828 228818
rect 293776 228754 293828 228760
rect 293776 227316 293828 227322
rect 293776 227258 293828 227264
rect 292672 223032 292724 223038
rect 292672 222974 292724 222980
rect 293224 222896 293276 222902
rect 293224 222838 293276 222844
rect 293236 218210 293264 222838
rect 293224 218204 293276 218210
rect 293224 218146 293276 218152
rect 293788 218074 293816 227258
rect 294340 227186 294368 231676
rect 294892 229094 294920 231676
rect 295444 229430 295472 231676
rect 295720 231662 296010 231690
rect 295432 229424 295484 229430
rect 295432 229366 295484 229372
rect 294800 229066 294920 229094
rect 294328 227180 294380 227186
rect 294328 227122 294380 227128
rect 294800 224262 294828 229066
rect 295156 228812 295208 228818
rect 295156 228754 295208 228760
rect 294972 225616 295024 225622
rect 294972 225558 295024 225564
rect 294788 224256 294840 224262
rect 294788 224198 294840 224204
rect 294984 218074 295012 225558
rect 292488 218068 292540 218074
rect 292488 218010 292540 218016
rect 293316 218068 293368 218074
rect 293316 218010 293368 218016
rect 293776 218068 293828 218074
rect 293776 218010 293828 218016
rect 294144 218068 294196 218074
rect 294144 218010 294196 218016
rect 294972 218068 295024 218074
rect 294972 218010 295024 218016
rect 292316 217246 292482 217274
rect 289142 217110 289216 217138
rect 289970 217110 290044 217138
rect 290798 217110 290872 217138
rect 291626 217110 291700 217138
rect 289142 216988 289170 217110
rect 289970 216988 289998 217110
rect 290798 216988 290826 217110
rect 291626 216988 291654 217110
rect 292454 216988 292482 217246
rect 293328 217138 293356 218010
rect 294156 217138 294184 218010
rect 295168 217274 295196 228754
rect 295720 221610 295748 231662
rect 296548 224534 296576 231676
rect 296824 231662 297114 231690
rect 296824 229094 296852 231662
rect 297652 230246 297680 231676
rect 297640 230240 297692 230246
rect 297640 230182 297692 230188
rect 297364 230104 297416 230110
rect 297364 230046 297416 230052
rect 296824 229066 297128 229094
rect 296536 224528 296588 224534
rect 296536 224470 296588 224476
rect 296628 224392 296680 224398
rect 296628 224334 296680 224340
rect 296444 224256 296496 224262
rect 296444 224198 296496 224204
rect 295708 221604 295760 221610
rect 295708 221546 295760 221552
rect 296456 219434 296484 224198
rect 296456 219406 296576 219434
rect 295800 219292 295852 219298
rect 295800 219234 295852 219240
rect 293282 217110 293356 217138
rect 294110 217110 294184 217138
rect 294938 217246 295196 217274
rect 293282 216988 293310 217110
rect 294110 216988 294138 217110
rect 294938 216988 294966 217246
rect 295812 217138 295840 219234
rect 296548 217274 296576 219406
rect 296640 219314 296668 224334
rect 296904 221604 296956 221610
rect 296904 221546 296956 221552
rect 296640 219298 296760 219314
rect 296640 219292 296772 219298
rect 296640 219286 296720 219292
rect 296720 219234 296772 219240
rect 296916 219162 296944 221546
rect 297100 220114 297128 229066
rect 297376 222018 297404 230046
rect 298204 227050 298232 231676
rect 298480 231662 298770 231690
rect 298192 227044 298244 227050
rect 298192 226986 298244 226992
rect 297364 222012 297416 222018
rect 297364 221954 297416 221960
rect 298480 221746 298508 231662
rect 298744 230376 298796 230382
rect 298744 230318 298796 230324
rect 298468 221740 298520 221746
rect 298468 221682 298520 221688
rect 297456 221468 297508 221474
rect 297456 221410 297508 221416
rect 297088 220108 297140 220114
rect 297088 220050 297140 220056
rect 296904 219156 296956 219162
rect 296904 219098 296956 219104
rect 297468 217274 297496 221410
rect 298284 220108 298336 220114
rect 298284 220050 298336 220056
rect 298296 217274 298324 220050
rect 298756 218890 298784 230318
rect 299308 230110 299336 231676
rect 299860 230382 299888 231676
rect 299848 230376 299900 230382
rect 299848 230318 299900 230324
rect 299296 230104 299348 230110
rect 299296 230046 299348 230052
rect 300412 228546 300440 231676
rect 300584 229832 300636 229838
rect 300584 229774 300636 229780
rect 300400 228540 300452 228546
rect 300400 228482 300452 228488
rect 300596 223174 300624 229774
rect 300964 228954 300992 231676
rect 301516 229838 301544 231676
rect 301792 231662 302082 231690
rect 302436 231662 302634 231690
rect 301504 229832 301556 229838
rect 301504 229774 301556 229780
rect 300952 228948 301004 228954
rect 300952 228890 301004 228896
rect 300768 228540 300820 228546
rect 300768 228482 300820 228488
rect 300584 223168 300636 223174
rect 300584 223110 300636 223116
rect 300584 223032 300636 223038
rect 300584 222974 300636 222980
rect 300596 219434 300624 222974
rect 300780 219434 300808 228482
rect 301792 221610 301820 231662
rect 301780 221604 301832 221610
rect 301780 221546 301832 221552
rect 302436 220658 302464 231662
rect 303172 225758 303200 231676
rect 303160 225752 303212 225758
rect 303160 225694 303212 225700
rect 303252 221740 303304 221746
rect 303252 221682 303304 221688
rect 302424 220652 302476 220658
rect 302424 220594 302476 220600
rect 299940 219428 299992 219434
rect 300596 219406 300716 219434
rect 300780 219428 300912 219434
rect 300780 219406 300860 219428
rect 299940 219370 299992 219376
rect 298744 218884 298796 218890
rect 298744 218826 298796 218832
rect 299112 218068 299164 218074
rect 299112 218010 299164 218016
rect 296548 217246 296622 217274
rect 295766 217110 295840 217138
rect 295766 216988 295794 217110
rect 296594 216988 296622 217246
rect 297422 217246 297496 217274
rect 298250 217246 298324 217274
rect 297422 216988 297450 217246
rect 298250 216988 298278 217246
rect 299124 217138 299152 218010
rect 299952 217138 299980 219370
rect 300688 217274 300716 219406
rect 300860 219370 300912 219376
rect 302424 219156 302476 219162
rect 302424 219098 302476 219104
rect 301596 219020 301648 219026
rect 301596 218962 301648 218968
rect 300688 217246 300762 217274
rect 299078 217110 299152 217138
rect 299906 217110 299980 217138
rect 299078 216988 299106 217110
rect 299906 216988 299934 217110
rect 300734 216988 300762 217246
rect 301608 217138 301636 218962
rect 302436 217138 302464 219098
rect 303264 217274 303292 221682
rect 303724 220386 303752 231676
rect 304276 229702 304304 231676
rect 304264 229696 304316 229702
rect 304264 229638 304316 229644
rect 304080 229152 304132 229158
rect 304080 229094 304132 229100
rect 304092 224398 304120 229094
rect 304828 228682 304856 231676
rect 304816 228676 304868 228682
rect 304816 228618 304868 228624
rect 305380 227322 305408 231676
rect 305644 229764 305696 229770
rect 305644 229706 305696 229712
rect 305368 227316 305420 227322
rect 305368 227258 305420 227264
rect 304632 227044 304684 227050
rect 304632 226986 304684 226992
rect 304080 224392 304132 224398
rect 304080 224334 304132 224340
rect 303712 220380 303764 220386
rect 303712 220322 303764 220328
rect 303436 220244 303488 220250
rect 303436 220186 303488 220192
rect 303448 218074 303476 220186
rect 304644 218074 304672 226986
rect 304908 221468 304960 221474
rect 304908 221410 304960 221416
rect 303436 218068 303488 218074
rect 303436 218010 303488 218016
rect 304080 218068 304132 218074
rect 304080 218010 304132 218016
rect 304632 218068 304684 218074
rect 304632 218010 304684 218016
rect 301562 217110 301636 217138
rect 302390 217110 302464 217138
rect 303218 217246 303292 217274
rect 301562 216988 301590 217110
rect 302390 216988 302418 217110
rect 303218 216988 303246 217246
rect 304092 217138 304120 218010
rect 304920 217274 304948 221410
rect 305656 219162 305684 229706
rect 305932 229094 305960 231676
rect 305932 229066 306144 229094
rect 305920 223576 305972 223582
rect 305920 223518 305972 223524
rect 305644 219156 305696 219162
rect 305644 219098 305696 219104
rect 305736 218884 305788 218890
rect 305736 218826 305788 218832
rect 304046 217110 304120 217138
rect 304874 217246 304948 217274
rect 304046 216988 304074 217110
rect 304874 216988 304902 217246
rect 305748 217138 305776 218826
rect 305932 218754 305960 223518
rect 306116 222902 306144 229066
rect 306484 223582 306512 231676
rect 307036 228818 307064 231676
rect 307312 231662 307602 231690
rect 307024 228812 307076 228818
rect 307024 228754 307076 228760
rect 307312 224262 307340 231662
rect 308140 225622 308168 231676
rect 308692 229158 308720 231676
rect 308680 229152 308732 229158
rect 308680 229094 308732 229100
rect 308772 227792 308824 227798
rect 308772 227734 308824 227740
rect 308128 225616 308180 225622
rect 308128 225558 308180 225564
rect 307300 224256 307352 224262
rect 307300 224198 307352 224204
rect 307484 224256 307536 224262
rect 307484 224198 307536 224204
rect 306472 223576 306524 223582
rect 306472 223518 306524 223524
rect 306104 222896 306156 222902
rect 306104 222838 306156 222844
rect 307496 219434 307524 224198
rect 307404 219406 307524 219434
rect 305920 218748 305972 218754
rect 305920 218690 305972 218696
rect 306564 218204 306616 218210
rect 306564 218146 306616 218152
rect 306576 217138 306604 218146
rect 307404 217274 307432 219406
rect 308784 218074 308812 227734
rect 308956 225616 309008 225622
rect 308956 225558 309008 225564
rect 308220 218068 308272 218074
rect 308220 218010 308272 218016
rect 308772 218068 308824 218074
rect 308772 218010 308824 218016
rect 305702 217110 305776 217138
rect 306530 217110 306604 217138
rect 307358 217246 307432 217274
rect 305702 216988 305730 217110
rect 306530 216988 306558 217110
rect 307358 216988 307386 217246
rect 308232 217138 308260 218010
rect 308968 217274 308996 225558
rect 309244 220114 309272 231676
rect 309796 228546 309824 231676
rect 310072 231662 310362 231690
rect 310808 231662 310914 231690
rect 311176 231662 311466 231690
rect 309784 228540 309836 228546
rect 309784 228482 309836 228488
rect 310072 221610 310100 231662
rect 310336 227928 310388 227934
rect 310336 227870 310388 227876
rect 310060 221604 310112 221610
rect 310060 221546 310112 221552
rect 309232 220108 309284 220114
rect 309232 220050 309284 220056
rect 310348 218074 310376 227870
rect 310520 220788 310572 220794
rect 310520 220730 310572 220736
rect 310532 219026 310560 220730
rect 310808 220250 310836 231662
rect 311176 220794 311204 231662
rect 312004 221746 312032 231676
rect 312556 223038 312584 231676
rect 313108 229770 313136 231676
rect 313464 230376 313516 230382
rect 313464 230318 313516 230324
rect 313096 229764 313148 229770
rect 313096 229706 313148 229712
rect 313188 229628 313240 229634
rect 313188 229570 313240 229576
rect 312544 223032 312596 223038
rect 312544 222974 312596 222980
rect 311992 221740 312044 221746
rect 311992 221682 312044 221688
rect 313004 220856 313056 220862
rect 313004 220798 313056 220804
rect 311164 220788 311216 220794
rect 311164 220730 311216 220736
rect 310796 220244 310848 220250
rect 310796 220186 310848 220192
rect 311532 219496 311584 219502
rect 311532 219438 311584 219444
rect 310520 219020 310572 219026
rect 310520 218962 310572 218968
rect 310704 218748 310756 218754
rect 310704 218690 310756 218696
rect 309876 218068 309928 218074
rect 309876 218010 309928 218016
rect 310336 218068 310388 218074
rect 310336 218010 310388 218016
rect 308968 217246 309042 217274
rect 308186 217110 308260 217138
rect 308186 216988 308214 217110
rect 309014 216988 309042 217246
rect 309888 217138 309916 218010
rect 310716 217138 310744 218690
rect 311544 217274 311572 219438
rect 313016 219434 313044 220798
rect 313016 219406 313136 219434
rect 312360 218068 312412 218074
rect 312360 218010 312412 218016
rect 309842 217110 309916 217138
rect 310670 217110 310744 217138
rect 311498 217246 311572 217274
rect 309842 216988 309870 217110
rect 310670 216988 310698 217110
rect 311498 216988 311526 217246
rect 312372 217138 312400 218010
rect 313108 217274 313136 219406
rect 313200 218090 313228 229570
rect 313476 218210 313504 230318
rect 313660 221474 313688 231676
rect 313936 231662 314226 231690
rect 313936 230382 313964 231662
rect 313924 230376 313976 230382
rect 313924 230318 313976 230324
rect 313924 230240 313976 230246
rect 313924 230182 313976 230188
rect 313648 221468 313700 221474
rect 313648 221410 313700 221416
rect 313936 219434 313964 230182
rect 314764 227050 314792 231676
rect 315316 230246 315344 231676
rect 315500 231662 315882 231690
rect 315304 230240 315356 230246
rect 315304 230182 315356 230188
rect 315500 227798 315528 231662
rect 315672 228676 315724 228682
rect 315672 228618 315724 228624
rect 315488 227792 315540 227798
rect 315488 227734 315540 227740
rect 314752 227044 314804 227050
rect 314752 226986 314804 226992
rect 315684 222194 315712 228618
rect 316420 227934 316448 231676
rect 316696 231662 316986 231690
rect 316408 227928 316460 227934
rect 316408 227870 316460 227876
rect 316696 224262 316724 231662
rect 317052 227792 317104 227798
rect 317052 227734 317104 227740
rect 316684 224256 316736 224262
rect 316684 224198 316736 224204
rect 313844 219406 313964 219434
rect 315592 222166 315712 222194
rect 313844 218890 313872 219406
rect 314016 219020 314068 219026
rect 314016 218962 314068 218968
rect 313832 218884 313884 218890
rect 313832 218826 313884 218832
rect 313464 218204 313516 218210
rect 313464 218146 313516 218152
rect 313200 218074 313320 218090
rect 313200 218068 313332 218074
rect 313200 218062 313280 218068
rect 313280 218010 313332 218016
rect 313108 217246 313182 217274
rect 312326 217110 312400 217138
rect 312326 216988 312354 217110
rect 313154 216988 313182 217246
rect 314028 217138 314056 218962
rect 315592 218074 315620 222166
rect 315764 221468 315816 221474
rect 315764 221410 315816 221416
rect 314844 218068 314896 218074
rect 314844 218010 314896 218016
rect 315580 218068 315632 218074
rect 315580 218010 315632 218016
rect 314856 217138 314884 218010
rect 315776 217274 315804 221410
rect 317064 218074 317092 227734
rect 317524 225622 317552 231676
rect 317708 231662 318090 231690
rect 318260 231662 318642 231690
rect 318812 231662 319194 231690
rect 317512 225616 317564 225622
rect 317512 225558 317564 225564
rect 317236 223780 317288 223786
rect 317236 223722 317288 223728
rect 316500 218068 316552 218074
rect 316500 218010 316552 218016
rect 317052 218068 317104 218074
rect 317052 218010 317104 218016
rect 313982 217110 314056 217138
rect 314810 217110 314884 217138
rect 315638 217246 315804 217274
rect 313982 216988 314010 217110
rect 314810 216988 314838 217110
rect 315638 216988 315666 217246
rect 316512 217138 316540 218010
rect 317248 217274 317276 223722
rect 317420 221672 317472 221678
rect 317420 221614 317472 221620
rect 317432 218754 317460 221614
rect 317708 219502 317736 231662
rect 318260 220862 318288 231662
rect 318812 221678 318840 231662
rect 319444 230376 319496 230382
rect 319444 230318 319496 230324
rect 318800 221672 318852 221678
rect 318800 221614 318852 221620
rect 318248 220856 318300 220862
rect 318248 220798 318300 220804
rect 318156 220720 318208 220726
rect 318156 220662 318208 220668
rect 317696 219496 317748 219502
rect 317696 219438 317748 219444
rect 317420 218748 317472 218754
rect 317420 218690 317472 218696
rect 318168 217274 318196 220662
rect 319456 219026 319484 230318
rect 319732 229634 319760 231676
rect 319720 229628 319772 229634
rect 319720 229570 319772 229576
rect 320284 228682 320312 231676
rect 320560 231662 320850 231690
rect 320272 228676 320324 228682
rect 320272 228618 320324 228624
rect 320560 227798 320588 231662
rect 321388 230382 321416 231676
rect 321376 230376 321428 230382
rect 321376 230318 321428 230324
rect 321940 230110 321968 231676
rect 322216 231662 322506 231690
rect 320824 230104 320876 230110
rect 320824 230046 320876 230052
rect 321928 230104 321980 230110
rect 321928 230046 321980 230052
rect 320548 227792 320600 227798
rect 320548 227734 320600 227740
rect 320836 221474 320864 230046
rect 321468 227792 321520 227798
rect 321468 227734 321520 227740
rect 320824 221468 320876 221474
rect 320824 221410 320876 221416
rect 320640 220856 320692 220862
rect 320640 220798 320692 220804
rect 319812 219428 319864 219434
rect 319812 219370 319864 219376
rect 319444 219020 319496 219026
rect 319444 218962 319496 218968
rect 318984 218204 319036 218210
rect 318984 218146 319036 218152
rect 317248 217246 317322 217274
rect 316466 217110 316540 217138
rect 316466 216988 316494 217110
rect 317294 216988 317322 217246
rect 318122 217246 318196 217274
rect 318122 216988 318150 217246
rect 318996 217138 319024 218146
rect 319824 217138 319852 219370
rect 320652 217274 320680 220798
rect 321480 217274 321508 227734
rect 322216 220726 322244 231662
rect 322756 229152 322808 229158
rect 322756 229094 322808 229100
rect 322204 220720 322256 220726
rect 322204 220662 322256 220668
rect 322768 218074 322796 229094
rect 323044 219502 323072 231676
rect 323596 223786 323624 231676
rect 323872 231662 324162 231690
rect 323584 223780 323636 223786
rect 323584 223722 323636 223728
rect 323032 219496 323084 219502
rect 323032 219438 323084 219444
rect 323872 219434 323900 231662
rect 324700 227798 324728 231676
rect 324976 231662 325266 231690
rect 324688 227792 324740 227798
rect 324688 227734 324740 227740
rect 324044 219496 324096 219502
rect 323320 219406 323900 219434
rect 323964 219444 324044 219450
rect 323964 219438 324096 219444
rect 323964 219422 324084 219438
rect 324976 219434 325004 231662
rect 325608 228540 325660 228546
rect 325608 228482 325660 228488
rect 323124 218748 323176 218754
rect 323124 218690 323176 218696
rect 322296 218068 322348 218074
rect 322296 218010 322348 218016
rect 322756 218068 322808 218074
rect 322756 218010 322808 218016
rect 318950 217110 319024 217138
rect 319778 217110 319852 217138
rect 320606 217246 320680 217274
rect 321434 217246 321508 217274
rect 318950 216988 318978 217110
rect 319778 216988 319806 217110
rect 320606 216988 320634 217246
rect 321434 216988 321462 217246
rect 322308 217138 322336 218010
rect 323136 217274 323164 218690
rect 323320 218210 323348 219406
rect 323308 218204 323360 218210
rect 323308 218146 323360 218152
rect 323964 217274 323992 219422
rect 324700 219406 325004 219434
rect 324700 218754 324728 219406
rect 324688 218748 324740 218754
rect 324688 218690 324740 218696
rect 324780 218612 324832 218618
rect 324780 218554 324832 218560
rect 322262 217110 322336 217138
rect 323090 217246 323164 217274
rect 323918 217246 323992 217274
rect 322262 216988 322290 217110
rect 323090 216988 323118 217246
rect 323918 216988 323946 217246
rect 324792 217138 324820 218554
rect 325620 217274 325648 228482
rect 325804 220862 325832 231676
rect 326356 229158 326384 231676
rect 326632 231662 326922 231690
rect 327474 231662 327672 231690
rect 326344 229152 326396 229158
rect 326344 229094 326396 229100
rect 325792 220856 325844 220862
rect 325792 220798 325844 220804
rect 326632 219434 326660 231662
rect 326080 219406 326660 219434
rect 326080 218618 326108 219406
rect 326068 218612 326120 218618
rect 326068 218554 326120 218560
rect 327264 218204 327316 218210
rect 327264 218146 327316 218152
rect 326436 218068 326488 218074
rect 326436 218010 326488 218016
rect 324746 217110 324820 217138
rect 325574 217246 325648 217274
rect 324746 216988 324774 217110
rect 325574 216988 325602 217246
rect 326448 217138 326476 218010
rect 327276 217138 327304 218146
rect 327644 218074 327672 231662
rect 327828 231662 328026 231690
rect 328472 231662 328578 231690
rect 328748 231662 329130 231690
rect 327828 219502 327856 231662
rect 328472 228562 328500 231662
rect 328748 230466 328776 231662
rect 328380 228546 328500 228562
rect 328368 228540 328500 228546
rect 328420 228534 328500 228540
rect 328564 230438 328776 230466
rect 328368 228482 328420 228488
rect 327816 219496 327868 219502
rect 327816 219438 327868 219444
rect 328564 218074 328592 230438
rect 329668 230382 329696 231676
rect 329944 231662 330234 231690
rect 330404 231662 330786 231690
rect 331338 231662 331628 231690
rect 328828 230376 328880 230382
rect 328828 230318 328880 230324
rect 329656 230376 329708 230382
rect 329656 230318 329708 230324
rect 328840 229094 328868 230318
rect 328840 229066 329696 229094
rect 327632 218068 327684 218074
rect 327632 218010 327684 218016
rect 328092 218068 328144 218074
rect 328092 218010 328144 218016
rect 328552 218068 328604 218074
rect 328552 218010 328604 218016
rect 328920 218068 328972 218074
rect 328920 218010 328972 218016
rect 328104 217138 328132 218010
rect 328932 217138 328960 218010
rect 329668 217274 329696 229066
rect 329944 218210 329972 231662
rect 330404 219434 330432 231662
rect 331220 224256 331272 224262
rect 331220 224198 331272 224204
rect 330128 219406 330432 219434
rect 329932 218204 329984 218210
rect 329932 218146 329984 218152
rect 330128 218074 330156 219406
rect 331232 218074 331260 224198
rect 331600 219434 331628 231662
rect 331876 230382 331904 231676
rect 332152 231662 332442 231690
rect 332704 231662 332994 231690
rect 331864 230376 331916 230382
rect 331864 230318 331916 230324
rect 332152 224262 332180 231662
rect 332140 224256 332192 224262
rect 332140 224198 332192 224204
rect 331416 219406 331628 219434
rect 330116 218068 330168 218074
rect 330116 218010 330168 218016
rect 330576 218068 330628 218074
rect 330576 218010 330628 218016
rect 331220 218068 331272 218074
rect 331220 218010 331272 218016
rect 329668 217246 329742 217274
rect 326402 217110 326476 217138
rect 327230 217110 327304 217138
rect 328058 217110 328132 217138
rect 328886 217110 328960 217138
rect 326402 216988 326430 217110
rect 327230 216988 327258 217110
rect 328058 216988 328086 217110
rect 328886 216988 328914 217110
rect 329714 216988 329742 217246
rect 330588 217138 330616 218010
rect 331416 217274 331444 219406
rect 332704 218074 332732 231662
rect 333532 230382 333560 231676
rect 333060 230376 333112 230382
rect 333060 230318 333112 230324
rect 333520 230376 333572 230382
rect 333520 230318 333572 230324
rect 332232 218068 332284 218074
rect 332232 218010 332284 218016
rect 332692 218068 332744 218074
rect 332692 218010 332744 218016
rect 330542 217110 330616 217138
rect 331370 217246 331444 217274
rect 330542 216988 330570 217110
rect 331370 216988 331398 217246
rect 332244 217138 332272 218010
rect 333072 217274 333100 230318
rect 334084 229294 334112 231676
rect 334360 231662 334650 231690
rect 334072 229288 334124 229294
rect 334072 229230 334124 229236
rect 334360 219434 334388 231662
rect 334532 230376 334584 230382
rect 334532 230318 334584 230324
rect 334544 229094 334572 230318
rect 335188 229158 335216 231676
rect 335740 230382 335768 231676
rect 336306 231662 336596 231690
rect 335728 230376 335780 230382
rect 335728 230318 335780 230324
rect 335728 229288 335780 229294
rect 335728 229230 335780 229236
rect 335176 229152 335228 229158
rect 335176 229094 335228 229100
rect 334544 229066 334664 229094
rect 333900 219406 334388 219434
rect 333900 217274 333928 219406
rect 332198 217110 332272 217138
rect 333026 217246 333100 217274
rect 333854 217246 333928 217274
rect 334636 217274 334664 229066
rect 335740 224262 335768 229230
rect 335912 229152 335964 229158
rect 335912 229094 335964 229100
rect 335728 224256 335780 224262
rect 335728 224198 335780 224204
rect 335924 219434 335952 229094
rect 336280 224256 336332 224262
rect 336280 224198 336332 224204
rect 335556 219406 335952 219434
rect 335556 217274 335584 219406
rect 334636 217246 334710 217274
rect 332198 216988 332226 217110
rect 333026 216988 333054 217246
rect 333854 216988 333882 217246
rect 334682 216988 334710 217246
rect 335510 217246 335584 217274
rect 336292 217274 336320 224198
rect 336568 218074 336596 231662
rect 336844 229094 336872 231676
rect 337396 230382 337424 231676
rect 337200 230376 337252 230382
rect 337200 230318 337252 230324
rect 337384 230376 337436 230382
rect 337384 230318 337436 230324
rect 336844 229066 337148 229094
rect 336556 218068 336608 218074
rect 336556 218010 336608 218016
rect 337120 217274 337148 229066
rect 337212 219434 337240 230318
rect 337948 220794 337976 231676
rect 338304 230376 338356 230382
rect 338304 230318 338356 230324
rect 338316 229094 338344 230318
rect 338500 229906 338528 231676
rect 339052 230314 339080 231676
rect 339604 230450 339632 231676
rect 340170 231662 340552 231690
rect 339592 230444 339644 230450
rect 339592 230386 339644 230392
rect 339040 230308 339092 230314
rect 339040 230250 339092 230256
rect 339868 230308 339920 230314
rect 339868 230250 339920 230256
rect 338488 229900 338540 229906
rect 338488 229842 338540 229848
rect 339316 229900 339368 229906
rect 339316 229842 339368 229848
rect 338316 229066 338804 229094
rect 337936 220788 337988 220794
rect 337936 220730 337988 220736
rect 337212 219406 337976 219434
rect 337948 217274 337976 219406
rect 338776 217274 338804 229066
rect 339328 218210 339356 229842
rect 339880 229094 339908 230250
rect 340524 229094 340552 231662
rect 340708 230110 340736 231676
rect 341064 230444 341116 230450
rect 341064 230386 341116 230392
rect 340696 230104 340748 230110
rect 340696 230046 340748 230052
rect 341076 229094 341104 230386
rect 341260 230246 341288 231676
rect 341826 231662 342208 231690
rect 341248 230240 341300 230246
rect 341248 230182 341300 230188
rect 339880 229066 340460 229094
rect 340524 229066 340644 229094
rect 341076 229066 342116 229094
rect 339316 218204 339368 218210
rect 339316 218146 339368 218152
rect 339592 218068 339644 218074
rect 339592 218010 339644 218016
rect 336292 217246 336366 217274
rect 337120 217246 337194 217274
rect 337948 217246 338022 217274
rect 338776 217246 338850 217274
rect 335510 216988 335538 217246
rect 336338 216988 336366 217246
rect 337166 216988 337194 217246
rect 337994 216988 338022 217246
rect 338822 216988 338850 217246
rect 339604 217138 339632 218010
rect 340432 217274 340460 229066
rect 340616 220658 340644 229066
rect 341248 220788 341300 220794
rect 341248 220730 341300 220736
rect 340604 220652 340656 220658
rect 340604 220594 340656 220600
rect 341260 217274 341288 220730
rect 342088 217274 342116 229066
rect 342180 222170 342208 231662
rect 342364 230382 342392 231676
rect 342352 230376 342404 230382
rect 342352 230318 342404 230324
rect 342916 229770 342944 231676
rect 343272 230376 343324 230382
rect 343272 230318 343324 230324
rect 342904 229764 342956 229770
rect 342904 229706 342956 229712
rect 342180 222142 342300 222170
rect 342272 219298 342300 222142
rect 343284 220250 343312 230318
rect 343468 220930 343496 231676
rect 344020 230382 344048 231676
rect 344008 230376 344060 230382
rect 344008 230318 344060 230324
rect 343824 230240 343876 230246
rect 343824 230182 343876 230188
rect 343456 220924 343508 220930
rect 343456 220866 343508 220872
rect 343272 220244 343324 220250
rect 343272 220186 343324 220192
rect 342260 219292 342312 219298
rect 342260 219234 342312 219240
rect 342904 218204 342956 218210
rect 342904 218146 342956 218152
rect 340432 217246 340506 217274
rect 341260 217246 341334 217274
rect 342088 217246 342162 217274
rect 339604 217110 339678 217138
rect 339650 216988 339678 217110
rect 340478 216988 340506 217246
rect 341306 216988 341334 217246
rect 342134 216988 342162 217246
rect 342916 217138 342944 218146
rect 343836 217274 343864 230182
rect 344572 230178 344600 231676
rect 344928 230376 344980 230382
rect 344928 230318 344980 230324
rect 344560 230172 344612 230178
rect 344560 230114 344612 230120
rect 344284 230104 344336 230110
rect 344284 230046 344336 230052
rect 344296 219502 344324 230046
rect 344940 221610 344968 230318
rect 345124 227798 345152 231676
rect 345690 231662 345888 231690
rect 345112 227792 345164 227798
rect 345112 227734 345164 227740
rect 344928 221604 344980 221610
rect 344928 221546 344980 221552
rect 345860 220794 345888 231662
rect 346044 231662 346242 231690
rect 346794 231662 347268 231690
rect 347346 231662 347636 231690
rect 345848 220788 345900 220794
rect 345848 220730 345900 220736
rect 344560 220652 344612 220658
rect 344560 220594 344612 220600
rect 344284 219496 344336 219502
rect 344284 219438 344336 219444
rect 343790 217246 343864 217274
rect 344572 217274 344600 220594
rect 345388 219292 345440 219298
rect 345388 219234 345440 219240
rect 344572 217246 344646 217274
rect 342916 217110 342990 217138
rect 342962 216988 342990 217110
rect 343790 216988 343818 217246
rect 344618 216988 344646 217246
rect 345400 217138 345428 219234
rect 346044 218210 346072 231662
rect 347044 220924 347096 220930
rect 347044 220866 347096 220872
rect 346400 220788 346452 220794
rect 346400 220730 346452 220736
rect 346216 219496 346268 219502
rect 346216 219438 346268 219444
rect 346032 218204 346084 218210
rect 346032 218146 346084 218152
rect 346228 217274 346256 219438
rect 346412 218074 346440 220730
rect 346400 218068 346452 218074
rect 346400 218010 346452 218016
rect 347056 217274 347084 220866
rect 347240 220658 347268 231662
rect 347608 221474 347636 231662
rect 347884 223582 347912 231676
rect 348450 231662 348832 231690
rect 348424 229764 348476 229770
rect 348424 229706 348476 229712
rect 347872 223576 347924 223582
rect 347872 223518 347924 223524
rect 347596 221468 347648 221474
rect 347596 221410 347648 221416
rect 348436 220794 348464 229706
rect 348804 222170 348832 231662
rect 348988 230382 349016 231676
rect 348976 230376 349028 230382
rect 348976 230318 349028 230324
rect 349540 228682 349568 231676
rect 350106 231662 350304 231690
rect 349804 230172 349856 230178
rect 349804 230114 349856 230120
rect 349528 228676 349580 228682
rect 349528 228618 349580 228624
rect 348804 222142 349200 222170
rect 348700 221604 348752 221610
rect 348700 221546 348752 221552
rect 348424 220788 348476 220794
rect 348424 220730 348476 220736
rect 347228 220652 347280 220658
rect 347228 220594 347280 220600
rect 347872 220244 347924 220250
rect 347872 220186 347924 220192
rect 347884 217274 347912 220186
rect 348712 217274 348740 221546
rect 349172 218618 349200 222142
rect 349816 220794 349844 230114
rect 349528 220788 349580 220794
rect 349528 220730 349580 220736
rect 349804 220788 349856 220794
rect 349804 220730 349856 220736
rect 349160 218612 349212 218618
rect 349160 218554 349212 218560
rect 349540 217274 349568 220730
rect 350276 219638 350304 231662
rect 350644 229294 350672 231676
rect 351210 231662 351684 231690
rect 350632 229288 350684 229294
rect 350632 229230 350684 229236
rect 351656 229094 351684 231662
rect 351564 229066 351684 229094
rect 351564 221882 351592 229066
rect 351748 227050 351776 231676
rect 351736 227044 351788 227050
rect 351736 226986 351788 226992
rect 352300 224262 352328 231676
rect 352564 230376 352616 230382
rect 352564 230318 352616 230324
rect 352288 224256 352340 224262
rect 352288 224198 352340 224204
rect 351552 221876 351604 221882
rect 351552 221818 351604 221824
rect 351184 220788 351236 220794
rect 351184 220730 351236 220736
rect 350264 219632 350316 219638
rect 350264 219574 350316 219580
rect 350356 218068 350408 218074
rect 350356 218010 350408 218016
rect 346228 217246 346302 217274
rect 347056 217246 347130 217274
rect 347884 217246 347958 217274
rect 348712 217246 348786 217274
rect 349540 217246 349614 217274
rect 345400 217110 345474 217138
rect 345446 216988 345474 217110
rect 346274 216988 346302 217246
rect 347102 216988 347130 217246
rect 347930 216988 347958 217246
rect 348758 216988 348786 217246
rect 349586 216988 349614 217246
rect 350368 217138 350396 218010
rect 351196 217274 351224 220730
rect 352576 220522 352604 230318
rect 352852 228818 352880 231676
rect 352840 228812 352892 228818
rect 352840 228754 352892 228760
rect 353404 228546 353432 231676
rect 353392 228540 353444 228546
rect 353392 228482 353444 228488
rect 352840 227792 352892 227798
rect 352840 227734 352892 227740
rect 352564 220516 352616 220522
rect 352564 220458 352616 220464
rect 352012 218204 352064 218210
rect 352012 218146 352064 218152
rect 351196 217246 351270 217274
rect 350368 217110 350442 217138
rect 350414 216988 350442 217110
rect 351242 216988 351270 217246
rect 352024 217138 352052 218146
rect 352852 217274 352880 227734
rect 353668 223576 353720 223582
rect 353668 223518 353720 223524
rect 353680 217274 353708 223518
rect 353956 223038 353984 231676
rect 354508 229094 354536 231676
rect 355060 230246 355088 231676
rect 355626 231662 356008 231690
rect 355048 230240 355100 230246
rect 355048 230182 355100 230188
rect 355324 229288 355376 229294
rect 355324 229230 355376 229236
rect 354324 229066 354536 229094
rect 353944 223032 353996 223038
rect 353944 222974 353996 222980
rect 354324 220386 354352 229066
rect 354496 220652 354548 220658
rect 354496 220594 354548 220600
rect 354312 220380 354364 220386
rect 354312 220322 354364 220328
rect 354508 217274 354536 220594
rect 355336 218754 355364 229230
rect 355980 220114 356008 231662
rect 356164 230382 356192 231676
rect 356730 231662 357112 231690
rect 356152 230376 356204 230382
rect 356152 230318 356204 230324
rect 357084 229094 357112 231662
rect 357268 230466 357296 231676
rect 357834 231662 358216 231690
rect 357268 230438 357480 230466
rect 357256 230376 357308 230382
rect 357256 230318 357308 230324
rect 357268 229094 357296 230318
rect 357452 230110 357480 230438
rect 357440 230104 357492 230110
rect 357440 230046 357492 230052
rect 358188 229094 358216 231662
rect 358372 229094 358400 231676
rect 358938 231662 359320 231690
rect 357084 229066 357204 229094
rect 357268 229066 357388 229094
rect 358188 229066 358308 229094
rect 358372 229066 358492 229094
rect 356152 221468 356204 221474
rect 356152 221410 356204 221416
rect 355968 220108 356020 220114
rect 355968 220050 356020 220056
rect 355324 218748 355376 218754
rect 355324 218690 355376 218696
rect 355324 218612 355376 218618
rect 355324 218554 355376 218560
rect 352852 217246 352926 217274
rect 353680 217246 353754 217274
rect 354508 217246 354582 217274
rect 352024 217110 352098 217138
rect 352070 216988 352098 217110
rect 352898 216988 352926 217246
rect 353726 216988 353754 217246
rect 354554 216988 354582 217246
rect 355336 217138 355364 218554
rect 356164 217274 356192 221410
rect 356980 219360 357032 219366
rect 356980 219302 357032 219308
rect 356164 217246 356238 217274
rect 355336 217110 355410 217138
rect 355382 216988 355410 217110
rect 356210 216988 356238 217246
rect 356992 217138 357020 219302
rect 357176 218618 357204 229066
rect 357360 221746 357388 229066
rect 358084 224256 358136 224262
rect 358084 224198 358136 224204
rect 357348 221740 357400 221746
rect 357348 221682 357400 221688
rect 357808 220516 357860 220522
rect 357808 220458 357860 220464
rect 357164 218612 357216 218618
rect 357164 218554 357216 218560
rect 357820 217274 357848 220458
rect 358096 218074 358124 224198
rect 358280 220250 358308 229066
rect 358464 224398 358492 229066
rect 359292 225622 359320 231662
rect 359476 229906 359504 231676
rect 359464 229900 359516 229906
rect 359464 229842 359516 229848
rect 359464 228676 359516 228682
rect 359464 228618 359516 228624
rect 359280 225616 359332 225622
rect 359280 225558 359332 225564
rect 358452 224392 358504 224398
rect 358452 224334 358504 224340
rect 358268 220244 358320 220250
rect 358268 220186 358320 220192
rect 358636 218748 358688 218754
rect 358636 218690 358688 218696
rect 358084 218068 358136 218074
rect 358084 218010 358136 218016
rect 357820 217246 357894 217274
rect 356992 217110 357066 217138
rect 357038 216988 357066 217110
rect 357866 216988 357894 217246
rect 358648 217138 358676 218690
rect 359476 217274 359504 228618
rect 360028 221610 360056 231676
rect 360580 230382 360608 231676
rect 360568 230376 360620 230382
rect 360568 230318 360620 230324
rect 360844 230240 360896 230246
rect 360844 230182 360896 230188
rect 360016 221604 360068 221610
rect 360016 221546 360068 221552
rect 360856 218754 360884 230182
rect 361132 229090 361160 231676
rect 361684 229770 361712 231676
rect 361672 229764 361724 229770
rect 361672 229706 361724 229712
rect 361120 229084 361172 229090
rect 361120 229026 361172 229032
rect 362236 228818 362264 231676
rect 362788 230466 362816 231676
rect 362788 230438 362908 230466
rect 362684 230376 362736 230382
rect 362684 230318 362736 230324
rect 361028 228812 361080 228818
rect 361028 228754 361080 228760
rect 362224 228812 362276 228818
rect 362224 228754 362276 228760
rect 360844 218748 360896 218754
rect 360844 218690 360896 218696
rect 361040 218210 361068 228754
rect 361580 227044 361632 227050
rect 361580 226986 361632 226992
rect 361212 221876 361264 221882
rect 361212 221818 361264 221824
rect 361028 218204 361080 218210
rect 361028 218146 361080 218152
rect 360292 218068 360344 218074
rect 360292 218010 360344 218016
rect 359476 217246 359550 217274
rect 358648 217110 358722 217138
rect 358694 216988 358722 217110
rect 359522 216988 359550 217246
rect 360304 217138 360332 218010
rect 361224 217274 361252 221818
rect 361178 217246 361252 217274
rect 361592 217258 361620 226986
rect 362696 222902 362724 230318
rect 362684 222896 362736 222902
rect 362684 222838 362736 222844
rect 362880 220522 362908 230438
rect 363340 225758 363368 231676
rect 363604 230104 363656 230110
rect 363604 230046 363656 230052
rect 363328 225752 363380 225758
rect 363328 225694 363380 225700
rect 362868 220516 362920 220522
rect 362868 220458 362920 220464
rect 361764 220380 361816 220386
rect 361764 220322 361816 220328
rect 361776 218074 361804 220322
rect 363616 219026 363644 230046
rect 363892 227186 363920 231676
rect 364444 230382 364472 231676
rect 364432 230376 364484 230382
rect 364432 230318 364484 230324
rect 364996 228546 365024 231676
rect 365548 230466 365576 231676
rect 366114 231662 366496 231690
rect 365548 230438 365760 230466
rect 365444 230376 365496 230382
rect 365444 230318 365496 230324
rect 364432 228540 364484 228546
rect 364432 228482 364484 228488
rect 364984 228540 365036 228546
rect 364984 228482 365036 228488
rect 363880 227180 363932 227186
rect 363880 227122 363932 227128
rect 363604 219020 363656 219026
rect 363604 218962 363656 218968
rect 361948 218204 362000 218210
rect 361948 218146 362000 218152
rect 361764 218068 361816 218074
rect 361764 218010 361816 218016
rect 361580 217252 361632 217258
rect 360304 217110 360378 217138
rect 360350 216988 360378 217110
rect 361178 216988 361206 217246
rect 361580 217194 361632 217200
rect 361960 217138 361988 218146
rect 363604 218068 363656 218074
rect 363604 218010 363656 218016
rect 362822 217252 362874 217258
rect 362822 217194 362874 217200
rect 361960 217110 362034 217138
rect 362006 216988 362034 217110
rect 362834 216988 362862 217194
rect 363616 217138 363644 218010
rect 364444 217274 364472 228482
rect 365456 220386 365484 230318
rect 365732 223174 365760 230438
rect 365720 223168 365772 223174
rect 365720 223110 365772 223116
rect 366088 223032 366140 223038
rect 366088 222974 366140 222980
rect 365444 220380 365496 220386
rect 365444 220322 365496 220328
rect 365260 218748 365312 218754
rect 365260 218690 365312 218696
rect 364444 217246 364518 217274
rect 363616 217110 363690 217138
rect 363662 216988 363690 217110
rect 364490 216988 364518 217246
rect 365272 217138 365300 218690
rect 366100 217274 366128 222974
rect 366468 219434 366496 231662
rect 366652 227050 366680 231676
rect 367204 230382 367232 231676
rect 367192 230376 367244 230382
rect 367192 230318 367244 230324
rect 367756 230042 367784 231676
rect 368124 231662 368322 231690
rect 367744 230036 367796 230042
rect 367744 229978 367796 229984
rect 366640 227044 366692 227050
rect 366640 226986 366692 226992
rect 367744 220108 367796 220114
rect 367744 220050 367796 220056
rect 366468 219406 366772 219434
rect 366744 218890 366772 219406
rect 366732 218884 366784 218890
rect 366732 218826 366784 218832
rect 366916 218612 366968 218618
rect 366916 218554 366968 218560
rect 366100 217246 366174 217274
rect 365272 217110 365346 217138
rect 365318 216988 365346 217110
rect 366146 216988 366174 217246
rect 366928 217138 366956 218554
rect 367756 217274 367784 220050
rect 368124 218754 368152 231662
rect 368860 230382 368888 231676
rect 368296 230376 368348 230382
rect 368296 230318 368348 230324
rect 368848 230376 368900 230382
rect 368848 230318 368900 230324
rect 368308 221474 368336 230318
rect 369412 230178 369440 231676
rect 369978 231662 370360 231690
rect 369768 230376 369820 230382
rect 369768 230318 369820 230324
rect 369400 230172 369452 230178
rect 369400 230114 369452 230120
rect 369124 229900 369176 229906
rect 369124 229842 369176 229848
rect 368296 221468 368348 221474
rect 368296 221410 368348 221416
rect 369136 220794 369164 229842
rect 369780 222018 369808 230318
rect 370332 228562 370360 231662
rect 370516 228682 370544 231676
rect 371068 230382 371096 231676
rect 371056 230376 371108 230382
rect 371056 230318 371108 230324
rect 370872 230036 370924 230042
rect 370872 229978 370924 229984
rect 370504 228676 370556 228682
rect 370504 228618 370556 228624
rect 370332 228534 370452 228562
rect 370228 225616 370280 225622
rect 370228 225558 370280 225564
rect 369768 222012 369820 222018
rect 369768 221954 369820 221960
rect 369400 221740 369452 221746
rect 369400 221682 369452 221688
rect 369124 220788 369176 220794
rect 369124 220730 369176 220736
rect 368572 219020 368624 219026
rect 368572 218962 368624 218968
rect 368112 218748 368164 218754
rect 368112 218690 368164 218696
rect 367756 217246 367830 217274
rect 366928 217110 367002 217138
rect 366974 216988 367002 217110
rect 367802 216988 367830 217246
rect 368584 217138 368612 218962
rect 369412 217274 369440 221682
rect 370240 217274 370268 225558
rect 370424 224262 370452 228534
rect 370884 224534 370912 229978
rect 371620 225622 371648 231676
rect 372186 231662 372568 231690
rect 372068 230376 372120 230382
rect 372068 230318 372120 230324
rect 371884 230172 371936 230178
rect 371884 230114 371936 230120
rect 371608 225616 371660 225622
rect 371608 225558 371660 225564
rect 370872 224528 370924 224534
rect 370872 224470 370924 224476
rect 370412 224256 370464 224262
rect 370412 224198 370464 224204
rect 371896 221762 371924 230114
rect 372080 221882 372108 230318
rect 372540 229430 372568 231662
rect 372724 230178 372752 231676
rect 372712 230172 372764 230178
rect 372712 230114 372764 230120
rect 372528 229424 372580 229430
rect 372528 229366 372580 229372
rect 373276 228954 373304 231676
rect 373736 231662 373842 231690
rect 373540 229084 373592 229090
rect 373540 229026 373592 229032
rect 373264 228948 373316 228954
rect 373264 228890 373316 228896
rect 372712 224392 372764 224398
rect 372712 224334 372764 224340
rect 372068 221876 372120 221882
rect 372068 221818 372120 221824
rect 371896 221734 372108 221762
rect 371884 220788 371936 220794
rect 371884 220730 371936 220736
rect 371056 220244 371108 220250
rect 371056 220186 371108 220192
rect 371068 217274 371096 220186
rect 371896 217274 371924 220730
rect 372080 220250 372108 221734
rect 372068 220244 372120 220250
rect 372068 220186 372120 220192
rect 372724 217274 372752 224334
rect 373552 217274 373580 229026
rect 373736 220114 373764 231662
rect 374380 230042 374408 231676
rect 374368 230036 374420 230042
rect 374368 229978 374420 229984
rect 374000 229764 374052 229770
rect 374000 229706 374052 229712
rect 373724 220108 373776 220114
rect 373724 220050 373776 220056
rect 369412 217246 369486 217274
rect 370240 217246 370314 217274
rect 371068 217246 371142 217274
rect 371896 217246 371970 217274
rect 372724 217246 372798 217274
rect 373552 217246 373626 217274
rect 374012 217258 374040 229706
rect 374932 229634 374960 231676
rect 374920 229628 374972 229634
rect 374920 229570 374972 229576
rect 374552 229424 374604 229430
rect 374552 229366 374604 229372
rect 374564 227458 374592 229366
rect 374552 227452 374604 227458
rect 374552 227394 374604 227400
rect 374644 227180 374696 227186
rect 374644 227122 374696 227128
rect 374368 221604 374420 221610
rect 374368 221546 374420 221552
rect 374380 217274 374408 221546
rect 374656 218074 374684 227122
rect 375484 223310 375512 231676
rect 375472 223304 375524 223310
rect 375472 223246 375524 223252
rect 376036 223038 376064 231676
rect 376392 228540 376444 228546
rect 376392 228482 376444 228488
rect 376404 228274 376432 228482
rect 376392 228268 376444 228274
rect 376392 228210 376444 228216
rect 376588 227322 376616 231676
rect 377140 229770 377168 231676
rect 377404 230036 377456 230042
rect 377404 229978 377456 229984
rect 377128 229764 377180 229770
rect 377128 229706 377180 229712
rect 376760 228812 376812 228818
rect 376760 228754 376812 228760
rect 376772 228546 376800 228754
rect 376760 228540 376812 228546
rect 376760 228482 376812 228488
rect 376576 227316 376628 227322
rect 376576 227258 376628 227264
rect 376852 225752 376904 225758
rect 376852 225694 376904 225700
rect 376024 223032 376076 223038
rect 376024 222974 376076 222980
rect 376024 222896 376076 222902
rect 376024 222838 376076 222844
rect 374644 218068 374696 218074
rect 374644 218010 374696 218016
rect 376036 217274 376064 222838
rect 376864 217274 376892 225694
rect 377416 222154 377444 229978
rect 377692 228818 377720 231676
rect 378244 230382 378272 231676
rect 378232 230376 378284 230382
rect 378232 230318 378284 230324
rect 378796 230246 378824 231676
rect 379164 231662 379362 231690
rect 378784 230240 378836 230246
rect 378784 230182 378836 230188
rect 379164 230042 379192 231662
rect 379336 230376 379388 230382
rect 379336 230318 379388 230324
rect 379152 230036 379204 230042
rect 379152 229978 379204 229984
rect 377680 228812 377732 228818
rect 377680 228754 377732 228760
rect 377680 228540 377732 228546
rect 377680 228482 377732 228488
rect 377404 222148 377456 222154
rect 377404 222090 377456 222096
rect 377692 217274 377720 228482
rect 379348 220794 379376 230318
rect 379900 224670 379928 231676
rect 380164 230240 380216 230246
rect 380164 230182 380216 230188
rect 379888 224664 379940 224670
rect 379888 224606 379940 224612
rect 380176 224482 380204 230182
rect 379992 224454 380204 224482
rect 379992 221746 380020 224454
rect 380164 223168 380216 223174
rect 380164 223110 380216 223116
rect 379980 221740 380032 221746
rect 379980 221682 380032 221688
rect 379336 220788 379388 220794
rect 379336 220730 379388 220736
rect 379336 220516 379388 220522
rect 379336 220458 379388 220464
rect 378508 218068 378560 218074
rect 378508 218010 378560 218016
rect 368584 217110 368658 217138
rect 368630 216988 368658 217110
rect 369458 216988 369486 217246
rect 370286 216988 370314 217246
rect 371114 216988 371142 217246
rect 371942 216988 371970 217246
rect 372770 216988 372798 217246
rect 373598 216988 373626 217246
rect 374000 217252 374052 217258
rect 374380 217246 374454 217274
rect 374000 217194 374052 217200
rect 374426 216988 374454 217246
rect 375242 217252 375294 217258
rect 376036 217246 376110 217274
rect 376864 217246 376938 217274
rect 377692 217246 377766 217274
rect 375242 217194 375294 217200
rect 375254 216988 375282 217194
rect 376082 216988 376110 217246
rect 376910 216988 376938 217246
rect 377738 216988 377766 217246
rect 378520 217138 378548 218010
rect 379348 217274 379376 220458
rect 380176 217274 380204 223110
rect 380452 222902 380480 231676
rect 381004 230246 381032 231676
rect 381570 231662 381952 231690
rect 380992 230240 381044 230246
rect 380992 230182 381044 230188
rect 380440 222896 380492 222902
rect 380440 222838 380492 222844
rect 380992 220380 381044 220386
rect 380992 220322 381044 220328
rect 381004 217274 381032 220322
rect 381924 219434 381952 231662
rect 382108 226166 382136 231676
rect 382674 231662 383056 231690
rect 382280 229900 382332 229906
rect 382280 229842 382332 229848
rect 382292 229090 382320 229842
rect 382280 229084 382332 229090
rect 382280 229026 382332 229032
rect 382648 228268 382700 228274
rect 382648 228210 382700 228216
rect 382096 226160 382148 226166
rect 382096 226102 382148 226108
rect 381924 219406 382228 219434
rect 382200 218890 382228 219406
rect 381820 218884 381872 218890
rect 381820 218826 381872 218832
rect 382188 218884 382240 218890
rect 382188 218826 382240 218832
rect 379348 217246 379422 217274
rect 380176 217246 380250 217274
rect 381004 217246 381078 217274
rect 378520 217110 378594 217138
rect 378566 216988 378594 217110
rect 379394 216988 379422 217246
rect 380222 216988 380250 217246
rect 381050 216988 381078 217246
rect 381832 217138 381860 218826
rect 382660 217274 382688 228210
rect 383028 224398 383056 231662
rect 383016 224392 383068 224398
rect 383016 224334 383068 224340
rect 383212 221610 383240 231676
rect 383778 231662 384160 231690
rect 383476 224528 383528 224534
rect 383476 224470 383528 224476
rect 383200 221604 383252 221610
rect 383200 221546 383252 221552
rect 383488 217274 383516 224470
rect 384132 223174 384160 231662
rect 384316 227186 384344 231676
rect 384684 231662 384882 231690
rect 384304 227180 384356 227186
rect 384304 227122 384356 227128
rect 384304 227044 384356 227050
rect 384304 226986 384356 226992
rect 384120 223168 384172 223174
rect 384120 223110 384172 223116
rect 384316 217274 384344 226986
rect 384684 220522 384712 231662
rect 385420 230382 385448 231676
rect 385408 230376 385460 230382
rect 385408 230318 385460 230324
rect 385972 229498 386000 231676
rect 386328 230376 386380 230382
rect 386328 230318 386380 230324
rect 385960 229492 386012 229498
rect 385960 229434 386012 229440
rect 386340 221474 386368 230318
rect 386524 228546 386552 231676
rect 387076 230382 387104 231676
rect 387064 230376 387116 230382
rect 387064 230318 387116 230324
rect 387064 228676 387116 228682
rect 387064 228618 387116 228624
rect 386512 228540 386564 228546
rect 386512 228482 386564 228488
rect 386788 224256 386840 224262
rect 386788 224198 386840 224204
rect 385960 221468 386012 221474
rect 385960 221410 386012 221416
rect 386328 221468 386380 221474
rect 386328 221410 386380 221416
rect 384672 220516 384724 220522
rect 384672 220458 384724 220464
rect 385132 218748 385184 218754
rect 385132 218690 385184 218696
rect 382660 217246 382734 217274
rect 383488 217246 383562 217274
rect 384316 217246 384390 217274
rect 381832 217110 381906 217138
rect 381878 216988 381906 217110
rect 382706 216988 382734 217246
rect 383534 216988 383562 217246
rect 384362 216988 384390 217246
rect 385144 217138 385172 218690
rect 385972 217274 386000 221410
rect 386800 217274 386828 224198
rect 387076 218074 387104 228618
rect 387628 224534 387656 231676
rect 388180 227050 388208 231676
rect 388444 230376 388496 230382
rect 388444 230318 388496 230324
rect 388456 229094 388484 230318
rect 388732 229094 388760 231676
rect 389284 229634 389312 231676
rect 389850 231662 390232 231690
rect 389732 230240 389784 230246
rect 389732 230182 389784 230188
rect 389272 229628 389324 229634
rect 389272 229570 389324 229576
rect 388456 229066 388668 229094
rect 388732 229066 388852 229094
rect 388444 228948 388496 228954
rect 388444 228890 388496 228896
rect 388456 228274 388484 228890
rect 388444 228268 388496 228274
rect 388444 228210 388496 228216
rect 388168 227044 388220 227050
rect 388168 226986 388220 226992
rect 387616 224528 387668 224534
rect 387616 224470 387668 224476
rect 387616 222012 387668 222018
rect 387616 221954 387668 221960
rect 387064 218068 387116 218074
rect 387064 218010 387116 218016
rect 387628 217274 387656 221954
rect 388640 219978 388668 229066
rect 388824 224262 388852 229066
rect 388812 224256 388864 224262
rect 388812 224198 388864 224204
rect 389744 221202 389772 230182
rect 390204 229294 390232 231662
rect 390388 230314 390416 231676
rect 390376 230308 390428 230314
rect 390376 230250 390428 230256
rect 390468 229628 390520 229634
rect 390468 229570 390520 229576
rect 390192 229288 390244 229294
rect 390192 229230 390244 229236
rect 390100 227452 390152 227458
rect 390100 227394 390152 227400
rect 389732 221196 389784 221202
rect 389732 221138 389784 221144
rect 389272 220244 389324 220250
rect 389272 220186 389324 220192
rect 388628 219972 388680 219978
rect 388628 219914 388680 219920
rect 388444 218068 388496 218074
rect 388444 218010 388496 218016
rect 385972 217246 386046 217274
rect 386800 217246 386874 217274
rect 387628 217246 387702 217274
rect 385144 217110 385218 217138
rect 385190 216988 385218 217110
rect 386018 216988 386046 217246
rect 386846 216988 386874 217246
rect 387674 216988 387702 217246
rect 388456 217138 388484 218010
rect 389284 217274 389312 220186
rect 390112 217274 390140 227394
rect 390480 220386 390508 229570
rect 390940 225894 390968 231676
rect 391492 229906 391520 231676
rect 392044 230042 392072 231676
rect 392610 231662 392992 231690
rect 392216 230172 392268 230178
rect 392216 230114 392268 230120
rect 392400 230172 392452 230178
rect 392400 230114 392452 230120
rect 392032 230036 392084 230042
rect 392032 229978 392084 229984
rect 391204 229900 391256 229906
rect 391204 229842 391256 229848
rect 391480 229900 391532 229906
rect 391480 229842 391532 229848
rect 391216 229090 391244 229842
rect 391664 229764 391716 229770
rect 391664 229706 391716 229712
rect 391204 229084 391256 229090
rect 391204 229026 391256 229032
rect 391676 226438 391704 229706
rect 391848 228948 391900 228954
rect 391848 228890 391900 228896
rect 391664 226432 391716 226438
rect 391664 226374 391716 226380
rect 390928 225888 390980 225894
rect 390928 225830 390980 225836
rect 390928 221876 390980 221882
rect 390928 221818 390980 221824
rect 390468 220380 390520 220386
rect 390468 220322 390520 220328
rect 390940 217274 390968 221818
rect 391860 219434 391888 228890
rect 392228 227458 392256 230114
rect 392412 229498 392440 230114
rect 392584 229900 392636 229906
rect 392584 229842 392636 229848
rect 392400 229492 392452 229498
rect 392400 229434 392452 229440
rect 392596 229094 392624 229842
rect 392964 229770 392992 231662
rect 392952 229764 393004 229770
rect 392952 229706 393004 229712
rect 392596 229066 392808 229094
rect 392216 227452 392268 227458
rect 392216 227394 392268 227400
rect 392584 225616 392636 225622
rect 392584 225558 392636 225564
rect 391768 219406 391888 219434
rect 391768 217274 391796 219406
rect 392596 217274 392624 225558
rect 392780 220658 392808 229066
rect 393148 228682 393176 231676
rect 393136 228676 393188 228682
rect 393136 228618 393188 228624
rect 393700 226302 393728 231676
rect 394252 229634 394280 231676
rect 394240 229628 394292 229634
rect 394240 229570 394292 229576
rect 393964 229288 394016 229294
rect 393964 229230 394016 229236
rect 393688 226296 393740 226302
rect 393688 226238 393740 226244
rect 393976 222154 394004 229230
rect 394240 228268 394292 228274
rect 394240 228210 394292 228216
rect 393412 222148 393464 222154
rect 393412 222090 393464 222096
rect 393964 222148 394016 222154
rect 393964 222090 394016 222096
rect 392768 220652 392820 220658
rect 392768 220594 392820 220600
rect 393424 217274 393452 222090
rect 394252 217274 394280 228210
rect 394804 227798 394832 231676
rect 394976 230172 395028 230178
rect 394976 230114 395028 230120
rect 394792 227792 394844 227798
rect 394792 227734 394844 227740
rect 394988 226522 395016 230114
rect 395356 227594 395384 231676
rect 395724 231662 395922 231690
rect 395344 227588 395396 227594
rect 395344 227530 395396 227536
rect 394988 226494 395292 226522
rect 395068 226432 395120 226438
rect 395068 226374 395120 226380
rect 395080 217274 395108 226374
rect 395264 222630 395292 226494
rect 395252 222624 395304 222630
rect 395252 222566 395304 222572
rect 395724 220250 395752 231662
rect 396460 229362 396488 231676
rect 396724 230036 396776 230042
rect 396724 229978 396776 229984
rect 396448 229356 396500 229362
rect 396448 229298 396500 229304
rect 396736 229094 396764 229978
rect 397012 229498 397040 231676
rect 397000 229492 397052 229498
rect 397000 229434 397052 229440
rect 397368 229356 397420 229362
rect 397368 229298 397420 229304
rect 396736 229066 396948 229094
rect 396724 227316 396776 227322
rect 396724 227258 396776 227264
rect 395712 220244 395764 220250
rect 395712 220186 395764 220192
rect 395896 220108 395948 220114
rect 395896 220050 395948 220056
rect 395908 217274 395936 220050
rect 396736 217274 396764 227258
rect 396920 222018 396948 229066
rect 396908 222012 396960 222018
rect 396908 221954 396960 221960
rect 397380 221882 397408 229298
rect 397564 228818 397592 231676
rect 398130 231662 398604 231690
rect 397736 229084 397788 229090
rect 397736 229026 397788 229032
rect 397552 228812 397604 228818
rect 397552 228754 397604 228760
rect 397748 228664 397776 229026
rect 397656 228636 397776 228664
rect 397368 221876 397420 221882
rect 397368 221818 397420 221824
rect 397656 217870 397684 228636
rect 397828 223304 397880 223310
rect 397828 223246 397880 223252
rect 397644 217864 397696 217870
rect 397644 217806 397696 217812
rect 397840 217546 397868 223246
rect 398576 220114 398604 231662
rect 398668 230058 398696 231676
rect 398668 230042 398788 230058
rect 398668 230036 398800 230042
rect 398668 230030 398748 230036
rect 398748 229978 398800 229984
rect 399220 229294 399248 231676
rect 399392 230308 399444 230314
rect 399392 230250 399444 230256
rect 399208 229288 399260 229294
rect 399208 229230 399260 229236
rect 399404 223582 399432 230250
rect 399576 229764 399628 229770
rect 399576 229706 399628 229712
rect 399392 223576 399444 223582
rect 399392 223518 399444 223524
rect 399588 223310 399616 229706
rect 399772 226030 399800 231676
rect 400324 228274 400352 231676
rect 400876 229906 400904 231676
rect 401336 231662 401442 231690
rect 400864 229900 400916 229906
rect 400864 229842 400916 229848
rect 400864 229628 400916 229634
rect 400864 229570 400916 229576
rect 400680 228948 400732 228954
rect 400680 228890 400732 228896
rect 400312 228268 400364 228274
rect 400312 228210 400364 228216
rect 399760 226024 399812 226030
rect 399760 225966 399812 225972
rect 399576 223304 399628 223310
rect 399576 223246 399628 223252
rect 399208 223032 399260 223038
rect 399208 222974 399260 222980
rect 398564 220108 398616 220114
rect 398564 220050 398616 220056
rect 398380 217864 398432 217870
rect 398380 217806 398432 217812
rect 397656 217518 397868 217546
rect 397656 217274 397684 217518
rect 389284 217246 389358 217274
rect 390112 217246 390186 217274
rect 390940 217246 391014 217274
rect 391768 217246 391842 217274
rect 392596 217246 392670 217274
rect 393424 217246 393498 217274
rect 394252 217246 394326 217274
rect 395080 217246 395154 217274
rect 395908 217246 395982 217274
rect 396736 217246 396810 217274
rect 388456 217110 388530 217138
rect 388502 216988 388530 217110
rect 389330 216988 389358 217246
rect 390158 216988 390186 217246
rect 390986 216988 391014 217246
rect 391814 216988 391842 217246
rect 392642 216988 392670 217246
rect 393470 216988 393498 217246
rect 394298 216988 394326 217246
rect 395126 216988 395154 217246
rect 395954 216988 395982 217246
rect 396782 216988 396810 217246
rect 397610 217246 397684 217274
rect 397610 216988 397638 217246
rect 398392 217138 398420 217806
rect 399220 217274 399248 222974
rect 400036 221740 400088 221746
rect 400036 221682 400088 221688
rect 400048 217274 400076 221682
rect 400692 219434 400720 228890
rect 400876 221338 400904 229570
rect 400864 221332 400916 221338
rect 400864 221274 400916 221280
rect 400692 219406 400904 219434
rect 400876 217274 400904 219406
rect 401336 218754 401364 231662
rect 401980 228954 402008 231676
rect 401968 228948 402020 228954
rect 401968 228890 402020 228896
rect 402244 227792 402296 227798
rect 402244 227734 402296 227740
rect 401692 227452 401744 227458
rect 401692 227394 401744 227400
rect 401324 218748 401376 218754
rect 401324 218690 401376 218696
rect 401704 217274 401732 227394
rect 402256 219298 402284 227734
rect 402532 225758 402560 231676
rect 403084 230382 403112 231676
rect 403072 230376 403124 230382
rect 403072 230318 403124 230324
rect 402520 225752 402572 225758
rect 402520 225694 402572 225700
rect 402980 224664 403032 224670
rect 402980 224606 403032 224612
rect 402520 220788 402572 220794
rect 402520 220730 402572 220736
rect 402244 219292 402296 219298
rect 402244 219234 402296 219240
rect 402532 217274 402560 220730
rect 399220 217246 399294 217274
rect 400048 217246 400122 217274
rect 400876 217246 400950 217274
rect 401704 217246 401778 217274
rect 402532 217246 402606 217274
rect 402992 217258 403020 224606
rect 403636 224398 403664 231676
rect 404096 231662 404202 231690
rect 404096 227458 404124 231662
rect 404268 230376 404320 230382
rect 404268 230318 404320 230324
rect 404084 227452 404136 227458
rect 404084 227394 404136 227400
rect 403440 224392 403492 224398
rect 403440 224334 403492 224340
rect 403624 224392 403676 224398
rect 403624 224334 403676 224340
rect 403452 224126 403480 224334
rect 403440 224120 403492 224126
rect 403440 224062 403492 224068
rect 404280 221746 404308 230318
rect 404740 230246 404768 231676
rect 404728 230240 404780 230246
rect 404728 230182 404780 230188
rect 405292 229498 405320 231676
rect 405844 230382 405872 231676
rect 405832 230376 405884 230382
rect 405832 230318 405884 230324
rect 405280 229492 405332 229498
rect 405280 229434 405332 229440
rect 404636 229424 404688 229430
rect 404636 229366 404688 229372
rect 404648 223038 404676 229366
rect 405004 229288 405056 229294
rect 405004 229230 405056 229236
rect 404636 223032 404688 223038
rect 404636 222974 404688 222980
rect 404268 221740 404320 221746
rect 404268 221682 404320 221688
rect 403348 221196 403400 221202
rect 403348 221138 403400 221144
rect 403360 217274 403388 221138
rect 405016 219162 405044 229230
rect 406396 225214 406424 231676
rect 406948 230466 406976 231676
rect 406948 230450 407252 230466
rect 406948 230444 407264 230450
rect 406948 230438 407212 230444
rect 407212 230386 407264 230392
rect 407028 230376 407080 230382
rect 407028 230318 407080 230324
rect 406384 225208 406436 225214
rect 406384 225150 406436 225156
rect 405372 224392 405424 224398
rect 405372 224334 405424 224340
rect 405004 219156 405056 219162
rect 405004 219098 405056 219104
rect 405384 218890 405412 224334
rect 405832 222896 405884 222902
rect 405832 222838 405884 222844
rect 405004 218884 405056 218890
rect 405004 218826 405056 218832
rect 405372 218884 405424 218890
rect 405372 218826 405424 218832
rect 405016 217274 405044 218826
rect 405844 217274 405872 222838
rect 406660 221604 406712 221610
rect 406660 221546 406712 221552
rect 406672 217274 406700 221546
rect 407040 219026 407068 230318
rect 407500 229634 407528 231676
rect 407488 229628 407540 229634
rect 407488 229570 407540 229576
rect 407764 229084 407816 229090
rect 407764 229026 407816 229032
rect 407776 228818 407804 229026
rect 407764 228812 407816 228818
rect 407764 228754 407816 228760
rect 407488 226160 407540 226166
rect 407488 226102 407540 226108
rect 407028 219020 407080 219026
rect 407028 218962 407080 218968
rect 407500 217274 407528 226102
rect 408052 222766 408080 231676
rect 408604 224806 408632 231676
rect 409170 231662 409552 231690
rect 408592 224800 408644 224806
rect 408592 224742 408644 224748
rect 409144 224120 409196 224126
rect 409144 224062 409196 224068
rect 408316 223168 408368 223174
rect 408316 223110 408368 223116
rect 408040 222760 408092 222766
rect 408040 222702 408092 222708
rect 408328 217274 408356 223110
rect 409156 217274 409184 224062
rect 409524 221202 409552 231662
rect 409708 224126 409736 231676
rect 409696 224120 409748 224126
rect 409696 224062 409748 224068
rect 410260 223446 410288 231676
rect 410616 227180 410668 227186
rect 410616 227122 410668 227128
rect 410248 223440 410300 223446
rect 410248 223382 410300 223388
rect 409972 221468 410024 221474
rect 409972 221410 410024 221416
rect 409512 221196 409564 221202
rect 409512 221138 409564 221144
rect 409984 217274 410012 221410
rect 410628 219434 410656 227122
rect 410812 224398 410840 231676
rect 411364 230178 411392 231676
rect 411930 231662 412312 231690
rect 411352 230172 411404 230178
rect 411352 230114 411404 230120
rect 410800 224392 410852 224398
rect 410800 224334 410852 224340
rect 411628 222624 411680 222630
rect 411628 222566 411680 222572
rect 410628 219406 410840 219434
rect 410812 217274 410840 219406
rect 411640 217274 411668 222566
rect 412284 221610 412312 231662
rect 412468 222902 412496 231676
rect 412824 230444 412876 230450
rect 412824 230386 412876 230392
rect 412836 229362 412864 230386
rect 412824 229356 412876 229362
rect 412824 229298 412876 229304
rect 413020 224670 413048 231676
rect 413572 230382 413600 231676
rect 413560 230376 413612 230382
rect 413560 230318 413612 230324
rect 413284 230308 413336 230314
rect 413284 230250 413336 230256
rect 413296 229094 413324 230250
rect 414124 230042 414152 231676
rect 414112 230036 414164 230042
rect 414112 229978 414164 229984
rect 413296 229066 413508 229094
rect 413008 224664 413060 224670
rect 413008 224606 413060 224612
rect 413284 224528 413336 224534
rect 413284 224470 413336 224476
rect 412456 222896 412508 222902
rect 412456 222838 412508 222844
rect 412272 221604 412324 221610
rect 412272 221546 412324 221552
rect 412456 220516 412508 220522
rect 412456 220458 412508 220464
rect 412468 217274 412496 220458
rect 413296 217274 413324 224470
rect 413480 220794 413508 229066
rect 414204 228540 414256 228546
rect 414204 228482 414256 228488
rect 413468 220788 413520 220794
rect 413468 220730 413520 220736
rect 414216 217274 414244 228482
rect 414676 224534 414704 231676
rect 415228 230178 415256 231676
rect 414848 230172 414900 230178
rect 414848 230114 414900 230120
rect 415216 230172 415268 230178
rect 415216 230114 415268 230120
rect 414860 228546 414888 230114
rect 415308 230036 415360 230042
rect 415308 229978 415360 229984
rect 414848 228540 414900 228546
rect 414848 228482 414900 228488
rect 414940 227044 414992 227050
rect 414940 226986 414992 226992
rect 414664 224528 414716 224534
rect 414664 224470 414716 224476
rect 398392 217110 398466 217138
rect 398438 216988 398466 217110
rect 399266 216988 399294 217246
rect 400094 216988 400122 217246
rect 400922 216988 400950 217246
rect 401750 216988 401778 217246
rect 402578 216988 402606 217246
rect 402980 217252 403032 217258
rect 403360 217246 403434 217274
rect 402980 217194 403032 217200
rect 403406 216988 403434 217246
rect 404222 217252 404274 217258
rect 405016 217246 405090 217274
rect 405844 217246 405918 217274
rect 406672 217246 406746 217274
rect 407500 217246 407574 217274
rect 408328 217246 408402 217274
rect 409156 217246 409230 217274
rect 409984 217246 410058 217274
rect 410812 217246 410886 217274
rect 411640 217246 411714 217274
rect 412468 217246 412542 217274
rect 413296 217246 413370 217274
rect 404222 217194 404274 217200
rect 404234 216988 404262 217194
rect 405062 216988 405090 217246
rect 405890 216988 405918 217246
rect 406718 216988 406746 217246
rect 407546 216988 407574 217246
rect 408374 216988 408402 217246
rect 409202 216988 409230 217246
rect 410030 216988 410058 217246
rect 410858 216988 410886 217246
rect 411686 216988 411714 217246
rect 412514 216988 412542 217246
rect 413342 216988 413370 217246
rect 414170 217246 414244 217274
rect 414952 217274 414980 226986
rect 415320 220522 415348 229978
rect 415780 226166 415808 231676
rect 416332 230042 416360 231676
rect 416898 231662 417280 231690
rect 416320 230036 416372 230042
rect 416320 229978 416372 229984
rect 416044 229900 416096 229906
rect 416044 229842 416096 229848
rect 415768 226160 415820 226166
rect 415768 226102 415820 226108
rect 416056 222290 416084 229842
rect 417252 223174 417280 231662
rect 417436 229094 417464 231676
rect 417436 229066 417648 229094
rect 417424 224256 417476 224262
rect 417424 224198 417476 224204
rect 417240 223168 417292 223174
rect 417240 223110 417292 223116
rect 416044 222284 416096 222290
rect 416044 222226 416096 222232
rect 416596 222148 416648 222154
rect 416596 222090 416648 222096
rect 415308 220516 415360 220522
rect 415308 220458 415360 220464
rect 415768 219972 415820 219978
rect 415768 219914 415820 219920
rect 415780 217274 415808 219914
rect 416608 217274 416636 222090
rect 417436 217274 417464 224198
rect 417620 223990 417648 229066
rect 417988 227322 418016 231676
rect 417976 227316 418028 227322
rect 417976 227258 418028 227264
rect 418540 225350 418568 231676
rect 418804 230376 418856 230382
rect 418804 230318 418856 230324
rect 418528 225344 418580 225350
rect 418528 225286 418580 225292
rect 417608 223984 417660 223990
rect 417608 223926 417660 223932
rect 418252 223576 418304 223582
rect 418252 223518 418304 223524
rect 418264 217274 418292 223518
rect 418816 219978 418844 230318
rect 419092 229906 419120 231676
rect 419658 231662 420040 231690
rect 419080 229900 419132 229906
rect 419080 229842 419132 229848
rect 419724 225888 419776 225894
rect 419724 225830 419776 225836
rect 419080 220380 419132 220386
rect 419080 220322 419132 220328
rect 418804 219972 418856 219978
rect 418804 219914 418856 219920
rect 419092 217274 419120 220322
rect 414952 217246 415026 217274
rect 415780 217246 415854 217274
rect 416608 217246 416682 217274
rect 417436 217246 417510 217274
rect 418264 217246 418338 217274
rect 419092 217246 419166 217274
rect 419736 217258 419764 225830
rect 420012 224942 420040 231662
rect 420196 230314 420224 231676
rect 420564 231662 420762 231690
rect 420184 230308 420236 230314
rect 420184 230250 420236 230256
rect 420184 229764 420236 229770
rect 420184 229706 420236 229712
rect 420000 224936 420052 224942
rect 420000 224878 420052 224884
rect 419908 222012 419960 222018
rect 419908 221954 419960 221960
rect 419920 217274 419948 221954
rect 420196 221066 420224 229706
rect 420184 221060 420236 221066
rect 420184 221002 420236 221008
rect 420564 220386 420592 231662
rect 421300 230450 421328 231676
rect 421288 230444 421340 230450
rect 421288 230386 421340 230392
rect 421852 229362 421880 231676
rect 422208 230444 422260 230450
rect 422208 230386 422260 230392
rect 421564 229356 421616 229362
rect 421564 229298 421616 229304
rect 421840 229356 421892 229362
rect 421840 229298 421892 229304
rect 421576 229094 421604 229298
rect 421392 229066 421604 229094
rect 420552 220380 420604 220386
rect 420552 220322 420604 220328
rect 421392 219706 421420 229066
rect 421840 224120 421892 224126
rect 421840 224062 421892 224068
rect 421564 223304 421616 223310
rect 421564 223246 421616 223252
rect 421380 219700 421432 219706
rect 421380 219642 421432 219648
rect 421576 217274 421604 223246
rect 421852 218618 421880 224062
rect 422220 221474 422248 230386
rect 422404 225894 422432 231676
rect 422956 229226 422984 231676
rect 422944 229220 422996 229226
rect 422944 229162 422996 229168
rect 423508 228818 423536 231676
rect 424060 230042 424088 231676
rect 424048 230036 424100 230042
rect 424048 229978 424100 229984
rect 424324 229628 424376 229634
rect 424324 229570 424376 229576
rect 423496 228812 423548 228818
rect 423496 228754 423548 228760
rect 424048 228676 424100 228682
rect 424048 228618 424100 228624
rect 422392 225888 422444 225894
rect 422392 225830 422444 225836
rect 422208 221468 422260 221474
rect 422208 221410 422260 221416
rect 423220 221332 423272 221338
rect 423220 221274 423272 221280
rect 422300 221196 422352 221202
rect 422300 221138 422352 221144
rect 422312 219434 422340 221138
rect 422484 220652 422536 220658
rect 422484 220594 422536 220600
rect 422300 219428 422352 219434
rect 422300 219370 422352 219376
rect 421840 218612 421892 218618
rect 421840 218554 421892 218560
rect 422496 217274 422524 220594
rect 414170 216988 414198 217246
rect 414998 216988 415026 217246
rect 415826 216988 415854 217246
rect 416654 216988 416682 217246
rect 417482 216988 417510 217246
rect 418310 216988 418338 217246
rect 419138 216988 419166 217246
rect 419724 217252 419776 217258
rect 419920 217246 419994 217274
rect 419724 217194 419776 217200
rect 419966 216988 419994 217246
rect 420782 217252 420834 217258
rect 421576 217246 421650 217274
rect 420782 217194 420834 217200
rect 420794 216988 420822 217194
rect 421622 216988 421650 217246
rect 422450 217246 422524 217274
rect 423232 217274 423260 221274
rect 424060 217274 424088 228618
rect 424336 222018 424364 229570
rect 424612 227186 424640 231676
rect 425178 231662 425376 231690
rect 424600 227180 424652 227186
rect 424600 227122 424652 227128
rect 425348 222630 425376 231662
rect 425716 229634 425744 231676
rect 425704 229628 425756 229634
rect 425704 229570 425756 229576
rect 426268 227050 426296 231676
rect 426820 228682 426848 231676
rect 427386 231662 427768 231690
rect 427084 229900 427136 229906
rect 427084 229842 427136 229848
rect 426808 228676 426860 228682
rect 426808 228618 426860 228624
rect 426256 227044 426308 227050
rect 426256 226986 426308 226992
rect 425704 226296 425756 226302
rect 425704 226238 425756 226244
rect 425336 222624 425388 222630
rect 425336 222566 425388 222572
rect 424324 222012 424376 222018
rect 424324 221954 424376 221960
rect 424876 219292 424928 219298
rect 424876 219234 424928 219240
rect 423232 217246 423306 217274
rect 424060 217246 424134 217274
rect 422450 216988 422478 217246
rect 423278 216988 423306 217246
rect 424106 216988 424134 217246
rect 424888 217138 424916 219234
rect 425716 217274 425744 226238
rect 425888 224528 425940 224534
rect 425888 224470 425940 224476
rect 425900 219162 425928 224470
rect 427096 221882 427124 229842
rect 427360 227588 427412 227594
rect 427360 227530 427412 227536
rect 426532 221876 426584 221882
rect 426532 221818 426584 221824
rect 427084 221876 427136 221882
rect 427084 221818 427136 221824
rect 425888 219156 425940 219162
rect 425888 219098 425940 219104
rect 426544 217274 426572 221818
rect 427372 217274 427400 227530
rect 427740 222494 427768 231662
rect 427924 230450 427952 231676
rect 427912 230444 427964 230450
rect 427912 230386 427964 230392
rect 428476 229906 428504 231676
rect 428844 231662 429042 231690
rect 428464 229900 428516 229906
rect 428464 229842 428516 229848
rect 428096 229764 428148 229770
rect 428096 229706 428148 229712
rect 428108 226302 428136 229706
rect 428844 229634 428872 231662
rect 429016 230444 429068 230450
rect 429016 230386 429068 230392
rect 429200 230444 429252 230450
rect 429200 230386 429252 230392
rect 428832 229628 428884 229634
rect 428832 229570 428884 229576
rect 428464 229492 428516 229498
rect 428464 229434 428516 229440
rect 428096 226296 428148 226302
rect 428096 226238 428148 226244
rect 428188 223032 428240 223038
rect 428188 222974 428240 222980
rect 427728 222488 427780 222494
rect 427728 222430 427780 222436
rect 428200 217274 428228 222974
rect 428476 221338 428504 229434
rect 429028 229094 429056 230386
rect 429212 230042 429240 230386
rect 429200 230036 429252 230042
rect 429200 229978 429252 229984
rect 429384 230036 429436 230042
rect 429384 229978 429436 229984
rect 429396 229226 429424 229978
rect 429384 229220 429436 229226
rect 429384 229162 429436 229168
rect 428844 229066 429056 229094
rect 428464 221332 428516 221338
rect 428464 221274 428516 221280
rect 428844 219842 428872 229066
rect 429580 227730 429608 231676
rect 429752 229492 429804 229498
rect 429752 229434 429804 229440
rect 429764 229226 429792 229434
rect 429752 229220 429804 229226
rect 429752 229162 429804 229168
rect 430132 229090 430160 231676
rect 429936 229084 429988 229090
rect 429936 229026 429988 229032
rect 430120 229084 430172 229090
rect 430120 229026 430172 229032
rect 429568 227724 429620 227730
rect 429568 227666 429620 227672
rect 429752 222148 429804 222154
rect 429752 222090 429804 222096
rect 429016 220244 429068 220250
rect 429016 220186 429068 220192
rect 428832 219836 428884 219842
rect 428832 219778 428884 219784
rect 429028 217274 429056 220186
rect 429764 217274 429792 222090
rect 429948 218074 429976 229026
rect 430684 223038 430712 231676
rect 431250 231662 431632 231690
rect 431224 223984 431276 223990
rect 431224 223926 431276 223932
rect 430672 223032 430724 223038
rect 430672 222974 430724 222980
rect 431236 219298 431264 223926
rect 431604 223310 431632 231662
rect 431788 223990 431816 231676
rect 432340 224262 432368 231676
rect 432604 228268 432656 228274
rect 432604 228210 432656 228216
rect 432328 224256 432380 224262
rect 432328 224198 432380 224204
rect 431776 223984 431828 223990
rect 431776 223926 431828 223932
rect 431592 223304 431644 223310
rect 431592 223246 431644 223252
rect 432328 220108 432380 220114
rect 432328 220050 432380 220056
rect 430856 219292 430908 219298
rect 430856 219234 430908 219240
rect 431224 219292 431276 219298
rect 431224 219234 431276 219240
rect 430868 218074 430896 219234
rect 429936 218068 429988 218074
rect 429936 218010 429988 218016
rect 430672 218068 430724 218074
rect 430672 218010 430724 218016
rect 430856 218068 430908 218074
rect 430856 218010 430908 218016
rect 431500 218068 431552 218074
rect 431500 218010 431552 218016
rect 425716 217246 425790 217274
rect 426544 217246 426618 217274
rect 427372 217246 427446 217274
rect 428200 217246 428274 217274
rect 429028 217246 429102 217274
rect 429764 217246 429930 217274
rect 424888 217110 424962 217138
rect 424934 216988 424962 217110
rect 425762 216988 425790 217246
rect 426590 216988 426618 217246
rect 427418 216988 427446 217246
rect 428246 216988 428274 217246
rect 429074 216988 429102 217246
rect 429902 216988 429930 217246
rect 430684 217138 430712 218010
rect 431512 217138 431540 218010
rect 432340 217274 432368 220050
rect 432616 218074 432644 228210
rect 432892 225486 432920 231676
rect 433458 231662 433840 231690
rect 432880 225480 432932 225486
rect 432880 225422 432932 225428
rect 433812 224126 433840 231662
rect 433996 229094 434024 231676
rect 433996 229066 434208 229094
rect 433984 226024 434036 226030
rect 433984 225966 434036 225972
rect 433800 224120 433852 224126
rect 433800 224062 433852 224068
rect 433156 221060 433208 221066
rect 433156 221002 433208 221008
rect 432604 218068 432656 218074
rect 432604 218010 432656 218016
rect 433168 217274 433196 221002
rect 433996 217274 434024 225966
rect 434180 224534 434208 229066
rect 434548 228274 434576 231676
rect 435100 230314 435128 231676
rect 434904 230308 434956 230314
rect 434904 230250 434956 230256
rect 435088 230308 435140 230314
rect 435088 230250 435140 230256
rect 434916 229498 434944 230250
rect 434904 229492 434956 229498
rect 434904 229434 434956 229440
rect 434536 228268 434588 228274
rect 434536 228210 434588 228216
rect 434168 224528 434220 224534
rect 434168 224470 434220 224476
rect 434168 224392 434220 224398
rect 434168 224334 434220 224340
rect 434180 218482 434208 224334
rect 435364 224256 435416 224262
rect 435364 224198 435416 224204
rect 434812 218748 434864 218754
rect 434812 218690 434864 218696
rect 434168 218476 434220 218482
rect 434168 218418 434220 218424
rect 432340 217246 432414 217274
rect 433168 217246 433242 217274
rect 433996 217246 434070 217274
rect 430684 217110 430758 217138
rect 431512 217110 431586 217138
rect 430730 216988 430758 217110
rect 431558 216988 431586 217110
rect 432386 216988 432414 217246
rect 433214 216988 433242 217246
rect 434042 216988 434070 217246
rect 434824 217138 434852 218690
rect 435376 218657 435404 224198
rect 435652 223582 435680 231676
rect 436218 231662 436600 231690
rect 436008 230308 436060 230314
rect 436008 230250 436060 230256
rect 435640 223576 435692 223582
rect 435640 223518 435692 223524
rect 436020 220250 436048 230250
rect 436572 226030 436600 231662
rect 436756 227866 436784 231676
rect 437112 228948 437164 228954
rect 437112 228890 437164 228896
rect 436744 227860 436796 227866
rect 436744 227802 436796 227808
rect 436560 226024 436612 226030
rect 436560 225966 436612 225972
rect 436468 221740 436520 221746
rect 436468 221682 436520 221688
rect 436008 220244 436060 220250
rect 436008 220186 436060 220192
rect 436284 219020 436336 219026
rect 436284 218962 436336 218968
rect 435362 218648 435418 218657
rect 435362 218583 435418 218592
rect 436296 218346 436324 218962
rect 436284 218340 436336 218346
rect 436284 218282 436336 218288
rect 435640 218068 435692 218074
rect 435640 218010 435692 218016
rect 435652 217138 435680 218010
rect 436480 217274 436508 221682
rect 437124 219434 437152 228890
rect 437308 220658 437336 231676
rect 437874 231662 438256 231690
rect 438228 224262 438256 231662
rect 438412 225622 438440 231676
rect 438964 229770 438992 231676
rect 439530 231662 439912 231690
rect 438952 229764 439004 229770
rect 438952 229706 439004 229712
rect 439504 229492 439556 229498
rect 439504 229434 439556 229440
rect 439516 228954 439544 229434
rect 439504 228948 439556 228954
rect 439504 228890 439556 228896
rect 439044 225752 439096 225758
rect 439044 225694 439096 225700
rect 438400 225616 438452 225622
rect 438400 225558 438452 225564
rect 438216 224256 438268 224262
rect 438216 224198 438268 224204
rect 438308 223984 438360 223990
rect 438308 223926 438360 223932
rect 437296 220652 437348 220658
rect 437296 220594 437348 220600
rect 437124 219406 437336 219434
rect 436928 219292 436980 219298
rect 436928 219234 436980 219240
rect 436940 219026 436968 219234
rect 436928 219020 436980 219026
rect 436928 218962 436980 218968
rect 437308 217274 437336 219406
rect 438124 218884 438176 218890
rect 438124 218826 438176 218832
rect 436480 217246 436554 217274
rect 437308 217246 437382 217274
rect 434824 217110 434898 217138
rect 435652 217110 435726 217138
rect 434870 216988 434898 217110
rect 435698 216988 435726 217110
rect 436526 216988 436554 217246
rect 437354 216988 437382 217246
rect 438136 217138 438164 218826
rect 438320 218754 438348 223926
rect 438308 218748 438360 218754
rect 438308 218690 438360 218696
rect 439056 217274 439084 225694
rect 439884 223530 439912 231662
rect 440068 223718 440096 231676
rect 440634 231662 441016 231690
rect 441186 231662 441568 231690
rect 440608 227452 440660 227458
rect 440608 227394 440660 227400
rect 440056 223712 440108 223718
rect 440056 223654 440108 223660
rect 439884 223502 440004 223530
rect 439780 221332 439832 221338
rect 439780 221274 439832 221280
rect 439010 217246 439084 217274
rect 439792 217274 439820 221274
rect 439976 221066 440004 223502
rect 439964 221060 440016 221066
rect 439964 221002 440016 221008
rect 440620 217274 440648 227394
rect 440988 225593 441016 231662
rect 440974 225584 441030 225593
rect 440974 225519 441030 225528
rect 441540 221746 441568 231662
rect 441724 230382 441752 231676
rect 442290 231662 442672 231690
rect 441896 230512 441948 230518
rect 441896 230454 441948 230460
rect 441712 230376 441764 230382
rect 441712 230318 441764 230324
rect 441908 230178 441936 230454
rect 441712 230172 441764 230178
rect 441712 230114 441764 230120
rect 441896 230172 441948 230178
rect 441896 230114 441948 230120
rect 441724 229498 441752 230114
rect 441896 229628 441948 229634
rect 441896 229570 441948 229576
rect 441712 229492 441764 229498
rect 441712 229434 441764 229440
rect 441908 226642 441936 229570
rect 442448 228268 442500 228274
rect 442448 228210 442500 228216
rect 441896 226636 441948 226642
rect 441896 226578 441948 226584
rect 441528 221740 441580 221746
rect 441528 221682 441580 221688
rect 442264 220788 442316 220794
rect 442264 220730 442316 220736
rect 441436 218340 441488 218346
rect 441436 218282 441488 218288
rect 439792 217246 439866 217274
rect 440620 217246 440694 217274
rect 438136 217110 438210 217138
rect 438182 216988 438210 217110
rect 439010 216988 439038 217246
rect 439838 216988 439866 217246
rect 440666 216988 440694 217246
rect 441448 217138 441476 218282
rect 442276 217274 442304 220730
rect 442460 218929 442488 228210
rect 442644 224126 442672 231662
rect 442828 230518 442856 231676
rect 442816 230512 442868 230518
rect 442816 230454 442868 230460
rect 443380 230382 443408 231676
rect 442908 230376 442960 230382
rect 442908 230318 442960 230324
rect 443368 230376 443420 230382
rect 443368 230318 443420 230324
rect 442632 224120 442684 224126
rect 442632 224062 442684 224068
rect 442920 220114 442948 230318
rect 443932 229094 443960 231676
rect 444196 230376 444248 230382
rect 444196 230318 444248 230324
rect 444208 229094 444236 230318
rect 444484 229634 444512 231676
rect 444760 231662 445050 231690
rect 444472 229628 444524 229634
rect 444472 229570 444524 229576
rect 444760 229094 444788 231662
rect 445588 229094 445616 231676
rect 446140 230314 446168 231676
rect 446324 231662 446706 231690
rect 447258 231662 447732 231690
rect 447810 231662 448192 231690
rect 446128 230308 446180 230314
rect 446128 230250 446180 230256
rect 446324 229094 446352 231662
rect 447508 230172 447560 230178
rect 447508 230114 447560 230120
rect 446772 230036 446824 230042
rect 446772 229978 446824 229984
rect 443932 229066 444144 229094
rect 444208 229066 444328 229094
rect 444760 229066 444972 229094
rect 443920 225208 443972 225214
rect 443920 225150 443972 225156
rect 443092 222012 443144 222018
rect 443092 221954 443144 221960
rect 442908 220108 442960 220114
rect 442908 220050 442960 220056
rect 442446 218920 442502 218929
rect 442446 218855 442502 218864
rect 443104 217274 443132 221954
rect 443932 217274 443960 225150
rect 444116 217598 444144 229066
rect 444300 221202 444328 229066
rect 444748 222760 444800 222766
rect 444748 222702 444800 222708
rect 444288 221196 444340 221202
rect 444288 221138 444340 221144
rect 444104 217592 444156 217598
rect 444104 217534 444156 217540
rect 444760 217274 444788 222702
rect 444944 221338 444972 229066
rect 445404 229066 445616 229094
rect 446232 229066 446352 229094
rect 444932 221332 444984 221338
rect 444932 221274 444984 221280
rect 445404 217734 445432 229066
rect 446232 220794 446260 229066
rect 446784 228274 446812 229978
rect 446956 229220 447008 229226
rect 446956 229162 447008 229168
rect 446772 228268 446824 228274
rect 446772 228210 446824 228216
rect 446968 227458 446996 229162
rect 446956 227452 447008 227458
rect 446956 227394 447008 227400
rect 447520 225758 447548 230114
rect 447508 225752 447560 225758
rect 447508 225694 447560 225700
rect 446404 225344 446456 225350
rect 446404 225286 446456 225292
rect 446220 220788 446272 220794
rect 446220 220730 446272 220736
rect 445576 219700 445628 219706
rect 445576 219642 445628 219648
rect 445392 217728 445444 217734
rect 445392 217670 445444 217676
rect 445588 217274 445616 219642
rect 446416 219026 446444 225286
rect 447232 224800 447284 224806
rect 447232 224742 447284 224748
rect 446956 221604 447008 221610
rect 446956 221546 447008 221552
rect 446404 219020 446456 219026
rect 446404 218962 446456 218968
rect 446404 218612 446456 218618
rect 446404 218554 446456 218560
rect 442276 217246 442350 217274
rect 443104 217246 443178 217274
rect 443932 217246 444006 217274
rect 444760 217246 444834 217274
rect 445588 217246 445662 217274
rect 441448 217110 441522 217138
rect 441494 216988 441522 217110
rect 442322 216988 442350 217246
rect 443150 216988 443178 217246
rect 443978 216988 444006 217246
rect 444806 216988 444834 217246
rect 445634 216988 445662 217246
rect 446416 217138 446444 218554
rect 446968 218074 446996 221546
rect 446956 218068 447008 218074
rect 446956 218010 447008 218016
rect 447244 217274 447272 224742
rect 447704 219570 447732 231662
rect 448164 230042 448192 231662
rect 448152 230036 448204 230042
rect 448152 229978 448204 229984
rect 448348 229226 448376 231676
rect 448914 231662 449296 231690
rect 448336 229220 448388 229226
rect 448336 229162 448388 229168
rect 449268 229094 449296 231662
rect 449452 229094 449480 231676
rect 449912 231662 450018 231690
rect 449268 229066 449388 229094
rect 449452 229066 449572 229094
rect 449164 226160 449216 226166
rect 449164 226102 449216 226108
rect 448060 223440 448112 223446
rect 448060 223382 448112 223388
rect 447692 219564 447744 219570
rect 447692 219506 447744 219512
rect 448072 217274 448100 223382
rect 449176 219434 449204 226102
rect 449360 219434 449388 229066
rect 449544 222873 449572 229066
rect 449530 222864 449586 222873
rect 449530 222799 449586 222808
rect 449912 222018 449940 231662
rect 450556 230654 450584 231676
rect 450544 230648 450596 230654
rect 450544 230590 450596 230596
rect 451108 230518 451136 231676
rect 451096 230512 451148 230518
rect 451096 230454 451148 230460
rect 450728 230444 450780 230450
rect 450728 230386 450780 230392
rect 450740 229498 450768 230386
rect 450544 229492 450596 229498
rect 450544 229434 450596 229440
rect 450728 229492 450780 229498
rect 450728 229434 450780 229440
rect 449900 222012 449952 222018
rect 449900 221954 449952 221960
rect 449900 221740 449952 221746
rect 449900 221682 449952 221688
rect 448888 219428 448940 219434
rect 448888 219370 448940 219376
rect 449164 219428 449216 219434
rect 449360 219406 449572 219434
rect 449164 219370 449216 219376
rect 447244 217246 447318 217274
rect 448072 217246 448146 217274
rect 446416 217110 446490 217138
rect 446462 216988 446490 217110
rect 447290 216988 447318 217246
rect 448118 216988 448146 217246
rect 448900 217138 448928 219370
rect 449544 217394 449572 219406
rect 449912 218210 449940 221682
rect 450556 218618 450584 229434
rect 451188 229356 451240 229362
rect 451188 229298 451240 229304
rect 451200 229106 451228 229298
rect 451200 229078 451320 229106
rect 451292 223446 451320 229078
rect 451660 228546 451688 231676
rect 452226 231662 452608 231690
rect 451464 228540 451516 228546
rect 451464 228482 451516 228488
rect 451648 228540 451700 228546
rect 451648 228482 451700 228488
rect 451280 223440 451332 223446
rect 451280 223382 451332 223388
rect 451476 223258 451504 228482
rect 451292 223230 451504 223258
rect 450544 218612 450596 218618
rect 450544 218554 450596 218560
rect 450544 218476 450596 218482
rect 450544 218418 450596 218424
rect 449900 218204 449952 218210
rect 449900 218146 449952 218152
rect 449716 218068 449768 218074
rect 449716 218010 449768 218016
rect 449532 217388 449584 217394
rect 449532 217330 449584 217336
rect 449728 217138 449756 218010
rect 450556 217138 450584 218418
rect 451292 217190 451320 223230
rect 451464 222896 451516 222902
rect 451464 222838 451516 222844
rect 451476 217274 451504 222838
rect 452580 222154 452608 231662
rect 452764 223854 452792 231676
rect 453316 229362 453344 231676
rect 453304 229356 453356 229362
rect 453304 229298 453356 229304
rect 453868 226166 453896 231676
rect 453856 226160 453908 226166
rect 453856 226102 453908 226108
rect 453856 224664 453908 224670
rect 453856 224606 453908 224612
rect 452752 223848 452804 223854
rect 452752 223790 452804 223796
rect 452568 222148 452620 222154
rect 452568 222090 452620 222096
rect 453028 220516 453080 220522
rect 453028 220458 453080 220464
rect 451430 217246 451504 217274
rect 453040 217274 453068 220458
rect 453868 217274 453896 224606
rect 454420 223990 454448 231676
rect 454972 228002 455000 231676
rect 455524 230178 455552 231676
rect 455512 230172 455564 230178
rect 455512 230114 455564 230120
rect 455878 229392 455934 229401
rect 456076 229362 456104 231676
rect 456536 231662 456642 231690
rect 455878 229327 455880 229336
rect 455932 229327 455934 229336
rect 456064 229356 456116 229362
rect 455880 229298 455932 229304
rect 456064 229298 456116 229304
rect 456536 228138 456564 231662
rect 457180 230178 457208 231676
rect 456708 230172 456760 230178
rect 456708 230114 456760 230120
rect 457168 230172 457220 230178
rect 457168 230114 457220 230120
rect 456524 228132 456576 228138
rect 456524 228074 456576 228080
rect 454960 227996 455012 228002
rect 454960 227938 455012 227944
rect 454868 224936 454920 224942
rect 454868 224878 454920 224884
rect 454408 223984 454460 223990
rect 454408 223926 454460 223932
rect 454684 219292 454736 219298
rect 454684 219234 454736 219240
rect 453040 217246 453114 217274
rect 453868 217246 453942 217274
rect 451280 217184 451332 217190
rect 448900 217110 448974 217138
rect 449728 217110 449802 217138
rect 450556 217110 450630 217138
rect 451280 217126 451332 217132
rect 448946 216988 448974 217110
rect 449774 216988 449802 217110
rect 450602 216988 450630 217110
rect 451430 216988 451458 217246
rect 452246 217184 452298 217190
rect 452246 217126 452298 217132
rect 452258 216988 452286 217126
rect 453086 216988 453114 217246
rect 453914 216988 453942 217246
rect 454696 217138 454724 219234
rect 454880 218890 454908 224878
rect 456720 221882 456748 230114
rect 457444 229084 457496 229090
rect 457444 229026 457496 229032
rect 456892 223168 456944 223174
rect 456892 223110 456944 223116
rect 456340 221876 456392 221882
rect 456340 221818 456392 221824
rect 456708 221876 456760 221882
rect 456708 221818 456760 221824
rect 455512 219972 455564 219978
rect 455512 219914 455564 219920
rect 454868 218884 454920 218890
rect 454868 218826 454920 218832
rect 455524 217274 455552 219914
rect 456064 217728 456116 217734
rect 456064 217670 456116 217676
rect 456076 217462 456104 217670
rect 456064 217456 456116 217462
rect 456064 217398 456116 217404
rect 456352 217274 456380 221818
rect 455524 217246 455598 217274
rect 456352 217246 456426 217274
rect 454696 217110 454770 217138
rect 454742 216988 454770 217110
rect 455570 216988 455598 217246
rect 456398 216988 456426 217246
rect 456904 217190 456932 223110
rect 457456 219434 457484 229026
rect 457732 224670 457760 231676
rect 458298 231662 458680 231690
rect 458850 231662 459232 231690
rect 458088 230172 458140 230178
rect 458088 230114 458140 230120
rect 458456 230172 458508 230178
rect 458456 230114 458508 230120
rect 457720 224664 457772 224670
rect 457720 224606 457772 224612
rect 458100 221746 458128 230114
rect 458468 229362 458496 230114
rect 458456 229356 458508 229362
rect 458456 229298 458508 229304
rect 458652 226778 458680 231662
rect 458822 229392 458878 229401
rect 458822 229327 458824 229336
rect 458876 229327 458878 229336
rect 458824 229298 458876 229304
rect 458640 226772 458692 226778
rect 458640 226714 458692 226720
rect 458640 225888 458692 225894
rect 458640 225830 458692 225836
rect 458088 221740 458140 221746
rect 458088 221682 458140 221688
rect 457444 219428 457496 219434
rect 457444 219370 457496 219376
rect 457168 218612 457220 218618
rect 457168 218554 457220 218560
rect 456892 217184 456944 217190
rect 456892 217126 456944 217132
rect 457180 217138 457208 218554
rect 458652 218482 458680 225830
rect 459008 222624 459060 222630
rect 459008 222566 459060 222572
rect 458824 219292 458876 219298
rect 458824 219234 458876 219240
rect 458640 218476 458692 218482
rect 458640 218418 458692 218424
rect 458042 217184 458094 217190
rect 457180 217110 457254 217138
rect 458042 217126 458094 217132
rect 458836 217138 458864 219234
rect 459020 218618 459048 222566
rect 459204 222358 459232 231662
rect 459388 225350 459416 231676
rect 459940 229090 459968 231676
rect 459928 229084 459980 229090
rect 459928 229026 459980 229032
rect 459376 225344 459428 225350
rect 459376 225286 459428 225292
rect 460492 223174 460520 231676
rect 461058 231662 461256 231690
rect 461228 229094 461256 231662
rect 461136 229066 461256 229094
rect 461136 225214 461164 229066
rect 461596 227594 461624 231676
rect 462148 229094 462176 231676
rect 461964 229066 462176 229094
rect 461584 227588 461636 227594
rect 461584 227530 461636 227536
rect 461308 226296 461360 226302
rect 461308 226238 461360 226244
rect 461124 225208 461176 225214
rect 461124 225150 461176 225156
rect 460480 223168 460532 223174
rect 460480 223110 460532 223116
rect 460204 222488 460256 222494
rect 460204 222430 460256 222436
rect 459192 222352 459244 222358
rect 459192 222294 459244 222300
rect 459836 220380 459888 220386
rect 459836 220322 459888 220328
rect 459652 219020 459704 219026
rect 459652 218962 459704 218968
rect 459008 218612 459060 218618
rect 459008 218554 459060 218560
rect 459664 217138 459692 218962
rect 459848 218346 459876 220322
rect 460216 219162 460244 222430
rect 460204 219156 460256 219162
rect 460204 219098 460256 219104
rect 460480 219020 460532 219026
rect 460480 218962 460532 218968
rect 459836 218340 459888 218346
rect 459836 218282 459888 218288
rect 460492 217138 460520 218962
rect 461320 217274 461348 226238
rect 461964 222494 461992 229066
rect 462136 227316 462188 227322
rect 462136 227258 462188 227264
rect 461952 222488 462004 222494
rect 461952 222430 462004 222436
rect 462148 217274 462176 227258
rect 462700 226302 462728 231676
rect 463266 231662 463556 231690
rect 463818 231662 464200 231690
rect 464370 231662 464752 231690
rect 462688 226296 462740 226302
rect 462688 226238 462740 226244
rect 462320 219836 462372 219842
rect 462320 219778 462372 219784
rect 462332 219434 462360 219778
rect 463528 219706 463556 231662
rect 464172 229226 464200 231662
rect 463700 229220 463752 229226
rect 463700 229162 463752 229168
rect 464160 229220 464212 229226
rect 464160 229162 464212 229168
rect 463712 220930 463740 229162
rect 464724 225486 464752 231662
rect 464908 229094 464936 231676
rect 465474 231662 465856 231690
rect 464908 229066 465028 229094
rect 464528 225480 464580 225486
rect 464528 225422 464580 225428
rect 464712 225480 464764 225486
rect 464712 225422 464764 225428
rect 464540 225298 464568 225422
rect 464540 225270 464844 225298
rect 464620 221468 464672 221474
rect 464620 221410 464672 221416
rect 463700 220924 463752 220930
rect 463700 220866 463752 220872
rect 463516 219700 463568 219706
rect 463516 219642 463568 219648
rect 462320 219428 462372 219434
rect 462320 219370 462372 219376
rect 463792 218884 463844 218890
rect 463792 218826 463844 218832
rect 462964 218340 463016 218346
rect 462964 218282 463016 218288
rect 461320 217246 461394 217274
rect 462148 217246 462222 217274
rect 457226 216988 457254 217110
rect 458054 216988 458082 217126
rect 458836 217110 458910 217138
rect 459664 217110 459738 217138
rect 460492 217110 460566 217138
rect 458882 216988 458910 217110
rect 459710 216988 459738 217110
rect 460538 216988 460566 217110
rect 461366 216988 461394 217246
rect 462194 216988 462222 217246
rect 462976 217138 463004 218282
rect 463804 217138 463832 218826
rect 464632 217274 464660 221410
rect 464816 218346 464844 225270
rect 465000 219842 465028 229066
rect 465264 228948 465316 228954
rect 465264 228890 465316 228896
rect 464988 219836 465040 219842
rect 464988 219778 465040 219784
rect 464804 218340 464856 218346
rect 464804 218282 464856 218288
rect 465276 217274 465304 228890
rect 465828 222766 465856 231662
rect 466012 225078 466040 231676
rect 466564 229226 466592 231676
rect 467130 231662 467512 231690
rect 466368 229220 466420 229226
rect 466368 229162 466420 229168
rect 466552 229220 466604 229226
rect 466552 229162 466604 229168
rect 466380 228274 466408 229162
rect 466184 228268 466236 228274
rect 466184 228210 466236 228216
rect 466368 228268 466420 228274
rect 466368 228210 466420 228216
rect 466000 225072 466052 225078
rect 466000 225014 466052 225020
rect 465816 222760 465868 222766
rect 465816 222702 465868 222708
rect 466196 219434 466224 228210
rect 467288 226024 467340 226030
rect 467288 225966 467340 225972
rect 467104 223440 467156 223446
rect 467104 223382 467156 223388
rect 466196 219406 466316 219434
rect 466288 217274 466316 219406
rect 467116 217274 467144 223382
rect 467300 219026 467328 225966
rect 467484 222630 467512 231662
rect 467668 225894 467696 231676
rect 468220 228818 468248 231676
rect 468024 228812 468076 228818
rect 468024 228754 468076 228760
rect 468208 228812 468260 228818
rect 468208 228754 468260 228760
rect 467656 225888 467708 225894
rect 467656 225830 467708 225836
rect 467472 222624 467524 222630
rect 467472 222566 467524 222572
rect 467288 219020 467340 219026
rect 467288 218962 467340 218968
rect 468036 217274 468064 228754
rect 468772 223446 468800 231676
rect 469324 226030 469352 231676
rect 469508 231662 469890 231690
rect 469312 226024 469364 226030
rect 469312 225966 469364 225972
rect 469312 225752 469364 225758
rect 469312 225694 469364 225700
rect 468760 223440 468812 223446
rect 468760 223382 468812 223388
rect 468760 218476 468812 218482
rect 468760 218418 468812 218424
rect 464632 217246 464706 217274
rect 465276 217246 465534 217274
rect 466288 217246 466362 217274
rect 467116 217246 467190 217274
rect 462976 217110 463050 217138
rect 463804 217110 463878 217138
rect 463022 216988 463050 217110
rect 463850 216988 463878 217110
rect 464678 216988 464706 217246
rect 465506 216988 465534 217246
rect 466334 216988 466362 217246
rect 467162 216988 467190 217246
rect 467990 217246 468064 217274
rect 467990 216988 468018 217246
rect 468772 217138 468800 218418
rect 469324 217190 469352 225694
rect 469508 219978 469536 231662
rect 470428 223310 470456 231676
rect 470784 229220 470836 229226
rect 470784 229162 470836 229168
rect 470796 226914 470824 229162
rect 470784 226908 470836 226914
rect 470784 226850 470836 226856
rect 470980 224942 471008 231676
rect 471244 227452 471296 227458
rect 471244 227394 471296 227400
rect 470968 224936 471020 224942
rect 470968 224878 471020 224884
rect 469864 223304 469916 223310
rect 469864 223246 469916 223252
rect 470416 223304 470468 223310
rect 470416 223246 470468 223252
rect 469496 219972 469548 219978
rect 469496 219914 469548 219920
rect 469876 218890 469904 223246
rect 471060 219292 471112 219298
rect 471060 219234 471112 219240
rect 469864 218884 469916 218890
rect 469864 218826 469916 218832
rect 469588 218612 469640 218618
rect 469588 218554 469640 218560
rect 469312 217184 469364 217190
rect 468772 217110 468846 217138
rect 469312 217126 469364 217132
rect 469600 217138 469628 218554
rect 471072 218074 471100 219234
rect 471060 218068 471112 218074
rect 471060 218010 471112 218016
rect 471256 217274 471284 227394
rect 471532 227322 471560 231676
rect 472084 229094 472112 231676
rect 471992 229066 472112 229094
rect 471520 227316 471572 227322
rect 471520 227258 471572 227264
rect 471428 223032 471480 223038
rect 471428 222974 471480 222980
rect 471440 219298 471468 222974
rect 471992 222902 472020 229066
rect 472164 227180 472216 227186
rect 472164 227122 472216 227128
rect 471980 222896 472032 222902
rect 471980 222838 472032 222844
rect 471428 219292 471480 219298
rect 471428 219234 471480 219240
rect 472176 217274 472204 227122
rect 472636 225758 472664 231676
rect 472624 225752 472676 225758
rect 472624 225694 472676 225700
rect 472624 225616 472676 225622
rect 472624 225558 472676 225564
rect 472636 218482 472664 225558
rect 473188 220522 473216 231676
rect 473452 229900 473504 229906
rect 473452 229842 473504 229848
rect 473464 229226 473492 229842
rect 473452 229220 473504 229226
rect 473452 229162 473504 229168
rect 473740 227458 473768 231676
rect 473728 227452 473780 227458
rect 473728 227394 473780 227400
rect 474292 227186 474320 231676
rect 474858 231662 475240 231690
rect 475212 230790 475240 231662
rect 475200 230784 475252 230790
rect 475200 230726 475252 230732
rect 475200 230172 475252 230178
rect 475200 230114 475252 230120
rect 475212 229906 475240 230114
rect 475200 229900 475252 229906
rect 475200 229842 475252 229848
rect 475396 228682 475424 231676
rect 475200 228676 475252 228682
rect 475200 228618 475252 228624
rect 475384 228676 475436 228682
rect 475384 228618 475436 228624
rect 474280 227180 474332 227186
rect 474280 227122 474332 227128
rect 473728 227044 473780 227050
rect 473728 226986 473780 226992
rect 473176 220516 473228 220522
rect 473176 220458 473228 220464
rect 472900 219156 472952 219162
rect 472900 219098 472952 219104
rect 472624 218476 472676 218482
rect 472624 218418 472676 218424
rect 471256 217246 471330 217274
rect 470462 217184 470514 217190
rect 469600 217110 469674 217138
rect 470462 217126 470514 217132
rect 468818 216988 468846 217110
rect 469646 216988 469674 217110
rect 470474 216988 470502 217126
rect 471302 216988 471330 217246
rect 472130 217246 472204 217274
rect 472130 216988 472158 217246
rect 472912 217138 472940 219098
rect 473740 217274 473768 226986
rect 474648 223576 474700 223582
rect 474648 223518 474700 223524
rect 474660 219586 474688 223518
rect 474660 219558 474780 219586
rect 474752 219434 474780 219558
rect 475212 219434 475240 228618
rect 475948 225622 475976 231676
rect 476500 230178 476528 231676
rect 476488 230172 476540 230178
rect 476488 230114 476540 230120
rect 476396 229220 476448 229226
rect 476396 229162 476448 229168
rect 476212 227724 476264 227730
rect 476212 227666 476264 227672
rect 475936 225616 475988 225622
rect 475936 225558 475988 225564
rect 474556 219428 474608 219434
rect 474556 219370 474608 219376
rect 474740 219428 474792 219434
rect 475212 219406 475424 219434
rect 474740 219370 474792 219376
rect 473740 217246 473814 217274
rect 472912 217110 472986 217138
rect 472958 216988 472986 217110
rect 473786 216988 473814 217246
rect 474568 217138 474596 219370
rect 475108 219156 475160 219162
rect 475108 219098 475160 219104
rect 474924 218884 474976 218890
rect 474924 218826 474976 218832
rect 474936 218346 474964 218826
rect 475120 218754 475148 219098
rect 475108 218748 475160 218754
rect 475108 218690 475160 218696
rect 474924 218340 474976 218346
rect 474924 218282 474976 218288
rect 475396 217274 475424 219406
rect 475752 219292 475804 219298
rect 475752 219234 475804 219240
rect 475764 218618 475792 219234
rect 475752 218612 475804 218618
rect 475752 218554 475804 218560
rect 476224 217274 476252 227666
rect 476408 219434 476436 229162
rect 477052 223582 477080 231676
rect 477604 228954 477632 231676
rect 477788 231662 478170 231690
rect 477592 228948 477644 228954
rect 477592 228890 477644 228896
rect 477592 226636 477644 226642
rect 477592 226578 477644 226584
rect 477040 223576 477092 223582
rect 477040 223518 477092 223524
rect 476408 219406 477080 219434
rect 477052 217274 477080 219406
rect 475396 217246 475470 217274
rect 476224 217246 476298 217274
rect 477052 217246 477126 217274
rect 474568 217110 474642 217138
rect 474614 216988 474642 217110
rect 475442 216988 475470 217246
rect 476270 216988 476298 217246
rect 477098 216988 477126 217246
rect 477604 217190 477632 226578
rect 477788 220386 477816 231662
rect 478708 223038 478736 231676
rect 479260 229226 479288 231676
rect 479524 230172 479576 230178
rect 479524 230114 479576 230120
rect 479248 229220 479300 229226
rect 479248 229162 479300 229168
rect 478696 223032 478748 223038
rect 478696 222974 478748 222980
rect 479536 220658 479564 230114
rect 479812 227050 479840 231676
rect 479984 230784 480036 230790
rect 479984 230726 480036 230732
rect 479996 230178 480024 230726
rect 479984 230172 480036 230178
rect 479984 230114 480036 230120
rect 480166 229392 480222 229401
rect 480166 229327 480168 229336
rect 480220 229327 480222 229336
rect 480168 229298 480220 229304
rect 479800 227044 479852 227050
rect 479800 226986 479852 226992
rect 480364 224806 480392 231676
rect 480930 231662 481312 231690
rect 481284 230790 481312 231662
rect 481272 230784 481324 230790
rect 481272 230726 481324 230732
rect 481468 230330 481496 231676
rect 481468 230302 481588 230330
rect 481364 230172 481416 230178
rect 481364 230114 481416 230120
rect 480534 229392 480590 229401
rect 480534 229327 480536 229336
rect 480588 229327 480590 229336
rect 480536 229298 480588 229304
rect 481376 227866 481404 230114
rect 481364 227860 481416 227866
rect 481364 227802 481416 227808
rect 480352 224800 480404 224806
rect 480352 224742 480404 224748
rect 478788 220652 478840 220658
rect 478788 220594 478840 220600
rect 479524 220652 479576 220658
rect 479524 220594 479576 220600
rect 477776 220380 477828 220386
rect 477776 220322 477828 220328
rect 478800 218385 478828 220594
rect 481560 220250 481588 230302
rect 481732 229356 481784 229362
rect 481732 229298 481784 229304
rect 481744 226642 481772 229298
rect 481732 226636 481784 226642
rect 481732 226578 481784 226584
rect 482020 224534 482048 231676
rect 482572 230178 482600 231676
rect 483138 231662 483336 231690
rect 482560 230172 482612 230178
rect 482560 230114 482612 230120
rect 481824 224528 481876 224534
rect 481824 224470 481876 224476
rect 482008 224528 482060 224534
rect 482008 224470 482060 224476
rect 481836 224233 481864 224470
rect 481822 224224 481878 224233
rect 481822 224159 481878 224168
rect 482650 224224 482706 224233
rect 482650 224159 482706 224168
rect 480260 220244 480312 220250
rect 480260 220186 480312 220192
rect 481548 220244 481600 220250
rect 481548 220186 481600 220192
rect 480272 219298 480300 220186
rect 480260 219292 480312 219298
rect 480260 219234 480312 219240
rect 482664 218754 482692 224159
rect 483018 223034 483074 223043
rect 483018 222969 483074 222978
rect 483308 220153 483336 231662
rect 483676 226273 483704 231676
rect 484228 229906 484256 231676
rect 484504 231662 484794 231690
rect 484032 229900 484084 229906
rect 484032 229842 484084 229848
rect 484216 229900 484268 229906
rect 484216 229842 484268 229848
rect 484044 226438 484072 229842
rect 484032 226432 484084 226438
rect 484032 226374 484084 226380
rect 483662 226264 483718 226273
rect 483662 226199 483718 226208
rect 484306 225992 484362 226001
rect 484306 225927 484362 225936
rect 483664 224800 483716 224806
rect 483662 224768 483664 224777
rect 483716 224768 483718 224777
rect 483662 224703 483718 224712
rect 484124 223576 484176 223582
rect 484124 223518 484176 223524
rect 484136 223038 484164 223518
rect 484124 223032 484176 223038
rect 484124 222974 484176 222980
rect 483294 220144 483350 220153
rect 483294 220079 483350 220088
rect 484320 219298 484348 225927
rect 484504 221474 484532 231662
rect 484860 229764 484912 229770
rect 484860 229706 484912 229712
rect 485044 229764 485096 229770
rect 485044 229706 485096 229712
rect 484872 229362 484900 229706
rect 484860 229356 484912 229362
rect 484860 229298 484912 229304
rect 485056 229226 485084 229706
rect 485044 229220 485096 229226
rect 485044 229162 485096 229168
rect 485332 227769 485360 231676
rect 485884 229226 485912 231676
rect 486068 231662 486450 231690
rect 485872 229220 485924 229226
rect 485872 229162 485924 229168
rect 485318 227760 485374 227769
rect 485318 227695 485374 227704
rect 486068 224954 486096 231662
rect 486068 224926 486648 224954
rect 485872 224800 485924 224806
rect 486240 224800 486292 224806
rect 485872 224742 485924 224748
rect 486238 224768 486240 224777
rect 486292 224768 486294 224777
rect 484860 224528 484912 224534
rect 484858 224496 484860 224505
rect 485884 224505 485912 224742
rect 486238 224703 486294 224712
rect 484912 224496 484914 224505
rect 484858 224431 484914 224440
rect 485870 224496 485926 224505
rect 485870 224431 485926 224440
rect 485044 224392 485096 224398
rect 485044 224334 485096 224340
rect 484676 224256 484728 224262
rect 484676 224198 484728 224204
rect 484688 222601 484716 224198
rect 484674 222592 484730 222601
rect 484674 222527 484730 222536
rect 484492 221468 484544 221474
rect 484492 221410 484544 221416
rect 483572 219292 483624 219298
rect 483572 219234 483624 219240
rect 483756 219292 483808 219298
rect 483756 219234 483808 219240
rect 484308 219292 484360 219298
rect 484308 219234 484360 219240
rect 482836 219156 482888 219162
rect 482836 219098 482888 219104
rect 481180 218748 481232 218754
rect 481180 218690 481232 218696
rect 482652 218748 482704 218754
rect 482652 218690 482704 218696
rect 480444 218612 480496 218618
rect 480444 218554 480496 218560
rect 478786 218376 478842 218385
rect 478786 218311 478842 218320
rect 477868 218068 477920 218074
rect 477868 218010 477920 218016
rect 479616 218068 479668 218074
rect 479616 218010 479668 218016
rect 477592 217184 477644 217190
rect 477592 217126 477644 217132
rect 477880 217138 477908 218010
rect 478742 217184 478794 217190
rect 477880 217110 477954 217138
rect 479628 217138 479656 218010
rect 480456 217274 480484 218554
rect 478742 217126 478794 217132
rect 477926 216988 477954 217110
rect 478754 216988 478782 217126
rect 479582 217110 479656 217138
rect 480410 217246 480484 217274
rect 481192 217274 481220 218690
rect 482190 218376 482246 218385
rect 482008 218340 482060 218346
rect 482190 218311 482192 218320
rect 482008 218282 482060 218288
rect 482244 218311 482246 218320
rect 482192 218282 482244 218288
rect 482020 217274 482048 218282
rect 482848 217274 482876 219098
rect 481192 217246 481266 217274
rect 482020 217246 482094 217274
rect 482848 217246 482922 217274
rect 479582 216988 479610 217110
rect 480410 216988 480438 217246
rect 481238 216988 481266 217246
rect 482066 216988 482094 217246
rect 482894 216988 482922 217246
rect 483584 217122 483612 219234
rect 483768 217274 483796 219234
rect 485056 219162 485084 224334
rect 485688 223984 485740 223990
rect 485872 223984 485924 223990
rect 485740 223932 485872 223938
rect 485688 223926 485924 223932
rect 485700 223910 485912 223926
rect 485688 223848 485740 223854
rect 485872 223848 485924 223854
rect 485740 223796 485872 223802
rect 485688 223790 485924 223796
rect 485700 223774 485912 223790
rect 486238 222592 486294 222601
rect 486238 222527 486294 222536
rect 485870 220144 485926 220153
rect 485734 220108 485786 220114
rect 485870 220079 485872 220088
rect 485734 220050 485786 220056
rect 485924 220079 485926 220088
rect 485872 220050 485924 220056
rect 485746 219994 485774 220050
rect 485746 219966 485912 219994
rect 485044 219156 485096 219162
rect 485044 219098 485096 219104
rect 485884 219026 485912 219966
rect 486252 219314 486280 222527
rect 486620 221610 486648 224926
rect 486792 224324 486844 224330
rect 486792 224266 486844 224272
rect 486804 223417 486832 224266
rect 486988 224262 487016 231676
rect 487540 229906 487568 231676
rect 487344 229900 487396 229906
rect 487344 229842 487396 229848
rect 487528 229900 487580 229906
rect 487528 229842 487580 229848
rect 487356 229401 487384 229842
rect 487342 229392 487398 229401
rect 487342 229327 487398 229336
rect 487620 227724 487672 227730
rect 487620 227666 487672 227672
rect 486976 224256 487028 224262
rect 486976 224198 487028 224204
rect 487068 223576 487120 223582
rect 487068 223518 487120 223524
rect 486790 223408 486846 223417
rect 486790 223343 486846 223352
rect 487080 223145 487108 223518
rect 487066 223136 487122 223145
rect 487066 223071 487122 223080
rect 486608 221604 486660 221610
rect 486608 221546 486660 221552
rect 486252 219286 486556 219314
rect 486148 219156 486200 219162
rect 486148 219098 486200 219104
rect 485412 219020 485464 219026
rect 485412 218962 485464 218968
rect 485872 219020 485924 219026
rect 485872 218962 485924 218968
rect 485424 218890 485452 218962
rect 485412 218884 485464 218890
rect 485412 218826 485464 218832
rect 484582 218648 484638 218657
rect 484582 218583 484638 218592
rect 484596 218113 484624 218583
rect 484582 218104 484638 218113
rect 484582 218039 484638 218048
rect 484596 217274 484624 218039
rect 485424 217274 485452 218826
rect 483722 217246 483796 217274
rect 484550 217246 484624 217274
rect 485378 217246 485452 217274
rect 483572 217116 483624 217122
rect 483572 217058 483624 217064
rect 483722 216988 483750 217246
rect 484550 216988 484578 217246
rect 485378 216988 485406 217246
rect 486160 217138 486188 219098
rect 486528 217938 486556 219286
rect 486976 218748 487028 218754
rect 486976 218690 487028 218696
rect 486516 217932 486568 217938
rect 486516 217874 486568 217880
rect 486988 217138 487016 218690
rect 487632 218521 487660 227666
rect 488092 226001 488120 231676
rect 489828 230784 489880 230790
rect 489828 230726 489880 230732
rect 489552 229356 489604 229362
rect 489552 229298 489604 229304
rect 489564 227730 489592 229298
rect 489840 229242 489868 230726
rect 495438 230344 495494 230353
rect 495438 230279 495494 230288
rect 499854 230344 499910 230353
rect 499854 230279 499910 230288
rect 505744 230308 505796 230314
rect 495452 229786 495480 230279
rect 499488 229900 499540 229906
rect 499488 229842 499540 229848
rect 495406 229770 495480 229786
rect 495394 229764 495480 229770
rect 495446 229758 495480 229764
rect 495394 229706 495446 229712
rect 499120 229696 499172 229702
rect 499120 229638 499172 229644
rect 495440 229628 495492 229634
rect 495440 229570 495492 229576
rect 490194 229528 490250 229537
rect 490024 229486 490194 229514
rect 490024 229362 490052 229486
rect 495452 229514 495480 229570
rect 495622 229528 495678 229537
rect 495452 229486 495622 229514
rect 490194 229463 490250 229472
rect 495622 229463 495678 229472
rect 495900 229492 495952 229498
rect 495900 229434 495952 229440
rect 490012 229356 490064 229362
rect 490012 229298 490064 229304
rect 490196 229356 490248 229362
rect 490196 229298 490248 229304
rect 489840 229226 489960 229242
rect 489840 229220 489972 229226
rect 489840 229214 489920 229220
rect 489920 229162 489972 229168
rect 490208 229129 490236 229298
rect 495912 229265 495940 229434
rect 499132 229378 499160 229638
rect 499500 229498 499528 229842
rect 499868 229634 499896 230279
rect 505744 230250 505796 230256
rect 499856 229628 499908 229634
rect 499856 229570 499908 229576
rect 502984 229628 503036 229634
rect 502984 229570 503036 229576
rect 504192 229622 504588 229650
rect 499670 229528 499726 229537
rect 499488 229492 499540 229498
rect 499670 229463 499672 229472
rect 499488 229434 499540 229440
rect 499724 229463 499726 229472
rect 502524 229492 502576 229498
rect 499672 229434 499724 229440
rect 502524 229434 502576 229440
rect 499132 229350 499620 229378
rect 495898 229256 495954 229265
rect 495898 229191 495954 229200
rect 490194 229120 490250 229129
rect 490194 229055 490250 229064
rect 495636 228954 496032 228970
rect 495394 228948 495446 228954
rect 495394 228890 495446 228896
rect 495636 228948 496044 228954
rect 495636 228942 495992 228948
rect 489918 228848 489974 228857
rect 495406 228834 495434 228890
rect 495406 228806 495480 228834
rect 489918 228783 489974 228792
rect 489932 227882 489960 228783
rect 495452 227905 495480 228806
rect 495636 228682 495664 228942
rect 495992 228890 496044 228896
rect 495806 228848 495862 228857
rect 495806 228783 495862 228792
rect 495820 228682 495848 228783
rect 495624 228676 495676 228682
rect 495624 228618 495676 228624
rect 495808 228676 495860 228682
rect 495808 228618 495860 228624
rect 489886 227866 489960 227882
rect 489874 227860 489960 227866
rect 489926 227854 489960 227860
rect 495438 227896 495494 227905
rect 495438 227831 495494 227840
rect 489874 227802 489926 227808
rect 490746 227760 490802 227769
rect 489552 227724 489604 227730
rect 490746 227695 490802 227704
rect 489552 227666 489604 227672
rect 488078 225992 488134 226001
rect 488078 225927 488134 225936
rect 487988 224528 488040 224534
rect 487988 224470 488040 224476
rect 488000 224126 488028 224470
rect 487988 224120 488040 224126
rect 487988 224062 488040 224068
rect 489368 219428 489420 219434
rect 489368 219370 489420 219376
rect 487894 218784 487950 218793
rect 487894 218719 487896 218728
rect 487948 218719 487950 218728
rect 487896 218690 487948 218696
rect 487618 218512 487674 218521
rect 487618 218447 487674 218456
rect 487908 217138 487936 218690
rect 489380 217274 489408 219370
rect 489564 219201 489592 227666
rect 489874 226296 489926 226302
rect 489926 226244 490052 226250
rect 489874 226238 490052 226244
rect 489886 226222 490052 226238
rect 490024 226030 490052 226222
rect 489874 226024 489926 226030
rect 489872 225992 489874 226001
rect 490012 226024 490064 226030
rect 489926 225992 489928 226001
rect 490012 225966 490064 225972
rect 489872 225927 489928 225936
rect 490760 224398 490788 227695
rect 491942 226264 491998 226273
rect 491942 226199 491998 226208
rect 491956 224534 491984 226199
rect 493874 225312 493930 225321
rect 493874 225247 493930 225256
rect 491944 224528 491996 224534
rect 491944 224470 491996 224476
rect 490748 224392 490800 224398
rect 490748 224334 490800 224340
rect 491208 221060 491260 221066
rect 491208 221002 491260 221008
rect 490196 219360 490248 219366
rect 490196 219302 490248 219308
rect 490380 219360 490432 219366
rect 490380 219302 490432 219308
rect 489828 219224 489880 219230
rect 489550 219192 489606 219201
rect 489828 219166 489880 219172
rect 489550 219127 489606 219136
rect 489840 218113 489868 219166
rect 489826 218104 489882 218113
rect 490208 218090 490236 219302
rect 490392 218754 490420 219302
rect 491220 219178 491248 221002
rect 491220 219150 491524 219178
rect 491496 219094 491524 219150
rect 491484 219088 491536 219094
rect 491484 219030 491536 219036
rect 491300 219020 491352 219026
rect 491300 218962 491352 218968
rect 491312 218754 491340 218962
rect 490380 218748 490432 218754
rect 490380 218690 490432 218696
rect 491300 218748 491352 218754
rect 491300 218690 491352 218696
rect 491114 218512 491170 218521
rect 490346 218482 490972 218498
rect 490334 218476 490972 218482
rect 490386 218470 490972 218476
rect 490334 218418 490386 218424
rect 490562 218240 490618 218249
rect 490944 218210 490972 218470
rect 491114 218447 491170 218456
rect 491300 218476 491352 218482
rect 490562 218175 490564 218184
rect 490616 218175 490618 218184
rect 490932 218204 490984 218210
rect 490564 218146 490616 218152
rect 490932 218146 490984 218152
rect 490378 218104 490434 218113
rect 490208 218062 490378 218090
rect 489826 218039 489882 218048
rect 490378 218039 490434 218048
rect 489380 217246 489546 217274
rect 486160 217110 486234 217138
rect 486988 217110 487062 217138
rect 486206 216988 486234 217110
rect 487034 216988 487062 217110
rect 487862 217110 487936 217138
rect 488678 217116 488730 217122
rect 487862 216988 487890 217110
rect 488678 217058 488730 217064
rect 488690 216988 488718 217058
rect 489518 216988 489546 217246
rect 490392 217138 490420 218039
rect 491128 217297 491156 218447
rect 491300 218418 491352 218424
rect 491312 218249 491340 218418
rect 491944 218340 491996 218346
rect 491944 218282 491996 218288
rect 491298 218240 491354 218249
rect 491298 218175 491354 218184
rect 491114 217288 491170 217297
rect 491114 217223 491170 217232
rect 490346 217110 490420 217138
rect 491128 217138 491156 217223
rect 491390 217152 491446 217161
rect 491128 217110 491202 217138
rect 490346 216988 490374 217110
rect 491174 216988 491202 217110
rect 491956 217138 491984 218282
rect 493888 218210 493916 225247
rect 499592 224954 499620 229350
rect 499592 224926 499988 224954
rect 496084 223712 496136 223718
rect 496084 223654 496136 223660
rect 494426 219192 494482 219201
rect 494426 219127 494482 219136
rect 493692 218204 493744 218210
rect 493692 218146 493744 218152
rect 493876 218204 493928 218210
rect 493876 218146 493928 218152
rect 493704 217977 493732 218146
rect 493690 217968 493746 217977
rect 492772 217932 492824 217938
rect 493690 217903 493746 217912
rect 492772 217874 492824 217880
rect 492784 217138 492812 217874
rect 493704 217138 493732 217903
rect 491956 217110 492030 217138
rect 492784 217110 492858 217138
rect 491390 217087 491392 217096
rect 491444 217087 491446 217096
rect 491392 217058 491444 217064
rect 492002 216988 492030 217110
rect 492830 216988 492858 217110
rect 493658 217110 493732 217138
rect 494440 217138 494468 219127
rect 495256 219088 495308 219094
rect 495256 219030 495308 219036
rect 495268 217297 495296 219030
rect 495254 217288 495310 217297
rect 496096 217274 496124 223654
rect 498198 223408 498254 223417
rect 498198 223343 498254 223352
rect 497740 218476 497792 218482
rect 497740 218418 497792 218424
rect 496912 218204 496964 218210
rect 496912 218146 496964 218152
rect 496096 217246 496170 217274
rect 495254 217223 495310 217232
rect 495268 217138 495296 217223
rect 494440 217110 494514 217138
rect 495268 217110 495342 217138
rect 493658 216988 493686 217110
rect 494486 216988 494514 217110
rect 495314 216988 495342 217110
rect 496142 216988 496170 217246
rect 496924 217138 496952 218146
rect 497752 217138 497780 218418
rect 498212 217190 498240 223343
rect 499960 219434 499988 224926
rect 502536 223145 502564 229434
rect 502522 223136 502578 223145
rect 502522 223071 502578 223080
rect 501052 221196 501104 221202
rect 501052 221138 501104 221144
rect 499592 219406 499988 219434
rect 499592 219065 499620 219406
rect 499578 219056 499634 219065
rect 498384 219020 498436 219026
rect 499578 218991 499634 219000
rect 500222 219056 500278 219065
rect 500222 218991 500278 219000
rect 498384 218962 498436 218968
rect 498396 218754 498424 218962
rect 498384 218748 498436 218754
rect 498752 218748 498804 218754
rect 498436 218708 498608 218736
rect 498384 218690 498436 218696
rect 498580 217274 498608 218708
rect 498752 218690 498804 218696
rect 498764 218482 498792 218690
rect 498752 218476 498804 218482
rect 498752 218418 498804 218424
rect 498580 217246 498654 217274
rect 498200 217184 498252 217190
rect 496924 217110 496998 217138
rect 497752 217110 497826 217138
rect 498200 217126 498252 217132
rect 496970 216988 496998 217110
rect 497798 216988 497826 217110
rect 498626 216988 498654 217246
rect 499442 217184 499494 217190
rect 499442 217126 499494 217132
rect 500236 217138 500264 218991
rect 501064 217308 501092 221138
rect 502536 219434 502564 223071
rect 502536 219406 502748 219434
rect 501880 217592 501932 217598
rect 501234 217560 501290 217569
rect 501880 217534 501932 217540
rect 501234 217495 501290 217504
rect 501248 217308 501276 217495
rect 501064 217280 501276 217308
rect 499454 216988 499482 217126
rect 500236 217110 500310 217138
rect 500282 216988 500310 217110
rect 501110 216988 501138 217280
rect 501892 217138 501920 217534
rect 502720 217308 502748 219406
rect 502996 218618 503024 229570
rect 504192 229498 504220 229622
rect 504180 229492 504232 229498
rect 504180 229434 504232 229440
rect 504364 229492 504416 229498
rect 504364 229434 504416 229440
rect 503536 221332 503588 221338
rect 503536 221274 503588 221280
rect 503548 220017 503576 221274
rect 503534 220008 503590 220017
rect 503534 219943 503590 219952
rect 502984 218612 503036 218618
rect 502984 218554 503036 218560
rect 503352 218340 503404 218346
rect 503352 218282 503404 218288
rect 503364 217569 503392 218282
rect 503350 217560 503406 217569
rect 503350 217495 503406 217504
rect 503548 217308 503576 219943
rect 504376 218074 504404 229434
rect 504560 221338 504588 229622
rect 505098 228848 505154 228857
rect 505098 228783 505154 228792
rect 505112 228698 505140 228783
rect 505066 228670 505140 228698
rect 505066 228546 505094 228670
rect 505054 228540 505106 228546
rect 505054 228482 505106 228488
rect 505192 228540 505244 228546
rect 505192 228482 505244 228488
rect 504914 227896 504970 227905
rect 505204 227882 505232 228482
rect 504970 227854 505232 227882
rect 504914 227831 504970 227840
rect 505098 226400 505154 226409
rect 505098 226335 505154 226344
rect 505112 226114 505140 226335
rect 505066 226086 505140 226114
rect 505066 226030 505094 226086
rect 505054 226024 505106 226030
rect 504914 225992 504970 226001
rect 505054 225966 505106 225972
rect 505192 226024 505244 226030
rect 505192 225966 505244 225972
rect 504914 225927 504970 225936
rect 504928 225842 504956 225927
rect 505204 225842 505232 225966
rect 504928 225814 505232 225842
rect 504732 225616 504784 225622
rect 504730 225584 504732 225593
rect 505192 225616 505244 225622
rect 504784 225584 504786 225593
rect 504730 225519 504786 225528
rect 505190 225584 505192 225593
rect 505244 225584 505246 225593
rect 505190 225519 505246 225528
rect 505008 223712 505060 223718
rect 505008 223654 505060 223660
rect 504548 221332 504600 221338
rect 504548 221274 504600 221280
rect 505020 220794 505048 223654
rect 505008 220788 505060 220794
rect 505008 220730 505060 220736
rect 505756 218657 505784 230250
rect 507124 230036 507176 230042
rect 507124 229978 507176 229984
rect 506020 220788 506072 220794
rect 506020 220730 506072 220736
rect 505742 218648 505798 218657
rect 505742 218583 505798 218592
rect 504364 218068 504416 218074
rect 504364 218010 504416 218016
rect 504364 217456 504416 217462
rect 504364 217398 504416 217404
rect 502720 217280 502794 217308
rect 503548 217280 503622 217308
rect 501892 217110 501966 217138
rect 501938 216988 501966 217110
rect 502766 216988 502794 217280
rect 503594 216988 503622 217280
rect 504376 217138 504404 217398
rect 505756 217308 505784 218583
rect 505250 217280 505784 217308
rect 506032 217308 506060 220730
rect 506848 219564 506900 219570
rect 506848 219506 506900 219512
rect 506860 217308 506888 219506
rect 507136 218113 507164 229978
rect 507504 229498 507532 232999
rect 510620 230648 510672 230654
rect 510620 230590 510672 230596
rect 507492 229492 507544 229498
rect 507492 229434 507544 229440
rect 507952 228948 508004 228954
rect 507952 228890 508004 228896
rect 508136 228948 508188 228954
rect 508136 228890 508188 228896
rect 507964 228682 507992 228890
rect 507952 228676 508004 228682
rect 507952 228618 508004 228624
rect 508148 228562 508176 228890
rect 507504 228546 508176 228562
rect 507492 228540 508176 228546
rect 507544 228534 508176 228540
rect 507492 228482 507544 228488
rect 509608 226432 509660 226438
rect 510160 226432 510212 226438
rect 509608 226374 509660 226380
rect 510158 226400 510160 226409
rect 510212 226400 510214 226409
rect 509620 226030 509648 226374
rect 510158 226335 510214 226344
rect 509608 226024 509660 226030
rect 509608 225966 509660 225972
rect 510158 222864 510214 222873
rect 510158 222799 510214 222808
rect 509194 222012 509246 222018
rect 509194 221954 509246 221960
rect 509206 221898 509234 221954
rect 509206 221870 509280 221898
rect 509252 221202 509280 221870
rect 509240 221196 509292 221202
rect 509240 221138 509292 221144
rect 508596 220924 508648 220930
rect 508596 220866 508648 220872
rect 508318 218648 508374 218657
rect 508318 218583 508374 218592
rect 508332 218113 508360 218583
rect 507122 218104 507178 218113
rect 507122 218039 507178 218048
rect 507674 218104 507730 218113
rect 507674 218039 507730 218048
rect 508318 218104 508374 218113
rect 508318 218039 508374 218048
rect 506032 217280 506106 217308
rect 506860 217280 506934 217308
rect 504376 217110 504450 217138
rect 504422 216988 504450 217110
rect 505250 216988 505278 217280
rect 506078 216988 506106 217280
rect 506906 216988 506934 217280
rect 507688 217138 507716 218039
rect 508608 217308 508636 220866
rect 510172 218657 510200 222799
rect 510158 218648 510214 218657
rect 510158 218583 510214 218592
rect 508562 217280 508636 217308
rect 507688 217110 507762 217138
rect 507734 216988 507762 217110
rect 508562 216988 508590 217280
rect 510172 217274 510200 218583
rect 509378 217252 509430 217258
rect 510172 217246 510246 217274
rect 510632 217258 510660 230590
rect 511276 229634 511304 238167
rect 512656 238066 512684 247114
rect 514036 238202 514064 259422
rect 567200 256760 567252 256766
rect 567200 256702 567252 256708
rect 559564 252612 559616 252618
rect 559564 252554 559616 252560
rect 514024 238196 514076 238202
rect 514024 238138 514076 238144
rect 512644 238060 512696 238066
rect 512644 238002 512696 238008
rect 512736 230512 512788 230518
rect 512736 230454 512788 230460
rect 511264 229628 511316 229634
rect 511264 229570 511316 229576
rect 511264 223576 511316 223582
rect 511264 223518 511316 223524
rect 511276 222222 511304 223518
rect 511264 222216 511316 222222
rect 511264 222158 511316 222164
rect 511080 221196 511132 221202
rect 511080 221138 511132 221144
rect 511092 219502 511120 221138
rect 511080 219496 511132 219502
rect 511080 219438 511132 219444
rect 511092 217274 511120 219438
rect 512748 218929 512776 230454
rect 541992 230172 542044 230178
rect 541992 230114 542044 230120
rect 536840 229356 536892 229362
rect 536840 229298 536892 229304
rect 533344 229220 533396 229226
rect 533344 229162 533396 229168
rect 525984 229084 526036 229090
rect 525984 229026 526036 229032
rect 513562 228848 513618 228857
rect 513562 228783 513618 228792
rect 513576 220998 513604 228783
rect 520924 228132 520976 228138
rect 520924 228074 520976 228080
rect 517796 227996 517848 228002
rect 517796 227938 517848 227944
rect 515956 226636 516008 226642
rect 515956 226578 516008 226584
rect 514576 226296 514628 226302
rect 514576 226238 514628 226244
rect 514588 226114 514616 226238
rect 514588 226086 514754 226114
rect 514726 226030 514754 226086
rect 514576 226024 514628 226030
rect 514574 225992 514576 226001
rect 514714 226024 514766 226030
rect 514628 225992 514630 226001
rect 514714 225966 514766 225972
rect 514574 225927 514630 225936
rect 515128 223848 515180 223854
rect 515128 223790 515180 223796
rect 514300 222080 514352 222086
rect 514300 222022 514352 222028
rect 513564 220992 513616 220998
rect 513564 220934 513616 220940
rect 512734 218920 512790 218929
rect 512734 218855 512790 218864
rect 512748 217274 512776 218855
rect 513576 217274 513604 220934
rect 509378 217194 509430 217200
rect 509390 216988 509418 217194
rect 510218 216988 510246 217246
rect 510620 217252 510672 217258
rect 510620 217194 510672 217200
rect 511046 217246 511120 217274
rect 511862 217252 511914 217258
rect 511046 216988 511074 217246
rect 511862 217194 511914 217200
rect 512702 217246 512776 217274
rect 513530 217246 513604 217274
rect 514312 217274 514340 222022
rect 515140 217274 515168 223790
rect 515968 221134 515996 226578
rect 516782 225992 516838 226001
rect 516782 225927 516838 225936
rect 515956 221128 516008 221134
rect 515956 221070 516008 221076
rect 515968 217274 515996 221070
rect 516796 217274 516824 225927
rect 517612 223984 517664 223990
rect 517612 223926 517664 223932
rect 517624 217274 517652 223926
rect 517808 222086 517836 227938
rect 518900 226160 518952 226166
rect 518900 226102 518952 226108
rect 518912 222601 518940 226102
rect 518898 222592 518954 222601
rect 518898 222527 518954 222536
rect 517796 222080 517848 222086
rect 517796 222022 517848 222028
rect 518440 222080 518492 222086
rect 518440 222022 518492 222028
rect 518452 217274 518480 222022
rect 514312 217246 514386 217274
rect 515140 217246 515214 217274
rect 515968 217246 516042 217274
rect 516796 217246 516870 217274
rect 517624 217246 517698 217274
rect 518452 217246 518526 217274
rect 518912 217258 518940 222527
rect 520936 221882 520964 228074
rect 523500 226772 523552 226778
rect 523500 226714 523552 226720
rect 522580 224120 522632 224126
rect 522580 224062 522632 224068
rect 522592 221882 522620 224062
rect 523224 223168 523276 223174
rect 523224 223110 523276 223116
rect 523236 222358 523264 223110
rect 523040 222352 523092 222358
rect 523040 222294 523092 222300
rect 523224 222352 523276 222358
rect 523224 222294 523276 222300
rect 519268 221876 519320 221882
rect 519268 221818 519320 221824
rect 520924 221876 520976 221882
rect 520924 221818 520976 221824
rect 522580 221876 522632 221882
rect 522580 221818 522632 221824
rect 519280 217274 519308 221818
rect 520936 217274 520964 221818
rect 521752 221740 521804 221746
rect 521752 221682 521804 221688
rect 521764 217274 521792 221682
rect 522592 217274 522620 221818
rect 511874 216988 511902 217194
rect 512702 216988 512730 217246
rect 513530 216988 513558 217246
rect 514358 216988 514386 217246
rect 515186 216988 515214 217246
rect 516014 216988 516042 217246
rect 516842 216988 516870 217246
rect 517670 216988 517698 217246
rect 518498 216988 518526 217246
rect 518900 217252 518952 217258
rect 519280 217246 519354 217274
rect 518900 217194 518952 217200
rect 519326 216988 519354 217246
rect 520142 217252 520194 217258
rect 520936 217246 521010 217274
rect 521764 217246 521838 217274
rect 522592 217246 522666 217274
rect 523052 217258 523080 222294
rect 523512 219434 523540 226714
rect 525064 225344 525116 225350
rect 525064 225286 525116 225292
rect 523684 223168 523736 223174
rect 523684 223110 523736 223116
rect 523696 222222 523724 223110
rect 524880 222488 524932 222494
rect 524880 222430 524932 222436
rect 523684 222216 523736 222222
rect 523684 222158 523736 222164
rect 523868 222216 523920 222222
rect 523868 222158 523920 222164
rect 523880 221882 523908 222158
rect 523868 221876 523920 221882
rect 523868 221818 523920 221824
rect 524326 220280 524382 220289
rect 524326 220215 524382 220224
rect 523512 219406 523724 219434
rect 520142 217194 520194 217200
rect 520154 216988 520182 217194
rect 520982 216988 521010 217246
rect 521810 216988 521838 217246
rect 522638 216988 522666 217246
rect 523040 217252 523092 217258
rect 523040 217194 523092 217200
rect 523696 217122 523724 219406
rect 524340 219026 524368 220215
rect 524328 219020 524380 219026
rect 524328 218962 524380 218968
rect 524892 217258 524920 222430
rect 525076 220969 525104 225286
rect 525996 221241 526024 229026
rect 531688 228268 531740 228274
rect 531688 228210 531740 228216
rect 527824 227588 527876 227594
rect 527824 227530 527876 227536
rect 526720 222420 526772 222426
rect 526720 222362 526772 222368
rect 527640 222420 527692 222426
rect 527640 222362 527692 222368
rect 525982 221232 526038 221241
rect 525982 221167 526038 221176
rect 525062 220960 525118 220969
rect 525062 220895 525118 220904
rect 525076 217274 525104 220895
rect 525996 217274 526024 221167
rect 526444 219972 526496 219978
rect 526444 219914 526496 219920
rect 526456 219094 526484 219914
rect 526444 219088 526496 219094
rect 526444 219030 526496 219036
rect 524282 217252 524334 217258
rect 524282 217194 524334 217200
rect 524880 217252 524932 217258
rect 525076 217246 525150 217274
rect 524880 217194 524932 217200
rect 523454 217116 523506 217122
rect 523454 217058 523506 217064
rect 523684 217116 523736 217122
rect 523684 217058 523736 217064
rect 523466 216988 523494 217058
rect 524294 216988 524322 217194
rect 525122 216988 525150 217246
rect 525950 217246 526024 217274
rect 525950 216988 525978 217246
rect 526732 217138 526760 222362
rect 527652 217274 527680 222362
rect 527836 218006 527864 227530
rect 530584 226296 530636 226302
rect 530584 226238 530636 226244
rect 528468 225208 528520 225214
rect 528468 225150 528520 225156
rect 528480 223530 528508 225150
rect 528480 223514 529428 223530
rect 528480 223508 529440 223514
rect 528480 223502 529388 223508
rect 528480 222426 528508 223502
rect 529388 223450 529440 223456
rect 529204 223440 529256 223446
rect 529204 223382 529256 223388
rect 529216 223174 529244 223382
rect 529020 223168 529072 223174
rect 529020 223110 529072 223116
rect 529204 223168 529256 223174
rect 529204 223110 529256 223116
rect 529032 222630 529060 223110
rect 529020 222624 529072 222630
rect 529020 222566 529072 222572
rect 528468 222420 528520 222426
rect 528468 222362 528520 222368
rect 529388 222148 529440 222154
rect 529388 222090 529440 222096
rect 529400 221338 529428 222090
rect 529756 221740 529808 221746
rect 529756 221682 529808 221688
rect 529388 221332 529440 221338
rect 529388 221274 529440 221280
rect 529572 221332 529624 221338
rect 529572 221274 529624 221280
rect 529388 219632 529440 219638
rect 529388 219574 529440 219580
rect 529400 219094 529428 219574
rect 529388 219088 529440 219094
rect 529388 219030 529440 219036
rect 529584 218890 529612 221274
rect 529768 221241 529796 221682
rect 529754 221232 529810 221241
rect 529754 221167 529810 221176
rect 530596 219094 530624 226238
rect 530860 219768 530912 219774
rect 530860 219710 530912 219716
rect 530124 219088 530176 219094
rect 530124 219030 530176 219036
rect 530584 219088 530636 219094
rect 530584 219030 530636 219036
rect 529572 218884 529624 218890
rect 529572 218826 529624 218832
rect 527824 218000 527876 218006
rect 527824 217942 527876 217948
rect 528376 218000 528428 218006
rect 528376 217942 528428 217948
rect 528388 217734 528416 217942
rect 528376 217728 528428 217734
rect 528376 217670 528428 217676
rect 527606 217246 527680 217274
rect 526732 217110 526806 217138
rect 526778 216988 526806 217110
rect 527606 216988 527634 217246
rect 528388 217138 528416 217670
rect 529250 217252 529302 217258
rect 529250 217194 529302 217200
rect 528388 217110 528462 217138
rect 528434 216988 528462 217110
rect 529262 216988 529290 217194
rect 530136 217138 530164 219030
rect 530596 218890 530624 219030
rect 530584 218884 530636 218890
rect 530584 218826 530636 218832
rect 530872 217870 530900 219710
rect 530860 217864 530912 217870
rect 530860 217806 530912 217812
rect 530090 217110 530164 217138
rect 530872 217138 530900 217806
rect 531700 217274 531728 228210
rect 533356 226302 533384 229162
rect 535920 226908 535972 226914
rect 535920 226850 535972 226856
rect 533344 226296 533396 226302
rect 533344 226238 533396 226244
rect 531964 225480 532016 225486
rect 531964 225422 532016 225428
rect 531976 219094 532004 225422
rect 535000 225072 535052 225078
rect 535000 225014 535052 225020
rect 533528 222760 533580 222766
rect 533528 222702 533580 222708
rect 533804 222760 533856 222766
rect 534172 222760 534224 222766
rect 533856 222720 534172 222748
rect 533804 222702 533856 222708
rect 534172 222702 534224 222708
rect 533540 222578 533568 222702
rect 533540 222550 534212 222578
rect 533528 222488 533580 222494
rect 533528 222430 533580 222436
rect 533540 221241 533568 222430
rect 533988 222420 534040 222426
rect 533988 222362 534040 222368
rect 533526 221232 533582 221241
rect 533526 221167 533582 221176
rect 534000 220969 534028 222362
rect 533986 220960 534042 220969
rect 533986 220895 534042 220904
rect 533344 219904 533396 219910
rect 533344 219846 533396 219852
rect 531964 219088 532016 219094
rect 531964 219030 532016 219036
rect 532516 219088 532568 219094
rect 532516 219030 532568 219036
rect 532528 218210 532556 219030
rect 532516 218204 532568 218210
rect 532516 218146 532568 218152
rect 531700 217246 531774 217274
rect 530872 217110 530946 217138
rect 530090 216988 530118 217110
rect 530918 216988 530946 217110
rect 531746 216988 531774 217246
rect 532528 217138 532556 218146
rect 533356 217138 533384 219846
rect 534184 217274 534212 222550
rect 535012 218346 535040 225014
rect 535932 219094 535960 226850
rect 536852 226166 536880 229298
rect 538404 228812 538456 228818
rect 538404 228754 538456 228760
rect 536840 226160 536892 226166
rect 536840 226102 536892 226108
rect 536840 225888 536892 225894
rect 536840 225830 536892 225836
rect 536852 224058 536880 225830
rect 536840 224052 536892 224058
rect 536840 223994 536892 224000
rect 537484 224052 537536 224058
rect 537484 223994 537536 224000
rect 536104 223508 536156 223514
rect 536104 223450 536156 223456
rect 536116 222562 536144 223450
rect 536104 222556 536156 222562
rect 536104 222498 536156 222504
rect 536654 221232 536710 221241
rect 536654 221167 536710 221176
rect 535920 219088 535972 219094
rect 535920 219030 535972 219036
rect 535000 218340 535052 218346
rect 535000 218282 535052 218288
rect 535012 217274 535040 218282
rect 535932 217274 535960 219030
rect 534184 217246 534258 217274
rect 535012 217246 535086 217274
rect 532528 217110 532602 217138
rect 533356 217110 533430 217138
rect 532574 216988 532602 217110
rect 533402 216988 533430 217110
rect 534230 216988 534258 217246
rect 535058 216988 535086 217246
rect 535886 217246 535960 217274
rect 535886 216988 535914 217246
rect 536668 217138 536696 221167
rect 537496 217274 537524 223994
rect 538416 220833 538444 228754
rect 540244 226024 540296 226030
rect 540244 225966 540296 225972
rect 540256 224954 540284 225966
rect 540072 224926 540284 224954
rect 539232 223168 539284 223174
rect 539232 223110 539284 223116
rect 538402 220824 538458 220833
rect 538402 220759 538458 220768
rect 538416 217274 538444 220759
rect 539048 220516 539100 220522
rect 539048 220458 539100 220464
rect 538680 219904 538732 219910
rect 538680 219846 538732 219852
rect 538692 219638 538720 219846
rect 539060 219774 539088 220458
rect 539048 219768 539100 219774
rect 539048 219710 539100 219716
rect 538680 219632 538732 219638
rect 538680 219574 538732 219580
rect 537496 217246 537570 217274
rect 536668 217110 536742 217138
rect 536714 216988 536742 217110
rect 537542 216988 537570 217246
rect 538370 217246 538444 217274
rect 538370 216988 538398 217246
rect 539244 217138 539272 223110
rect 540072 218482 540100 224926
rect 542004 223310 542032 230114
rect 551928 229900 551980 229906
rect 551928 229842 551980 229848
rect 548340 228676 548392 228682
rect 548340 228618 548392 228624
rect 546592 227452 546644 227458
rect 546592 227394 546644 227400
rect 543464 227316 543516 227322
rect 543464 227258 543516 227264
rect 543476 224954 543504 227258
rect 543740 225752 543792 225758
rect 543740 225694 543792 225700
rect 542360 224936 542412 224942
rect 542360 224878 542412 224884
rect 543384 224926 543504 224954
rect 543752 224942 543780 225694
rect 543740 224936 543792 224942
rect 541624 223304 541676 223310
rect 541624 223246 541676 223252
rect 541992 223304 542044 223310
rect 541992 223246 542044 223252
rect 540796 220516 540848 220522
rect 540796 220458 540848 220464
rect 540808 219910 540836 220458
rect 540796 219904 540848 219910
rect 540796 219846 540848 219852
rect 540980 219904 541032 219910
rect 540980 219846 541032 219852
rect 540060 218476 540112 218482
rect 540060 218418 540112 218424
rect 540072 217274 540100 218418
rect 539198 217110 539272 217138
rect 540026 217246 540100 217274
rect 539198 216988 539226 217110
rect 540026 216988 540054 217246
rect 540808 217138 540836 219846
rect 540992 219094 541020 219846
rect 540980 219088 541032 219094
rect 540980 219030 541032 219036
rect 541636 217138 541664 223246
rect 542372 218618 542400 224878
rect 543384 220561 543412 224926
rect 543740 224878 543792 224884
rect 545028 224936 545080 224942
rect 545028 224878 545080 224884
rect 544384 224052 544436 224058
rect 544384 223994 544436 224000
rect 544396 223938 544424 223994
rect 544028 223922 544424 223938
rect 544016 223916 544424 223922
rect 544068 223910 544424 223916
rect 544016 223858 544068 223864
rect 544200 222896 544252 222902
rect 544200 222838 544252 222844
rect 544212 222194 544240 222838
rect 544212 222166 544608 222194
rect 543554 221096 543610 221105
rect 543554 221031 543610 221040
rect 543568 220658 543596 221031
rect 543556 220652 543608 220658
rect 544384 220652 544436 220658
rect 543556 220594 543608 220600
rect 543936 220612 544384 220640
rect 543370 220552 543426 220561
rect 543370 220487 543426 220496
rect 542360 218612 542412 218618
rect 542360 218554 542412 218560
rect 542372 217274 542400 218554
rect 543384 217274 543412 220487
rect 543936 220402 543964 220612
rect 544384 220594 544436 220600
rect 543844 220386 543964 220402
rect 543832 220380 543964 220386
rect 543884 220374 543964 220380
rect 543832 220322 543884 220328
rect 543832 219768 543884 219774
rect 543832 219710 543884 219716
rect 543844 218006 543872 219710
rect 543832 218000 543884 218006
rect 543832 217942 543884 217948
rect 542372 217246 542538 217274
rect 540808 217110 540882 217138
rect 541636 217110 541710 217138
rect 540854 216988 540882 217110
rect 541682 216988 541710 217110
rect 542510 216988 542538 217246
rect 543338 217246 543412 217274
rect 544580 217258 544608 222166
rect 544154 217252 544206 217258
rect 543338 216988 543366 217246
rect 544154 217194 544206 217200
rect 544568 217252 544620 217258
rect 544568 217194 544620 217200
rect 544166 216988 544194 217194
rect 545040 217138 545068 224878
rect 545210 220824 545266 220833
rect 545210 220759 545266 220768
rect 545224 219774 545252 220759
rect 545762 220552 545818 220561
rect 545762 220487 545818 220496
rect 545776 220386 545804 220487
rect 545764 220380 545816 220386
rect 545764 220322 545816 220328
rect 545212 219768 545264 219774
rect 545212 219710 545264 219716
rect 545856 218000 545908 218006
rect 545856 217942 545908 217948
rect 545868 217138 545896 217942
rect 546604 217274 546632 227394
rect 547512 227180 547564 227186
rect 547512 227122 547564 227128
rect 547524 219366 547552 227122
rect 548352 223174 548380 228618
rect 548524 228540 548576 228546
rect 548524 228482 548576 228488
rect 548340 223168 548392 223174
rect 548340 223110 548392 223116
rect 548536 222986 548564 228482
rect 549904 225616 549956 225622
rect 549904 225558 549956 225564
rect 549076 223168 549128 223174
rect 549076 223110 549128 223116
rect 548352 222958 548748 222986
rect 547512 219360 547564 219366
rect 547512 219302 547564 219308
rect 547524 217274 547552 219302
rect 548156 217864 548208 217870
rect 548156 217806 548208 217812
rect 548168 217598 548196 217806
rect 548156 217592 548208 217598
rect 548156 217534 548208 217540
rect 548352 217274 548380 222958
rect 548720 222873 548748 222958
rect 548706 222864 548762 222873
rect 548706 222799 548762 222808
rect 546604 217246 546678 217274
rect 544994 217110 545068 217138
rect 545822 217110 545896 217138
rect 544994 216988 545022 217110
rect 545822 216988 545850 217110
rect 546650 216988 546678 217246
rect 547478 217246 547552 217274
rect 548306 217246 548380 217274
rect 547478 216988 547506 217246
rect 548306 216988 548334 217246
rect 549088 217138 549116 223110
rect 549916 222426 549944 225558
rect 551940 223446 551968 229842
rect 558184 229764 558236 229770
rect 558184 229706 558236 229712
rect 552204 228948 552256 228954
rect 552204 228890 552256 228896
rect 551928 223440 551980 223446
rect 551928 223382 551980 223388
rect 550640 223168 550692 223174
rect 550640 223110 550692 223116
rect 549904 222420 549956 222426
rect 549904 222362 549956 222368
rect 549444 219360 549496 219366
rect 549444 219302 549496 219308
rect 549456 218074 549484 219302
rect 549444 218068 549496 218074
rect 549444 218010 549496 218016
rect 549916 217274 549944 222362
rect 550652 219094 550680 223110
rect 551560 223032 551612 223038
rect 551560 222974 551612 222980
rect 551744 223032 551796 223038
rect 551744 222974 551796 222980
rect 550822 221096 550878 221105
rect 550822 221031 550878 221040
rect 550640 219088 550692 219094
rect 550640 219030 550692 219036
rect 549916 217246 549990 217274
rect 549088 217110 549162 217138
rect 549134 216988 549162 217110
rect 549962 216988 549990 217246
rect 550836 217138 550864 221031
rect 551572 217274 551600 222974
rect 551756 219230 551784 222974
rect 551744 219224 551796 219230
rect 551744 219166 551796 219172
rect 552216 219026 552244 228890
rect 555700 227044 555752 227050
rect 555700 226986 555752 226992
rect 553400 225072 553452 225078
rect 553400 225014 553452 225020
rect 552756 224936 552808 224942
rect 552756 224878 552808 224884
rect 552768 224670 552796 224878
rect 552756 224664 552808 224670
rect 552756 224606 552808 224612
rect 552940 224664 552992 224670
rect 552940 224606 552992 224612
rect 552952 223922 552980 224606
rect 553412 223922 553440 225014
rect 555712 224954 555740 226986
rect 556712 226296 556764 226302
rect 556712 226238 556764 226244
rect 555620 224926 555740 224954
rect 552940 223916 552992 223922
rect 552940 223858 552992 223864
rect 553400 223916 553452 223922
rect 553400 223858 553452 223864
rect 555422 223408 555478 223417
rect 555422 223343 555478 223352
rect 554044 222896 554096 222902
rect 554044 222838 554096 222844
rect 554688 222896 554740 222902
rect 554688 222838 554740 222844
rect 553308 222148 553360 222154
rect 553308 222090 553360 222096
rect 553320 222034 553348 222090
rect 553320 222006 553532 222034
rect 553504 221241 553532 222006
rect 553490 221232 553546 221241
rect 553490 221167 553546 221176
rect 553306 221096 553362 221105
rect 553306 221031 553362 221040
rect 553320 220810 553348 221031
rect 553320 220782 553394 220810
rect 553366 220726 553394 220782
rect 553354 220720 553406 220726
rect 553122 220688 553178 220697
rect 553354 220662 553406 220668
rect 553122 220623 553124 220632
rect 553176 220623 553178 220632
rect 553504 220646 553900 220674
rect 553124 220594 553176 220600
rect 552940 220244 552992 220250
rect 552940 220186 552992 220192
rect 552204 219020 552256 219026
rect 552204 218962 552256 218968
rect 552388 219020 552440 219026
rect 552388 218962 552440 218968
rect 551572 217246 551646 217274
rect 550790 217110 550864 217138
rect 550790 216988 550818 217110
rect 551618 216988 551646 217246
rect 552400 217138 552428 218962
rect 552952 217258 552980 220186
rect 553136 217274 553164 220594
rect 553504 220561 553532 220646
rect 553490 220552 553546 220561
rect 553490 220487 553546 220496
rect 553674 220552 553730 220561
rect 553674 220487 553730 220496
rect 553688 220266 553716 220487
rect 553872 220386 553900 220646
rect 553860 220380 553912 220386
rect 553860 220322 553912 220328
rect 553412 220238 553716 220266
rect 553412 220114 553440 220238
rect 553400 220108 553452 220114
rect 553400 220050 553452 220056
rect 552940 217252 552992 217258
rect 553136 217246 553302 217274
rect 552940 217194 552992 217200
rect 552400 217110 552474 217138
rect 552446 216988 552474 217110
rect 553274 216988 553302 217246
rect 554056 217138 554084 222838
rect 554700 218754 554728 222838
rect 555436 222766 555464 223343
rect 555424 222760 555476 222766
rect 555424 222702 555476 222708
rect 554870 221232 554926 221241
rect 554870 221167 554926 221176
rect 554884 219162 554912 221167
rect 555620 220096 555648 224926
rect 556724 224806 556752 226238
rect 558196 224954 558224 229706
rect 558196 224926 558408 224954
rect 556528 224800 556580 224806
rect 556528 224742 556580 224748
rect 556712 224800 556764 224806
rect 556712 224742 556764 224748
rect 557356 224800 557408 224806
rect 557356 224742 557408 224748
rect 557816 224800 557868 224806
rect 557816 224742 557868 224748
rect 556342 222864 556398 222873
rect 556342 222799 556398 222808
rect 555976 222148 556028 222154
rect 555976 222090 556028 222096
rect 555988 221610 556016 222090
rect 555976 221604 556028 221610
rect 555976 221546 556028 221552
rect 556356 221474 556384 222799
rect 556344 221468 556396 221474
rect 556344 221410 556396 221416
rect 555620 220068 555740 220096
rect 554872 219156 554924 219162
rect 554872 219098 554924 219104
rect 554688 218748 554740 218754
rect 554688 218690 554740 218696
rect 554884 217138 554912 219098
rect 555712 217462 555740 220068
rect 555700 217456 555752 217462
rect 555700 217398 555752 217404
rect 555712 217274 555740 217398
rect 556540 217274 556568 224742
rect 557368 224505 557396 224742
rect 557828 224534 557856 224742
rect 557816 224528 557868 224534
rect 557354 224496 557410 224505
rect 557816 224470 557868 224476
rect 558000 224528 558052 224534
rect 558000 224470 558052 224476
rect 557354 224431 557410 224440
rect 557368 217274 557396 224431
rect 558012 224262 558040 224470
rect 558000 224256 558052 224262
rect 558000 224198 558052 224204
rect 558000 223304 558052 223310
rect 558000 223246 558052 223252
rect 558012 222873 558040 223246
rect 557998 222864 558054 222873
rect 557998 222799 558054 222808
rect 558380 220726 558408 224926
rect 559012 224936 559064 224942
rect 559012 224878 559064 224884
rect 558550 224496 558606 224505
rect 558550 224431 558606 224440
rect 558564 224058 558592 224431
rect 558552 224052 558604 224058
rect 558552 223994 558604 224000
rect 558550 223408 558606 223417
rect 558550 223343 558606 223352
rect 558564 223038 558592 223343
rect 558552 223032 558604 223038
rect 558552 222974 558604 222980
rect 558368 220720 558420 220726
rect 558368 220662 558420 220668
rect 558000 220516 558052 220522
rect 558000 220458 558052 220464
rect 558012 220250 558040 220458
rect 557816 220244 557868 220250
rect 557816 220186 557868 220192
rect 558000 220244 558052 220250
rect 558000 220186 558052 220192
rect 557828 219910 557856 220186
rect 557816 219904 557868 219910
rect 557816 219846 557868 219852
rect 558184 219020 558236 219026
rect 558184 218962 558236 218968
rect 558196 218754 558224 218962
rect 558184 218748 558236 218754
rect 558184 218690 558236 218696
rect 555712 217246 555786 217274
rect 556540 217246 556614 217274
rect 557368 217246 557442 217274
rect 554056 217110 554130 217138
rect 554884 217110 554958 217138
rect 554102 216988 554130 217110
rect 554930 216988 554958 217110
rect 555758 216988 555786 217246
rect 556586 216988 556614 217246
rect 557414 216988 557442 217246
rect 558230 217252 558282 217258
rect 558230 217194 558282 217200
rect 558242 216988 558270 217194
rect 559024 217138 559052 224878
rect 559576 222902 559604 252554
rect 567212 229094 567240 256702
rect 567212 229066 568160 229094
rect 561772 226160 561824 226166
rect 561772 226102 561824 226108
rect 561496 224800 561548 224806
rect 561496 224742 561548 224748
rect 559564 222896 559616 222902
rect 559564 222838 559616 222844
rect 559838 222864 559894 222873
rect 559838 222799 559894 222808
rect 559852 219366 559880 222799
rect 560666 220552 560722 220561
rect 560666 220487 560722 220496
rect 559840 219360 559892 219366
rect 559840 219302 559892 219308
rect 559852 217138 559880 219302
rect 560680 217138 560708 220487
rect 561508 217138 561536 224742
rect 561784 219162 561812 226102
rect 568132 224954 568160 229066
rect 568132 224926 568528 224954
rect 566464 224528 566516 224534
rect 566464 224470 566516 224476
rect 563980 224392 564032 224398
rect 563980 224334 564032 224340
rect 563244 221604 563296 221610
rect 563244 221546 563296 221552
rect 562782 220960 562838 220969
rect 562782 220895 562838 220904
rect 562796 220726 562824 220895
rect 562784 220720 562836 220726
rect 562968 220720 563020 220726
rect 562784 220662 562836 220668
rect 562966 220688 562968 220697
rect 563020 220688 563022 220697
rect 562966 220623 563022 220632
rect 561772 219156 561824 219162
rect 561772 219098 561824 219104
rect 562324 219156 562376 219162
rect 562324 219098 562376 219104
rect 562336 217138 562364 219098
rect 563256 217138 563284 221546
rect 559024 217110 559098 217138
rect 559852 217110 559926 217138
rect 560680 217110 560754 217138
rect 561508 217110 561582 217138
rect 562336 217110 562410 217138
rect 559070 216988 559098 217110
rect 559898 216988 559926 217110
rect 560726 216988 560754 217110
rect 561554 216988 561582 217110
rect 562382 216988 562410 217110
rect 563210 217110 563284 217138
rect 563992 217138 564020 224334
rect 564808 223440 564860 223446
rect 564808 223382 564860 223388
rect 564622 220552 564678 220561
rect 564622 220487 564678 220496
rect 564636 220250 564664 220487
rect 564624 220244 564676 220250
rect 564624 220186 564676 220192
rect 564820 217841 564848 223382
rect 565728 222148 565780 222154
rect 565728 222090 565780 222096
rect 565358 220552 565414 220561
rect 565358 220487 565414 220496
rect 565372 220046 565400 220487
rect 565360 220040 565412 220046
rect 565360 219982 565412 219988
rect 564806 217832 564862 217841
rect 564806 217767 564862 217776
rect 564820 217138 564848 217767
rect 565740 217138 565768 222090
rect 563992 217110 564066 217138
rect 564820 217110 564894 217138
rect 563210 216988 563238 217110
rect 564038 216988 564066 217110
rect 564866 216988 564894 217110
rect 565694 217110 565768 217138
rect 566476 217138 566504 224470
rect 567752 223032 567804 223038
rect 567804 222980 568160 222986
rect 567752 222974 568160 222980
rect 567764 222958 568160 222974
rect 568132 222902 568160 222958
rect 568120 222896 568172 222902
rect 568120 222838 568172 222844
rect 567672 222278 568068 222306
rect 567672 222154 567700 222278
rect 567660 222148 567712 222154
rect 567660 222090 567712 222096
rect 567844 222148 567896 222154
rect 567844 222090 567896 222096
rect 567856 221474 567884 222090
rect 568040 221762 568068 222278
rect 568040 221734 568344 221762
rect 568316 221610 568344 221734
rect 568304 221604 568356 221610
rect 568304 221546 568356 221552
rect 567844 221468 567896 221474
rect 567844 221410 567896 221416
rect 567290 220824 567346 220833
rect 567290 220759 567346 220768
rect 567304 217841 567332 220759
rect 568028 219360 568080 219366
rect 568028 219302 568080 219308
rect 568212 219360 568264 219366
rect 568212 219302 568264 219308
rect 567474 219192 567530 219201
rect 567474 219127 567476 219136
rect 567528 219127 567530 219136
rect 567660 219156 567712 219162
rect 567476 219098 567528 219104
rect 567660 219098 567712 219104
rect 567672 218754 567700 219098
rect 568040 219026 568068 219302
rect 567844 219020 567896 219026
rect 567844 218962 567896 218968
rect 568028 219020 568080 219026
rect 568028 218962 568080 218968
rect 567856 218754 567884 218962
rect 567660 218748 567712 218754
rect 567660 218690 567712 218696
rect 567844 218748 567896 218754
rect 567844 218690 567896 218696
rect 568224 218090 568252 219302
rect 567672 218074 568252 218090
rect 567660 218068 568252 218074
rect 567712 218062 568252 218068
rect 567660 218010 567712 218016
rect 567844 218000 567896 218006
rect 567844 217942 567896 217948
rect 567290 217832 567346 217841
rect 567290 217767 567346 217776
rect 567304 217138 567332 217767
rect 567856 217258 567884 217942
rect 568500 217410 568528 224926
rect 568224 217382 568528 217410
rect 568224 217274 568252 217382
rect 567844 217252 567896 217258
rect 567844 217194 567896 217200
rect 568178 217246 568252 217274
rect 568592 217258 568620 261462
rect 571340 250504 571392 250510
rect 571340 250446 571392 250452
rect 570052 246356 570104 246362
rect 570052 246298 570104 246304
rect 568764 238196 568816 238202
rect 568764 238138 568816 238144
rect 568776 229094 568804 238138
rect 570064 229094 570092 246298
rect 568776 229066 568988 229094
rect 570064 229066 570644 229094
rect 568960 217274 568988 229066
rect 570144 218000 570196 218006
rect 570144 217942 570196 217948
rect 570156 217462 570184 217942
rect 570144 217456 570196 217462
rect 570144 217398 570196 217404
rect 570616 217274 570644 229066
rect 571352 224954 571380 250446
rect 632704 242208 632756 242214
rect 632704 242150 632756 242156
rect 629944 240780 629996 240786
rect 629944 240722 629996 240728
rect 577504 234048 577556 234054
rect 577504 233990 577556 233996
rect 571352 224926 572300 224954
rect 571432 223032 571484 223038
rect 571432 222974 571484 222980
rect 568580 217252 568632 217258
rect 566476 217110 566550 217138
rect 567304 217110 567378 217138
rect 565694 216988 565722 217110
rect 566522 216988 566550 217110
rect 567350 216988 567378 217110
rect 568178 216988 568206 217246
rect 568960 217246 569034 217274
rect 568580 217194 568632 217200
rect 569006 216988 569034 217246
rect 569822 217252 569874 217258
rect 570616 217246 570690 217274
rect 569822 217194 569874 217200
rect 569834 216988 569862 217194
rect 570662 216988 570690 217246
rect 571444 217138 571472 222974
rect 572272 217274 572300 224926
rect 572536 220720 572588 220726
rect 572536 220662 572588 220668
rect 572548 220561 572576 220662
rect 572674 220652 572726 220658
rect 572674 220594 572726 220600
rect 574560 220652 574612 220658
rect 574560 220594 574612 220600
rect 574744 220652 574796 220658
rect 574744 220594 574796 220600
rect 572534 220552 572590 220561
rect 572534 220487 572590 220496
rect 572686 220402 572714 220594
rect 572548 220374 572714 220402
rect 572548 219201 572576 220374
rect 572534 219192 572590 219201
rect 572534 219127 572590 219136
rect 574190 219192 574246 219201
rect 574190 219127 574246 219136
rect 574204 218074 574232 219127
rect 574192 218068 574244 218074
rect 574192 218010 574244 218016
rect 574282 217832 574338 217841
rect 574282 217767 574338 217776
rect 572272 217246 572346 217274
rect 571444 217110 571518 217138
rect 571490 216988 571518 217110
rect 572318 216988 572346 217246
rect 574296 216986 574324 217767
rect 574284 216980 574336 216986
rect 574284 216922 574336 216928
rect 574374 216472 574430 216481
rect 574374 216407 574430 216416
rect 574388 213246 574416 216407
rect 574572 215966 574600 220594
rect 574756 220046 574784 220594
rect 574926 220552 574982 220561
rect 574926 220487 574982 220496
rect 574940 220046 574968 220487
rect 574744 220040 574796 220046
rect 574744 219982 574796 219988
rect 574928 220040 574980 220046
rect 574928 219982 574980 219988
rect 574744 219292 574796 219298
rect 574744 219234 574796 219240
rect 574560 215960 574612 215966
rect 574560 215902 574612 215908
rect 574756 214606 574784 219234
rect 575110 219192 575166 219201
rect 574928 219156 574980 219162
rect 575110 219127 575166 219136
rect 574928 219098 574980 219104
rect 574940 216374 574968 219098
rect 574928 216368 574980 216374
rect 574928 216310 574980 216316
rect 574928 216096 574980 216102
rect 574926 216064 574928 216073
rect 574980 216064 574982 216073
rect 574926 215999 574982 216008
rect 575124 214742 575152 219127
rect 575296 219020 575348 219026
rect 575296 218962 575348 218968
rect 575308 216238 575336 218962
rect 575478 216744 575534 216753
rect 575478 216679 575534 216688
rect 575296 216232 575348 216238
rect 575296 216174 575348 216180
rect 575112 214736 575164 214742
rect 575112 214678 575164 214684
rect 574744 214600 574796 214606
rect 574744 214542 574796 214548
rect 575492 213382 575520 216679
rect 575480 213376 575532 213382
rect 575480 213318 575532 213324
rect 574376 213240 574428 213246
rect 574376 213182 574428 213188
rect 50988 212696 51040 212702
rect 50988 212638 51040 212644
rect 50344 203040 50396 203046
rect 50344 202982 50396 202988
rect 44548 191820 44600 191826
rect 44548 191762 44600 191768
rect 44364 191684 44416 191690
rect 44364 191626 44416 191632
rect 42432 183524 42484 183530
rect 42432 183466 42484 183472
rect 44180 183524 44232 183530
rect 44180 183466 44232 183472
rect 41786 183424 41842 183433
rect 41786 183359 41842 183368
rect 41800 183124 41828 183359
rect 42444 182491 42472 183466
rect 42182 182463 42472 182491
rect 577516 97986 577544 233990
rect 613290 225312 613346 225321
rect 613290 225247 613346 225256
rect 590936 224460 590988 224466
rect 590936 224402 590988 224408
rect 597560 224460 597612 224466
rect 597560 224402 597612 224408
rect 590948 223650 590976 224402
rect 591120 224188 591172 224194
rect 591120 224130 591172 224136
rect 591132 223650 591160 224130
rect 590936 223644 590988 223650
rect 590936 223586 590988 223592
rect 591120 223644 591172 223650
rect 591120 223586 591172 223592
rect 596824 222896 596876 222902
rect 596824 222838 596876 222844
rect 596836 222630 596864 222838
rect 596640 222624 596692 222630
rect 596640 222566 596692 222572
rect 596824 222624 596876 222630
rect 596824 222566 596876 222572
rect 596652 222442 596680 222566
rect 596652 222414 597048 222442
rect 597020 222358 597048 222414
rect 597008 222352 597060 222358
rect 597008 222294 597060 222300
rect 591304 222148 591356 222154
rect 591304 222090 591356 222096
rect 591488 222148 591540 222154
rect 591488 222090 591540 222096
rect 591316 220862 591344 222090
rect 591120 220856 591172 220862
rect 591120 220798 591172 220804
rect 591304 220856 591356 220862
rect 591304 220798 591356 220804
rect 591132 220674 591160 220798
rect 591500 220674 591528 222090
rect 591994 222012 592046 222018
rect 591994 221954 592046 221960
rect 592006 221898 592034 221954
rect 592006 221870 592080 221898
rect 592052 221241 592080 221870
rect 593972 221332 594024 221338
rect 593972 221274 594024 221280
rect 592038 221232 592094 221241
rect 592038 221167 592094 221176
rect 591132 220646 591528 220674
rect 578882 215384 578938 215393
rect 578882 215319 578938 215328
rect 578330 212936 578386 212945
rect 578330 212871 578386 212880
rect 578344 211342 578372 212871
rect 578332 211336 578384 211342
rect 578332 211278 578384 211284
rect 578896 208282 578924 215319
rect 580632 211336 580684 211342
rect 580632 211278 580684 211284
rect 579526 210352 579582 210361
rect 579526 210287 579582 210296
rect 579540 210118 579568 210287
rect 579528 210112 579580 210118
rect 579528 210054 579580 210060
rect 579526 208584 579582 208593
rect 579582 208542 579752 208570
rect 579526 208519 579582 208528
rect 578884 208276 578936 208282
rect 578884 208218 578936 208224
rect 579526 205864 579582 205873
rect 579526 205799 579528 205808
rect 579580 205799 579582 205808
rect 579528 205770 579580 205776
rect 579724 204270 579752 208542
rect 580644 206990 580672 211278
rect 593984 210202 594012 221274
rect 594156 221264 594208 221270
rect 594154 221232 594156 221241
rect 594208 221232 594210 221241
rect 594154 221167 594210 221176
rect 597008 220652 597060 220658
rect 597008 220594 597060 220600
rect 596270 220280 596326 220289
rect 596270 220215 596326 220224
rect 596640 220244 596692 220250
rect 596088 218884 596140 218890
rect 596088 218826 596140 218832
rect 595166 217560 595222 217569
rect 595166 217495 595222 217504
rect 594800 213376 594852 213382
rect 594800 213318 594852 213324
rect 594812 210202 594840 213318
rect 595180 210202 595208 217495
rect 595718 217288 595774 217297
rect 595718 217223 595774 217232
rect 595732 210202 595760 217223
rect 596100 216714 596128 218826
rect 596088 216708 596140 216714
rect 596088 216650 596140 216656
rect 596284 215294 596312 220215
rect 596640 220186 596692 220192
rect 596456 220176 596508 220182
rect 596456 220118 596508 220124
rect 596468 219502 596496 220118
rect 596652 219774 596680 220186
rect 597020 219910 597048 220594
rect 597008 219904 597060 219910
rect 597008 219846 597060 219852
rect 596640 219768 596692 219774
rect 596640 219710 596692 219716
rect 596456 219496 596508 219502
rect 596456 219438 596508 219444
rect 597192 218204 597244 218210
rect 597192 218146 597244 218152
rect 596652 217790 597048 217818
rect 596652 217734 596680 217790
rect 596640 217728 596692 217734
rect 596640 217670 596692 217676
rect 596824 217728 596876 217734
rect 596824 217670 596876 217676
rect 596836 217462 596864 217670
rect 597020 217462 597048 217790
rect 596824 217456 596876 217462
rect 596824 217398 596876 217404
rect 597008 217456 597060 217462
rect 597008 217398 597060 217404
rect 597008 217184 597060 217190
rect 597008 217126 597060 217132
rect 596822 217016 596878 217025
rect 596822 216951 596878 216960
rect 596284 215266 596588 215294
rect 596560 210202 596588 215266
rect 596836 210202 596864 216951
rect 597020 216918 597048 217126
rect 597008 216912 597060 216918
rect 597008 216854 597060 216860
rect 597204 216850 597232 218146
rect 597192 216844 597244 216850
rect 597192 216786 597244 216792
rect 593984 210174 594412 210202
rect 594812 210174 594964 210202
rect 595180 210174 595516 210202
rect 595732 210174 596068 210202
rect 596560 210174 596620 210202
rect 596836 210174 597172 210202
rect 597572 210118 597600 224402
rect 610440 224324 610492 224330
rect 610440 224266 610492 224272
rect 610452 223650 610480 224266
rect 611634 224224 611690 224233
rect 610808 224188 610860 224194
rect 611634 224159 611690 224168
rect 610808 224130 610860 224136
rect 610820 223786 610848 224130
rect 610808 223780 610860 223786
rect 610808 223722 610860 223728
rect 610440 223644 610492 223650
rect 610440 223586 610492 223592
rect 597836 222080 597888 222086
rect 597836 222022 597888 222028
rect 597848 214470 597876 222022
rect 600320 221876 600372 221882
rect 600320 221818 600372 221824
rect 598940 220992 598992 220998
rect 598940 220934 598992 220940
rect 598018 220008 598074 220017
rect 598018 219943 598074 219952
rect 597836 214464 597888 214470
rect 597836 214406 597888 214412
rect 598032 210202 598060 219943
rect 598952 214470 598980 220934
rect 599124 219360 599176 219366
rect 599124 219302 599176 219308
rect 598480 214464 598532 214470
rect 598480 214406 598532 214412
rect 598940 214464 598992 214470
rect 598940 214406 598992 214412
rect 597724 210174 598060 210202
rect 598492 210202 598520 214406
rect 599136 210202 599164 219302
rect 600332 214470 600360 221818
rect 602252 221740 602304 221746
rect 602252 221682 602304 221688
rect 601056 221264 601108 221270
rect 601056 221206 601108 221212
rect 600872 221128 600924 221134
rect 600872 221070 600924 221076
rect 599584 214464 599636 214470
rect 599584 214406 599636 214412
rect 600320 214464 600372 214470
rect 600320 214406 600372 214412
rect 599596 210202 599624 214406
rect 600884 210338 600912 221070
rect 601068 215294 601096 221206
rect 601700 218476 601752 218482
rect 601700 218418 601752 218424
rect 601712 217598 601740 218418
rect 601976 217864 602028 217870
rect 601976 217806 602028 217812
rect 601516 217592 601568 217598
rect 601514 217560 601516 217569
rect 601700 217592 601752 217598
rect 601568 217560 601570 217569
rect 601700 217534 601752 217540
rect 601514 217495 601570 217504
rect 601332 217456 601384 217462
rect 601654 217456 601706 217462
rect 601332 217398 601384 217404
rect 601620 217404 601654 217410
rect 601620 217398 601706 217404
rect 601344 217297 601372 217398
rect 601620 217382 601694 217398
rect 601330 217288 601386 217297
rect 601330 217223 601386 217232
rect 601620 216714 601648 217382
rect 601792 217048 601844 217054
rect 601792 216990 601844 216996
rect 601608 216708 601660 216714
rect 601608 216650 601660 216656
rect 600700 210310 600912 210338
rect 600976 215266 601096 215294
rect 600700 210202 600728 210310
rect 598492 210174 598828 210202
rect 599136 210174 599380 210202
rect 599596 210174 599932 210202
rect 600484 210174 600728 210202
rect 600976 210202 601004 215266
rect 601240 214464 601292 214470
rect 601240 214406 601292 214412
rect 601252 210202 601280 214406
rect 601804 210202 601832 216990
rect 601988 216714 602016 217806
rect 601976 216708 602028 216714
rect 601976 216650 602028 216656
rect 602264 210202 602292 221682
rect 611360 221604 611412 221610
rect 611360 221546 611412 221552
rect 609980 221468 610032 221474
rect 609980 221410 610032 221416
rect 607220 220856 607272 220862
rect 607220 220798 607272 220804
rect 605012 220244 605064 220250
rect 605012 220186 605064 220192
rect 603908 219632 603960 219638
rect 603908 219574 603960 219580
rect 603446 217560 603502 217569
rect 603446 217495 603502 217504
rect 603078 217288 603134 217297
rect 603078 217223 603134 217232
rect 603092 210202 603120 217223
rect 603460 210202 603488 217495
rect 603920 210202 603948 219574
rect 604552 219496 604604 219502
rect 604552 219438 604604 219444
rect 604564 210202 604592 219438
rect 605024 210202 605052 220186
rect 605932 219904 605984 219910
rect 605932 219846 605984 219852
rect 605944 210202 605972 219846
rect 606116 219768 606168 219774
rect 606116 219710 606168 219716
rect 606128 210202 606156 219710
rect 606760 216708 606812 216714
rect 606760 216650 606812 216656
rect 606772 210202 606800 216650
rect 607232 210202 607260 220798
rect 607772 220516 607824 220522
rect 607772 220458 607824 220464
rect 607784 210202 607812 220458
rect 608876 220380 608928 220386
rect 608876 220322 608928 220328
rect 608508 218340 608560 218346
rect 608508 218282 608560 218288
rect 608520 217734 608548 218282
rect 608324 217728 608376 217734
rect 608324 217670 608376 217676
rect 608508 217728 608560 217734
rect 608508 217670 608560 217676
rect 608336 213790 608364 217670
rect 608324 213784 608376 213790
rect 608324 213726 608376 213732
rect 608888 210202 608916 220322
rect 609610 218376 609666 218385
rect 609610 218311 609666 218320
rect 609060 217320 609112 217326
rect 609060 217262 609112 217268
rect 600976 210174 601036 210202
rect 601252 210174 601588 210202
rect 601804 210174 602140 210202
rect 602264 210174 602692 210202
rect 603092 210174 603244 210202
rect 603460 210174 603796 210202
rect 603920 210174 604348 210202
rect 604564 210174 604900 210202
rect 605024 210174 605452 210202
rect 605944 210174 606004 210202
rect 606128 210174 606556 210202
rect 606772 210174 607108 210202
rect 607232 210174 607660 210202
rect 607784 210174 608212 210202
rect 608764 210174 608916 210202
rect 609072 210202 609100 217262
rect 609624 216850 609652 218311
rect 609612 216844 609664 216850
rect 609612 216786 609664 216792
rect 609992 214606 610020 221410
rect 610164 220040 610216 220046
rect 610164 219982 610216 219988
rect 609980 214600 610032 214606
rect 609980 214542 610032 214548
rect 609520 213784 609572 213790
rect 609520 213726 609572 213732
rect 609532 210202 609560 213726
rect 610176 210202 610204 219982
rect 610624 214600 610676 214606
rect 610624 214542 610676 214548
rect 610636 210202 610664 214542
rect 611372 210202 611400 221546
rect 611648 210202 611676 224159
rect 612830 216744 612886 216753
rect 612830 216679 612886 216688
rect 612280 214736 612332 214742
rect 612280 214678 612332 214684
rect 612292 210202 612320 214678
rect 612844 210202 612872 216679
rect 613304 210202 613332 225247
rect 617708 224188 617760 224194
rect 617708 224130 617760 224136
rect 617064 223644 617116 223650
rect 617064 223586 617116 223592
rect 614394 223136 614450 223145
rect 614394 223071 614450 223080
rect 614120 218068 614172 218074
rect 614120 218010 614172 218016
rect 614132 210202 614160 218010
rect 614408 210202 614436 223071
rect 616878 218920 616934 218929
rect 616878 218855 616934 218864
rect 616142 218648 616198 218657
rect 616142 218583 616198 218592
rect 615038 218104 615094 218113
rect 615038 218039 615094 218048
rect 615052 210202 615080 218039
rect 615684 216844 615736 216850
rect 615684 216786 615736 216792
rect 615696 210202 615724 216786
rect 616156 210202 616184 218583
rect 616892 210202 616920 218855
rect 617076 210338 617104 223586
rect 617076 210310 617196 210338
rect 617168 210202 617196 210310
rect 617720 210202 617748 224130
rect 626724 224052 626776 224058
rect 626724 223994 626776 224000
rect 623780 223916 623832 223922
rect 623780 223858 623832 223864
rect 622584 223780 622636 223786
rect 622584 223722 622636 223728
rect 620468 223032 620520 223038
rect 620468 222974 620520 222980
rect 619180 222896 619232 222902
rect 619180 222838 619232 222844
rect 620284 222896 620336 222902
rect 620284 222838 620336 222844
rect 619192 222630 619220 222838
rect 618720 222624 618772 222630
rect 618534 222592 618590 222601
rect 618720 222566 618772 222572
rect 619180 222624 619232 222630
rect 619180 222566 619232 222572
rect 618534 222527 618590 222536
rect 618352 222216 618404 222222
rect 618352 222158 618404 222164
rect 618364 214606 618392 222158
rect 618352 214600 618404 214606
rect 618352 214542 618404 214548
rect 618548 210202 618576 222527
rect 618732 222222 618760 222566
rect 620296 222494 620324 222838
rect 620480 222494 620508 222974
rect 620284 222488 620336 222494
rect 620284 222430 620336 222436
rect 620468 222488 620520 222494
rect 620468 222430 620520 222436
rect 619732 222352 619784 222358
rect 619732 222294 619784 222300
rect 618720 222216 618772 222222
rect 618720 222158 618772 222164
rect 618904 214600 618956 214606
rect 618904 214542 618956 214548
rect 618916 210202 618944 214542
rect 619744 210202 619772 222294
rect 619916 222216 619968 222222
rect 619916 222158 619968 222164
rect 619928 210202 619956 222158
rect 621664 217728 621716 217734
rect 621664 217670 621716 217676
rect 620560 217456 620612 217462
rect 620560 217398 620612 217404
rect 620572 210202 620600 217398
rect 621112 216980 621164 216986
rect 621112 216922 621164 216928
rect 621124 210202 621152 216922
rect 621676 210202 621704 217670
rect 622596 210202 622624 223722
rect 623320 218612 623372 218618
rect 623320 218554 623372 218560
rect 622768 217592 622820 217598
rect 622768 217534 622820 217540
rect 609072 210174 609316 210202
rect 609532 210174 609868 210202
rect 610176 210174 610420 210202
rect 610636 210174 610972 210202
rect 611372 210174 611524 210202
rect 611648 210174 612076 210202
rect 612292 210174 612628 210202
rect 612844 210174 613180 210202
rect 613304 210174 613732 210202
rect 614132 210174 614284 210202
rect 614408 210174 614836 210202
rect 615052 210174 615388 210202
rect 615696 210174 615940 210202
rect 616156 210174 616492 210202
rect 616892 210174 617044 210202
rect 617168 210174 617596 210202
rect 617720 210174 618148 210202
rect 618548 210174 618700 210202
rect 618916 210174 619252 210202
rect 619744 210174 619804 210202
rect 619928 210174 620356 210202
rect 620572 210174 620908 210202
rect 621124 210174 621460 210202
rect 621676 210174 622012 210202
rect 622564 210174 622624 210202
rect 622780 210202 622808 217534
rect 623332 210202 623360 218554
rect 623792 210202 623820 223858
rect 625344 222896 625396 222902
rect 625344 222838 625396 222844
rect 625068 218748 625120 218754
rect 625068 218690 625120 218696
rect 625080 215234 625108 218690
rect 625080 215206 625200 215234
rect 624424 214464 624476 214470
rect 624424 214406 624476 214412
rect 624436 210202 624464 214406
rect 625172 213994 625200 215206
rect 625160 213988 625212 213994
rect 625160 213930 625212 213936
rect 625356 210202 625384 222838
rect 625528 216368 625580 216374
rect 625528 216310 625580 216316
rect 622780 210174 623116 210202
rect 623332 210174 623668 210202
rect 623792 210174 624220 210202
rect 624436 210174 624772 210202
rect 625324 210174 625384 210202
rect 625540 210202 625568 216310
rect 626080 213988 626132 213994
rect 626080 213930 626132 213936
rect 626092 210202 626120 213930
rect 626736 210202 626764 223994
rect 629300 222624 629352 222630
rect 629300 222566 629352 222572
rect 628840 217320 628892 217326
rect 628840 217262 628892 217268
rect 627184 216232 627236 216238
rect 627184 216174 627236 216180
rect 627196 210202 627224 216174
rect 628288 216096 628340 216102
rect 628288 216038 628340 216044
rect 627920 215960 627972 215966
rect 627920 215902 627972 215908
rect 627932 210202 627960 215902
rect 628300 210202 628328 216038
rect 628852 210202 628880 217262
rect 629312 210202 629340 222566
rect 629956 213450 629984 240722
rect 631324 233912 631376 233918
rect 631324 233854 631376 233860
rect 631336 229094 631364 233854
rect 631336 229066 631456 229094
rect 630680 227792 630732 227798
rect 630680 227734 630732 227740
rect 629944 213444 629996 213450
rect 629944 213386 629996 213392
rect 629944 213240 629996 213246
rect 629944 213182 629996 213188
rect 629956 210202 629984 213182
rect 630692 210202 630720 227734
rect 630956 222760 631008 222766
rect 630956 222702 631008 222708
rect 630968 210202 630996 222702
rect 631232 222488 631284 222494
rect 631232 222430 631284 222436
rect 631244 210338 631272 222430
rect 631428 212770 631456 229066
rect 632716 213926 632744 242150
rect 633440 238060 633492 238066
rect 633440 238002 633492 238008
rect 633452 229094 633480 238002
rect 641904 231804 641956 231810
rect 641904 231746 641956 231752
rect 641720 231668 641772 231674
rect 641720 231610 641772 231616
rect 633452 229066 634308 229094
rect 632704 213920 632756 213926
rect 632704 213862 632756 213868
rect 633440 213920 633492 213926
rect 633440 213862 633492 213868
rect 631416 212764 631468 212770
rect 631416 212706 631468 212712
rect 632704 212764 632756 212770
rect 632704 212706 632756 212712
rect 631244 210310 631548 210338
rect 631520 210202 631548 210310
rect 632716 210202 632744 212706
rect 633452 210202 633480 213862
rect 633808 213444 633860 213450
rect 633808 213386 633860 213392
rect 633820 210202 633848 213386
rect 634280 210202 634308 229066
rect 637212 213920 637264 213926
rect 637212 213862 637264 213868
rect 636660 213376 636712 213382
rect 636660 213318 636712 213324
rect 635556 213240 635608 213246
rect 635556 213182 635608 213188
rect 635568 210202 635596 213182
rect 636672 210202 636700 213318
rect 637224 210202 637252 213862
rect 638868 213784 638920 213790
rect 638868 213726 638920 213732
rect 638316 213512 638368 213518
rect 638316 213454 638368 213460
rect 638328 210202 638356 213454
rect 638880 210202 638908 213726
rect 639972 213648 640024 213654
rect 639972 213590 640024 213596
rect 639984 210202 640012 213590
rect 641536 213104 641588 213110
rect 641536 213046 641588 213052
rect 640248 212968 640300 212974
rect 640248 212910 640300 212916
rect 640260 210202 640288 212910
rect 641548 210202 641576 213046
rect 625540 210174 625876 210202
rect 626092 210174 626428 210202
rect 626736 210174 626980 210202
rect 627196 210174 627532 210202
rect 627932 210174 628084 210202
rect 628300 210174 628636 210202
rect 628852 210174 629188 210202
rect 629312 210174 629740 210202
rect 629956 210174 630292 210202
rect 630692 210174 630844 210202
rect 630968 210174 631396 210202
rect 631520 210174 631948 210202
rect 632716 210174 633052 210202
rect 633452 210174 633604 210202
rect 633820 210174 634156 210202
rect 634280 210174 634708 210202
rect 635260 210174 635596 210202
rect 636364 210174 636700 210202
rect 636916 210174 637252 210202
rect 638020 210174 638356 210202
rect 638572 210174 638908 210202
rect 639676 210174 640012 210202
rect 640228 210174 640288 210202
rect 641332 210174 641576 210202
rect 641732 210202 641760 231610
rect 641916 229094 641944 231746
rect 643100 231532 643152 231538
rect 643100 231474 643152 231480
rect 641916 229066 642588 229094
rect 642560 210202 642588 229066
rect 643112 210202 643140 231474
rect 644480 231124 644532 231130
rect 644480 231066 644532 231072
rect 644492 229094 644520 231066
rect 644492 229066 644612 229094
rect 644584 212534 644612 229066
rect 644492 212506 644612 212534
rect 644492 211070 644520 212506
rect 644480 211064 644532 211070
rect 644480 211006 644532 211012
rect 644676 210746 644704 278015
rect 645136 274718 645164 277780
rect 645872 277766 646346 277794
rect 647252 277766 647542 277794
rect 645124 274712 645176 274718
rect 645124 274654 645176 274660
rect 645872 268666 645900 277766
rect 647252 269822 647280 277766
rect 648724 277394 648752 277780
rect 648632 277366 648752 277394
rect 647240 269816 647292 269822
rect 647240 269758 647292 269764
rect 645860 268660 645912 268666
rect 645860 268602 645912 268608
rect 648632 265674 648660 277366
rect 648620 265668 648672 265674
rect 648620 265610 648672 265616
rect 645860 231396 645912 231402
rect 645860 231338 645912 231344
rect 644848 211064 644900 211070
rect 644848 211006 644900 211012
rect 644584 210718 644704 210746
rect 644584 210202 644612 210718
rect 644860 210202 644888 211006
rect 645872 210202 645900 231338
rect 648618 229800 648674 229809
rect 648618 229735 648674 229744
rect 648632 229094 648660 229735
rect 648632 229066 649212 229094
rect 647238 228576 647294 228585
rect 647238 228511 647294 228520
rect 646410 226672 646466 226681
rect 646410 226607 646466 226616
rect 646424 210202 646452 226607
rect 647252 212430 647280 228511
rect 647514 227488 647570 227497
rect 647514 227423 647570 227432
rect 647240 212424 647292 212430
rect 647240 212366 647292 212372
rect 647528 210202 647556 227423
rect 648160 212424 648212 212430
rect 648160 212366 648212 212372
rect 648172 210202 648200 212366
rect 649184 210202 649212 229066
rect 650104 213246 650132 990082
rect 650736 988780 650788 988786
rect 650736 988722 650788 988728
rect 650368 231260 650420 231266
rect 650368 231202 650420 231208
rect 650092 213240 650144 213246
rect 650092 213182 650144 213188
rect 650380 210202 650408 231202
rect 650550 228304 650606 228313
rect 650550 228239 650606 228248
rect 650564 219434 650592 228239
rect 650564 219406 650684 219434
rect 650656 210338 650684 219406
rect 650748 213466 650776 988722
rect 650932 213926 650960 991578
rect 651472 991500 651524 991506
rect 651472 991442 651524 991448
rect 651104 987420 651156 987426
rect 651104 987362 651156 987368
rect 650920 213920 650972 213926
rect 650920 213862 650972 213868
rect 650748 213438 650868 213466
rect 650840 213382 650868 213438
rect 650828 213376 650880 213382
rect 650828 213318 650880 213324
rect 651116 212974 651144 987362
rect 651484 213518 651512 991442
rect 651840 984632 651892 984638
rect 651840 984574 651892 984580
rect 651654 975896 651710 975905
rect 651654 975831 651710 975840
rect 651668 975730 651696 975831
rect 651656 975724 651708 975730
rect 651656 975666 651708 975672
rect 651654 962568 651710 962577
rect 651654 962503 651710 962512
rect 651668 961926 651696 962503
rect 651656 961920 651708 961926
rect 651656 961862 651708 961868
rect 651654 949376 651710 949385
rect 651654 949311 651710 949320
rect 651668 948122 651696 949311
rect 651656 948116 651708 948122
rect 651656 948058 651708 948064
rect 651656 937032 651708 937038
rect 651656 936974 651708 936980
rect 651668 936193 651696 936974
rect 651654 936184 651710 936193
rect 651654 936119 651710 936128
rect 651654 922720 651710 922729
rect 651654 922655 651710 922664
rect 651668 921874 651696 922655
rect 651656 921868 651708 921874
rect 651656 921810 651708 921816
rect 651654 909528 651710 909537
rect 651654 909463 651656 909472
rect 651708 909463 651710 909472
rect 651656 909434 651708 909440
rect 651654 896200 651710 896209
rect 651654 896135 651710 896144
rect 651668 895694 651696 896135
rect 651656 895688 651708 895694
rect 651656 895630 651708 895636
rect 651654 882872 651710 882881
rect 651654 882807 651710 882816
rect 651668 881890 651696 882807
rect 651656 881884 651708 881890
rect 651656 881826 651708 881832
rect 651654 869680 651710 869689
rect 651654 869615 651710 869624
rect 651668 869446 651696 869615
rect 651656 869440 651708 869446
rect 651656 869382 651708 869388
rect 651654 856352 651710 856361
rect 651654 856287 651710 856296
rect 651668 855642 651696 856287
rect 651656 855636 651708 855642
rect 651656 855578 651708 855584
rect 651654 843024 651710 843033
rect 651654 842959 651710 842968
rect 651668 841838 651696 842959
rect 651656 841832 651708 841838
rect 651656 841774 651708 841780
rect 651654 829832 651710 829841
rect 651654 829767 651710 829776
rect 651668 829462 651696 829767
rect 651656 829456 651708 829462
rect 651656 829398 651708 829404
rect 651654 816504 651710 816513
rect 651654 816439 651710 816448
rect 651668 815658 651696 816439
rect 651656 815652 651708 815658
rect 651656 815594 651708 815600
rect 651654 803312 651710 803321
rect 651654 803247 651656 803256
rect 651708 803247 651710 803256
rect 651656 803218 651708 803224
rect 651654 789984 651710 789993
rect 651654 789919 651710 789928
rect 651668 789410 651696 789919
rect 651656 789404 651708 789410
rect 651656 789346 651708 789352
rect 651654 776656 651710 776665
rect 651654 776591 651710 776600
rect 651668 775606 651696 776591
rect 651656 775600 651708 775606
rect 651656 775542 651708 775548
rect 651654 763328 651710 763337
rect 651654 763263 651656 763272
rect 651708 763263 651710 763272
rect 651656 763234 651708 763240
rect 651654 736808 651710 736817
rect 651654 736743 651710 736752
rect 651668 735622 651696 736743
rect 651656 735616 651708 735622
rect 651656 735558 651708 735564
rect 651654 723480 651710 723489
rect 651654 723415 651710 723424
rect 651668 723178 651696 723415
rect 651656 723172 651708 723178
rect 651656 723114 651708 723120
rect 651654 710288 651710 710297
rect 651654 710223 651710 710232
rect 651668 709374 651696 710223
rect 651656 709368 651708 709374
rect 651656 709310 651708 709316
rect 651656 696992 651708 696998
rect 651654 696960 651656 696969
rect 651708 696960 651710 696969
rect 651654 696895 651710 696904
rect 651654 683632 651710 683641
rect 651654 683567 651710 683576
rect 651668 683194 651696 683567
rect 651656 683188 651708 683194
rect 651656 683130 651708 683136
rect 651654 670440 651710 670449
rect 651654 670375 651710 670384
rect 651668 669390 651696 670375
rect 651656 669384 651708 669390
rect 651656 669326 651708 669332
rect 651654 657112 651710 657121
rect 651654 657047 651710 657056
rect 651668 656946 651696 657047
rect 651656 656940 651708 656946
rect 651656 656882 651708 656888
rect 651654 643784 651710 643793
rect 651654 643719 651710 643728
rect 651668 643142 651696 643719
rect 651656 643136 651708 643142
rect 651656 643078 651708 643084
rect 651654 617264 651710 617273
rect 651654 617199 651710 617208
rect 651668 616894 651696 617199
rect 651656 616888 651708 616894
rect 651656 616830 651708 616836
rect 651654 590744 651710 590753
rect 651654 590679 651656 590688
rect 651708 590679 651710 590688
rect 651656 590650 651708 590656
rect 651654 577416 651710 577425
rect 651654 577351 651710 577360
rect 651668 576910 651696 577351
rect 651656 576904 651708 576910
rect 651656 576846 651708 576852
rect 651654 564088 651710 564097
rect 651654 564023 651710 564032
rect 651668 563106 651696 564023
rect 651656 563100 651708 563106
rect 651656 563042 651708 563048
rect 651654 550896 651710 550905
rect 651654 550831 651710 550840
rect 651668 550662 651696 550831
rect 651656 550656 651708 550662
rect 651656 550598 651708 550604
rect 651654 524240 651710 524249
rect 651654 524175 651710 524184
rect 651668 523054 651696 524175
rect 651656 523048 651708 523054
rect 651656 522990 651708 522996
rect 651654 511048 651710 511057
rect 651654 510983 651710 510992
rect 651668 510678 651696 510983
rect 651656 510672 651708 510678
rect 651656 510614 651708 510620
rect 651654 497720 651710 497729
rect 651654 497655 651710 497664
rect 651668 496874 651696 497655
rect 651656 496868 651708 496874
rect 651656 496810 651708 496816
rect 651654 484528 651710 484537
rect 651654 484463 651656 484472
rect 651708 484463 651710 484472
rect 651656 484434 651708 484440
rect 651654 471200 651710 471209
rect 651654 471135 651710 471144
rect 651668 470626 651696 471135
rect 651656 470620 651708 470626
rect 651656 470562 651708 470568
rect 651654 457872 651710 457881
rect 651654 457807 651710 457816
rect 651668 456822 651696 457807
rect 651656 456816 651708 456822
rect 651656 456758 651708 456764
rect 651654 444544 651710 444553
rect 651654 444479 651656 444488
rect 651708 444479 651710 444488
rect 651656 444450 651708 444456
rect 651654 418024 651710 418033
rect 651654 417959 651710 417968
rect 651668 416838 651696 417959
rect 651656 416832 651708 416838
rect 651656 416774 651708 416780
rect 651654 404696 651710 404705
rect 651654 404631 651710 404640
rect 651668 404394 651696 404631
rect 651656 404388 651708 404394
rect 651656 404330 651708 404336
rect 651654 391504 651710 391513
rect 651654 391439 651710 391448
rect 651668 390590 651696 391439
rect 651656 390584 651708 390590
rect 651656 390526 651708 390532
rect 651656 378208 651708 378214
rect 651654 378176 651656 378185
rect 651708 378176 651710 378185
rect 651654 378111 651710 378120
rect 651654 364848 651710 364857
rect 651654 364783 651710 364792
rect 651668 364410 651696 364783
rect 651656 364404 651708 364410
rect 651656 364346 651708 364352
rect 651654 351656 651710 351665
rect 651654 351591 651710 351600
rect 651668 350606 651696 351591
rect 651656 350600 651708 350606
rect 651656 350542 651708 350548
rect 651654 338328 651710 338337
rect 651654 338263 651710 338272
rect 651668 338162 651696 338263
rect 651656 338156 651708 338162
rect 651656 338098 651708 338104
rect 651654 325000 651710 325009
rect 651654 324935 651710 324944
rect 651668 324358 651696 324935
rect 651656 324352 651708 324358
rect 651656 324294 651708 324300
rect 651654 285288 651710 285297
rect 651654 285223 651710 285232
rect 651668 284374 651696 285223
rect 651656 284368 651708 284374
rect 651656 284310 651708 284316
rect 651654 226944 651710 226953
rect 651654 226879 651710 226888
rect 651472 213512 651524 213518
rect 651472 213454 651524 213460
rect 651104 212968 651156 212974
rect 651104 212910 651156 212916
rect 650656 210310 650868 210338
rect 641732 210174 641884 210202
rect 642560 210174 642988 210202
rect 643112 210174 643540 210202
rect 644584 210174 644644 210202
rect 644860 210174 645196 210202
rect 645872 210174 646300 210202
rect 646424 210174 646852 210202
rect 647528 210174 647956 210202
rect 648172 210174 648508 210202
rect 649184 210174 649612 210202
rect 650164 210174 650408 210202
rect 650840 210202 650868 210310
rect 651668 210202 651696 226879
rect 651852 213110 651880 984574
rect 652022 750136 652078 750145
rect 652022 750071 652078 750080
rect 652036 749426 652064 750071
rect 652024 749420 652076 749426
rect 652024 749362 652076 749368
rect 652022 630592 652078 630601
rect 652022 630527 652078 630536
rect 652036 629338 652064 630527
rect 652024 629332 652076 629338
rect 652024 629274 652076 629280
rect 652022 603936 652078 603945
rect 652022 603871 652078 603880
rect 652036 603158 652064 603871
rect 652024 603152 652076 603158
rect 652024 603094 652076 603100
rect 652022 537568 652078 537577
rect 652022 537503 652078 537512
rect 652036 536858 652064 537503
rect 652024 536852 652076 536858
rect 652024 536794 652076 536800
rect 652022 431352 652078 431361
rect 652022 431287 652078 431296
rect 652036 430642 652064 431287
rect 652024 430636 652076 430642
rect 652024 430578 652076 430584
rect 652022 311808 652078 311817
rect 652022 311743 652078 311752
rect 651840 213104 651892 213110
rect 651840 213046 651892 213052
rect 652036 210458 652064 311743
rect 652206 298480 652262 298489
rect 652206 298415 652262 298424
rect 652220 210594 652248 298415
rect 652496 213790 652524 992870
rect 652484 213784 652536 213790
rect 652484 213726 652536 213732
rect 652772 213654 652800 993006
rect 658924 987692 658976 987698
rect 658924 987634 658976 987640
rect 658936 937242 658964 987634
rect 664444 984904 664496 984910
rect 664444 984846 664496 984852
rect 661684 975724 661736 975730
rect 661684 975666 661736 975672
rect 660304 957772 660356 957778
rect 660304 957714 660356 957720
rect 658924 937236 658976 937242
rect 658924 937178 658976 937184
rect 660316 937038 660344 957714
rect 661696 938466 661724 975666
rect 663064 961920 663116 961926
rect 663064 961862 663116 961868
rect 663076 941866 663104 961862
rect 663064 941860 663116 941866
rect 663064 941802 663116 941808
rect 661684 938460 661736 938466
rect 661684 938402 661736 938408
rect 660304 937032 660356 937038
rect 660304 936974 660356 936980
rect 663064 921868 663116 921874
rect 663064 921810 663116 921816
rect 658924 869440 658976 869446
rect 658924 869382 658976 869388
rect 658936 714882 658964 869382
rect 659108 855636 659160 855642
rect 659108 855578 659160 855584
rect 659120 716310 659148 855578
rect 661868 841832 661920 841838
rect 661868 841774 661920 841780
rect 660304 829456 660356 829462
rect 660304 829398 660356 829404
rect 660316 779006 660344 829398
rect 661684 815652 661736 815658
rect 661684 815594 661736 815600
rect 660488 789404 660540 789410
rect 660488 789346 660540 789352
rect 660304 779000 660356 779006
rect 660304 778942 660356 778948
rect 660304 763224 660356 763230
rect 660304 763166 660356 763172
rect 659292 749420 659344 749426
rect 659292 749362 659344 749368
rect 659108 716304 659160 716310
rect 659108 716246 659160 716252
rect 658924 714876 658976 714882
rect 658924 714818 658976 714824
rect 658924 683188 658976 683194
rect 658924 683130 658976 683136
rect 658936 579698 658964 683130
rect 659108 629332 659160 629338
rect 659108 629274 659160 629280
rect 658924 579692 658976 579698
rect 658924 579634 658976 579640
rect 658924 563100 658976 563106
rect 658924 563042 658976 563048
rect 658936 554062 658964 563042
rect 658924 554056 658976 554062
rect 658924 553998 658976 554004
rect 659120 534274 659148 629274
rect 659304 625462 659332 749362
rect 659476 723172 659528 723178
rect 659476 723114 659528 723120
rect 659488 689314 659516 723114
rect 659476 689308 659528 689314
rect 659476 689250 659528 689256
rect 659292 625456 659344 625462
rect 659292 625398 659344 625404
rect 660316 625190 660344 763166
rect 660500 669526 660528 789346
rect 661696 670750 661724 815594
rect 661880 715154 661908 841774
rect 663076 760442 663104 921810
rect 663248 803276 663300 803282
rect 663248 803218 663300 803224
rect 663064 760436 663116 760442
rect 663064 760378 663116 760384
rect 661868 715148 661920 715154
rect 661868 715090 661920 715096
rect 663064 709368 663116 709374
rect 663064 709310 663116 709316
rect 661868 696992 661920 696998
rect 661868 696934 661920 696940
rect 661684 670744 661736 670750
rect 661684 670686 661736 670692
rect 660488 669520 660540 669526
rect 660488 669462 660540 669468
rect 661684 656940 661736 656946
rect 661684 656882 661736 656888
rect 660304 625184 660356 625190
rect 660304 625126 660356 625132
rect 660488 616888 660540 616894
rect 660488 616830 660540 616836
rect 660304 603152 660356 603158
rect 660304 603094 660356 603100
rect 659292 550656 659344 550662
rect 659292 550598 659344 550604
rect 659108 534268 659160 534274
rect 659108 534210 659160 534216
rect 659108 510672 659160 510678
rect 659108 510614 659160 510620
rect 658924 430636 658976 430642
rect 658924 430578 658976 430584
rect 654140 278180 654192 278186
rect 654140 278122 654192 278128
rect 653034 276992 653090 277001
rect 653034 276927 653090 276936
rect 652760 213648 652812 213654
rect 652760 213590 652812 213596
rect 652208 210588 652260 210594
rect 652208 210530 652260 210536
rect 652024 210452 652076 210458
rect 652024 210394 652076 210400
rect 653048 210202 653076 276927
rect 653220 228404 653272 228410
rect 653220 228346 653272 228352
rect 650840 210174 651268 210202
rect 651668 210174 651820 210202
rect 652924 210174 653076 210202
rect 653232 210202 653260 228346
rect 654152 210202 654180 278122
rect 658280 278044 658332 278050
rect 658280 277986 658332 277992
rect 656898 276720 656954 276729
rect 656898 276655 656954 276664
rect 655520 264240 655572 264246
rect 655520 264182 655572 264188
rect 654322 230072 654378 230081
rect 654322 230007 654378 230016
rect 654336 229094 654364 230007
rect 655532 229094 655560 264182
rect 656912 229094 656940 276655
rect 654336 229066 654732 229094
rect 655532 229066 655652 229094
rect 656912 229066 657492 229094
rect 654704 210202 654732 229066
rect 655624 210338 655652 229066
rect 656346 227216 656402 227225
rect 656346 227151 656402 227160
rect 655624 210310 655836 210338
rect 655808 210202 655836 210310
rect 656360 210202 656388 227151
rect 657464 210202 657492 229066
rect 658292 210202 658320 277986
rect 658936 268054 658964 430578
rect 659120 357474 659148 510614
rect 659304 403306 659332 550598
rect 660316 491366 660344 603094
rect 660500 599622 660528 616830
rect 660488 599616 660540 599622
rect 660488 599558 660540 599564
rect 660488 536852 660540 536858
rect 660488 536794 660540 536800
rect 660304 491360 660356 491366
rect 660304 491302 660356 491308
rect 660304 416832 660356 416838
rect 660304 416774 660356 416780
rect 659292 403300 659344 403306
rect 659292 403242 659344 403248
rect 659108 357468 659160 357474
rect 659108 357410 659160 357416
rect 659660 278316 659712 278322
rect 659660 278258 659712 278264
rect 658924 268048 658976 268054
rect 658924 267990 658976 267996
rect 658462 265568 658518 265577
rect 658462 265503 658518 265512
rect 658476 229094 658504 265503
rect 658476 229066 659148 229094
rect 659120 210202 659148 229066
rect 659672 212430 659700 278258
rect 659844 276684 659896 276690
rect 659844 276626 659896 276632
rect 659660 212424 659712 212430
rect 659660 212366 659712 212372
rect 659856 210202 659884 276626
rect 660316 267918 660344 416774
rect 660500 403170 660528 536794
rect 661696 535498 661724 656882
rect 661880 581058 661908 696934
rect 662052 669384 662104 669390
rect 662052 669326 662104 669332
rect 662064 643754 662092 669326
rect 662052 643748 662104 643754
rect 662052 643690 662104 643696
rect 661868 581052 661920 581058
rect 661868 580994 661920 581000
rect 663076 579834 663104 709310
rect 663260 670886 663288 803218
rect 663432 775600 663484 775606
rect 663432 775542 663484 775548
rect 663444 734874 663472 775542
rect 663432 734868 663484 734874
rect 663432 734810 663484 734816
rect 663248 670880 663300 670886
rect 663248 670822 663300 670828
rect 663708 614168 663760 614174
rect 663708 614110 663760 614116
rect 663248 590708 663300 590714
rect 663248 590650 663300 590656
rect 663064 579828 663116 579834
rect 663064 579770 663116 579776
rect 661684 535492 661736 535498
rect 661684 535434 661736 535440
rect 661684 523048 661736 523054
rect 661684 522990 661736 522996
rect 660672 444440 660724 444446
rect 660672 444382 660724 444388
rect 660488 403164 660540 403170
rect 660488 403106 660540 403112
rect 660684 312050 660712 444382
rect 661696 403034 661724 522990
rect 661868 496868 661920 496874
rect 661868 496810 661920 496816
rect 661684 403028 661736 403034
rect 661684 402970 661736 402976
rect 661684 378208 661736 378214
rect 661684 378150 661736 378156
rect 660672 312044 660724 312050
rect 660672 311986 660724 311992
rect 661040 278452 661092 278458
rect 661040 278394 661092 278400
rect 660304 267912 660356 267918
rect 660304 267854 660356 267860
rect 660304 212424 660356 212430
rect 660304 212366 660356 212372
rect 660316 210202 660344 212366
rect 661052 210202 661080 278394
rect 661316 230988 661368 230994
rect 661316 230930 661368 230936
rect 661328 212430 661356 230930
rect 661696 222630 661724 378150
rect 661880 357610 661908 496810
rect 663260 491502 663288 590650
rect 663248 491496 663300 491502
rect 663248 491438 663300 491444
rect 663248 470620 663300 470626
rect 663248 470562 663300 470568
rect 663064 390584 663116 390590
rect 663064 390526 663116 390532
rect 661868 357604 661920 357610
rect 661868 357546 661920 357552
rect 661868 350600 661920 350606
rect 661868 350542 661920 350548
rect 661684 222624 661736 222630
rect 661684 222566 661736 222572
rect 661498 222048 661554 222057
rect 661498 221983 661554 221992
rect 661316 212424 661368 212430
rect 661316 212366 661368 212372
rect 661512 210202 661540 221983
rect 661880 215294 661908 350542
rect 662052 284368 662104 284374
rect 662052 284310 662104 284316
rect 661788 215266 661908 215294
rect 662064 215294 662092 284310
rect 662418 223952 662474 223961
rect 662418 223887 662474 223896
rect 662064 215266 662184 215294
rect 661788 210730 661816 215266
rect 661960 212424 662012 212430
rect 661960 212366 662012 212372
rect 661776 210724 661828 210730
rect 661776 210666 661828 210672
rect 661972 210202 662000 212366
rect 662156 210322 662184 215266
rect 662432 212430 662460 223887
rect 663076 222222 663104 390526
rect 663260 313478 663288 470562
rect 663432 456816 663484 456822
rect 663432 456758 663484 456764
rect 663248 313472 663300 313478
rect 663248 313414 663300 313420
rect 663444 313342 663472 456758
rect 663432 313336 663484 313342
rect 663432 313278 663484 313284
rect 663720 244934 663748 614110
rect 664260 550656 664312 550662
rect 664260 550598 664312 550604
rect 664272 484566 664300 550598
rect 664260 484560 664312 484566
rect 664260 484502 664312 484508
rect 664260 309392 664312 309398
rect 664260 309334 664312 309340
rect 664272 265130 664300 309334
rect 664260 265124 664312 265130
rect 664260 265066 664312 265072
rect 664260 264988 664312 264994
rect 664260 264930 664312 264936
rect 663708 244928 663760 244934
rect 663708 244870 663760 244876
rect 663064 222216 663116 222222
rect 663064 222158 663116 222164
rect 662602 221776 662658 221785
rect 662602 221711 662658 221720
rect 662420 212424 662472 212430
rect 662420 212366 662472 212372
rect 662144 210316 662196 210322
rect 662144 210258 662196 210264
rect 662616 210202 662644 221711
rect 663798 221504 663854 221513
rect 663798 221439 663854 221448
rect 663812 219434 663840 221439
rect 664272 221270 664300 264930
rect 664260 221264 664312 221270
rect 664260 221206 664312 221212
rect 663982 219736 664038 219745
rect 663982 219671 664038 219680
rect 663812 219406 663932 219434
rect 663904 212534 663932 219406
rect 663812 212506 663932 212534
rect 663064 212424 663116 212430
rect 663064 212366 663116 212372
rect 663076 210202 663104 212366
rect 663812 211070 663840 212506
rect 663800 211064 663852 211070
rect 663800 211006 663852 211012
rect 663996 210712 664024 219671
rect 664168 211064 664220 211070
rect 664168 211006 664220 211012
rect 663996 210684 664116 210712
rect 664088 210202 664116 210684
rect 653232 210174 653476 210202
rect 654152 210174 654580 210202
rect 654704 210174 655132 210202
rect 655808 210174 656236 210202
rect 656360 210174 656788 210202
rect 657464 210174 657892 210202
rect 658292 210174 658444 210202
rect 659120 210174 659548 210202
rect 659856 210174 660100 210202
rect 660316 210174 660652 210202
rect 661052 210174 661204 210202
rect 661512 210174 661756 210202
rect 661972 210174 662308 210202
rect 662616 210174 662860 210202
rect 663076 210174 663412 210202
rect 663964 210174 664116 210202
rect 664180 210202 664208 211006
rect 664456 210905 664484 984846
rect 665824 984768 665876 984774
rect 665824 984710 665876 984716
rect 664628 895688 664680 895694
rect 664628 895630 664680 895636
rect 664640 760578 664668 895630
rect 664628 760572 664680 760578
rect 664628 760514 664680 760520
rect 664628 735616 664680 735622
rect 664628 735558 664680 735564
rect 664640 625326 664668 735558
rect 665456 654288 665508 654294
rect 665456 654230 665508 654236
rect 665272 647760 665324 647766
rect 665272 647702 665324 647708
rect 664812 643136 664864 643142
rect 664812 643078 664864 643084
rect 664628 625320 664680 625326
rect 664628 625262 664680 625268
rect 664628 576904 664680 576910
rect 664628 576846 664680 576852
rect 664640 491638 664668 576846
rect 664824 535702 664852 643078
rect 665284 574122 665312 647702
rect 665468 574258 665496 654230
rect 665640 603152 665692 603158
rect 665640 603094 665692 603100
rect 665456 574252 665508 574258
rect 665456 574194 665508 574200
rect 665272 574116 665324 574122
rect 665272 574058 665324 574064
rect 665088 564460 665140 564466
rect 665088 564402 665140 564408
rect 664812 535696 664864 535702
rect 664812 535638 664864 535644
rect 664628 491632 664680 491638
rect 664628 491574 664680 491580
rect 665100 485858 665128 564402
rect 665652 529990 665680 603094
rect 665640 529984 665692 529990
rect 665640 529926 665692 529932
rect 665088 485852 665140 485858
rect 665088 485794 665140 485800
rect 664996 484424 665048 484430
rect 664996 484366 665048 484372
rect 664812 404388 664864 404394
rect 664812 404330 664864 404336
rect 664628 364404 664680 364410
rect 664628 364346 664680 364352
rect 664640 222902 664668 364346
rect 664824 267782 664852 404330
rect 665008 357746 665036 484366
rect 664996 357740 665048 357746
rect 664996 357682 665048 357688
rect 665088 309188 665140 309194
rect 665088 309130 665140 309136
rect 664812 267776 664864 267782
rect 664812 267718 664864 267724
rect 664812 266416 664864 266422
rect 664812 266358 664864 266364
rect 664628 222896 664680 222902
rect 664628 222838 664680 222844
rect 664824 222766 664852 266358
rect 665100 265266 665128 309130
rect 665272 265464 665324 265470
rect 665272 265406 665324 265412
rect 665088 265260 665140 265266
rect 665088 265202 665140 265208
rect 665284 265146 665312 265406
rect 665100 265118 665312 265146
rect 664812 222760 664864 222766
rect 664812 222702 664864 222708
rect 665100 219638 665128 265118
rect 665088 219632 665140 219638
rect 665088 219574 665140 219580
rect 665836 211177 665864 984710
rect 666100 742484 666152 742490
rect 666100 742426 666152 742432
rect 666112 665242 666140 742426
rect 666284 692844 666336 692850
rect 666284 692786 666336 692792
rect 666100 665236 666152 665242
rect 666100 665178 666152 665184
rect 666100 641776 666152 641782
rect 666100 641718 666152 641724
rect 666112 570178 666140 641718
rect 666296 619682 666324 692786
rect 666284 619676 666336 619682
rect 666284 619618 666336 619624
rect 666376 610020 666428 610026
rect 666376 609962 666428 609968
rect 666100 570172 666152 570178
rect 666100 570114 666152 570120
rect 666192 560380 666244 560386
rect 666192 560322 666244 560328
rect 666204 557682 666232 560322
rect 666204 557654 666324 557682
rect 666100 557592 666152 557598
rect 666100 557534 666152 557540
rect 666112 485994 666140 557534
rect 666100 485988 666152 485994
rect 666100 485930 666152 485936
rect 666296 483138 666324 557654
rect 666388 538214 666416 609962
rect 666572 538214 666600 994230
rect 666744 993336 666796 993342
rect 666744 993278 666796 993284
rect 666388 538186 666508 538214
rect 666572 538186 666692 538214
rect 666480 528630 666508 538186
rect 666468 528624 666520 528630
rect 666468 528566 666520 528572
rect 666664 509234 666692 538186
rect 666572 509206 666692 509234
rect 666284 483132 666336 483138
rect 666284 483074 666336 483080
rect 666376 313608 666428 313614
rect 666376 313550 666428 313556
rect 666388 313342 666416 313550
rect 666376 313336 666428 313342
rect 666376 313278 666428 313284
rect 666192 311908 666244 311914
rect 666192 311850 666244 311856
rect 666204 266830 666232 311850
rect 666376 310548 666428 310554
rect 666376 310490 666428 310496
rect 666192 266824 666244 266830
rect 666192 266766 666244 266772
rect 666388 266558 666416 310490
rect 666376 266552 666428 266558
rect 666376 266494 666428 266500
rect 666192 263628 666244 263634
rect 666192 263570 666244 263576
rect 666204 219774 666232 263570
rect 666376 262540 666428 262546
rect 666376 262482 666428 262488
rect 666388 241466 666416 262482
rect 666376 241460 666428 241466
rect 666376 241402 666428 241408
rect 666192 219768 666244 219774
rect 666192 219710 666244 219716
rect 665822 211168 665878 211177
rect 665822 211103 665878 211112
rect 664442 210896 664498 210905
rect 664442 210831 664498 210840
rect 664180 210174 664516 210202
rect 582288 210112 582340 210118
rect 582288 210054 582340 210060
rect 597560 210112 597612 210118
rect 597560 210054 597612 210060
rect 597928 210112 597980 210118
rect 597980 210060 598276 210066
rect 597928 210054 598276 210060
rect 580632 206984 580684 206990
rect 580632 206926 580684 206932
rect 581000 205828 581052 205834
rect 581000 205770 581052 205776
rect 579712 204264 579764 204270
rect 579712 204206 579764 204212
rect 578330 203280 578386 203289
rect 578330 203215 578386 203224
rect 578344 202910 578372 203215
rect 578332 202904 578384 202910
rect 578332 202846 578384 202852
rect 580264 202904 580316 202910
rect 580264 202846 580316 202852
rect 579158 200696 579214 200705
rect 579158 200631 579214 200640
rect 579172 200190 579200 200631
rect 579160 200184 579212 200190
rect 579160 200126 579212 200132
rect 580276 200054 580304 202846
rect 581012 202842 581040 205770
rect 582300 205562 582328 210054
rect 597940 210038 598276 210054
rect 591304 209840 591356 209846
rect 591304 209782 591356 209788
rect 632152 209840 632204 209846
rect 632204 209788 632500 209794
rect 632152 209782 632500 209788
rect 589462 208312 589518 208321
rect 589462 208247 589464 208256
rect 589516 208247 589518 208256
rect 589464 208218 589516 208224
rect 589556 206984 589608 206990
rect 589554 206952 589556 206961
rect 589608 206952 589610 206961
rect 589554 206887 589610 206896
rect 582288 205556 582340 205562
rect 582288 205498 582340 205504
rect 589464 205556 589516 205562
rect 589464 205498 589516 205504
rect 589476 205193 589504 205498
rect 589462 205184 589518 205193
rect 589462 205119 589518 205128
rect 589464 204264 589516 204270
rect 589464 204206 589516 204212
rect 589476 203697 589504 204206
rect 589462 203688 589518 203697
rect 589462 203623 589518 203632
rect 581000 202836 581052 202842
rect 581000 202778 581052 202784
rect 589464 202836 589516 202842
rect 589464 202778 589516 202784
rect 589476 202201 589504 202778
rect 589462 202192 589518 202201
rect 589462 202127 589518 202136
rect 590568 200184 590620 200190
rect 590568 200126 590620 200132
rect 580264 200048 580316 200054
rect 580264 199990 580316 199996
rect 589464 200048 589516 200054
rect 589464 199990 589516 199996
rect 589476 199889 589504 199990
rect 589462 199880 589518 199889
rect 589462 199815 589518 199824
rect 590580 198665 590608 200126
rect 590566 198656 590622 198665
rect 590566 198591 590622 198600
rect 578882 198112 578938 198121
rect 578882 198047 578938 198056
rect 578896 197402 578924 198047
rect 578884 197396 578936 197402
rect 578884 197338 578936 197344
rect 589464 197396 589516 197402
rect 589464 197338 589516 197344
rect 589476 197033 589504 197338
rect 589462 197024 589518 197033
rect 589462 196959 589518 196968
rect 579526 196072 579582 196081
rect 579526 196007 579528 196016
rect 579580 196007 579582 196016
rect 589556 196036 589608 196042
rect 579528 195978 579580 195984
rect 589556 195978 589608 195984
rect 589568 195537 589596 195978
rect 589554 195528 589610 195537
rect 589554 195463 589610 195472
rect 579526 193896 579582 193905
rect 579526 193831 579528 193840
rect 579580 193831 579582 193840
rect 589556 193860 589608 193866
rect 579528 193802 579580 193808
rect 589556 193802 589608 193808
rect 589568 193633 589596 193802
rect 589554 193624 589610 193633
rect 589554 193559 589610 193568
rect 589462 191720 589518 191729
rect 589462 191655 589518 191664
rect 579526 191176 579582 191185
rect 589476 191146 589504 191655
rect 579526 191111 579528 191120
rect 579580 191111 579582 191120
rect 589464 191140 589516 191146
rect 579528 191082 579580 191088
rect 589464 191082 589516 191088
rect 589462 190088 589518 190097
rect 589462 190023 589518 190032
rect 589476 189038 589504 190023
rect 579528 189032 579580 189038
rect 579526 189000 579528 189009
rect 589464 189032 589516 189038
rect 579580 189000 579582 189009
rect 589464 188974 589516 188980
rect 579526 188935 579582 188944
rect 589646 188456 589702 188465
rect 589646 188391 589702 188400
rect 579528 186992 579580 186998
rect 579528 186934 579580 186940
rect 589464 186992 589516 186998
rect 589464 186934 589516 186940
rect 579540 186697 579568 186934
rect 589476 186833 589504 186934
rect 589462 186824 589518 186833
rect 589462 186759 589518 186768
rect 579526 186688 579582 186697
rect 579526 186623 579582 186632
rect 589462 185192 589518 185201
rect 589462 185127 589518 185136
rect 589476 184958 589504 185127
rect 579436 184952 579488 184958
rect 579436 184894 579488 184900
rect 589464 184952 589516 184958
rect 589464 184894 589516 184900
rect 578516 184816 578568 184822
rect 578516 184758 578568 184764
rect 578528 184385 578556 184758
rect 578514 184376 578570 184385
rect 578514 184311 578570 184320
rect 579448 182073 579476 184894
rect 589660 184822 589688 188391
rect 589648 184816 589700 184822
rect 589648 184758 589700 184764
rect 589462 183560 589518 183569
rect 589462 183495 589518 183504
rect 589476 182238 589504 183495
rect 580908 182232 580960 182238
rect 580908 182174 580960 182180
rect 589464 182232 589516 182238
rect 589464 182174 589516 182180
rect 579434 182064 579490 182073
rect 579434 181999 579490 182008
rect 580920 179382 580948 182174
rect 589462 181928 589518 181937
rect 589462 181863 589518 181872
rect 589476 180878 589504 181863
rect 583116 180872 583168 180878
rect 583116 180814 583168 180820
rect 589464 180872 589516 180878
rect 589464 180814 589516 180820
rect 581736 179444 581788 179450
rect 581736 179386 581788 179392
rect 578332 179376 578384 179382
rect 578332 179318 578384 179324
rect 580908 179376 580960 179382
rect 580908 179318 580960 179324
rect 578344 179217 578372 179318
rect 578330 179208 578386 179217
rect 578330 179143 578386 179152
rect 579712 178084 579764 178090
rect 579712 178026 579764 178032
rect 579528 176656 579580 176662
rect 579528 176598 579580 176604
rect 579540 176497 579568 176598
rect 579526 176488 579582 176497
rect 579526 176423 579582 176432
rect 578700 174888 578752 174894
rect 578700 174830 578752 174836
rect 578712 174729 578740 174830
rect 578698 174720 578754 174729
rect 578698 174655 578754 174664
rect 579526 172136 579582 172145
rect 579724 172122 579752 178026
rect 581748 174894 581776 179386
rect 583128 176662 583156 180814
rect 589462 180296 589518 180305
rect 589462 180231 589518 180240
rect 589476 179450 589504 180231
rect 589464 179444 589516 179450
rect 589464 179386 589516 179392
rect 589462 178664 589518 178673
rect 589462 178599 589518 178608
rect 589476 178090 589504 178599
rect 589464 178084 589516 178090
rect 589464 178026 589516 178032
rect 589462 177032 589518 177041
rect 589462 176967 589518 176976
rect 583116 176656 583168 176662
rect 583116 176598 583168 176604
rect 589278 175400 589334 175409
rect 587164 175364 587216 175370
rect 589278 175335 589280 175344
rect 587164 175306 587216 175312
rect 589332 175335 589334 175344
rect 589280 175306 589332 175312
rect 581736 174888 581788 174894
rect 581736 174830 581788 174836
rect 581736 173188 581788 173194
rect 581736 173130 581788 173136
rect 579582 172094 579752 172122
rect 579526 172071 579582 172080
rect 579804 171148 579856 171154
rect 579804 171090 579856 171096
rect 578884 170400 578936 170406
rect 578884 170342 578936 170348
rect 578896 166977 578924 170342
rect 579252 169584 579304 169590
rect 579250 169552 579252 169561
rect 579304 169552 579306 169561
rect 579250 169487 579306 169496
rect 578882 166968 578938 166977
rect 578882 166903 578938 166912
rect 579816 166818 579844 171090
rect 581748 169590 581776 173130
rect 587176 170406 587204 175306
rect 589476 173194 589504 176967
rect 589738 173768 589794 173777
rect 589738 173703 589794 173712
rect 589464 173188 589516 173194
rect 589464 173130 589516 173136
rect 589462 172136 589518 172145
rect 589462 172071 589518 172080
rect 589476 171154 589504 172071
rect 589464 171148 589516 171154
rect 589464 171090 589516 171096
rect 588542 170504 588598 170513
rect 588542 170439 588598 170448
rect 587164 170400 587216 170406
rect 587164 170342 587216 170348
rect 581736 169584 581788 169590
rect 581736 169526 581788 169532
rect 583024 168428 583076 168434
rect 583024 168370 583076 168376
rect 581644 167068 581696 167074
rect 581644 167010 581696 167016
rect 579724 166790 579844 166818
rect 579528 166320 579580 166326
rect 579528 166262 579580 166268
rect 579540 164529 579568 166262
rect 579526 164520 579582 164529
rect 579526 164455 579582 164464
rect 579724 164234 579752 166790
rect 579540 164206 579752 164234
rect 580264 164280 580316 164286
rect 580264 164222 580316 164228
rect 579540 162489 579568 164206
rect 579526 162480 579582 162489
rect 579526 162415 579582 162424
rect 579528 159996 579580 160002
rect 579528 159938 579580 159944
rect 579540 159769 579568 159938
rect 579526 159760 579582 159769
rect 579526 159695 579582 159704
rect 579252 157344 579304 157350
rect 579252 157286 579304 157292
rect 579264 157185 579292 157286
rect 579250 157176 579306 157185
rect 579250 157111 579306 157120
rect 578700 155508 578752 155514
rect 578700 155450 578752 155456
rect 578712 155145 578740 155450
rect 578698 155136 578754 155145
rect 578698 155071 578754 155080
rect 580276 153474 580304 164222
rect 581656 155514 581684 167010
rect 583036 157350 583064 168370
rect 587348 162920 587400 162926
rect 587348 162862 587400 162868
rect 585968 160132 586020 160138
rect 585968 160074 586020 160080
rect 584404 157412 584456 157418
rect 584404 157354 584456 157360
rect 583024 157344 583076 157350
rect 583024 157286 583076 157292
rect 581644 155508 581696 155514
rect 581644 155450 581696 155456
rect 583208 154624 583260 154630
rect 583208 154566 583260 154572
rect 578332 153468 578384 153474
rect 578332 153410 578384 153416
rect 580264 153468 580316 153474
rect 580264 153410 580316 153416
rect 578344 152697 578372 153410
rect 581828 153264 581880 153270
rect 581828 153206 581880 153212
rect 578330 152688 578386 152697
rect 578330 152623 578386 152632
rect 578424 152516 578476 152522
rect 578424 152458 578476 152464
rect 578436 147665 578464 152458
rect 580632 151088 580684 151094
rect 580632 151030 580684 151036
rect 579528 150408 579580 150414
rect 579528 150350 579580 150356
rect 579540 150113 579568 150350
rect 579526 150104 579582 150113
rect 579526 150039 579582 150048
rect 578422 147656 578478 147665
rect 578422 147591 578478 147600
rect 578792 145444 578844 145450
rect 578792 145386 578844 145392
rect 578804 144673 578832 145386
rect 578790 144664 578846 144673
rect 578790 144599 578846 144608
rect 578884 144220 578936 144226
rect 578884 144162 578936 144168
rect 578332 137896 578384 137902
rect 578332 137838 578384 137844
rect 578344 137737 578372 137838
rect 578330 137728 578386 137737
rect 578330 137663 578386 137672
rect 578332 133816 578384 133822
rect 578332 133758 578384 133764
rect 578344 133113 578372 133758
rect 578330 133104 578386 133113
rect 578330 133039 578386 133048
rect 578896 125361 578924 144162
rect 579252 143472 579304 143478
rect 579252 143414 579304 143420
rect 579264 142905 579292 143414
rect 579250 142896 579306 142905
rect 579250 142831 579306 142840
rect 579528 140616 579580 140622
rect 579528 140558 579580 140564
rect 579540 140321 579568 140558
rect 579526 140312 579582 140321
rect 579526 140247 579582 140256
rect 580264 140072 580316 140078
rect 580264 140014 580316 140020
rect 579068 138712 579120 138718
rect 579068 138654 579120 138660
rect 579080 130665 579108 138654
rect 579344 135176 579396 135182
rect 579342 135144 579344 135153
rect 579396 135144 579398 135153
rect 579342 135079 579398 135088
rect 579252 133476 579304 133482
rect 579252 133418 579304 133424
rect 579066 130656 579122 130665
rect 579066 130591 579122 130600
rect 578882 125352 578938 125361
rect 578882 125287 578938 125296
rect 578424 124908 578476 124914
rect 578424 124850 578476 124856
rect 578436 120873 578464 124850
rect 578884 122664 578936 122670
rect 578882 122632 578884 122641
rect 578936 122632 578938 122641
rect 578882 122567 578938 122576
rect 578422 120864 578478 120873
rect 578422 120799 578478 120808
rect 578516 118312 578568 118318
rect 578514 118280 578516 118289
rect 578568 118280 578570 118289
rect 578514 118215 578570 118224
rect 579068 117360 579120 117366
rect 579068 117302 579120 117308
rect 578884 116000 578936 116006
rect 578884 115942 578936 115948
rect 578332 106820 578384 106826
rect 578332 106762 578384 106768
rect 578344 105913 578372 106762
rect 578330 105904 578386 105913
rect 578330 105839 578386 105848
rect 577504 97980 577556 97986
rect 577504 97922 577556 97928
rect 578608 96620 578660 96626
rect 578608 96562 578660 96568
rect 578620 96257 578648 96562
rect 578606 96248 578662 96257
rect 578606 96183 578662 96192
rect 578516 89616 578568 89622
rect 578516 89558 578568 89564
rect 578528 89049 578556 89558
rect 578514 89040 578570 89049
rect 578514 88975 578570 88984
rect 577504 77308 577556 77314
rect 577504 77250 577556 77256
rect 392564 53230 392624 53258
rect 78476 53094 78628 53122
rect 130824 53094 131068 53122
rect 78600 50289 78628 53094
rect 78586 50280 78642 50289
rect 78586 50215 78642 50224
rect 131040 49745 131068 53094
rect 145380 53100 145432 53106
rect 183172 53094 183508 53122
rect 235520 53094 235856 53122
rect 287868 53094 288204 53122
rect 340216 53094 340552 53122
rect 145380 53042 145432 53048
rect 145392 50810 145420 53042
rect 145084 50782 145420 50810
rect 183480 50386 183508 53094
rect 235828 51066 235856 53094
rect 288176 52358 288204 53094
rect 288164 52352 288216 52358
rect 288164 52294 288216 52300
rect 288176 51066 288204 52294
rect 340524 51066 340552 53094
rect 392596 52494 392624 53230
rect 444912 53094 445248 53122
rect 497260 53094 497596 53122
rect 391940 52488 391992 52494
rect 391940 52430 391992 52436
rect 392584 52488 392636 52494
rect 392584 52430 392636 52436
rect 391952 51066 391980 52430
rect 405096 51740 405148 51746
rect 405096 51682 405148 51688
rect 235816 51060 235868 51066
rect 235816 51002 235868 51008
rect 288164 51060 288216 51066
rect 288164 51002 288216 51008
rect 340512 51060 340564 51066
rect 340512 51002 340564 51008
rect 391940 51060 391992 51066
rect 391940 51002 391992 51008
rect 183468 50380 183520 50386
rect 183468 50322 183520 50328
rect 131026 49736 131082 49745
rect 131026 49671 131082 49680
rect 151910 47288 151966 47297
rect 151910 47223 151966 47232
rect 142172 46702 142370 46730
rect 142172 40338 142200 46702
rect 151924 45937 151952 47223
rect 151910 45928 151966 45937
rect 151910 45863 151966 45872
rect 194048 44872 194100 44878
rect 194048 44814 194100 44820
rect 187514 42120 187570 42129
rect 187358 42078 187514 42106
rect 194060 42092 194088 44814
rect 315948 43444 316000 43450
rect 315948 43386 316000 43392
rect 306976 42392 307032 42401
rect 306976 42327 307032 42336
rect 310104 42392 310160 42401
rect 310104 42327 310160 42336
rect 306990 42092 307018 42327
rect 310118 42092 310146 42327
rect 315960 42231 315988 43386
rect 315948 42225 316000 42231
rect 315948 42167 316000 42173
rect 361946 42120 362002 42129
rect 361790 42078 361946 42106
rect 187514 42055 187570 42064
rect 365166 42120 365222 42129
rect 364918 42078 365166 42106
rect 361946 42055 362002 42064
rect 405108 42106 405136 51682
rect 445220 50522 445248 53094
rect 497568 50561 497596 53094
rect 549272 53094 549608 53122
rect 549272 50561 549300 53094
rect 577516 52494 577544 77250
rect 578896 76809 578924 115942
rect 579080 79257 579108 117302
rect 579264 115705 579292 133418
rect 579528 128240 579580 128246
rect 579528 128182 579580 128188
rect 579540 127945 579568 128182
rect 579526 127936 579582 127945
rect 579526 127871 579582 127880
rect 580276 118318 580304 140014
rect 580448 133952 580500 133958
rect 580448 133894 580500 133900
rect 580264 118312 580316 118318
rect 580264 118254 580316 118260
rect 579250 115696 579306 115705
rect 579250 115631 579306 115640
rect 579528 113144 579580 113150
rect 579526 113112 579528 113121
rect 579580 113112 579582 113121
rect 579526 113047 579582 113056
rect 579528 111240 579580 111246
rect 579528 111182 579580 111188
rect 579540 111081 579568 111182
rect 579526 111072 579582 111081
rect 579526 111007 579582 111016
rect 579252 108792 579304 108798
rect 579252 108734 579304 108740
rect 579264 108497 579292 108734
rect 579250 108488 579306 108497
rect 579250 108423 579306 108432
rect 579252 107228 579304 107234
rect 579252 107170 579304 107176
rect 579264 100609 579292 107170
rect 580460 106826 580488 133894
rect 580644 133822 580672 151030
rect 581644 135312 581696 135318
rect 581644 135254 581696 135260
rect 580632 133816 580684 133822
rect 580632 133758 580684 133764
rect 580632 115252 580684 115258
rect 580632 115194 580684 115200
rect 580448 106820 580500 106826
rect 580448 106762 580500 106768
rect 580264 106344 580316 106350
rect 580264 106286 580316 106292
rect 579526 103456 579582 103465
rect 579526 103391 579528 103400
rect 579580 103391 579582 103400
rect 579528 103362 579580 103368
rect 579250 100600 579306 100609
rect 579250 100535 579306 100544
rect 579528 99340 579580 99346
rect 579528 99282 579580 99288
rect 579540 98841 579568 99282
rect 579526 98832 579582 98841
rect 579526 98767 579582 98776
rect 579528 93832 579580 93838
rect 579528 93774 579580 93780
rect 579540 93673 579568 93774
rect 579526 93664 579582 93673
rect 579526 93599 579582 93608
rect 579526 91080 579582 91089
rect 579526 91015 579528 91024
rect 579580 91015 579582 91024
rect 579528 90986 579580 90992
rect 579528 86964 579580 86970
rect 579528 86906 579580 86912
rect 579540 86465 579568 86906
rect 579526 86456 579582 86465
rect 579526 86391 579582 86400
rect 579344 84040 579396 84046
rect 579344 83982 579396 83988
rect 579356 83881 579384 83982
rect 579342 83872 579398 83881
rect 579342 83807 579398 83816
rect 579526 81424 579582 81433
rect 579526 81359 579528 81368
rect 579580 81359 579582 81368
rect 579528 81330 579580 81336
rect 579252 80096 579304 80102
rect 579252 80038 579304 80044
rect 579066 79248 579122 79257
rect 579066 79183 579122 79192
rect 578882 76800 578938 76809
rect 578882 76735 578938 76744
rect 578516 69012 578568 69018
rect 578516 68954 578568 68960
rect 578528 68785 578556 68954
rect 578514 68776 578570 68785
rect 578514 68711 578570 68720
rect 579264 64569 579292 80038
rect 579528 74520 579580 74526
rect 579528 74462 579580 74468
rect 579540 74225 579568 74462
rect 579526 74216 579582 74225
rect 579526 74151 579582 74160
rect 579528 71528 579580 71534
rect 579526 71496 579528 71505
rect 579580 71496 579582 71505
rect 579526 71431 579582 71440
rect 579528 67516 579580 67522
rect 579528 67458 579580 67464
rect 579540 67017 579568 67458
rect 579526 67008 579582 67017
rect 579526 66943 579582 66952
rect 579250 64560 579306 64569
rect 579250 64495 579306 64504
rect 580276 62014 580304 106286
rect 580644 89622 580672 115194
rect 581656 108798 581684 135254
rect 581840 135182 581868 153206
rect 583220 137902 583248 154566
rect 583760 140820 583812 140826
rect 583760 140762 583812 140768
rect 583208 137896 583260 137902
rect 583208 137838 583260 137844
rect 583024 137284 583076 137290
rect 583024 137226 583076 137232
rect 581828 135176 581880 135182
rect 581828 135118 581880 135124
rect 581828 121508 581880 121514
rect 581828 121450 581880 121456
rect 581644 108792 581696 108798
rect 581644 108734 581696 108740
rect 581644 103556 581696 103562
rect 581644 103498 581696 103504
rect 580632 89616 580684 89622
rect 580632 89558 580684 89564
rect 578516 62008 578568 62014
rect 578516 61950 578568 61956
rect 580264 62008 580316 62014
rect 580264 61950 580316 61956
rect 578528 61849 578556 61950
rect 578514 61840 578570 61849
rect 578514 61775 578570 61784
rect 579528 59016 579580 59022
rect 579526 58984 579528 58993
rect 579580 58984 579582 58993
rect 579526 58919 579582 58928
rect 581656 57934 581684 103498
rect 581840 84046 581868 121450
rect 583036 113150 583064 137226
rect 583772 133482 583800 140762
rect 584416 140622 584444 157354
rect 585980 145450 586008 160074
rect 587360 150414 587388 162862
rect 588556 160002 588584 170439
rect 589462 168872 589518 168881
rect 589462 168807 589518 168816
rect 589476 168434 589504 168807
rect 589464 168428 589516 168434
rect 589464 168370 589516 168376
rect 589462 167240 589518 167249
rect 589462 167175 589518 167184
rect 589476 167074 589504 167175
rect 589464 167068 589516 167074
rect 589464 167010 589516 167016
rect 589752 166326 589780 173703
rect 589740 166320 589792 166326
rect 589740 166262 589792 166268
rect 589462 165608 589518 165617
rect 589462 165543 589518 165552
rect 589476 164286 589504 165543
rect 589464 164280 589516 164286
rect 589464 164222 589516 164228
rect 589738 163976 589794 163985
rect 589738 163911 589794 163920
rect 589752 162926 589780 163911
rect 589740 162920 589792 162926
rect 589740 162862 589792 162868
rect 590106 162344 590162 162353
rect 590106 162279 590162 162288
rect 589462 160712 589518 160721
rect 589462 160647 589518 160656
rect 589476 160138 589504 160647
rect 589464 160132 589516 160138
rect 589464 160074 589516 160080
rect 588544 159996 588596 160002
rect 588544 159938 588596 159944
rect 588726 159080 588782 159089
rect 588726 159015 588782 159024
rect 587348 150408 587400 150414
rect 587348 150350 587400 150356
rect 587164 149116 587216 149122
rect 587164 149058 587216 149064
rect 586888 146328 586940 146334
rect 586888 146270 586940 146276
rect 585968 145444 586020 145450
rect 585968 145386 586020 145392
rect 585784 144968 585836 144974
rect 585784 144910 585836 144916
rect 584404 140616 584456 140622
rect 584404 140558 584456 140564
rect 583760 133476 583812 133482
rect 583760 133418 583812 133424
rect 584772 132524 584824 132530
rect 584772 132466 584824 132472
rect 584588 118720 584640 118726
rect 584588 118662 584640 118668
rect 583024 113144 583076 113150
rect 583024 113086 583076 113092
rect 584404 109064 584456 109070
rect 584404 109006 584456 109012
rect 583208 107704 583260 107710
rect 583208 107646 583260 107652
rect 583024 104916 583076 104922
rect 583024 104858 583076 104864
rect 581828 84040 581880 84046
rect 581828 83982 581880 83988
rect 583036 59022 583064 104858
rect 583220 80102 583248 107646
rect 583208 80096 583260 80102
rect 583208 80038 583260 80044
rect 584416 71534 584444 109006
rect 584600 81394 584628 118662
rect 584784 107234 584812 132466
rect 585796 122670 585824 144910
rect 586900 144226 586928 146270
rect 586888 144220 586940 144226
rect 586888 144162 586940 144168
rect 585968 128376 586020 128382
rect 585968 128318 586020 128324
rect 585784 122664 585836 122670
rect 585784 122606 585836 122612
rect 585784 113212 585836 113218
rect 585784 113154 585836 113160
rect 584772 107228 584824 107234
rect 584772 107170 584824 107176
rect 584588 81388 584640 81394
rect 584588 81330 584640 81336
rect 584588 75948 584640 75954
rect 584588 75890 584640 75896
rect 584404 71528 584456 71534
rect 584404 71470 584456 71476
rect 583024 59016 583076 59022
rect 583024 58958 583076 58964
rect 579068 57928 579120 57934
rect 579068 57870 579120 57876
rect 581644 57928 581696 57934
rect 581644 57870 581696 57876
rect 579080 57225 579108 57870
rect 579066 57216 579122 57225
rect 579066 57151 579122 57160
rect 578516 55208 578568 55214
rect 578516 55150 578568 55156
rect 578528 54777 578556 55150
rect 578514 54768 578570 54777
rect 578514 54703 578570 54712
rect 584600 53106 584628 75890
rect 585796 67522 585824 113154
rect 585980 91050 586008 128318
rect 587176 128246 587204 149058
rect 588542 144392 588598 144401
rect 588542 144327 588598 144336
rect 587164 128240 587216 128246
rect 587164 128182 587216 128188
rect 587348 125656 587400 125662
rect 587348 125598 587400 125604
rect 586152 120760 586204 120766
rect 586152 120702 586204 120708
rect 586164 111246 586192 120702
rect 586152 111240 586204 111246
rect 586152 111182 586204 111188
rect 587164 110492 587216 110498
rect 587164 110434 587216 110440
rect 586520 96076 586572 96082
rect 586520 96018 586572 96024
rect 586532 93838 586560 96018
rect 586520 93832 586572 93838
rect 586520 93774 586572 93780
rect 585968 91044 586020 91050
rect 585968 90986 586020 90992
rect 587176 69018 587204 110434
rect 587360 96626 587388 125598
rect 588556 124914 588584 144327
rect 588740 143478 588768 159015
rect 589462 157448 589518 157457
rect 589462 157383 589464 157392
rect 589516 157383 589518 157392
rect 589464 157354 589516 157360
rect 589370 155816 589426 155825
rect 589370 155751 589426 155760
rect 589384 154630 589412 155751
rect 589372 154624 589424 154630
rect 589372 154566 589424 154572
rect 589462 154184 589518 154193
rect 589462 154119 589518 154128
rect 589476 153270 589504 154119
rect 589464 153264 589516 153270
rect 589464 153206 589516 153212
rect 589738 152552 589794 152561
rect 590120 152522 590148 162279
rect 589738 152487 589794 152496
rect 590108 152516 590160 152522
rect 589752 151094 589780 152487
rect 590108 152458 590160 152464
rect 589740 151088 589792 151094
rect 589740 151030 589792 151036
rect 589922 150920 589978 150929
rect 589922 150855 589978 150864
rect 589278 149288 589334 149297
rect 589278 149223 589334 149232
rect 589292 149122 589320 149223
rect 589280 149116 589332 149122
rect 589280 149058 589332 149064
rect 589462 147656 589518 147665
rect 589462 147591 589518 147600
rect 589476 146334 589504 147591
rect 589464 146328 589516 146334
rect 589464 146270 589516 146276
rect 589462 146024 589518 146033
rect 589462 145959 589518 145968
rect 589476 144974 589504 145959
rect 589464 144968 589516 144974
rect 589464 144910 589516 144916
rect 588728 143472 588780 143478
rect 588728 143414 588780 143420
rect 589462 141128 589518 141137
rect 589462 141063 589518 141072
rect 589476 140826 589504 141063
rect 589464 140820 589516 140826
rect 589464 140762 589516 140768
rect 589462 139496 589518 139505
rect 589462 139431 589518 139440
rect 589476 137290 589504 139431
rect 589936 138718 589964 150855
rect 590290 142760 590346 142769
rect 590290 142695 590346 142704
rect 590304 140078 590332 142695
rect 590292 140072 590344 140078
rect 590292 140014 590344 140020
rect 589924 138712 589976 138718
rect 589924 138654 589976 138660
rect 589922 137864 589978 137873
rect 589922 137799 589978 137808
rect 589464 137284 589516 137290
rect 589464 137226 589516 137232
rect 589462 136232 589518 136241
rect 589462 136167 589518 136176
rect 589476 135318 589504 136167
rect 589464 135312 589516 135318
rect 589464 135254 589516 135260
rect 589462 134600 589518 134609
rect 589462 134535 589518 134544
rect 589476 133958 589504 134535
rect 589464 133952 589516 133958
rect 589464 133894 589516 133900
rect 589462 132968 589518 132977
rect 589462 132903 589518 132912
rect 589476 132530 589504 132903
rect 589464 132524 589516 132530
rect 589464 132466 589516 132472
rect 588910 131336 588966 131345
rect 588910 131271 588966 131280
rect 588544 124908 588596 124914
rect 588544 124850 588596 124856
rect 588726 124808 588782 124817
rect 588726 124743 588782 124752
rect 588544 98048 588596 98054
rect 588544 97990 588596 97996
rect 587348 96620 587400 96626
rect 587348 96562 587400 96568
rect 587164 69012 587216 69018
rect 587164 68954 587216 68960
rect 585784 67516 585836 67522
rect 585784 67458 585836 67464
rect 588556 55214 588584 97990
rect 588740 86970 588768 124743
rect 588924 99346 588952 131271
rect 589462 129704 589518 129713
rect 589462 129639 589518 129648
rect 589476 128382 589504 129639
rect 589464 128376 589516 128382
rect 589464 128318 589516 128324
rect 589278 126440 589334 126449
rect 589278 126375 589334 126384
rect 589292 125662 589320 126375
rect 589280 125656 589332 125662
rect 589280 125598 589332 125604
rect 589462 121544 589518 121553
rect 589462 121479 589464 121488
rect 589516 121479 589518 121488
rect 589464 121450 589516 121456
rect 589936 120766 589964 137799
rect 590106 128072 590162 128081
rect 590106 128007 590162 128016
rect 589924 120760 589976 120766
rect 589924 120702 589976 120708
rect 589462 119912 589518 119921
rect 589462 119847 589518 119856
rect 589476 118726 589504 119847
rect 589464 118720 589516 118726
rect 589464 118662 589516 118668
rect 589462 118280 589518 118289
rect 589462 118215 589518 118224
rect 589476 117366 589504 118215
rect 589464 117360 589516 117366
rect 589464 117302 589516 117308
rect 589462 116648 589518 116657
rect 589462 116583 589518 116592
rect 589476 116006 589504 116583
rect 589464 116000 589516 116006
rect 589464 115942 589516 115948
rect 589922 115016 589978 115025
rect 589922 114951 589978 114960
rect 589462 113384 589518 113393
rect 589462 113319 589518 113328
rect 589476 113218 589504 113319
rect 589464 113212 589516 113218
rect 589464 113154 589516 113160
rect 589646 111752 589702 111761
rect 589646 111687 589702 111696
rect 589660 110498 589688 111687
rect 589648 110492 589700 110498
rect 589648 110434 589700 110440
rect 589462 110120 589518 110129
rect 589462 110055 589518 110064
rect 589476 109070 589504 110055
rect 589464 109064 589516 109070
rect 589464 109006 589516 109012
rect 589462 108488 589518 108497
rect 589462 108423 589518 108432
rect 589476 107710 589504 108423
rect 589464 107704 589516 107710
rect 589464 107646 589516 107652
rect 589462 106856 589518 106865
rect 589462 106791 589518 106800
rect 589476 106350 589504 106791
rect 589464 106344 589516 106350
rect 589464 106286 589516 106292
rect 589462 105224 589518 105233
rect 589462 105159 589518 105168
rect 589476 104922 589504 105159
rect 589464 104916 589516 104922
rect 589464 104858 589516 104864
rect 589462 103592 589518 103601
rect 589462 103527 589464 103536
rect 589516 103527 589518 103536
rect 589464 103498 589516 103504
rect 589370 101960 589426 101969
rect 589370 101895 589426 101904
rect 588912 99340 588964 99346
rect 588912 99282 588964 99288
rect 589384 98054 589412 101895
rect 589372 98048 589424 98054
rect 589372 97990 589424 97996
rect 588728 86964 588780 86970
rect 588728 86906 588780 86912
rect 589936 74526 589964 114951
rect 590120 96082 590148 128007
rect 590290 123176 590346 123185
rect 590290 123111 590346 123120
rect 590304 115258 590332 123111
rect 590292 115252 590344 115258
rect 590292 115194 590344 115200
rect 591316 103426 591344 209782
rect 632164 209766 632500 209782
rect 666572 184793 666600 509206
rect 666756 245993 666784 993278
rect 667388 993200 667440 993206
rect 667388 993142 667440 993148
rect 666928 991772 666980 991778
rect 666928 991714 666980 991720
rect 666742 245984 666798 245993
rect 666742 245919 666798 245928
rect 666940 245721 666968 991714
rect 667204 403436 667256 403442
rect 667204 403378 667256 403384
rect 667216 403170 667244 403378
rect 667204 403164 667256 403170
rect 667204 403106 667256 403112
rect 667112 338156 667164 338162
rect 667112 338098 667164 338104
rect 666926 245712 666982 245721
rect 666926 245647 666982 245656
rect 666742 222320 666798 222329
rect 666742 222255 666798 222264
rect 666558 184784 666614 184793
rect 666558 184719 666614 184728
rect 666756 109381 666784 222255
rect 666928 196716 666980 196722
rect 666928 196658 666980 196664
rect 666940 192681 666968 196658
rect 666926 192672 666982 192681
rect 666926 192607 666982 192616
rect 666928 192296 666980 192302
rect 666928 192238 666980 192244
rect 666940 160041 666968 192238
rect 667124 178090 667152 338098
rect 667400 246129 667428 993142
rect 667664 985040 667716 985046
rect 667664 984982 667716 984988
rect 667386 246120 667442 246129
rect 667386 246055 667442 246064
rect 667480 220856 667532 220862
rect 667480 220798 667532 220804
rect 667492 210610 667520 220798
rect 667676 215294 667704 984982
rect 667952 215294 667980 994366
rect 672724 990276 672776 990282
rect 672724 990218 672776 990224
rect 668308 988916 668360 988922
rect 668308 988858 668360 988864
rect 668124 987556 668176 987562
rect 668124 987498 668176 987504
rect 668136 245993 668164 987498
rect 668122 245984 668178 245993
rect 668122 245919 668178 245928
rect 668320 245721 668348 988858
rect 669964 985992 670016 985998
rect 669964 985934 670016 985940
rect 669976 935950 670004 985934
rect 671344 985176 671396 985182
rect 671344 985118 671396 985124
rect 671356 937378 671384 985118
rect 671528 948116 671580 948122
rect 671528 948058 671580 948064
rect 671540 938738 671568 948058
rect 671528 938732 671580 938738
rect 671528 938674 671580 938680
rect 672736 938602 672764 990218
rect 675404 966521 675432 966723
rect 675390 966512 675446 966521
rect 675390 966447 675446 966456
rect 673276 966340 673328 966346
rect 673276 966282 673328 966288
rect 675116 966340 675168 966346
rect 675116 966282 675168 966288
rect 672906 959168 672962 959177
rect 672906 959103 672962 959112
rect 672724 938596 672776 938602
rect 672724 938538 672776 938544
rect 672724 937576 672776 937582
rect 672724 937518 672776 937524
rect 671344 937372 671396 937378
rect 671344 937314 671396 937320
rect 672540 937100 672592 937106
rect 672540 937042 672592 937048
rect 669964 935944 670016 935950
rect 669964 935886 670016 935892
rect 670976 935808 671028 935814
rect 670976 935750 671028 935756
rect 670608 927444 670660 927450
rect 670608 927386 670660 927392
rect 670424 879096 670476 879102
rect 670424 879038 670476 879044
rect 670056 865292 670108 865298
rect 670056 865234 670108 865240
rect 669780 789404 669832 789410
rect 669780 789346 669832 789352
rect 669044 782536 669096 782542
rect 669044 782478 669096 782484
rect 668582 728784 668638 728793
rect 668582 728719 668638 728728
rect 668596 663814 668624 728719
rect 669056 709782 669084 782478
rect 669410 775024 669466 775033
rect 669410 774959 669466 774968
rect 669228 743844 669280 743850
rect 669228 743786 669280 743792
rect 669044 709776 669096 709782
rect 669044 709718 669096 709724
rect 668766 688664 668822 688673
rect 668766 688599 668822 688608
rect 668584 663808 668636 663814
rect 668584 663750 668636 663756
rect 668780 615806 668808 688599
rect 669042 685128 669098 685137
rect 669042 685063 669098 685072
rect 669056 617273 669084 685063
rect 669240 663950 669268 743786
rect 669424 710705 669452 774959
rect 669596 745272 669648 745278
rect 669596 745214 669648 745220
rect 669608 743850 669636 745214
rect 669596 743844 669648 743850
rect 669596 743786 669648 743792
rect 669594 735176 669650 735185
rect 669594 735111 669650 735120
rect 669410 710696 669466 710705
rect 669410 710631 669466 710640
rect 669608 666126 669636 735111
rect 669792 709646 669820 789346
rect 670068 755070 670096 865234
rect 670240 783760 670292 783766
rect 670240 783702 670292 783708
rect 670056 755064 670108 755070
rect 670056 755006 670108 755012
rect 669964 750100 670016 750106
rect 669964 750042 670016 750048
rect 669780 709640 669832 709646
rect 669780 709582 669832 709588
rect 669780 685908 669832 685914
rect 669780 685850 669832 685856
rect 669596 666120 669648 666126
rect 669596 666062 669648 666068
rect 669228 663944 669280 663950
rect 669228 663886 669280 663892
rect 669228 650072 669280 650078
rect 669228 650014 669280 650020
rect 669042 617264 669098 617273
rect 669042 617199 669098 617208
rect 668768 615800 668820 615806
rect 668768 615742 668820 615748
rect 668584 610156 668636 610162
rect 668584 610098 668636 610104
rect 668306 245712 668362 245721
rect 668306 245647 668362 245656
rect 668400 222624 668452 222630
rect 668400 222566 668452 222572
rect 668412 222222 668440 222566
rect 668400 222216 668452 222222
rect 668400 222158 668452 222164
rect 668398 219464 668454 219473
rect 668398 219399 668454 219408
rect 667676 215266 667888 215294
rect 667952 215266 668164 215294
rect 667296 210588 667348 210594
rect 667492 210582 667796 210610
rect 667296 210530 667348 210536
rect 667112 178084 667164 178090
rect 667112 178026 667164 178032
rect 666926 160032 666982 160041
rect 666926 159967 666982 159976
rect 667308 132530 667336 210530
rect 667480 210316 667532 210322
rect 667480 210258 667532 210264
rect 667492 132802 667520 210258
rect 667768 202874 667796 210582
rect 667584 202846 667796 202874
rect 667584 201494 667612 202846
rect 667584 201466 667704 201494
rect 667676 196586 667704 201466
rect 667860 196722 667888 215266
rect 667848 196716 667900 196722
rect 667848 196658 667900 196664
rect 667664 196580 667716 196586
rect 667664 196522 667716 196528
rect 667848 196376 667900 196382
rect 667848 196318 667900 196324
rect 667860 179414 667888 196318
rect 668136 187785 668164 215266
rect 668122 187776 668178 187785
rect 668122 187711 668178 187720
rect 668216 183524 668268 183530
rect 668216 183466 668268 183472
rect 667768 179386 667888 179414
rect 667768 176866 667796 179386
rect 667938 177984 667994 177993
rect 667938 177919 667940 177928
rect 667992 177919 667994 177928
rect 667940 177890 667992 177896
rect 667756 176860 667808 176866
rect 667756 176802 667808 176808
rect 667940 174752 667992 174758
rect 667938 174720 667940 174729
rect 667992 174720 667994 174729
rect 667938 174655 667994 174664
rect 667940 169720 667992 169726
rect 667938 169688 667940 169697
rect 667992 169688 667994 169697
rect 667938 169623 667994 169632
rect 668032 164960 668084 164966
rect 668030 164928 668032 164937
rect 668084 164928 668086 164937
rect 668030 164863 668086 164872
rect 667480 132796 667532 132802
rect 667480 132738 667532 132744
rect 667296 132524 667348 132530
rect 667296 132466 667348 132472
rect 667940 130960 667992 130966
rect 667940 130902 667992 130908
rect 667952 130665 667980 130902
rect 667938 130656 667994 130665
rect 667938 130591 667994 130600
rect 667940 126200 667992 126206
rect 667940 126142 667992 126148
rect 667952 125769 667980 126142
rect 667938 125760 667994 125769
rect 667938 125695 667994 125704
rect 668228 120873 668256 183466
rect 668412 132494 668440 219399
rect 668596 168201 668624 610098
rect 668860 598800 668912 598806
rect 668860 598742 668912 598748
rect 668872 525842 668900 598742
rect 669042 593600 669098 593609
rect 669042 593535 669098 593544
rect 669056 529378 669084 593535
rect 669240 571402 669268 650014
rect 669594 642152 669650 642161
rect 669594 642087 669650 642096
rect 669608 572966 669636 642087
rect 669792 619886 669820 685850
rect 669780 619880 669832 619886
rect 669780 619822 669832 619828
rect 669596 572960 669648 572966
rect 669596 572902 669648 572908
rect 669228 571396 669280 571402
rect 669228 571338 669280 571344
rect 669780 554804 669832 554810
rect 669780 554746 669832 554752
rect 669044 529372 669096 529378
rect 669044 529314 669096 529320
rect 668860 525836 668912 525842
rect 668860 525778 668912 525784
rect 669792 484022 669820 554746
rect 669780 484016 669832 484022
rect 669780 483958 669832 483964
rect 668768 474088 668820 474094
rect 668768 474030 668820 474036
rect 668582 168192 668638 168201
rect 668582 168127 668638 168136
rect 668582 165744 668638 165753
rect 668582 165679 668638 165688
rect 668596 163305 668624 165679
rect 668582 163296 668638 163305
rect 668582 163231 668638 163240
rect 668780 158409 668808 474030
rect 669780 353320 669832 353326
rect 669780 353262 669832 353268
rect 669596 350736 669648 350742
rect 669596 350678 669648 350684
rect 669226 342136 669282 342145
rect 669226 342071 669282 342080
rect 669240 325514 669268 342071
rect 669608 335646 669636 350678
rect 669596 335640 669648 335646
rect 669596 335582 669648 335588
rect 669792 325650 669820 353262
rect 669780 325644 669832 325650
rect 669780 325586 669832 325592
rect 669228 325508 669280 325514
rect 669228 325450 669280 325456
rect 669780 300824 669832 300830
rect 669780 300766 669832 300772
rect 669320 268524 669372 268530
rect 669320 268466 669372 268472
rect 669332 267918 669360 268466
rect 669320 267912 669372 267918
rect 669320 267854 669372 267860
rect 669320 265600 669372 265606
rect 669320 265542 669372 265548
rect 669332 264926 669360 265542
rect 669320 264920 669372 264926
rect 669320 264862 669372 264868
rect 669412 262132 669464 262138
rect 669412 262074 669464 262080
rect 669136 259888 669188 259894
rect 669136 259830 669188 259836
rect 669148 242049 669176 259830
rect 669424 250442 669452 262074
rect 669596 253224 669648 253230
rect 669596 253166 669648 253172
rect 669412 250436 669464 250442
rect 669412 250378 669464 250384
rect 669320 244928 669372 244934
rect 669320 244870 669372 244876
rect 669134 242040 669190 242049
rect 669134 241975 669190 241984
rect 669134 225040 669190 225049
rect 669134 224975 669190 224984
rect 669148 224890 669176 224975
rect 669148 224862 669268 224890
rect 668950 223680 669006 223689
rect 668950 223615 669006 223624
rect 668964 223530 668992 223615
rect 668872 223502 668992 223530
rect 668872 219434 668900 223502
rect 669044 221060 669096 221066
rect 669044 221002 669096 221008
rect 668872 219406 668992 219434
rect 668766 158400 668822 158409
rect 668584 158364 668636 158370
rect 668766 158335 668822 158344
rect 668584 158306 668636 158312
rect 668596 143721 668624 158306
rect 668768 150272 668820 150278
rect 668766 150240 668768 150249
rect 668820 150240 668822 150249
rect 668766 150175 668822 150184
rect 668768 145580 668820 145586
rect 668768 145522 668820 145528
rect 668780 145353 668808 145522
rect 668766 145344 668822 145353
rect 668766 145279 668822 145288
rect 668582 143712 668638 143721
rect 668582 143647 668638 143656
rect 668676 140480 668728 140486
rect 668674 140448 668676 140457
rect 668728 140448 668730 140457
rect 668674 140383 668730 140392
rect 668766 138680 668822 138689
rect 668766 138615 668822 138624
rect 668780 138446 668808 138615
rect 668768 138440 668820 138446
rect 668768 138382 668820 138388
rect 668768 136536 668820 136542
rect 668768 136478 668820 136484
rect 668780 135561 668808 136478
rect 668766 135552 668822 135561
rect 668766 135487 668822 135496
rect 668412 132466 668808 132494
rect 668780 131170 668808 132466
rect 668768 131164 668820 131170
rect 668768 131106 668820 131112
rect 668584 129804 668636 129810
rect 668584 129746 668636 129752
rect 668214 120864 668270 120873
rect 668214 120799 668270 120808
rect 667940 117836 667992 117842
rect 667940 117778 667992 117784
rect 667952 117609 667980 117778
rect 667938 117600 667994 117609
rect 667938 117535 667994 117544
rect 668400 115864 668452 115870
rect 668398 115832 668400 115841
rect 668452 115832 668454 115841
rect 668398 115767 668454 115776
rect 668400 114368 668452 114374
rect 668398 114336 668400 114345
rect 668452 114336 668454 114345
rect 668398 114271 668454 114280
rect 668032 112940 668084 112946
rect 668032 112882 668084 112888
rect 668044 112713 668072 112882
rect 668030 112704 668086 112713
rect 668030 112639 668086 112648
rect 666742 109372 666798 109381
rect 666742 109307 666798 109316
rect 591304 103420 591356 103426
rect 591304 103362 591356 103368
rect 668596 102921 668624 129746
rect 668780 113174 668808 131106
rect 668964 128382 668992 219406
rect 669056 179414 669084 221002
rect 669240 195974 669268 224862
rect 669148 195946 669268 195974
rect 669148 190454 669176 195946
rect 669332 192302 669360 244870
rect 669320 192296 669372 192302
rect 669320 192238 669372 192244
rect 669148 190426 669268 190454
rect 669240 189074 669268 190426
rect 669240 189046 669544 189074
rect 669228 182912 669280 182918
rect 669226 182880 669228 182889
rect 669280 182880 669282 182889
rect 669226 182815 669282 182824
rect 669056 179386 669176 179414
rect 669148 176633 669176 179386
rect 669134 176624 669190 176633
rect 669134 176559 669190 176568
rect 669516 173894 669544 189046
rect 669148 173866 669544 173894
rect 669148 166994 669176 173866
rect 669412 171964 669464 171970
rect 669412 171906 669464 171912
rect 669148 166966 669268 166994
rect 669240 161474 669268 166966
rect 669148 161446 669268 161474
rect 669148 129946 669176 161446
rect 669424 149054 669452 171906
rect 669412 149048 669464 149054
rect 669412 148990 669464 148996
rect 669136 129940 669188 129946
rect 669136 129882 669188 129888
rect 669148 129810 669176 129882
rect 669136 129804 669188 129810
rect 669136 129746 669188 129752
rect 669228 129056 669280 129062
rect 669226 129024 669228 129033
rect 669280 129024 669282 129033
rect 669226 128959 669282 128968
rect 668952 128376 669004 128382
rect 668952 128318 669004 128324
rect 668964 113174 668992 128318
rect 669608 126206 669636 253166
rect 669792 130966 669820 300766
rect 669976 174758 670004 750042
rect 670252 708830 670280 783702
rect 670436 754662 670464 879038
rect 670424 754656 670476 754662
rect 670424 754598 670476 754604
rect 670422 734496 670478 734505
rect 670422 734431 670478 734440
rect 670240 708824 670292 708830
rect 670240 708766 670292 708772
rect 670148 705084 670200 705090
rect 670148 705026 670200 705032
rect 669964 174752 670016 174758
rect 669964 174694 670016 174700
rect 670160 169726 670188 705026
rect 670436 662862 670464 734431
rect 670424 662856 670476 662862
rect 670424 662798 670476 662804
rect 670332 659932 670384 659938
rect 670332 659874 670384 659880
rect 670148 169720 670200 169726
rect 670148 169662 670200 169668
rect 669964 167884 670016 167890
rect 669964 167826 670016 167832
rect 669780 130960 669832 130966
rect 669780 130902 669832 130908
rect 669596 126200 669648 126206
rect 669596 126142 669648 126148
rect 669228 124160 669280 124166
rect 669226 124128 669228 124137
rect 669280 124128 669282 124137
rect 669226 124063 669282 124072
rect 669136 119264 669188 119270
rect 669134 119232 669136 119241
rect 669188 119232 669190 119241
rect 669134 119167 669190 119176
rect 669976 117842 670004 167826
rect 670344 164966 670372 659874
rect 670620 217977 670648 927386
rect 670792 788044 670844 788050
rect 670792 787986 670844 787992
rect 670804 711278 670832 787986
rect 670988 758742 671016 935750
rect 671804 935672 671856 935678
rect 671804 935614 671856 935620
rect 671344 909492 671396 909498
rect 671344 909434 671396 909440
rect 671160 866720 671212 866726
rect 671160 866662 671212 866668
rect 670976 758736 671028 758742
rect 670976 758678 671028 758684
rect 671172 753438 671200 866662
rect 671356 761598 671384 909434
rect 671528 881884 671580 881890
rect 671528 881826 671580 881832
rect 671540 869038 671568 881826
rect 671528 869032 671580 869038
rect 671528 868974 671580 868980
rect 671528 777028 671580 777034
rect 671528 776970 671580 776976
rect 671344 761592 671396 761598
rect 671344 761534 671396 761540
rect 671344 757444 671396 757450
rect 671344 757386 671396 757392
rect 671356 756254 671384 757386
rect 671356 756226 671476 756254
rect 671160 753432 671212 753438
rect 671160 753374 671212 753380
rect 671250 734224 671306 734233
rect 671250 734159 671306 734168
rect 671264 727274 671292 734159
rect 671448 727274 671476 756226
rect 671540 746594 671568 776970
rect 671816 758402 671844 935614
rect 672354 868048 672410 868057
rect 672354 867983 672410 867992
rect 672172 786684 672224 786690
rect 672172 786626 672224 786632
rect 671988 759892 672040 759898
rect 671988 759834 672040 759840
rect 671804 758396 671856 758402
rect 671804 758338 671856 758344
rect 671804 758260 671856 758266
rect 671804 758202 671856 758208
rect 671540 746566 671660 746594
rect 671264 727246 671384 727274
rect 671448 727246 671568 727274
rect 670976 715012 671028 715018
rect 670976 714954 671028 714960
rect 670792 711272 670844 711278
rect 670792 711214 670844 711220
rect 670988 669798 671016 714954
rect 671160 714060 671212 714066
rect 671160 714002 671212 714008
rect 670976 669792 671028 669798
rect 670976 669734 671028 669740
rect 671172 669662 671200 714002
rect 671160 669656 671212 669662
rect 671160 669598 671212 669604
rect 671160 669384 671212 669390
rect 671160 669326 671212 669332
rect 670976 667276 671028 667282
rect 670976 667218 671028 667224
rect 670792 647760 670844 647766
rect 670792 647702 670844 647708
rect 670804 647465 670832 647702
rect 670790 647456 670846 647465
rect 670790 647391 670846 647400
rect 670792 643680 670844 643686
rect 670792 643622 670844 643628
rect 670804 641918 670832 643622
rect 670792 641912 670844 641918
rect 670792 641854 670844 641860
rect 670792 641776 670844 641782
rect 670792 641718 670844 641724
rect 670804 640082 670832 641718
rect 670792 640076 670844 640082
rect 670792 640018 670844 640024
rect 670792 623824 670844 623830
rect 670792 623766 670844 623772
rect 670804 580038 670832 623766
rect 670988 622470 671016 667218
rect 671172 624102 671200 669326
rect 671356 669066 671384 727246
rect 671540 712910 671568 727246
rect 671632 712994 671660 746566
rect 671816 713726 671844 758202
rect 672000 715358 672028 759834
rect 671988 715352 672040 715358
rect 671988 715294 672040 715300
rect 671804 713720 671856 713726
rect 671804 713662 671856 713668
rect 671896 713244 671948 713250
rect 671896 713186 671948 713192
rect 671632 712966 671752 712994
rect 671528 712904 671580 712910
rect 671528 712846 671580 712852
rect 671724 712722 671752 712966
rect 671540 712694 671752 712722
rect 671540 708422 671568 712694
rect 671712 712428 671764 712434
rect 671712 712370 671764 712376
rect 671528 708416 671580 708422
rect 671528 708358 671580 708364
rect 671724 673454 671752 712370
rect 671908 673454 671936 713186
rect 672184 712094 672212 786626
rect 672368 751806 672396 867983
rect 672552 760306 672580 937042
rect 672540 760300 672592 760306
rect 672540 760242 672592 760248
rect 672736 759558 672764 937518
rect 672920 932958 672948 959103
rect 673092 956412 673144 956418
rect 673092 956354 673144 956360
rect 672908 932952 672960 932958
rect 672908 932894 672960 932900
rect 673104 930170 673132 956354
rect 673288 933094 673316 966282
rect 675128 966090 675156 966282
rect 675128 966062 675418 966090
rect 675772 965161 675800 965435
rect 675758 965152 675814 965161
rect 675758 965087 675814 965096
rect 675220 963581 675418 963609
rect 675220 963393 675248 963581
rect 675206 963384 675262 963393
rect 675206 963319 675262 963328
rect 675312 963070 675432 963098
rect 675312 963030 675340 963070
rect 674668 963002 675340 963030
rect 675404 963016 675432 963070
rect 674288 961920 674340 961926
rect 674288 961862 674340 961868
rect 674104 957908 674156 957914
rect 674104 957850 674156 957856
rect 673276 933088 673328 933094
rect 673276 933030 673328 933036
rect 674116 931462 674144 957850
rect 674300 932249 674328 961862
rect 674470 952232 674526 952241
rect 674470 952167 674526 952176
rect 674484 933473 674512 952167
rect 674470 933464 674526 933473
rect 674470 933399 674526 933408
rect 674668 932657 674696 963002
rect 675128 962390 675418 962418
rect 675128 961926 675156 962390
rect 675758 962024 675814 962033
rect 675758 961959 675814 961968
rect 675116 961920 675168 961926
rect 675116 961862 675168 961868
rect 675772 961755 675800 961959
rect 674930 959440 674986 959449
rect 674930 959375 674986 959384
rect 674944 954530 674972 959375
rect 675128 959262 675418 959290
rect 675128 959177 675156 959262
rect 675114 959168 675170 959177
rect 675114 959103 675170 959112
rect 675772 958361 675800 958732
rect 675758 958352 675814 958361
rect 675758 958287 675814 958296
rect 675312 958174 675432 958202
rect 675312 958066 675340 958174
rect 675128 958038 675340 958066
rect 675404 958052 675432 958174
rect 675128 957914 675156 958038
rect 675116 957908 675168 957914
rect 675116 957850 675168 957856
rect 675128 957426 675418 957454
rect 675128 956418 675156 957426
rect 675300 957364 675352 957370
rect 675300 957306 675352 957312
rect 675116 956412 675168 956418
rect 675116 956354 675168 956360
rect 675312 955482 675340 957306
rect 675758 956448 675814 956457
rect 675758 956383 675814 956392
rect 675772 956216 675800 956383
rect 675312 955454 675524 955482
rect 675496 955060 675524 955454
rect 674944 954502 675064 954530
rect 675036 954258 675064 954502
rect 675036 954230 675156 954258
rect 674930 948968 674986 948977
rect 674930 948903 674986 948912
rect 674944 941905 674972 948903
rect 675128 946694 675156 954230
rect 675680 954009 675708 954380
rect 675666 954000 675722 954009
rect 675666 953935 675722 953944
rect 675220 953754 675340 953782
rect 675220 949454 675248 953754
rect 675312 953714 675340 953754
rect 675404 953714 675432 953768
rect 675312 953686 675432 953714
rect 675404 952241 675432 952544
rect 675390 952232 675446 952241
rect 675390 952167 675446 952176
rect 677506 951552 677562 951561
rect 677506 951487 677562 951496
rect 675852 949476 675904 949482
rect 675220 949426 675852 949454
rect 675852 949418 675904 949424
rect 675942 949240 675998 949249
rect 675942 949175 675998 949184
rect 675956 948802 675984 949175
rect 675944 948796 675996 948802
rect 675944 948738 675996 948744
rect 675128 946666 675248 946694
rect 674930 941896 674986 941905
rect 675220 941848 675248 946666
rect 675850 941896 675906 941905
rect 674930 941831 674986 941840
rect 675128 941820 675248 941848
rect 675484 941860 675536 941866
rect 674930 938360 674986 938369
rect 674930 938295 674986 938304
rect 674944 937106 674972 938295
rect 674932 937100 674984 937106
rect 674932 937042 674984 937048
rect 675128 934153 675156 941820
rect 675850 941831 675906 941840
rect 675484 941802 675536 941808
rect 675496 940001 675524 941802
rect 675482 939992 675538 940001
rect 675482 939927 675538 939936
rect 675666 939584 675722 939593
rect 675666 939519 675722 939528
rect 675298 939176 675354 939185
rect 675298 939111 675354 939120
rect 675312 938738 675340 939111
rect 675482 938768 675538 938777
rect 675300 938732 675352 938738
rect 675482 938703 675538 938712
rect 675300 938674 675352 938680
rect 675496 938602 675524 938703
rect 675484 938596 675536 938602
rect 675484 938538 675536 938544
rect 675680 938482 675708 939519
rect 675496 938466 675708 938482
rect 675484 938460 675708 938466
rect 675536 938454 675708 938460
rect 675484 938402 675536 938408
rect 675298 937952 675354 937961
rect 675298 937887 675354 937896
rect 675312 937242 675340 937887
rect 675484 937576 675536 937582
rect 675482 937544 675484 937553
rect 675536 937544 675538 937553
rect 675482 937479 675538 937488
rect 675484 937372 675536 937378
rect 675484 937314 675536 937320
rect 675300 937236 675352 937242
rect 675300 937178 675352 937184
rect 675496 937145 675524 937314
rect 675482 937136 675538 937145
rect 675482 937071 675538 937080
rect 675666 936728 675722 936737
rect 675666 936663 675722 936672
rect 675482 936320 675538 936329
rect 675482 936255 675538 936264
rect 675496 935950 675524 936255
rect 675484 935944 675536 935950
rect 675298 935912 675354 935921
rect 675484 935886 675536 935892
rect 675298 935847 675354 935856
rect 675312 935678 675340 935847
rect 675484 935808 675536 935814
rect 675680 935762 675708 936663
rect 675536 935756 675708 935762
rect 675484 935750 675708 935756
rect 675496 935734 675708 935750
rect 675300 935672 675352 935678
rect 675300 935614 675352 935620
rect 675864 934697 675892 941831
rect 675850 934688 675906 934697
rect 675850 934623 675906 934632
rect 675114 934144 675170 934153
rect 675114 934079 675170 934088
rect 675298 933872 675354 933881
rect 675298 933807 675354 933816
rect 675312 932958 675340 933807
rect 675484 933088 675536 933094
rect 675482 933056 675484 933065
rect 675536 933056 675538 933065
rect 675482 932991 675538 933000
rect 675300 932952 675352 932958
rect 675300 932894 675352 932900
rect 674654 932648 674710 932657
rect 674654 932583 674710 932592
rect 674286 932240 674342 932249
rect 674286 932175 674342 932184
rect 674104 931456 674156 931462
rect 675484 931456 675536 931462
rect 674104 931398 674156 931404
rect 675482 931424 675484 931433
rect 675536 931424 675538 931433
rect 675482 931359 675538 931368
rect 677520 931161 677548 951487
rect 683302 950056 683358 950065
rect 683302 949991 683358 950000
rect 678244 949476 678296 949482
rect 678244 949418 678296 949424
rect 677506 931152 677562 931161
rect 677506 931087 677562 931096
rect 675482 930200 675538 930209
rect 673092 930164 673144 930170
rect 675482 930135 675484 930144
rect 673092 930106 673144 930112
rect 675536 930135 675538 930144
rect 675484 930106 675536 930112
rect 678256 930102 678284 949418
rect 682384 948796 682436 948802
rect 682384 948738 682436 948744
rect 682396 935241 682424 948738
rect 683316 935649 683344 949991
rect 703694 940508 703722 940644
rect 704154 940508 704182 940644
rect 704614 940508 704642 940644
rect 705074 940508 705102 940644
rect 705534 940508 705562 940644
rect 705994 940508 706022 940644
rect 706454 940508 706482 940644
rect 706914 940508 706942 940644
rect 707374 940508 707402 940644
rect 707834 940508 707862 940644
rect 708294 940508 708322 940644
rect 708754 940508 708782 940644
rect 709214 940508 709242 940644
rect 683302 935640 683358 935649
rect 683302 935575 683358 935584
rect 682382 935232 682438 935241
rect 682382 935167 682438 935176
rect 678244 930096 678296 930102
rect 678244 930038 678296 930044
rect 683120 930096 683172 930102
rect 683120 930038 683172 930044
rect 675482 929792 675538 929801
rect 675482 929727 675538 929736
rect 675496 928810 675524 929727
rect 683132 929529 683160 930038
rect 683118 929520 683174 929529
rect 683118 929455 683174 929464
rect 673276 928804 673328 928810
rect 673276 928746 673328 928752
rect 675484 928804 675536 928810
rect 675484 928746 675536 928752
rect 672998 864240 673054 864249
rect 672998 864175 673054 864184
rect 672724 759552 672776 759558
rect 672724 759494 672776 759500
rect 672632 759076 672684 759082
rect 672632 759018 672684 759024
rect 672356 751800 672408 751806
rect 672356 751742 672408 751748
rect 672356 751324 672408 751330
rect 672356 751266 672408 751272
rect 672368 727274 672396 751266
rect 672368 727246 672580 727274
rect 672552 724514 672580 727246
rect 672460 724486 672580 724514
rect 672460 715714 672488 724486
rect 672644 715834 672672 759018
rect 673012 752321 673040 864175
rect 673288 775574 673316 928746
rect 675482 928568 675538 928577
rect 675482 928503 675538 928512
rect 675496 927450 675524 928503
rect 675484 927444 675536 927450
rect 675484 927386 675536 927392
rect 675300 879096 675352 879102
rect 675300 879038 675352 879044
rect 675312 877146 675340 879038
rect 675772 877169 675800 877540
rect 675758 877160 675814 877169
rect 675312 877118 675432 877146
rect 675404 876860 675432 877118
rect 675758 877095 675814 877104
rect 675298 876480 675354 876489
rect 675298 876415 675354 876424
rect 675312 876262 675340 876415
rect 675312 876234 675418 876262
rect 675404 874041 675432 874412
rect 675390 874032 675446 874041
rect 675390 873967 675446 873976
rect 674484 873854 675340 873882
rect 673828 868080 673880 868086
rect 673828 868022 673880 868028
rect 673104 775546 673316 775574
rect 673104 754474 673132 775546
rect 673274 773664 673330 773673
rect 673274 773599 673330 773608
rect 673288 765914 673316 773599
rect 673288 765886 673408 765914
rect 673104 754446 673224 754474
rect 672998 752312 673054 752321
rect 672998 752247 673054 752256
rect 673000 752140 673052 752146
rect 673000 752082 673052 752088
rect 673012 750734 673040 752082
rect 673196 752026 673224 754446
rect 673380 752146 673408 765886
rect 673644 765332 673696 765338
rect 673644 765274 673696 765280
rect 673656 761462 673684 765274
rect 673840 761938 673868 868022
rect 674484 854321 674512 873854
rect 675312 873746 675340 873854
rect 675404 873746 675432 873868
rect 675312 873718 675432 873746
rect 675772 872817 675800 873188
rect 675758 872808 675814 872817
rect 675758 872743 675814 872752
rect 675404 872273 675432 872576
rect 675390 872264 675446 872273
rect 675390 872199 675446 872208
rect 674668 869774 675064 869802
rect 674470 854312 674526 854321
rect 674470 854247 674526 854256
rect 674472 783896 674524 783902
rect 674472 783838 674524 783844
rect 674012 782672 674064 782678
rect 674012 782614 674064 782620
rect 674024 778546 674052 782614
rect 674288 779204 674340 779210
rect 674288 779146 674340 779152
rect 673932 778518 674052 778546
rect 673932 765082 673960 778518
rect 674104 778388 674156 778394
rect 674104 778330 674156 778336
rect 674116 775574 674144 778330
rect 674024 775546 674144 775574
rect 674024 772814 674052 775546
rect 674024 772786 674236 772814
rect 674208 771434 674236 772786
rect 674116 771406 674236 771434
rect 674116 765338 674144 771406
rect 674104 765332 674156 765338
rect 674104 765274 674156 765280
rect 673932 765054 674236 765082
rect 673828 761932 673880 761938
rect 673828 761874 673880 761880
rect 673828 761796 673880 761802
rect 673828 761738 673880 761744
rect 673644 761456 673696 761462
rect 673644 761398 673696 761404
rect 673840 753030 673868 761738
rect 674012 761456 674064 761462
rect 674012 761398 674064 761404
rect 673828 753024 673880 753030
rect 673828 752966 673880 752972
rect 673368 752140 673420 752146
rect 673368 752082 673420 752088
rect 673196 751998 673408 752026
rect 673380 750734 673408 751998
rect 674024 750734 674052 761398
rect 674208 760394 674236 765054
rect 673012 750706 673224 750734
rect 673000 738472 673052 738478
rect 673000 738414 673052 738420
rect 672814 730144 672870 730153
rect 672814 730079 672870 730088
rect 672632 715828 672684 715834
rect 672632 715770 672684 715776
rect 672460 715686 672580 715714
rect 672356 715624 672408 715630
rect 672356 715566 672408 715572
rect 672368 714542 672396 715566
rect 672356 714536 672408 714542
rect 672356 714478 672408 714484
rect 672172 712088 672224 712094
rect 672172 712030 672224 712036
rect 672264 706308 672316 706314
rect 672264 706250 672316 706256
rect 672080 698488 672132 698494
rect 672080 698430 672132 698436
rect 672092 698294 672120 698430
rect 672276 698294 672304 706250
rect 671264 669038 671384 669066
rect 671540 673426 671752 673454
rect 671816 673426 671936 673454
rect 672000 698266 672120 698294
rect 672184 698266 672304 698294
rect 671264 664170 671292 669038
rect 671540 667758 671568 673426
rect 671816 668574 671844 673426
rect 671804 668568 671856 668574
rect 671804 668510 671856 668516
rect 672000 668250 672028 698266
rect 672184 678974 672212 698266
rect 672552 692774 672580 715686
rect 672276 692746 672580 692774
rect 672276 688634 672304 692746
rect 672276 688606 672396 688634
rect 671908 668222 672028 668250
rect 672092 678946 672212 678974
rect 671908 667978 671936 668222
rect 671908 667950 672028 667978
rect 671802 667856 671858 667865
rect 671802 667791 671858 667800
rect 671528 667752 671580 667758
rect 671528 667694 671580 667700
rect 671620 667616 671672 667622
rect 671620 667558 671672 667564
rect 671632 666618 671660 667558
rect 671632 666590 671752 666618
rect 671264 664142 671384 664170
rect 671356 661638 671384 664142
rect 671344 661632 671396 661638
rect 671344 661574 671396 661580
rect 671344 661156 671396 661162
rect 671344 661098 671396 661104
rect 671160 624096 671212 624102
rect 671160 624038 671212 624044
rect 671160 623960 671212 623966
rect 671160 623902 671212 623908
rect 670976 622464 671028 622470
rect 670976 622406 671028 622412
rect 670976 616140 671028 616146
rect 670976 616082 671028 616088
rect 670792 580032 670844 580038
rect 670792 579974 670844 579980
rect 670792 569628 670844 569634
rect 670792 569570 670844 569576
rect 670606 217968 670662 217977
rect 670606 217903 670662 217912
rect 670608 216980 670660 216986
rect 670608 216922 670660 216928
rect 670620 193361 670648 216922
rect 670804 211177 670832 569570
rect 670988 345001 671016 616082
rect 671172 601694 671200 623902
rect 671356 610162 671384 661098
rect 671724 659654 671752 666590
rect 671816 666554 671844 667791
rect 671816 666526 671936 666554
rect 671540 659626 671752 659654
rect 671540 624306 671568 659626
rect 671712 649120 671764 649126
rect 671712 649062 671764 649068
rect 671528 624300 671580 624306
rect 671528 624242 671580 624248
rect 671724 624186 671752 649062
rect 671448 624158 671752 624186
rect 671448 617250 671476 624158
rect 671908 623914 671936 666526
rect 671632 623886 671936 623914
rect 671632 622878 671660 623886
rect 671620 622872 671672 622878
rect 671620 622814 671672 622820
rect 672000 622690 672028 667950
rect 671908 622662 672028 622690
rect 671712 622600 671764 622606
rect 671712 622542 671764 622548
rect 671724 621014 671752 622542
rect 671908 621246 671936 622662
rect 671896 621240 671948 621246
rect 671896 621182 671948 621188
rect 671540 620986 671752 621014
rect 671896 621036 671948 621042
rect 671540 618202 671568 620986
rect 671896 620978 671948 620984
rect 671540 618174 671752 618202
rect 671448 617222 671660 617250
rect 671632 616706 671660 617222
rect 671540 616690 671660 616706
rect 671528 616684 671660 616690
rect 671580 616678 671660 616684
rect 671528 616626 671580 616632
rect 671724 616554 671752 618174
rect 671908 616865 671936 620978
rect 671894 616856 671950 616865
rect 671894 616791 671950 616800
rect 671896 616684 671948 616690
rect 671896 616626 671948 616632
rect 671712 616548 671764 616554
rect 671712 616490 671764 616496
rect 671712 616412 671764 616418
rect 671712 616354 671764 616360
rect 671344 610156 671396 610162
rect 671344 610098 671396 610104
rect 671526 608696 671582 608705
rect 671526 608631 671582 608640
rect 671172 601666 671384 601694
rect 671160 579420 671212 579426
rect 671160 579362 671212 579368
rect 671172 565078 671200 579362
rect 671356 579086 671384 601666
rect 671344 579080 671396 579086
rect 671344 579022 671396 579028
rect 671540 578898 671568 608631
rect 671724 608594 671752 616354
rect 671356 578870 671568 578898
rect 671632 608566 671752 608594
rect 671356 577454 671384 578870
rect 671632 578066 671660 608566
rect 671908 601694 671936 616626
rect 671816 601666 671936 601694
rect 671620 578060 671672 578066
rect 671620 578002 671672 578008
rect 671528 577788 671580 577794
rect 671528 577730 671580 577736
rect 671344 577448 671396 577454
rect 671344 577390 671396 577396
rect 671344 576972 671396 576978
rect 671344 576914 671396 576920
rect 671356 572714 671384 576914
rect 671356 572686 671476 572714
rect 671448 569954 671476 572686
rect 671356 569926 671476 569954
rect 671356 565282 671384 569926
rect 671344 565276 671396 565282
rect 671344 565218 671396 565224
rect 671160 565072 671212 565078
rect 671160 565014 671212 565020
rect 671160 564936 671212 564942
rect 671160 564878 671212 564884
rect 671172 560368 671200 564878
rect 671344 564800 671396 564806
rect 671396 564748 671476 564754
rect 671344 564742 671476 564748
rect 671356 564726 671476 564742
rect 671172 560340 671292 560368
rect 671264 538214 671292 560340
rect 671448 560294 671476 564726
rect 671172 538186 671292 538214
rect 671356 560266 671476 560294
rect 671172 531486 671200 538186
rect 671356 534410 671384 560266
rect 671344 534404 671396 534410
rect 671344 534346 671396 534352
rect 671540 532914 671568 577730
rect 671816 573782 671844 601666
rect 671804 573776 671856 573782
rect 671804 573718 671856 573724
rect 671712 570852 671764 570858
rect 671712 570794 671764 570800
rect 671528 532908 671580 532914
rect 671528 532850 671580 532856
rect 671160 531480 671212 531486
rect 671160 531422 671212 531428
rect 671252 524476 671304 524482
rect 671252 524418 671304 524424
rect 670974 344992 671030 345001
rect 670974 344927 671030 344936
rect 670974 278760 671030 278769
rect 670974 278695 671030 278704
rect 670988 216617 671016 278695
rect 670974 216608 671030 216617
rect 670974 216543 671030 216552
rect 670976 212084 671028 212090
rect 670976 212026 671028 212032
rect 670790 211168 670846 211177
rect 670790 211103 670846 211112
rect 670790 210896 670846 210905
rect 670790 210831 670846 210840
rect 670804 201521 670832 210831
rect 670790 201512 670846 201521
rect 670790 201447 670846 201456
rect 670606 193352 670662 193361
rect 670606 193287 670662 193296
rect 670988 183530 671016 212026
rect 670976 183524 671028 183530
rect 670976 183466 671028 183472
rect 670608 170332 670660 170338
rect 670608 170274 670660 170280
rect 670332 164960 670384 164966
rect 670332 164902 670384 164908
rect 670620 147626 670648 170274
rect 670976 166932 671028 166938
rect 670976 166874 671028 166880
rect 670608 147620 670660 147626
rect 670608 147562 670660 147568
rect 670148 121508 670200 121514
rect 670148 121450 670200 121456
rect 669964 117836 670016 117842
rect 669964 117778 670016 117784
rect 668780 113146 668900 113174
rect 668964 113146 669084 113174
rect 668872 111738 668900 113146
rect 668872 111710 668992 111738
rect 668768 111648 668820 111654
rect 668768 111590 668820 111596
rect 668780 111081 668808 111590
rect 668766 111072 668822 111081
rect 668766 111007 668822 111016
rect 668964 106049 668992 111710
rect 669056 106162 669084 113146
rect 670160 112946 670188 121450
rect 670988 115870 671016 166874
rect 671264 150278 671292 524418
rect 671436 480684 671488 480690
rect 671436 480626 671488 480632
rect 671252 150272 671304 150278
rect 671252 150214 671304 150220
rect 671448 145586 671476 480626
rect 671724 474094 671752 570794
rect 671896 553512 671948 553518
rect 671896 553454 671948 553460
rect 671908 482390 671936 553454
rect 671896 482384 671948 482390
rect 671896 482326 671948 482332
rect 671712 474088 671764 474094
rect 671712 474030 671764 474036
rect 671804 396364 671856 396370
rect 671804 396306 671856 396312
rect 671620 392012 671672 392018
rect 671620 391954 671672 391960
rect 671632 350534 671660 391954
rect 671816 382362 671844 396306
rect 671804 382356 671856 382362
rect 671804 382298 671856 382304
rect 671896 351960 671948 351966
rect 671896 351902 671948 351908
rect 671908 350690 671936 351902
rect 671908 350662 672028 350690
rect 671804 350600 671856 350606
rect 671804 350542 671856 350548
rect 671540 350506 671660 350534
rect 671540 340874 671568 350506
rect 671816 347774 671844 350542
rect 671816 347746 671936 347774
rect 671908 346394 671936 347746
rect 671816 346366 671936 346394
rect 671816 345273 671844 346366
rect 671802 345264 671858 345273
rect 671802 345199 671858 345208
rect 671712 345024 671764 345030
rect 671712 344966 671764 344972
rect 671540 340846 671660 340874
rect 671632 211154 671660 340846
rect 671724 211290 671752 344966
rect 672000 341578 672028 350662
rect 671908 341550 672028 341578
rect 671908 333946 671936 341550
rect 671896 333940 671948 333946
rect 671896 333882 671948 333888
rect 671896 259684 671948 259690
rect 671896 259626 671948 259632
rect 671908 245721 671936 259626
rect 671894 245712 671950 245721
rect 671894 245647 671950 245656
rect 671896 219496 671948 219502
rect 671816 219444 671896 219450
rect 671816 219438 671948 219444
rect 671816 219406 671936 219438
rect 671908 216209 671936 219406
rect 671894 216200 671950 216209
rect 671894 216135 671950 216144
rect 672092 216050 672120 678946
rect 672368 538214 672396 688606
rect 672632 687268 672684 687274
rect 672632 687210 672684 687216
rect 672644 618254 672672 687210
rect 672828 673454 672856 730079
rect 673012 717614 673040 738414
rect 673196 717614 673224 750706
rect 672736 673426 672856 673454
rect 672920 717586 673040 717614
rect 673104 717586 673224 717614
rect 673288 750706 673408 750734
rect 673932 750706 674052 750734
rect 674116 760366 674236 760394
rect 674116 750734 674144 760366
rect 674116 750706 674236 750734
rect 672736 663898 672764 673426
rect 672920 664086 672948 717586
rect 673104 710054 673132 717586
rect 673092 710048 673144 710054
rect 673092 709990 673144 709996
rect 673092 697128 673144 697134
rect 673092 697070 673144 697076
rect 672908 664080 672960 664086
rect 672908 664022 672960 664028
rect 672736 663870 672948 663898
rect 672920 663513 672948 663870
rect 672906 663504 672962 663513
rect 672906 663439 672962 663448
rect 672908 651432 672960 651438
rect 672908 651374 672960 651380
rect 672632 618248 672684 618254
rect 672632 618190 672684 618196
rect 672540 605872 672592 605878
rect 672540 605814 672592 605820
rect 672552 538214 672580 605814
rect 672724 578604 672776 578610
rect 672724 578546 672776 578552
rect 672736 563054 672764 578546
rect 672920 578270 672948 651374
rect 673104 619478 673132 697070
rect 673092 619472 673144 619478
rect 673092 619414 673144 619420
rect 673092 607640 673144 607646
rect 673092 607582 673144 607588
rect 672908 578264 672960 578270
rect 672908 578206 672960 578212
rect 672276 538186 672396 538214
rect 672460 538186 672580 538214
rect 672644 563026 672764 563054
rect 672276 528554 672304 538186
rect 672460 531622 672488 538186
rect 672644 534614 672672 563026
rect 672814 554024 672870 554033
rect 672814 553959 672870 553968
rect 672632 534608 672684 534614
rect 672632 534550 672684 534556
rect 672632 534132 672684 534138
rect 672632 534074 672684 534080
rect 672448 531616 672500 531622
rect 672448 531558 672500 531564
rect 672644 531434 672672 534074
rect 672644 531406 672764 531434
rect 672540 531344 672592 531350
rect 672540 531286 672592 531292
rect 672276 528526 672396 528554
rect 672368 297770 672396 528526
rect 672552 487354 672580 531286
rect 672736 490074 672764 531406
rect 672828 505094 672856 553959
rect 673104 530126 673132 607582
rect 673092 530120 673144 530126
rect 673092 530062 673144 530068
rect 672828 505066 672948 505094
rect 672724 490068 672776 490074
rect 672724 490010 672776 490016
rect 672540 487348 672592 487354
rect 672540 487290 672592 487296
rect 672920 483614 672948 505066
rect 672908 483608 672960 483614
rect 672908 483550 672960 483556
rect 672724 400580 672776 400586
rect 672724 400522 672776 400528
rect 672540 396092 672592 396098
rect 672540 396034 672592 396040
rect 672552 378049 672580 396034
rect 672538 378040 672594 378049
rect 672538 377975 672594 377984
rect 672736 355230 672764 400522
rect 673092 399764 673144 399770
rect 673092 399706 673144 399712
rect 672908 393372 672960 393378
rect 672908 393314 672960 393320
rect 672920 376514 672948 393314
rect 672908 376508 672960 376514
rect 672908 376450 672960 376456
rect 672724 355224 672776 355230
rect 672724 355166 672776 355172
rect 673104 354890 673132 399706
rect 673288 394641 673316 750706
rect 673736 748876 673788 748882
rect 673736 748818 673788 748824
rect 673748 741074 673776 748818
rect 673932 748746 673960 750706
rect 674208 748898 674236 750706
rect 674116 748882 674236 748898
rect 674104 748876 674236 748882
rect 674156 748870 674236 748876
rect 674104 748818 674156 748824
rect 673920 748740 673972 748746
rect 673920 748682 673972 748688
rect 674104 748400 674156 748406
rect 674104 748342 674156 748348
rect 674116 741074 674144 748342
rect 673748 741046 673960 741074
rect 674116 741046 674236 741074
rect 673458 734904 673514 734913
rect 673458 734839 673514 734848
rect 673472 682825 673500 734839
rect 673932 734174 673960 741046
rect 673932 734146 674144 734174
rect 673826 732728 673882 732737
rect 673826 732663 673882 732672
rect 673642 725928 673698 725937
rect 673642 725863 673698 725872
rect 673656 683097 673684 725863
rect 673642 683088 673698 683097
rect 673642 683023 673698 683032
rect 673458 682816 673514 682825
rect 673458 682751 673514 682760
rect 673840 663270 673868 732663
rect 674116 732034 674144 734146
rect 673932 732006 674144 732034
rect 673932 727274 673960 732006
rect 673932 727246 674144 727274
rect 674116 707606 674144 727246
rect 674208 726730 674236 741046
rect 674300 730266 674328 779146
rect 674484 775574 674512 783838
rect 674668 775574 674696 869774
rect 674838 869680 674894 869689
rect 674838 869615 674894 869624
rect 674852 865434 674880 869615
rect 675036 869530 675064 869774
rect 675680 869689 675708 870060
rect 675666 869680 675722 869689
rect 675666 869615 675722 869624
rect 675036 869502 675418 869530
rect 675024 869032 675076 869038
rect 674944 868980 675024 868986
rect 674944 868974 675076 868980
rect 674944 868958 675064 868974
rect 674944 866266 674972 868958
rect 675128 868861 675418 868889
rect 675128 868086 675156 868861
rect 675116 868080 675168 868086
rect 675496 868057 675524 868224
rect 675116 868022 675168 868028
rect 675482 868048 675538 868057
rect 675482 867983 675538 867992
rect 675128 867021 675418 867049
rect 675128 866726 675156 867021
rect 675116 866720 675168 866726
rect 675116 866662 675168 866668
rect 674944 866238 675432 866266
rect 675404 865844 675432 866238
rect 674840 865428 674892 865434
rect 674840 865370 674892 865376
rect 674840 865292 674892 865298
rect 674840 865234 674892 865240
rect 674852 863841 674880 865234
rect 675220 865181 675418 865209
rect 675220 865178 675248 865181
rect 675128 865150 675248 865178
rect 674838 863832 674894 863841
rect 674838 863767 674894 863776
rect 675128 859754 675156 865150
rect 675300 865088 675352 865094
rect 675300 865030 675352 865036
rect 675036 859726 675156 859754
rect 675036 856994 675064 859726
rect 675036 856966 675156 856994
rect 674932 789404 674984 789410
rect 674932 789346 674984 789352
rect 674944 788730 674972 789346
rect 674932 788724 674984 788730
rect 674932 788666 674984 788672
rect 675128 788610 675156 856966
rect 675312 789374 675340 865030
rect 675496 864249 675524 864552
rect 675482 864240 675538 864249
rect 675482 864175 675538 864184
rect 675482 863832 675538 863841
rect 675482 863767 675538 863776
rect 675496 863328 675524 863767
rect 674852 788582 675156 788610
rect 675220 789346 675340 789374
rect 674852 782474 674880 788582
rect 675220 788474 675248 789346
rect 674760 782446 674880 782474
rect 674944 788446 675248 788474
rect 674760 776506 674788 782446
rect 674944 780337 674972 788446
rect 675128 788310 675418 788338
rect 675128 788050 675156 788310
rect 675300 788248 675352 788254
rect 675300 788190 675352 788196
rect 675116 788044 675168 788050
rect 675116 787986 675168 787992
rect 675312 787693 675340 788190
rect 675312 787665 675418 787693
rect 675128 787018 675418 787046
rect 675128 786690 675156 787018
rect 675116 786684 675168 786690
rect 675116 786626 675168 786632
rect 675220 785182 675418 785210
rect 675220 783902 675248 785182
rect 675404 784281 675432 784652
rect 675390 784272 675446 784281
rect 675390 784207 675446 784216
rect 675208 783896 675260 783902
rect 675496 783850 675524 783972
rect 675208 783838 675260 783844
rect 675404 783822 675524 783850
rect 675404 783766 675432 783822
rect 675392 783760 675444 783766
rect 675392 783702 675444 783708
rect 675220 783346 675418 783374
rect 675220 782678 675248 783346
rect 675208 782672 675260 782678
rect 675208 782614 675260 782620
rect 675300 782536 675352 782542
rect 675300 782478 675352 782484
rect 675312 781402 675340 782478
rect 675312 781374 675432 781402
rect 675404 780844 675432 781374
rect 674930 780328 674986 780337
rect 674930 780263 674986 780272
rect 675496 779929 675524 780300
rect 675482 779920 675538 779929
rect 675482 779855 675538 779864
rect 675312 779674 675418 779702
rect 675312 779210 675340 779674
rect 675300 779204 675352 779210
rect 675300 779146 675352 779152
rect 675312 779062 675432 779090
rect 675116 779000 675168 779006
rect 675116 778942 675168 778948
rect 675128 776642 675156 778942
rect 675312 778394 675340 779062
rect 675404 779008 675432 779062
rect 675300 778388 675352 778394
rect 675300 778330 675352 778336
rect 675404 777322 675432 777852
rect 675312 777294 675432 777322
rect 675312 777034 675340 777294
rect 675300 777028 675352 777034
rect 675300 776970 675352 776976
rect 675128 776614 675418 776642
rect 674760 776478 675156 776506
rect 674392 775546 674512 775574
rect 674576 775546 674696 775574
rect 674392 730365 674420 775546
rect 674576 772721 674604 775546
rect 674932 775464 674984 775470
rect 674746 775432 674802 775441
rect 674932 775406 674984 775412
rect 674746 775367 674802 775376
rect 674562 772712 674618 772721
rect 674562 772647 674618 772656
rect 674760 756254 674788 775367
rect 674484 756226 674788 756254
rect 674484 732306 674512 756226
rect 674944 751097 674972 775406
rect 675128 771769 675156 776478
rect 675404 775554 675432 776016
rect 675312 775526 675432 775554
rect 675312 775470 675340 775526
rect 675300 775464 675352 775470
rect 675300 775406 675352 775412
rect 675404 775033 675432 775336
rect 675390 775024 675446 775033
rect 675390 774959 675446 774968
rect 675404 773673 675432 774180
rect 675390 773664 675446 773673
rect 675390 773599 675446 773608
rect 675390 773392 675446 773401
rect 675390 773327 675446 773336
rect 675114 771760 675170 771769
rect 675114 771695 675170 771704
rect 675404 765914 675432 773327
rect 675850 772712 675906 772721
rect 675850 772647 675906 772656
rect 679622 772712 679678 772721
rect 679622 772647 679678 772656
rect 675864 772138 675892 772647
rect 675852 772132 675904 772138
rect 675852 772074 675904 772080
rect 675850 771760 675906 771769
rect 675850 771695 675906 771704
rect 675864 771322 675892 771695
rect 675852 771316 675904 771322
rect 675852 771258 675904 771264
rect 675404 765886 675892 765914
rect 675484 761592 675536 761598
rect 675482 761560 675484 761569
rect 675536 761560 675538 761569
rect 675482 761495 675538 761504
rect 675298 761152 675354 761161
rect 675298 761087 675354 761096
rect 675312 760442 675340 761087
rect 675482 760744 675538 760753
rect 675482 760679 675538 760688
rect 675496 760578 675524 760679
rect 675484 760572 675536 760578
rect 675484 760514 675536 760520
rect 675300 760436 675352 760442
rect 675300 760378 675352 760384
rect 675482 760336 675538 760345
rect 675482 760271 675484 760280
rect 675536 760271 675538 760280
rect 675484 760242 675536 760248
rect 675482 759928 675538 759937
rect 675482 759863 675484 759872
rect 675536 759863 675538 759872
rect 675484 759834 675536 759840
rect 675484 759552 675536 759558
rect 675482 759520 675484 759529
rect 675536 759520 675538 759529
rect 675482 759455 675538 759464
rect 675482 759112 675538 759121
rect 675482 759047 675484 759056
rect 675536 759047 675538 759056
rect 675484 759018 675536 759024
rect 675484 758736 675536 758742
rect 675482 758704 675484 758713
rect 675536 758704 675538 758713
rect 675482 758639 675538 758648
rect 675300 758396 675352 758402
rect 675300 758338 675352 758344
rect 675312 757897 675340 758338
rect 675482 758296 675538 758305
rect 675482 758231 675484 758240
rect 675536 758231 675538 758240
rect 675484 758202 675536 758208
rect 675298 757888 675354 757897
rect 675298 757823 675354 757832
rect 675482 757480 675538 757489
rect 675482 757415 675484 757424
rect 675536 757415 675538 757424
rect 675484 757386 675536 757392
rect 675864 755857 675892 765886
rect 676954 761832 677010 761841
rect 676954 761767 677010 761776
rect 676968 757081 676996 761767
rect 676954 757072 677010 757081
rect 676954 757007 677010 757016
rect 679636 756265 679664 772647
rect 683394 772440 683450 772449
rect 683394 772375 683450 772384
rect 683212 772132 683264 772138
rect 683212 772074 683264 772080
rect 682382 771352 682438 771361
rect 681004 771316 681056 771322
rect 682382 771287 682438 771296
rect 681004 771258 681056 771264
rect 681016 756673 681044 771258
rect 681002 756664 681058 756673
rect 681002 756599 681058 756608
rect 679622 756256 679678 756265
rect 679622 756191 679678 756200
rect 675850 755848 675906 755857
rect 675850 755783 675906 755792
rect 682396 755449 682424 771287
rect 682382 755440 682438 755449
rect 682382 755375 682438 755384
rect 675484 755064 675536 755070
rect 675482 755032 675484 755041
rect 675536 755032 675538 755041
rect 675482 754967 675538 754976
rect 675484 754656 675536 754662
rect 675482 754624 675484 754633
rect 675536 754624 675538 754633
rect 675482 754559 675538 754568
rect 675484 753432 675536 753438
rect 675482 753400 675484 753409
rect 675536 753400 675538 753409
rect 675482 753335 675538 753344
rect 675484 753024 675536 753030
rect 675482 752992 675484 753001
rect 675536 752992 675538 753001
rect 675482 752927 675538 752936
rect 675850 752312 675906 752321
rect 675850 752247 675906 752256
rect 675484 751800 675536 751806
rect 675482 751768 675484 751777
rect 675536 751768 675538 751777
rect 675482 751703 675538 751712
rect 675482 751360 675538 751369
rect 675482 751295 675484 751304
rect 675536 751295 675538 751304
rect 675484 751266 675536 751272
rect 675864 751126 675892 752247
rect 683224 752185 683252 772074
rect 683408 752593 683436 772375
rect 684038 772032 684094 772041
rect 684038 771967 684094 771976
rect 684052 754225 684080 771967
rect 703694 762076 703722 762212
rect 704154 762076 704182 762212
rect 704614 762076 704642 762212
rect 705074 762076 705102 762212
rect 705534 762076 705562 762212
rect 705994 762076 706022 762212
rect 706454 762076 706482 762212
rect 706914 762076 706942 762212
rect 707374 762076 707402 762212
rect 707834 762076 707862 762212
rect 708294 762076 708322 762212
rect 708754 762076 708782 762212
rect 709214 762076 709242 762212
rect 684038 754216 684094 754225
rect 684038 754151 684094 754160
rect 683394 752584 683450 752593
rect 683394 752519 683450 752528
rect 683210 752176 683266 752185
rect 683210 752111 683266 752120
rect 675852 751120 675904 751126
rect 674930 751088 674986 751097
rect 675852 751062 675904 751068
rect 683120 751120 683172 751126
rect 683120 751062 683172 751068
rect 674930 751023 674986 751032
rect 683132 750757 683160 751062
rect 683118 750748 683174 750757
rect 683118 750683 683174 750692
rect 675482 750136 675538 750145
rect 675482 750071 675484 750080
rect 675536 750071 675538 750080
rect 675484 750042 675536 750048
rect 675300 745272 675352 745278
rect 675300 745214 675352 745220
rect 675312 742642 675340 745214
rect 675588 743073 675616 743308
rect 675574 743064 675630 743073
rect 675574 742999 675630 743008
rect 675404 742642 675432 742696
rect 675312 742614 675432 742642
rect 675300 742484 675352 742490
rect 675300 742426 675352 742432
rect 674840 741668 674892 741674
rect 674840 741610 674892 741616
rect 674484 732278 674788 732306
rect 674392 730337 674604 730365
rect 674300 730238 674420 730266
rect 674392 728414 674420 730238
rect 674380 728408 674432 728414
rect 674380 728350 674432 728356
rect 674576 728113 674604 730337
rect 674760 728226 674788 732278
rect 674852 729314 674880 741610
rect 675312 740194 675340 742426
rect 675496 741674 675524 742016
rect 675484 741668 675536 741674
rect 675484 741610 675536 741616
rect 675312 740166 675418 740194
rect 675128 739622 675418 739650
rect 675128 738478 675156 739622
rect 675404 738721 675432 739024
rect 675390 738712 675446 738721
rect 675390 738647 675446 738656
rect 675116 738472 675168 738478
rect 675116 738414 675168 738420
rect 675128 738330 675418 738358
rect 675128 738177 675156 738330
rect 675114 738168 675170 738177
rect 675114 738103 675170 738112
rect 675404 735842 675432 735896
rect 675312 735814 675432 735842
rect 675312 734806 675340 735814
rect 675496 734913 675524 735319
rect 675482 734904 675538 734913
rect 675482 734839 675538 734848
rect 675300 734800 675352 734806
rect 675300 734742 675352 734748
rect 675024 734732 675076 734738
rect 675024 734674 675076 734680
rect 675036 731626 675064 734674
rect 675300 734596 675352 734602
rect 675300 734538 675352 734544
rect 675312 733689 675340 734538
rect 675496 734505 675524 734672
rect 675482 734496 675538 734505
rect 675482 734431 675538 734440
rect 675482 734224 675538 734233
rect 675482 734159 675538 734168
rect 675496 734031 675524 734159
rect 675298 733680 675354 733689
rect 675298 733615 675354 733624
rect 675404 732737 675432 732836
rect 675390 732728 675446 732737
rect 675390 732663 675446 732672
rect 675312 731734 675432 731762
rect 675312 731626 675340 731734
rect 675036 731598 675340 731626
rect 675404 731612 675432 731734
rect 675220 730986 675418 731014
rect 674852 729286 675064 729314
rect 675036 728906 675064 729286
rect 675220 729026 675248 730986
rect 675404 730153 675432 730351
rect 675390 730144 675446 730153
rect 675390 730079 675446 730088
rect 675208 729020 675260 729026
rect 675208 728962 675260 728968
rect 675036 728878 675248 728906
rect 675024 728816 675076 728822
rect 675024 728758 675076 728764
rect 674760 728198 674880 728226
rect 674562 728104 674618 728113
rect 674562 728039 674618 728048
rect 674208 726702 674328 726730
rect 674300 723217 674328 726702
rect 674852 724514 674880 728198
rect 674484 724486 674880 724514
rect 674286 723208 674342 723217
rect 674286 723143 674342 723152
rect 674104 707600 674156 707606
rect 674104 707542 674156 707548
rect 674484 707169 674512 724486
rect 674840 715352 674892 715358
rect 674838 715320 674840 715329
rect 674892 715320 674894 715329
rect 674838 715255 674894 715264
rect 674470 707160 674526 707169
rect 674470 707095 674526 707104
rect 675036 698294 675064 728758
rect 675220 721585 675248 728878
rect 675404 728793 675432 729164
rect 675390 728784 675446 728793
rect 675390 728719 675446 728728
rect 675484 728408 675536 728414
rect 675484 728350 675536 728356
rect 675496 728090 675524 728350
rect 676034 728104 676090 728113
rect 675496 728062 675892 728090
rect 675864 726578 675892 728062
rect 676034 728039 676090 728048
rect 676048 726850 676076 728039
rect 676036 726844 676088 726850
rect 676036 726786 676088 726792
rect 683120 726844 683172 726850
rect 683120 726786 683172 726792
rect 675852 726572 675904 726578
rect 675852 726514 675904 726520
rect 675850 723208 675906 723217
rect 675850 723143 675906 723152
rect 675206 721576 675262 721585
rect 675206 721511 675262 721520
rect 675864 719710 675892 723143
rect 675852 719704 675904 719710
rect 675852 719646 675904 719652
rect 675482 716544 675538 716553
rect 675482 716479 675538 716488
rect 675496 716310 675524 716479
rect 675484 716304 675536 716310
rect 675484 716246 675536 716252
rect 675298 716136 675354 716145
rect 675298 716071 675354 716080
rect 675312 714882 675340 716071
rect 675482 715728 675538 715737
rect 675482 715663 675538 715672
rect 675496 715154 675524 715663
rect 675484 715148 675536 715154
rect 675484 715090 675536 715096
rect 675482 714912 675538 714921
rect 675300 714876 675352 714882
rect 675482 714847 675484 714856
rect 675300 714818 675352 714824
rect 675536 714847 675538 714856
rect 675484 714818 675536 714824
rect 675484 714536 675536 714542
rect 675482 714504 675484 714513
rect 675536 714504 675538 714513
rect 675482 714439 675538 714448
rect 675482 714096 675538 714105
rect 675482 714031 675484 714040
rect 675536 714031 675538 714040
rect 675484 714002 675536 714008
rect 675484 713720 675536 713726
rect 675482 713688 675484 713697
rect 675536 713688 675538 713697
rect 675482 713623 675538 713632
rect 677690 713488 677746 713497
rect 676036 713448 676088 713454
rect 677690 713423 677692 713432
rect 676036 713390 676088 713396
rect 677744 713423 677746 713432
rect 677692 713390 677744 713396
rect 675482 713280 675538 713289
rect 675482 713215 675484 713224
rect 675536 713215 675538 713224
rect 675484 713186 675536 713192
rect 675484 712904 675536 712910
rect 675482 712872 675484 712881
rect 675536 712872 675538 712881
rect 675482 712807 675538 712816
rect 675482 712464 675538 712473
rect 675482 712399 675484 712408
rect 675536 712399 675538 712408
rect 675484 712370 675536 712376
rect 675484 712088 675536 712094
rect 675482 712056 675484 712065
rect 675536 712056 675538 712065
rect 675482 711991 675538 712000
rect 676048 711657 676076 713390
rect 676034 711648 676090 711657
rect 676034 711583 676090 711592
rect 675484 711272 675536 711278
rect 675482 711240 675484 711249
rect 675536 711240 675538 711249
rect 675482 711175 675538 711184
rect 683132 710841 683160 726786
rect 683488 726572 683540 726578
rect 683488 726514 683540 726520
rect 683304 719704 683356 719710
rect 683304 719646 683356 719652
rect 683118 710832 683174 710841
rect 683118 710767 683174 710776
rect 675850 710696 675906 710705
rect 675850 710631 675906 710640
rect 675482 710424 675538 710433
rect 675482 710359 675538 710368
rect 675300 710048 675352 710054
rect 675298 710016 675300 710025
rect 675352 710016 675354 710025
rect 675298 709951 675354 709960
rect 675496 709782 675524 710359
rect 675484 709776 675536 709782
rect 675484 709718 675536 709724
rect 675484 709640 675536 709646
rect 675482 709608 675484 709617
rect 675536 709608 675538 709617
rect 675482 709543 675538 709552
rect 675484 708824 675536 708830
rect 675482 708792 675484 708801
rect 675536 708792 675538 708801
rect 675482 708727 675538 708736
rect 675484 708416 675536 708422
rect 675482 708384 675484 708393
rect 675536 708384 675538 708393
rect 675482 708319 675538 708328
rect 675484 707600 675536 707606
rect 675482 707568 675484 707577
rect 675536 707568 675538 707577
rect 675482 707503 675538 707512
rect 675482 706344 675538 706353
rect 675482 706279 675484 706288
rect 675536 706279 675538 706288
rect 675484 706250 675536 706256
rect 675864 705362 675892 710631
rect 683316 706761 683344 719646
rect 683500 707985 683528 726514
rect 703694 717196 703722 717264
rect 704154 717196 704182 717264
rect 704614 717196 704642 717264
rect 705074 717196 705102 717264
rect 705534 717196 705562 717264
rect 705994 717196 706022 717264
rect 706454 717196 706482 717264
rect 706914 717196 706942 717264
rect 707374 717196 707402 717264
rect 707834 717196 707862 717264
rect 708294 717196 708322 717264
rect 708754 717196 708782 717264
rect 709214 717196 709242 717264
rect 683486 707976 683542 707985
rect 683486 707911 683542 707920
rect 683302 706752 683358 706761
rect 683302 706687 683358 706696
rect 683118 705528 683174 705537
rect 683118 705463 683174 705472
rect 683132 705362 683160 705463
rect 675852 705356 675904 705362
rect 675852 705298 675904 705304
rect 683120 705356 683172 705362
rect 683120 705298 683172 705304
rect 675482 705120 675538 705129
rect 675482 705055 675484 705064
rect 675536 705055 675538 705064
rect 675484 705026 675536 705032
rect 675208 698488 675260 698494
rect 675208 698430 675260 698436
rect 675220 698337 675248 698430
rect 675220 698309 675418 698337
rect 674944 698266 675064 698294
rect 674288 694816 674340 694822
rect 674288 694758 674340 694764
rect 674104 689172 674156 689178
rect 674104 689114 674156 689120
rect 674116 688634 674144 689114
rect 674116 688606 674236 688634
rect 674012 670404 674064 670410
rect 674012 670346 674064 670352
rect 674024 669526 674052 670346
rect 674012 669520 674064 669526
rect 674012 669462 674064 669468
rect 674010 668944 674066 668953
rect 674010 668879 674066 668888
rect 674024 667622 674052 668879
rect 674012 667616 674064 667622
rect 674012 667558 674064 667564
rect 673828 663264 673880 663270
rect 673828 663206 673880 663212
rect 674010 644736 674066 644745
rect 674010 644671 674066 644680
rect 674024 644489 674052 644671
rect 674024 644461 674144 644489
rect 673734 644328 673790 644337
rect 673734 644263 673790 644272
rect 673460 639056 673512 639062
rect 673380 639004 673460 639010
rect 673380 638998 673512 639004
rect 673380 638982 673500 638998
rect 673380 576994 673408 638982
rect 673550 599856 673606 599865
rect 673550 599791 673606 599800
rect 673564 577266 673592 599791
rect 673748 577590 673776 644263
rect 673918 643512 673974 643521
rect 673918 643447 673974 643456
rect 673932 640334 673960 643447
rect 673932 640306 674052 640334
rect 674024 611354 674052 640306
rect 673840 611326 674052 611354
rect 673840 592034 673868 611326
rect 674116 608594 674144 644461
rect 674208 630674 674236 688606
rect 674300 645854 674328 694758
rect 674472 694204 674524 694210
rect 674472 694146 674524 694152
rect 674484 645854 674512 694146
rect 674944 694113 674972 698266
rect 675128 697666 675418 697694
rect 675128 697134 675156 697666
rect 675116 697128 675168 697134
rect 675116 697070 675168 697076
rect 675404 696833 675432 697035
rect 675390 696824 675446 696833
rect 675390 696759 675446 696768
rect 675128 695181 675418 695209
rect 675128 694822 675156 695181
rect 675116 694816 675168 694822
rect 675116 694758 675168 694764
rect 675312 694742 675432 694770
rect 675114 694648 675170 694657
rect 675312 694634 675340 694742
rect 675170 694606 675340 694634
rect 675404 694620 675432 694742
rect 675114 694583 675170 694592
rect 675392 694204 675444 694210
rect 675392 694146 675444 694152
rect 674930 694104 674986 694113
rect 674930 694039 674986 694048
rect 675404 694008 675432 694146
rect 675312 693382 675432 693410
rect 675312 693342 675340 693382
rect 675128 693314 675340 693342
rect 675404 693328 675432 693382
rect 675128 693025 675156 693314
rect 675114 693016 675170 693025
rect 675114 692951 675170 692960
rect 675116 692844 675168 692850
rect 675116 692786 675168 692792
rect 675128 690894 675156 692786
rect 675128 690866 675418 690894
rect 674668 690322 675340 690350
rect 674300 645826 674420 645854
rect 674484 645826 674604 645854
rect 674392 636954 674420 645826
rect 674380 636948 674432 636954
rect 674380 636890 674432 636896
rect 674576 636194 674604 645826
rect 674484 636166 674604 636194
rect 674208 630646 674328 630674
rect 674300 617817 674328 630646
rect 674484 618633 674512 636166
rect 674470 618624 674526 618633
rect 674470 618559 674526 618568
rect 674286 617808 674342 617817
rect 674286 617743 674342 617752
rect 674668 617001 674696 690322
rect 675312 690282 675340 690322
rect 675404 690282 675432 690336
rect 675312 690254 675432 690282
rect 675312 689710 675432 689738
rect 675312 689670 675340 689710
rect 675128 689642 675340 689670
rect 675404 689656 675432 689710
rect 674932 689308 674984 689314
rect 674932 689250 674984 689256
rect 674944 686678 674972 689250
rect 675128 689178 675156 689642
rect 675116 689172 675168 689178
rect 675116 689114 675168 689120
rect 675128 689030 675418 689058
rect 675128 688673 675156 689030
rect 675114 688664 675170 688673
rect 675114 688599 675170 688608
rect 675128 687806 675418 687834
rect 675128 687274 675156 687806
rect 675116 687268 675168 687274
rect 675116 687210 675168 687216
rect 674944 686650 675340 686678
rect 675312 686610 675340 686650
rect 675404 686610 675432 686664
rect 675312 686582 675432 686610
rect 675036 685970 675418 685998
rect 674840 685908 674892 685914
rect 674840 685850 674892 685856
rect 674852 684321 674880 685850
rect 674838 684312 674894 684321
rect 674838 684247 674894 684256
rect 674838 669760 674894 669769
rect 674838 669695 674894 669704
rect 674852 669390 674880 669695
rect 674840 669384 674892 669390
rect 674840 669326 674892 669332
rect 674840 664080 674892 664086
rect 674838 664048 674840 664057
rect 674892 664048 674894 664057
rect 674838 663983 674894 663992
rect 674840 650072 674892 650078
rect 674840 650014 674892 650020
rect 674852 648650 674880 650014
rect 674840 648644 674892 648650
rect 674840 648586 674892 648592
rect 675036 647234 675064 685970
rect 675298 685672 675354 685681
rect 675298 685607 675354 685616
rect 675312 676214 675340 685607
rect 675496 685137 675524 685372
rect 675482 685128 675538 685137
rect 675482 685063 675538 685072
rect 675482 684312 675538 684321
rect 675482 684247 675538 684256
rect 675496 684148 675524 684247
rect 675850 683088 675906 683097
rect 675850 683023 675906 683032
rect 675864 682446 675892 683023
rect 676034 682816 676090 682825
rect 676034 682751 676090 682760
rect 675852 682440 675904 682446
rect 675852 682382 675904 682388
rect 676048 682310 676076 682751
rect 683212 682440 683264 682446
rect 683212 682382 683264 682388
rect 676036 682304 676088 682310
rect 676036 682246 676088 682252
rect 681002 681864 681058 681873
rect 681002 681799 681058 681808
rect 675220 676186 675340 676214
rect 675220 650185 675248 676186
rect 675482 671392 675538 671401
rect 675482 671327 675538 671336
rect 675496 671158 675524 671327
rect 675484 671152 675536 671158
rect 675484 671094 675536 671100
rect 675482 670984 675538 670993
rect 675482 670919 675538 670928
rect 675496 670750 675524 670919
rect 675484 670744 675536 670750
rect 675484 670686 675536 670692
rect 675482 670576 675538 670585
rect 675482 670511 675538 670520
rect 675496 670410 675524 670511
rect 675484 670404 675536 670410
rect 675484 670346 675536 670352
rect 675482 670168 675538 670177
rect 675482 670103 675538 670112
rect 675496 669798 675524 670103
rect 675484 669792 675536 669798
rect 675484 669734 675536 669740
rect 675484 669656 675536 669662
rect 675484 669598 675536 669604
rect 675496 669361 675524 669598
rect 675482 669352 675538 669361
rect 675482 669287 675538 669296
rect 675484 668568 675536 668574
rect 675482 668536 675484 668545
rect 675536 668536 675538 668545
rect 675482 668471 675538 668480
rect 675484 667752 675536 667758
rect 675482 667720 675484 667729
rect 675536 667720 675538 667729
rect 675482 667655 675538 667664
rect 675482 667312 675538 667321
rect 675482 667247 675484 667256
rect 675536 667247 675538 667256
rect 675484 667218 675536 667224
rect 681016 667049 681044 681799
rect 681002 667040 681058 667049
rect 681002 666975 681058 666984
rect 675484 666120 675536 666126
rect 675482 666088 675484 666097
rect 675536 666088 675538 666097
rect 675482 666023 675538 666032
rect 675482 665680 675538 665689
rect 675482 665615 675538 665624
rect 675496 665242 675524 665615
rect 675484 665236 675536 665242
rect 675484 665178 675536 665184
rect 675666 664864 675722 664873
rect 675666 664799 675722 664808
rect 675482 664456 675538 664465
rect 675482 664391 675538 664400
rect 675496 663950 675524 664391
rect 675484 663944 675536 663950
rect 675484 663886 675536 663892
rect 675484 663808 675536 663814
rect 675680 663762 675708 664799
rect 675536 663756 675708 663762
rect 675484 663750 675708 663756
rect 675496 663734 675708 663750
rect 675850 663504 675906 663513
rect 675850 663439 675906 663448
rect 675484 663264 675536 663270
rect 675482 663232 675484 663241
rect 675536 663232 675538 663241
rect 675482 663167 675538 663176
rect 675484 662856 675536 662862
rect 675482 662824 675484 662833
rect 675536 662824 675538 662833
rect 675482 662759 675538 662768
rect 675484 661632 675536 661638
rect 675482 661600 675484 661609
rect 675536 661600 675538 661609
rect 675482 661535 675538 661544
rect 675482 661192 675538 661201
rect 675482 661127 675484 661136
rect 675536 661127 675538 661136
rect 675484 661098 675536 661104
rect 675482 659968 675538 659977
rect 675482 659903 675484 659912
rect 675536 659903 675538 659912
rect 675484 659874 675536 659880
rect 675864 659870 675892 663439
rect 683224 662561 683252 682382
rect 683396 682304 683448 682310
rect 683396 682246 683448 682252
rect 683210 662552 683266 662561
rect 683210 662487 683266 662496
rect 683408 662153 683436 682246
rect 684038 674112 684094 674121
rect 684038 674047 684094 674056
rect 684052 663785 684080 674047
rect 703694 671908 703722 672044
rect 704154 671908 704182 672044
rect 704614 671908 704642 672044
rect 705074 671908 705102 672044
rect 705534 671908 705562 672044
rect 705994 671908 706022 672044
rect 706454 671908 706482 672044
rect 706914 671908 706942 672044
rect 707374 671908 707402 672044
rect 707834 671908 707862 672044
rect 708294 671908 708322 672044
rect 708754 671908 708782 672044
rect 709214 671908 709242 672044
rect 684038 663776 684094 663785
rect 684038 663711 684094 663720
rect 683394 662144 683450 662153
rect 683394 662079 683450 662088
rect 683118 660104 683174 660113
rect 683118 660039 683174 660048
rect 683132 659870 683160 660039
rect 675852 659864 675904 659870
rect 675852 659806 675904 659812
rect 683120 659864 683172 659870
rect 683120 659806 683172 659812
rect 675392 654288 675444 654294
rect 675312 654236 675392 654242
rect 675312 654230 675444 654236
rect 675312 654214 675432 654230
rect 675312 653018 675340 654214
rect 675312 652990 675432 653018
rect 675404 652460 675432 652990
rect 675588 652905 675616 653140
rect 675574 652896 675630 652905
rect 675574 652831 675630 652840
rect 675404 651438 675432 651848
rect 675392 651432 675444 651438
rect 675392 651374 675444 651380
rect 675206 650176 675262 650185
rect 675206 650111 675262 650120
rect 675404 649890 675432 650012
rect 674944 647206 675064 647234
rect 675128 649862 675432 649890
rect 674944 643929 674972 647206
rect 674930 643920 674986 643929
rect 674930 643855 674986 643864
rect 675128 642410 675156 649862
rect 675404 649126 675432 649468
rect 675392 649120 675444 649126
rect 675392 649062 675444 649068
rect 675390 648952 675446 648961
rect 675390 648887 675446 648896
rect 675404 648788 675432 648887
rect 675392 648644 675444 648650
rect 675392 648586 675444 648592
rect 675404 648530 675432 648586
rect 675404 648502 675524 648530
rect 675496 648176 675524 648502
rect 675390 648000 675446 648009
rect 674944 642382 675156 642410
rect 675220 647958 675390 647986
rect 674944 642274 674972 642382
rect 674852 642246 674972 642274
rect 674852 631258 674880 642246
rect 675220 642138 675248 647958
rect 675390 647935 675446 647944
rect 675666 647456 675722 647465
rect 675666 647391 675722 647400
rect 675680 647234 675708 647391
rect 675312 647206 675708 647234
rect 675312 645674 675340 647206
rect 675312 645646 675418 645674
rect 675404 644745 675432 645116
rect 675390 644736 675446 644745
rect 675390 644671 675446 644680
rect 675404 644337 675432 644475
rect 675390 644328 675446 644337
rect 675390 644263 675446 644272
rect 675404 643521 675432 643824
rect 675390 643512 675446 643521
rect 675390 643447 675446 643456
rect 675404 642161 675432 642635
rect 675128 642110 675248 642138
rect 675390 642152 675446 642161
rect 675128 638874 675156 642110
rect 675390 642087 675446 642096
rect 675300 641912 675352 641918
rect 675300 641854 675352 641860
rect 675312 641458 675340 641854
rect 675312 641430 675418 641458
rect 675680 640393 675708 640795
rect 675666 640384 675722 640393
rect 675666 640319 675722 640328
rect 675312 640138 675418 640166
rect 675312 640082 675340 640138
rect 675300 640076 675352 640082
rect 675300 640018 675352 640024
rect 675300 639056 675352 639062
rect 675352 639004 675432 639010
rect 675300 638998 675432 639004
rect 675312 638982 675432 638998
rect 675404 638928 675432 638982
rect 675128 638846 675340 638874
rect 675312 637945 675340 638846
rect 675482 638208 675538 638217
rect 675482 638143 675538 638152
rect 675298 637936 675354 637945
rect 675298 637871 675354 637880
rect 675206 637664 675262 637673
rect 675206 637599 675262 637608
rect 675220 631417 675248 637599
rect 675496 637378 675524 638143
rect 675850 637936 675906 637945
rect 675850 637871 675906 637880
rect 675864 637498 675892 637871
rect 675852 637492 675904 637498
rect 675852 637434 675904 637440
rect 679624 637492 679676 637498
rect 679624 637434 679676 637440
rect 675496 637350 675892 637378
rect 675484 636880 675536 636886
rect 675484 636822 675536 636828
rect 675496 636585 675524 636822
rect 675482 636576 675538 636585
rect 675482 636511 675538 636520
rect 675864 636206 675892 637350
rect 675852 636200 675904 636206
rect 675852 636142 675904 636148
rect 675206 631408 675262 631417
rect 675206 631343 675262 631352
rect 675390 631408 675446 631417
rect 675390 631343 675446 631352
rect 675404 631258 675432 631343
rect 674852 631230 675432 631258
rect 675298 626376 675354 626385
rect 675298 626311 675354 626320
rect 675114 625968 675170 625977
rect 675114 625903 675170 625912
rect 675128 625190 675156 625903
rect 675312 625462 675340 626311
rect 675482 625560 675538 625569
rect 675482 625495 675538 625504
rect 675300 625456 675352 625462
rect 675300 625398 675352 625404
rect 675496 625326 675524 625495
rect 675484 625320 675536 625326
rect 675484 625262 675536 625268
rect 675116 625184 675168 625190
rect 675116 625126 675168 625132
rect 675298 625152 675354 625161
rect 675298 625087 675354 625096
rect 675114 624744 675170 624753
rect 675114 624679 675170 624688
rect 675128 623830 675156 624679
rect 675312 624102 675340 625087
rect 675482 624336 675538 624345
rect 675482 624271 675484 624280
rect 675536 624271 675538 624280
rect 675484 624242 675536 624248
rect 675300 624096 675352 624102
rect 675300 624038 675352 624044
rect 675484 623960 675536 623966
rect 675482 623928 675484 623937
rect 675536 623928 675538 623937
rect 675482 623863 675538 623872
rect 675116 623824 675168 623830
rect 675116 623766 675168 623772
rect 675298 623656 675354 623665
rect 676402 623656 676458 623665
rect 675354 623614 676402 623642
rect 675298 623591 675354 623600
rect 676402 623591 676458 623600
rect 675482 623520 675538 623529
rect 675482 623455 675538 623464
rect 675298 623112 675354 623121
rect 675298 623047 675354 623056
rect 675312 622606 675340 623047
rect 675496 622878 675524 623455
rect 675484 622872 675536 622878
rect 675484 622814 675536 622820
rect 675482 622704 675538 622713
rect 675482 622639 675538 622648
rect 675300 622600 675352 622606
rect 675300 622542 675352 622548
rect 675496 622470 675524 622639
rect 675484 622464 675536 622470
rect 675484 622406 675536 622412
rect 675298 622296 675354 622305
rect 675298 622231 675354 622240
rect 675312 621042 675340 622231
rect 679636 622033 679664 637434
rect 683394 636848 683450 636857
rect 683394 636783 683450 636792
rect 683210 636576 683266 636585
rect 683210 636511 683266 636520
rect 682384 636200 682436 636206
rect 682384 636142 682436 636148
rect 679622 622024 679678 622033
rect 679622 621959 679678 621968
rect 682396 621625 682424 636142
rect 682382 621616 682438 621625
rect 682382 621551 682438 621560
rect 675484 621240 675536 621246
rect 675484 621182 675536 621188
rect 675496 621081 675524 621182
rect 675482 621072 675538 621081
rect 675300 621036 675352 621042
rect 675482 621007 675538 621016
rect 675300 620978 675352 620984
rect 683224 620809 683252 636511
rect 683408 634814 683436 636783
rect 683408 634786 683620 634814
rect 683394 623656 683450 623665
rect 683394 623591 683450 623600
rect 683210 620800 683266 620809
rect 683210 620735 683266 620744
rect 675482 620256 675538 620265
rect 675482 620191 675538 620200
rect 675300 619880 675352 619886
rect 675298 619848 675300 619857
rect 675352 619848 675354 619857
rect 675298 619783 675354 619792
rect 675496 619682 675524 620191
rect 675484 619676 675536 619682
rect 675484 619618 675536 619624
rect 675484 619472 675536 619478
rect 675482 619440 675484 619449
rect 675536 619440 675538 619449
rect 675482 619375 675538 619384
rect 675484 618248 675536 618254
rect 675482 618216 675484 618225
rect 675536 618216 675538 618225
rect 675482 618151 675538 618160
rect 683408 617545 683436 623591
rect 683592 619177 683620 634786
rect 703694 626892 703722 627028
rect 704154 626892 704182 627028
rect 704614 626892 704642 627028
rect 705074 626892 705102 627028
rect 705534 626892 705562 627028
rect 705994 626892 706022 627028
rect 706454 626892 706482 627028
rect 706914 626892 706942 627028
rect 707374 626892 707402 627028
rect 707834 626892 707862 627028
rect 708294 626892 708322 627028
rect 708754 626892 708782 627028
rect 709214 626892 709242 627028
rect 683578 619168 683634 619177
rect 683578 619103 683634 619112
rect 683394 617536 683450 617545
rect 683394 617471 683450 617480
rect 675850 617264 675906 617273
rect 675850 617199 675906 617208
rect 674654 616992 674710 617001
rect 674654 616927 674710 616936
rect 675482 616584 675538 616593
rect 675482 616519 675538 616528
rect 675298 616176 675354 616185
rect 675298 616111 675300 616120
rect 675352 616111 675354 616120
rect 675300 616082 675352 616088
rect 675496 615806 675524 616519
rect 675484 615800 675536 615806
rect 675484 615742 675536 615748
rect 675864 615670 675892 617199
rect 675852 615664 675904 615670
rect 675852 615606 675904 615612
rect 683120 615664 683172 615670
rect 683120 615606 683172 615612
rect 683132 615505 683160 615606
rect 683118 615496 683174 615505
rect 683118 615431 683174 615440
rect 675482 614952 675538 614961
rect 675482 614887 675538 614896
rect 675496 614174 675524 614887
rect 675484 614168 675536 614174
rect 675484 614110 675536 614116
rect 675116 610020 675168 610026
rect 675116 609962 675168 609968
rect 674116 608566 674328 608594
rect 674012 601384 674064 601390
rect 674012 601326 674064 601332
rect 674024 599978 674052 601326
rect 673932 599950 674052 599978
rect 673932 592770 673960 599950
rect 674300 599706 674328 608566
rect 675128 607493 675156 609962
rect 675312 608110 675418 608138
rect 675312 607646 675340 608110
rect 675300 607640 675352 607646
rect 675300 607582 675352 607588
rect 675128 607465 675418 607493
rect 675128 606818 675418 606846
rect 675128 605878 675156 606818
rect 675116 605872 675168 605878
rect 675116 605814 675168 605820
rect 674852 604982 675418 605010
rect 674656 603356 674708 603362
rect 674656 603298 674708 603304
rect 674668 601390 674696 603298
rect 674656 601384 674708 601390
rect 674656 601326 674708 601332
rect 674024 599678 674328 599706
rect 674024 598934 674052 599678
rect 674288 599548 674340 599554
rect 674288 599490 674340 599496
rect 674024 598906 674144 598934
rect 674116 592929 674144 598906
rect 674102 592920 674158 592929
rect 674102 592855 674158 592864
rect 673932 592742 674236 592770
rect 673840 592006 673960 592034
rect 673932 591598 673960 592006
rect 674208 591682 674236 592742
rect 674116 591654 674236 591682
rect 673920 591592 673972 591598
rect 673920 591534 673972 591540
rect 674116 589274 674144 591654
rect 674116 589246 674236 589274
rect 674208 582374 674236 589246
rect 673932 582346 674236 582374
rect 673736 577584 673788 577590
rect 673736 577526 673788 577532
rect 673564 577238 673868 577266
rect 673380 576966 673684 576994
rect 673656 574569 673684 576966
rect 673642 574560 673698 574569
rect 673642 574495 673698 574504
rect 673840 569954 673868 577238
rect 673564 569926 673868 569954
rect 673564 547097 673592 569926
rect 673736 561740 673788 561746
rect 673736 561682 673788 561688
rect 673550 547088 673606 547097
rect 673550 547023 673606 547032
rect 673552 531820 673604 531826
rect 673552 531762 673604 531768
rect 673564 531486 673592 531762
rect 673552 531480 673604 531486
rect 673552 531422 673604 531428
rect 673748 485518 673776 561682
rect 673932 528358 673960 582346
rect 674104 577584 674156 577590
rect 674104 577526 674156 577532
rect 674116 572558 674144 577526
rect 674104 572552 674156 572558
rect 674104 572494 674156 572500
rect 674104 557728 674156 557734
rect 674104 557670 674156 557676
rect 673920 528352 673972 528358
rect 673920 528294 673972 528300
rect 674116 528154 674144 557670
rect 674104 528148 674156 528154
rect 674104 528090 674156 528096
rect 674300 528034 674328 599490
rect 674564 597508 674616 597514
rect 674564 597450 674616 597456
rect 674576 563054 674604 597450
rect 674852 586265 674880 604982
rect 675114 604480 675170 604489
rect 675170 604438 675418 604466
rect 675114 604415 675170 604424
rect 675496 603378 675524 603772
rect 675404 603362 675524 603378
rect 675392 603356 675524 603362
rect 675444 603350 675524 603356
rect 675392 603298 675444 603304
rect 675128 603146 675418 603174
rect 675128 602993 675156 603146
rect 675300 603084 675352 603090
rect 675300 603026 675352 603032
rect 675114 602984 675170 602993
rect 675114 602919 675170 602928
rect 675312 601694 675340 603026
rect 675220 601666 675340 601694
rect 675220 601202 675248 601666
rect 675220 601174 675432 601202
rect 675404 600644 675432 601174
rect 675496 599865 675524 600100
rect 675482 599856 675538 599865
rect 675482 599791 675538 599800
rect 675116 599548 675168 599554
rect 675168 599496 675418 599502
rect 675116 599490 675418 599496
rect 675128 599474 675418 599490
rect 675116 599412 675168 599418
rect 675116 599354 675168 599360
rect 675128 596442 675156 599354
rect 675312 598862 675432 598890
rect 675312 598738 675340 598862
rect 675404 598808 675432 598862
rect 675300 598732 675352 598738
rect 675300 598674 675352 598680
rect 675404 597530 675432 597652
rect 675312 597514 675432 597530
rect 675300 597508 675432 597514
rect 675352 597502 675432 597508
rect 675300 597450 675352 597456
rect 675128 596414 675418 596442
rect 675036 595802 675340 595830
rect 674838 586256 674894 586265
rect 674838 586191 674894 586200
rect 675036 582374 675064 595802
rect 675312 595762 675340 595802
rect 675404 595762 675432 595816
rect 675312 595734 675432 595762
rect 674944 582346 675064 582374
rect 675128 595122 675418 595150
rect 674748 580032 674800 580038
rect 674748 579974 674800 579980
rect 674760 579873 674788 579974
rect 674746 579864 674802 579873
rect 674746 579799 674802 579808
rect 674944 571577 674972 582346
rect 674930 571568 674986 571577
rect 674930 571503 674986 571512
rect 675128 563054 675156 595122
rect 675404 593609 675432 593980
rect 675390 593600 675446 593609
rect 675390 593535 675446 593544
rect 675850 592920 675906 592929
rect 675850 592855 675906 592864
rect 678242 592920 678298 592929
rect 678242 592855 678298 592864
rect 675484 591592 675536 591598
rect 675484 591534 675536 591540
rect 675496 591274 675524 591534
rect 675864 591462 675892 592855
rect 676034 592648 676090 592657
rect 676034 592583 676090 592592
rect 675852 591456 675904 591462
rect 675852 591398 675904 591404
rect 675852 591320 675904 591326
rect 675496 591268 675852 591274
rect 675496 591262 675904 591268
rect 675496 591246 675892 591262
rect 675482 581088 675538 581097
rect 675482 581023 675484 581032
rect 675536 581023 675538 581032
rect 675484 580994 675536 581000
rect 675298 580680 675354 580689
rect 675298 580615 675354 580624
rect 675312 579834 675340 580615
rect 675482 580272 675538 580281
rect 675482 580207 675538 580216
rect 675300 579828 675352 579834
rect 675300 579770 675352 579776
rect 675496 579698 675524 580207
rect 675484 579692 675536 579698
rect 675484 579634 675536 579640
rect 675482 579456 675538 579465
rect 675482 579391 675484 579400
rect 675536 579391 675538 579400
rect 675484 579362 675536 579368
rect 675484 579080 675536 579086
rect 675482 579048 675484 579057
rect 675536 579048 675538 579057
rect 675482 578983 675538 578992
rect 675482 578640 675538 578649
rect 675482 578575 675484 578584
rect 675536 578575 675538 578584
rect 675484 578546 675536 578552
rect 675484 578264 675536 578270
rect 675298 578232 675354 578241
rect 675484 578206 675536 578212
rect 675298 578167 675354 578176
rect 675312 578066 675340 578167
rect 675300 578060 675352 578066
rect 675300 578002 675352 578008
rect 675298 577824 675354 577833
rect 675298 577759 675300 577768
rect 675352 577759 675354 577768
rect 675300 577730 675352 577736
rect 675300 577448 675352 577454
rect 675298 577416 675300 577425
rect 675352 577416 675354 577425
rect 675298 577351 675354 577360
rect 675298 577008 675354 577017
rect 675298 576943 675300 576952
rect 675352 576943 675354 576952
rect 675300 576914 675352 576920
rect 675496 576609 675524 578206
rect 675482 576600 675538 576609
rect 675482 576535 675538 576544
rect 676048 575793 676076 592583
rect 676034 575784 676090 575793
rect 676034 575719 676090 575728
rect 678256 575657 678284 592855
rect 683212 591456 683264 591462
rect 683212 591398 683264 591404
rect 678242 575648 678298 575657
rect 678242 575583 678298 575592
rect 675298 574968 675354 574977
rect 675298 574903 675354 574912
rect 675312 574122 675340 574903
rect 675484 574320 675536 574326
rect 675484 574262 675536 574268
rect 675496 574161 675524 574262
rect 675482 574152 675538 574161
rect 675300 574116 675352 574122
rect 675482 574087 675538 574096
rect 675300 574058 675352 574064
rect 675484 573776 675536 573782
rect 675482 573744 675484 573753
rect 675536 573744 675538 573753
rect 675482 573679 675538 573688
rect 675484 572960 675536 572966
rect 675482 572928 675484 572937
rect 675536 572928 675538 572937
rect 675482 572863 675538 572872
rect 675484 572552 675536 572558
rect 675482 572520 675484 572529
rect 675536 572520 675538 572529
rect 675482 572455 675538 572464
rect 675482 572112 675538 572121
rect 675482 572047 675538 572056
rect 675496 571402 675524 572047
rect 683224 571985 683252 591398
rect 683396 591320 683448 591326
rect 683396 591262 683448 591268
rect 683210 571976 683266 571985
rect 683210 571911 683266 571920
rect 675484 571396 675536 571402
rect 675484 571338 675536 571344
rect 683408 571169 683436 591262
rect 703694 581740 703722 581876
rect 704154 581740 704182 581876
rect 704614 581740 704642 581876
rect 705074 581740 705102 581876
rect 705534 581740 705562 581876
rect 705994 581740 706022 581876
rect 706454 581740 706482 581876
rect 706914 581740 706942 581876
rect 707374 581740 707402 581876
rect 707834 581740 707862 581876
rect 708294 581740 708322 581876
rect 708754 581740 708782 581876
rect 709214 581740 709242 581876
rect 683394 571160 683450 571169
rect 683394 571095 683450 571104
rect 675482 570888 675538 570897
rect 675482 570823 675484 570832
rect 675536 570823 675538 570832
rect 675484 570794 675536 570800
rect 683118 570344 683174 570353
rect 683118 570279 683174 570288
rect 675496 570178 675892 570194
rect 675484 570172 675892 570178
rect 675536 570166 675892 570172
rect 675484 570114 675536 570120
rect 675864 570110 675892 570166
rect 683132 570110 683160 570279
rect 675852 570104 675904 570110
rect 675852 570046 675904 570052
rect 683120 570104 683172 570110
rect 683120 570046 683172 570052
rect 675482 569664 675538 569673
rect 675482 569599 675484 569608
rect 675536 569599 675538 569608
rect 675484 569570 675536 569576
rect 675300 564460 675352 564466
rect 675300 564402 675352 564408
rect 674484 563026 674604 563054
rect 674944 563026 675156 563054
rect 675312 563054 675340 564402
rect 675312 563026 675432 563054
rect 674484 554826 674512 563026
rect 674484 554798 674696 554826
rect 674472 554328 674524 554334
rect 673932 528006 674328 528034
rect 674392 554276 674472 554282
rect 674392 554270 674524 554276
rect 674392 554254 674512 554270
rect 673932 527678 673960 528006
rect 674104 527944 674156 527950
rect 674104 527886 674156 527892
rect 673920 527672 673972 527678
rect 673920 527614 673972 527620
rect 673736 485512 673788 485518
rect 673736 485454 673788 485460
rect 674116 483177 674144 527886
rect 674102 483168 674158 483177
rect 674102 483103 674158 483112
rect 674392 482769 674420 554254
rect 674668 554044 674696 554798
rect 674576 554016 674696 554044
rect 674576 546825 674604 554016
rect 674944 553874 674972 563026
rect 675404 562904 675432 563026
rect 675128 562278 675418 562306
rect 675128 561746 675156 562278
rect 675390 561912 675446 561921
rect 675390 561847 675446 561856
rect 675116 561740 675168 561746
rect 675116 561682 675168 561688
rect 675404 561612 675432 561847
rect 675300 560380 675352 560386
rect 675300 560322 675352 560328
rect 675312 558498 675340 560322
rect 675496 559473 675524 559776
rect 675482 559464 675538 559473
rect 675482 559399 675538 559408
rect 675772 559065 675800 559232
rect 675758 559056 675814 559065
rect 675758 558991 675814 559000
rect 675404 558498 675432 558620
rect 675312 558470 675432 558498
rect 675128 557926 675418 557954
rect 675128 557734 675156 557926
rect 675116 557728 675168 557734
rect 675116 557670 675168 557676
rect 675300 557592 675352 557598
rect 675300 557534 675352 557540
rect 675312 555370 675340 557534
rect 675404 555370 675432 555492
rect 675312 555342 675432 555370
rect 675128 554905 675418 554933
rect 675128 554334 675156 554905
rect 675300 554804 675352 554810
rect 675300 554746 675352 554752
rect 675116 554328 675168 554334
rect 675116 554270 675168 554276
rect 675116 554056 675168 554062
rect 674760 553846 674972 553874
rect 675036 554004 675116 554010
rect 675036 553998 675168 554004
rect 675036 553982 675156 553998
rect 674760 547369 674788 553846
rect 675036 551253 675064 553982
rect 675312 553738 675340 554746
rect 675496 554033 675524 554268
rect 675482 554024 675538 554033
rect 675482 553959 675538 553968
rect 675128 553710 675340 553738
rect 675128 552446 675156 553710
rect 675404 553602 675432 553656
rect 675312 553574 675432 553602
rect 675312 553518 675340 553574
rect 675300 553512 675352 553518
rect 675300 553454 675352 553460
rect 675128 552418 675418 552446
rect 675036 551225 675418 551253
rect 675024 550656 675076 550662
rect 675024 550598 675076 550604
rect 675036 549817 675064 550598
rect 675404 550361 675432 550596
rect 675390 550352 675446 550361
rect 675390 550287 675446 550296
rect 675220 549937 675418 549965
rect 675022 549808 675078 549817
rect 675022 549743 675078 549752
rect 675220 548978 675248 549937
rect 675482 549264 675538 549273
rect 675482 549199 675538 549208
rect 674944 548950 675248 548978
rect 674746 547360 674802 547369
rect 674746 547295 674802 547304
rect 674562 546816 674618 546825
rect 674562 546751 674618 546760
rect 674562 535120 674618 535129
rect 674562 535055 674618 535064
rect 674576 534274 674604 535055
rect 674748 534608 674800 534614
rect 674748 534550 674800 534556
rect 674564 534268 674616 534274
rect 674564 534210 674616 534216
rect 674760 534177 674788 534550
rect 674746 534168 674802 534177
rect 674746 534103 674802 534112
rect 674562 533624 674618 533633
rect 674562 533559 674618 533568
rect 674576 528554 674604 533559
rect 674746 531992 674802 532001
rect 674746 531927 674802 531936
rect 674760 531350 674788 531927
rect 674748 531344 674800 531350
rect 674748 531286 674800 531292
rect 674576 528526 674696 528554
rect 674668 495434 674696 528526
rect 674576 495406 674696 495434
rect 674576 490113 674604 495406
rect 674746 492144 674802 492153
rect 674746 492079 674802 492088
rect 674760 491502 674788 492079
rect 674748 491496 674800 491502
rect 674748 491438 674800 491444
rect 674562 490104 674618 490113
rect 674562 490039 674618 490048
rect 674748 485512 674800 485518
rect 674748 485454 674800 485460
rect 674760 485217 674788 485454
rect 674746 485208 674802 485217
rect 674746 485143 674802 485152
rect 674378 482760 674434 482769
rect 674378 482695 674434 482704
rect 673736 481908 673788 481914
rect 673736 481850 673788 481856
rect 673274 394632 673330 394641
rect 673274 394567 673330 394576
rect 673460 394324 673512 394330
rect 673460 394266 673512 394272
rect 673472 393258 673500 394266
rect 673380 393230 673500 393258
rect 673380 377874 673408 393230
rect 673368 377868 673420 377874
rect 673368 377810 673420 377816
rect 673092 354884 673144 354890
rect 673092 354826 673144 354832
rect 673092 354748 673144 354754
rect 673092 354690 673144 354696
rect 672816 353456 672868 353462
rect 672816 353398 672868 353404
rect 672632 348900 672684 348906
rect 672632 348842 672684 348848
rect 672644 332450 672672 348842
rect 672632 332444 672684 332450
rect 672632 332386 672684 332392
rect 672828 310078 672856 353398
rect 673104 310894 673132 354690
rect 673368 353592 673420 353598
rect 673368 353534 673420 353540
rect 673380 340746 673408 353534
rect 673552 349308 673604 349314
rect 673552 349250 673604 349256
rect 673368 340740 673420 340746
rect 673368 340682 673420 340688
rect 673274 340504 673330 340513
rect 673274 340439 673330 340448
rect 673288 338026 673316 340439
rect 673276 338020 673328 338026
rect 673276 337962 673328 337968
rect 673564 335510 673592 349250
rect 673552 335504 673604 335510
rect 673552 335446 673604 335452
rect 673552 324352 673604 324358
rect 673552 324294 673604 324300
rect 673092 310888 673144 310894
rect 673092 310830 673144 310836
rect 672816 310072 672868 310078
rect 672816 310014 672868 310020
rect 673092 305516 673144 305522
rect 673092 305458 673144 305464
rect 672540 303476 672592 303482
rect 672540 303418 672592 303424
rect 672552 302234 672580 303418
rect 672460 302206 672580 302234
rect 672460 299474 672488 302206
rect 672460 299446 672580 299474
rect 672356 297764 672408 297770
rect 672356 297706 672408 297712
rect 672552 294794 672580 299446
rect 672724 297764 672776 297770
rect 672724 297706 672776 297712
rect 672000 216034 672120 216050
rect 671988 216028 672120 216034
rect 672040 216022 672120 216028
rect 672184 294766 672580 294794
rect 672184 216050 672212 294766
rect 672736 289882 672764 297706
rect 672356 289876 672408 289882
rect 672356 289818 672408 289824
rect 672724 289876 672776 289882
rect 672724 289818 672776 289824
rect 672368 217394 672396 289818
rect 673104 285569 673132 305458
rect 673368 303884 673420 303890
rect 673368 303826 673420 303832
rect 673380 286521 673408 303826
rect 673366 286512 673422 286521
rect 673366 286447 673422 286456
rect 673090 285560 673146 285569
rect 673090 285495 673146 285504
rect 672538 278760 672594 278769
rect 672538 278695 672594 278704
rect 672356 217388 672408 217394
rect 672356 217330 672408 217336
rect 672184 216022 672304 216050
rect 671988 215970 672040 215976
rect 672276 215626 672304 216022
rect 672264 215620 672316 215626
rect 672264 215562 672316 215568
rect 671986 215520 672042 215529
rect 671986 215455 672042 215464
rect 672172 215484 672224 215490
rect 672000 215294 672028 215455
rect 672172 215426 672224 215432
rect 672184 215370 672212 215426
rect 671908 215266 672028 215294
rect 672092 215342 672212 215370
rect 671908 214146 671936 215266
rect 671908 214118 672028 214146
rect 671724 211262 671844 211290
rect 671540 211126 671660 211154
rect 671540 201494 671568 211126
rect 671816 209774 671844 211262
rect 671724 209746 671844 209774
rect 671724 206786 671752 209746
rect 671712 206780 671764 206786
rect 671712 206722 671764 206728
rect 671712 206644 671764 206650
rect 671712 206586 671764 206592
rect 671724 204049 671752 206586
rect 671632 204021 671752 204049
rect 671632 202722 671660 204021
rect 671632 202694 671752 202722
rect 671540 201466 671660 201494
rect 671436 145580 671488 145586
rect 671436 145522 671488 145528
rect 671632 140486 671660 201466
rect 671724 166994 671752 202694
rect 672000 201346 672028 214118
rect 672092 209250 672120 215342
rect 672264 215280 672316 215286
rect 672184 215228 672264 215234
rect 672184 215222 672316 215228
rect 672184 215206 672304 215222
rect 672184 209522 672212 215206
rect 672356 215144 672408 215150
rect 672356 215086 672408 215092
rect 672368 210497 672396 215086
rect 672552 212673 672580 278695
rect 673368 260500 673420 260506
rect 673368 260442 673420 260448
rect 673092 258868 673144 258874
rect 673092 258810 673144 258816
rect 672724 258460 672776 258466
rect 672724 258402 672776 258408
rect 672538 212664 672594 212673
rect 672538 212599 672594 212608
rect 672540 210724 672592 210730
rect 672540 210666 672592 210672
rect 672354 210488 672410 210497
rect 672354 210423 672410 210432
rect 672184 209494 672304 209522
rect 672276 209438 672304 209494
rect 672264 209432 672316 209438
rect 672264 209374 672316 209380
rect 672354 209264 672410 209273
rect 672092 209222 672354 209250
rect 672354 209199 672410 209208
rect 672264 208956 672316 208962
rect 672264 208898 672316 208904
rect 672276 208162 672304 208898
rect 672092 208134 672304 208162
rect 672092 207890 672120 208134
rect 672092 207862 672212 207890
rect 671988 201340 672040 201346
rect 671988 201282 672040 201288
rect 671988 168700 672040 168706
rect 671988 168642 672040 168648
rect 671724 166966 671844 166994
rect 671620 140480 671672 140486
rect 671620 140422 671672 140428
rect 671816 136542 671844 166966
rect 672000 151774 672028 168642
rect 672184 168337 672212 207862
rect 672354 183560 672410 183569
rect 672354 183495 672410 183504
rect 672368 182918 672396 183495
rect 672356 182912 672408 182918
rect 672356 182854 672408 182860
rect 672552 178294 672580 210666
rect 672540 178288 672592 178294
rect 672540 178230 672592 178236
rect 672356 169108 672408 169114
rect 672356 169050 672408 169056
rect 672170 168328 672226 168337
rect 672170 168263 672226 168272
rect 672368 153202 672396 169050
rect 672540 168292 672592 168298
rect 672540 168234 672592 168240
rect 672356 153196 672408 153202
rect 672356 153138 672408 153144
rect 671988 151768 672040 151774
rect 671988 151710 672040 151716
rect 671804 136536 671856 136542
rect 671804 136478 671856 136484
rect 671344 122868 671396 122874
rect 671344 122810 671396 122816
rect 670976 115864 671028 115870
rect 670976 115806 671028 115812
rect 671356 114374 671384 122810
rect 671528 120760 671580 120766
rect 671528 120702 671580 120708
rect 671344 114368 671396 114374
rect 671344 114310 671396 114316
rect 670148 112940 670200 112946
rect 670148 112882 670200 112888
rect 671540 111654 671568 120702
rect 672552 119270 672580 168234
rect 672736 129062 672764 258402
rect 672908 250436 672960 250442
rect 672908 250378 672960 250384
rect 672920 241777 672948 250378
rect 672906 241768 672962 241777
rect 673104 241738 673132 258810
rect 672906 241703 672962 241712
rect 673092 241732 673144 241738
rect 673092 241674 673144 241680
rect 673380 241602 673408 260442
rect 673368 241596 673420 241602
rect 673368 241538 673420 241544
rect 672908 217388 672960 217394
rect 672908 217330 672960 217336
rect 672920 215150 672948 217330
rect 673368 216164 673420 216170
rect 673368 216106 673420 216112
rect 672908 215144 672960 215150
rect 672908 215086 672960 215092
rect 673092 213716 673144 213722
rect 673092 213658 673144 213664
rect 672908 213308 672960 213314
rect 672908 213250 672960 213256
rect 672724 129056 672776 129062
rect 672724 128998 672776 129004
rect 672724 125656 672776 125662
rect 672724 125598 672776 125604
rect 672540 119264 672592 119270
rect 672540 119206 672592 119212
rect 671528 111648 671580 111654
rect 671528 111590 671580 111596
rect 672736 111178 672764 125598
rect 672920 124166 672948 213250
rect 673104 200530 673132 213658
rect 673380 201890 673408 216106
rect 673368 201884 673420 201890
rect 673368 201826 673420 201832
rect 673092 200524 673144 200530
rect 673092 200466 673144 200472
rect 673564 190097 673592 324294
rect 673748 210497 673776 481850
rect 674944 481545 674972 548950
rect 675496 548760 675524 549199
rect 675482 547904 675538 547913
rect 675482 547839 675538 547848
rect 675206 545864 675262 545873
rect 675206 545799 675262 545808
rect 675220 511994 675248 545799
rect 675496 543734 675524 547839
rect 675758 547632 675814 547641
rect 675758 547567 675814 547576
rect 675128 511966 675248 511994
rect 675312 543706 675524 543734
rect 675128 508881 675156 511966
rect 675114 508872 675170 508881
rect 675114 508807 675170 508816
rect 675114 491736 675170 491745
rect 675114 491671 675170 491680
rect 675128 491366 675156 491671
rect 675116 491360 675168 491366
rect 675116 491302 675168 491308
rect 675312 487234 675340 543706
rect 675482 536072 675538 536081
rect 675482 536007 675538 536016
rect 675496 535702 675524 536007
rect 675484 535696 675536 535702
rect 675484 535638 675536 535644
rect 675482 535528 675538 535537
rect 675482 535463 675484 535472
rect 675536 535463 675538 535472
rect 675484 535434 675536 535440
rect 675482 534848 675538 534857
rect 675482 534783 675538 534792
rect 675496 534614 675524 534783
rect 675484 534608 675536 534614
rect 675484 534550 675536 534556
rect 675482 534440 675538 534449
rect 675482 534375 675538 534384
rect 675496 534138 675524 534375
rect 675484 534132 675536 534138
rect 675484 534074 675536 534080
rect 675482 533216 675538 533225
rect 675482 533151 675538 533160
rect 675496 532914 675524 533151
rect 675484 532908 675536 532914
rect 675484 532850 675536 532856
rect 675482 532400 675538 532409
rect 675482 532335 675538 532344
rect 675496 531826 675524 532335
rect 675484 531820 675536 531826
rect 675484 531762 675536 531768
rect 675484 531616 675536 531622
rect 675482 531584 675484 531593
rect 675536 531584 675538 531593
rect 675482 531519 675538 531528
rect 675482 530768 675538 530777
rect 675482 530703 675538 530712
rect 675496 530126 675524 530703
rect 675484 530120 675536 530126
rect 675484 530062 675536 530068
rect 675484 529984 675536 529990
rect 675482 529952 675484 529961
rect 675536 529952 675538 529961
rect 675482 529887 675538 529896
rect 675482 529408 675538 529417
rect 675482 529343 675484 529352
rect 675536 529343 675538 529352
rect 675484 529314 675536 529320
rect 675482 529136 675538 529145
rect 675482 529071 675538 529080
rect 675496 528630 675524 529071
rect 675484 528624 675536 528630
rect 675484 528566 675536 528572
rect 675484 528352 675536 528358
rect 675482 528320 675484 528329
rect 675536 528320 675538 528329
rect 675482 528255 675538 528264
rect 675484 527672 675536 527678
rect 675482 527640 675484 527649
rect 675536 527640 675538 527649
rect 675482 527575 675538 527584
rect 675482 526144 675538 526153
rect 675482 526079 675538 526088
rect 675496 525842 675524 526079
rect 675484 525836 675536 525842
rect 675484 525778 675536 525784
rect 675482 524648 675538 524657
rect 675482 524583 675538 524592
rect 675496 524482 675524 524583
rect 675484 524476 675536 524482
rect 675484 524418 675536 524424
rect 675484 491632 675536 491638
rect 675484 491574 675536 491580
rect 675496 491337 675524 491574
rect 675482 491328 675538 491337
rect 675482 491263 675538 491272
rect 675482 490920 675538 490929
rect 675482 490855 675538 490864
rect 675496 490074 675524 490855
rect 675484 490068 675536 490074
rect 675484 490010 675536 490016
rect 675482 488472 675538 488481
rect 675482 488407 675538 488416
rect 675496 487354 675524 488407
rect 675772 487665 675800 547567
rect 675942 547360 675998 547369
rect 675942 547295 675944 547304
rect 675996 547295 675998 547304
rect 678244 547324 678296 547330
rect 675944 547266 675996 547272
rect 678244 547266 678296 547272
rect 676128 547188 676180 547194
rect 676128 547130 676180 547136
rect 675942 547088 675998 547097
rect 675942 547023 675998 547032
rect 675956 545766 675984 547023
rect 676140 546825 676168 547130
rect 676126 546816 676182 546825
rect 676126 546751 676182 546760
rect 675944 545760 675996 545766
rect 675944 545702 675996 545708
rect 675942 532876 675998 532885
rect 675942 532811 675998 532820
rect 675956 489297 675984 532811
rect 678256 525774 678284 547266
rect 683396 547188 683448 547194
rect 683396 547130 683448 547136
rect 683212 545760 683264 545766
rect 683212 545702 683264 545708
rect 682382 545184 682438 545193
rect 682382 545119 682438 545128
rect 682396 530641 682424 545119
rect 682382 530632 682438 530641
rect 682382 530567 682438 530576
rect 683224 526969 683252 545702
rect 683408 528193 683436 547130
rect 703694 536724 703722 536860
rect 704154 536724 704182 536860
rect 704614 536724 704642 536860
rect 705074 536724 705102 536860
rect 705534 536724 705562 536860
rect 705994 536724 706022 536860
rect 706454 536724 706482 536860
rect 706914 536724 706942 536860
rect 707374 536724 707402 536860
rect 707834 536724 707862 536860
rect 708294 536724 708322 536860
rect 708754 536724 708782 536860
rect 709214 536724 709242 536860
rect 683394 528184 683450 528193
rect 683394 528119 683450 528128
rect 683210 526960 683266 526969
rect 683210 526895 683266 526904
rect 678244 525768 678296 525774
rect 683120 525768 683172 525774
rect 678244 525710 678296 525716
rect 683118 525736 683120 525745
rect 683172 525736 683174 525745
rect 683118 525671 683174 525680
rect 676126 508872 676182 508881
rect 676126 508807 676182 508816
rect 676140 503538 676168 508807
rect 676128 503532 676180 503538
rect 676128 503474 676180 503480
rect 679624 503532 679676 503538
rect 679624 503474 679676 503480
rect 677414 490512 677470 490521
rect 677414 490447 677470 490456
rect 677230 489696 677286 489705
rect 677230 489631 677286 489640
rect 675942 489288 675998 489297
rect 675942 489223 675998 489232
rect 676034 488880 676090 488889
rect 676034 488815 676090 488824
rect 676048 488186 676076 488815
rect 676048 488158 676168 488186
rect 675942 488064 675998 488073
rect 675942 487999 675998 488008
rect 675758 487656 675814 487665
rect 675758 487591 675814 487600
rect 675484 487348 675536 487354
rect 675484 487290 675536 487296
rect 675312 487206 675524 487234
rect 675298 486840 675354 486849
rect 675298 486775 675354 486784
rect 675312 485858 675340 486775
rect 675496 486441 675524 487206
rect 675482 486432 675538 486441
rect 675482 486367 675538 486376
rect 675482 486024 675538 486033
rect 675482 485959 675484 485968
rect 675536 485959 675538 485968
rect 675484 485930 675536 485936
rect 675300 485852 675352 485858
rect 675300 485794 675352 485800
rect 675482 485616 675538 485625
rect 675482 485551 675538 485560
rect 675496 484566 675524 485551
rect 675484 484560 675536 484566
rect 675484 484502 675536 484508
rect 675482 484392 675538 484401
rect 675482 484327 675538 484336
rect 675300 484016 675352 484022
rect 675298 483984 675300 483993
rect 675352 483984 675354 483993
rect 675298 483919 675354 483928
rect 675300 483608 675352 483614
rect 675298 483576 675300 483585
rect 675352 483576 675354 483585
rect 675298 483511 675354 483520
rect 675496 483138 675524 484327
rect 675484 483132 675536 483138
rect 675484 483074 675536 483080
rect 675484 482384 675536 482390
rect 675482 482352 675484 482361
rect 675536 482352 675538 482361
rect 675482 482287 675538 482296
rect 675482 481944 675538 481953
rect 675482 481879 675484 481888
rect 675536 481879 675538 481888
rect 675484 481850 675536 481856
rect 674930 481536 674986 481545
rect 674930 481471 674986 481480
rect 675482 480720 675538 480729
rect 675482 480655 675484 480664
rect 675536 480655 675538 480664
rect 675484 480626 675536 480632
rect 675956 408494 675984 487999
rect 676140 476114 676168 488158
rect 676048 476086 676168 476114
rect 676048 470594 676076 476086
rect 676048 470566 676168 470594
rect 676140 412634 676168 470566
rect 675864 408466 675984 408494
rect 676048 412606 676168 412634
rect 675298 403880 675354 403889
rect 675298 403815 675354 403824
rect 675312 403442 675340 403815
rect 675482 403472 675538 403481
rect 675300 403436 675352 403442
rect 675482 403407 675538 403416
rect 675300 403378 675352 403384
rect 675496 403238 675524 403407
rect 675484 403232 675536 403238
rect 675484 403174 675536 403180
rect 675482 403064 675538 403073
rect 675482 402999 675484 403008
rect 675536 402999 675538 403008
rect 675484 402970 675536 402976
rect 674654 402248 674710 402257
rect 674654 402183 674710 402192
rect 673920 401396 673972 401402
rect 673920 401338 673972 401344
rect 673932 357338 673960 401338
rect 674286 396128 674342 396137
rect 674286 396063 674342 396072
rect 674102 393680 674158 393689
rect 674102 393615 674158 393624
rect 673920 357332 673972 357338
rect 673920 357274 673972 357280
rect 673920 357060 673972 357066
rect 673920 357002 673972 357008
rect 673932 312526 673960 357002
rect 673920 312520 673972 312526
rect 673920 312462 673972 312468
rect 673918 249792 673974 249801
rect 673918 249727 673974 249736
rect 673932 214033 673960 249727
rect 673918 214024 673974 214033
rect 673918 213959 673974 213968
rect 673734 210488 673790 210497
rect 673734 210423 673790 210432
rect 673920 210452 673972 210458
rect 673920 210394 673972 210400
rect 673550 190088 673606 190097
rect 673550 190023 673606 190032
rect 673182 183560 673238 183569
rect 673182 183495 673238 183504
rect 673196 177954 673224 183495
rect 673184 177948 673236 177954
rect 673184 177890 673236 177896
rect 673276 176724 673328 176730
rect 673276 176666 673328 176672
rect 673092 175228 673144 175234
rect 673092 175170 673144 175176
rect 673104 130286 673132 175170
rect 673288 171850 673316 176666
rect 673196 171822 673316 171850
rect 673196 147674 673224 171822
rect 673368 171216 673420 171222
rect 673288 171164 673368 171170
rect 673288 171158 673420 171164
rect 673288 171142 673408 171158
rect 673288 166994 673316 171142
rect 673288 166966 673408 166994
rect 673380 157010 673408 166966
rect 673368 157004 673420 157010
rect 673368 156946 673420 156952
rect 673196 147646 673408 147674
rect 673380 131306 673408 147646
rect 673932 133006 673960 210394
rect 674116 158370 674144 393615
rect 674300 382226 674328 396063
rect 674470 395720 674526 395729
rect 674470 395655 674526 395664
rect 674288 382220 674340 382226
rect 674288 382162 674340 382168
rect 674484 375358 674512 395655
rect 674472 375352 674524 375358
rect 674472 375294 674524 375300
rect 674668 357513 674696 402183
rect 675482 401432 675538 401441
rect 675482 401367 675484 401376
rect 675536 401367 675538 401376
rect 675484 401338 675536 401344
rect 675482 400616 675538 400625
rect 675482 400551 675484 400560
rect 675536 400551 675538 400560
rect 675484 400522 675536 400528
rect 675864 400217 675892 408466
rect 676048 401033 676076 412606
rect 677244 402121 677272 489631
rect 677428 402937 677456 490447
rect 679636 487257 679664 503474
rect 683302 500984 683358 500993
rect 683302 500919 683358 500928
rect 679622 487248 679678 487257
rect 679622 487183 679678 487192
rect 683316 484809 683344 500919
rect 703694 492796 703722 492864
rect 704154 492796 704182 492864
rect 704614 492796 704642 492864
rect 705074 492796 705102 492864
rect 705534 492796 705562 492864
rect 705994 492796 706022 492864
rect 706454 492796 706482 492864
rect 706914 492796 706942 492864
rect 707374 492796 707402 492864
rect 707834 492796 707862 492864
rect 708294 492796 708322 492864
rect 708754 492796 708782 492864
rect 709214 492796 709242 492864
rect 683302 484800 683358 484809
rect 683302 484735 683358 484744
rect 703694 404532 703722 404668
rect 704154 404532 704182 404668
rect 704614 404532 704642 404668
rect 705074 404532 705102 404668
rect 705534 404532 705562 404668
rect 705994 404532 706022 404668
rect 706454 404532 706482 404668
rect 706914 404532 706942 404668
rect 707374 404532 707402 404668
rect 707834 404532 707862 404668
rect 708294 404532 708322 404668
rect 708754 404532 708782 404668
rect 709214 404532 709242 404668
rect 677414 402928 677470 402937
rect 677414 402863 677470 402872
rect 677230 402112 677286 402121
rect 677230 402047 677286 402056
rect 676034 401024 676090 401033
rect 676034 400959 676090 400968
rect 675850 400208 675906 400217
rect 675850 400143 675906 400152
rect 675482 399800 675538 399809
rect 675482 399735 675484 399744
rect 675536 399735 675538 399744
rect 675484 399706 675536 399712
rect 675666 399392 675722 399401
rect 675666 399327 675722 399336
rect 675114 398168 675170 398177
rect 675114 398103 675170 398112
rect 675128 382582 675156 398103
rect 675298 397352 675354 397361
rect 675298 397287 675354 397296
rect 675312 396098 675340 397287
rect 675482 396536 675538 396545
rect 675482 396471 675538 396480
rect 675496 396370 675524 396471
rect 675484 396364 675536 396370
rect 675484 396306 675536 396312
rect 675300 396092 675352 396098
rect 675300 396034 675352 396040
rect 675680 395978 675708 399327
rect 676218 398440 676274 398449
rect 676218 398375 676274 398384
rect 675220 395950 675708 395978
rect 675220 384449 675248 395950
rect 676232 394618 676260 398375
rect 681002 397624 681058 397633
rect 681002 397559 681058 397568
rect 675312 394590 676260 394618
rect 675312 386186 675340 394590
rect 675482 394496 675538 394505
rect 675482 394431 675538 394440
rect 675496 394330 675524 394431
rect 675484 394324 675536 394330
rect 675484 394266 675536 394272
rect 675482 394088 675538 394097
rect 675482 394023 675538 394032
rect 675496 393378 675524 394023
rect 675484 393372 675536 393378
rect 675484 393314 675536 393320
rect 675482 392456 675538 392465
rect 675482 392391 675538 392400
rect 675496 392018 675524 392391
rect 675484 392012 675536 392018
rect 675484 391954 675536 391960
rect 681016 388521 681044 397559
rect 683026 392728 683082 392737
rect 683026 392663 683082 392672
rect 683040 389881 683068 392663
rect 683026 389872 683082 389881
rect 683026 389807 683082 389816
rect 681002 388512 681058 388521
rect 681002 388447 681058 388456
rect 675312 386158 675432 386186
rect 675404 385696 675432 386158
rect 675772 384985 675800 385084
rect 675758 384976 675814 384985
rect 675758 384911 675814 384920
rect 675220 384421 675418 384449
rect 675312 382622 675432 382650
rect 675312 382582 675340 382622
rect 675128 382554 675340 382582
rect 675404 382568 675432 382622
rect 675392 382356 675444 382362
rect 675392 382298 675444 382304
rect 675116 382220 675168 382226
rect 675116 382162 675168 382168
rect 675128 381426 675156 382162
rect 675404 382024 675432 382298
rect 675128 381398 675418 381426
rect 675772 380633 675800 380732
rect 675758 380624 675814 380633
rect 675758 380559 675814 380568
rect 675758 378720 675814 378729
rect 675758 378655 675814 378664
rect 675772 378284 675800 378655
rect 675300 377868 675352 377874
rect 675300 377810 675352 377816
rect 675312 377618 675340 377810
rect 675404 377618 675432 377740
rect 675312 377590 675432 377618
rect 675758 377360 675814 377369
rect 675758 377295 675814 377304
rect 675772 377060 675800 377295
rect 675116 376508 675168 376514
rect 675168 376456 675340 376462
rect 675116 376450 675340 376456
rect 675128 376434 675340 376450
rect 675312 376394 675340 376434
rect 675404 376394 675432 376448
rect 675312 376366 675432 376394
rect 675116 375352 675168 375358
rect 675116 375294 675168 375300
rect 675128 375238 675156 375294
rect 675128 375210 675418 375238
rect 675298 375048 675354 375057
rect 675298 374983 675354 374992
rect 675312 373402 675340 374983
rect 675312 373374 675418 373402
rect 675666 373008 675722 373017
rect 675666 372943 675722 372952
rect 675680 372776 675708 372943
rect 675114 372600 675170 372609
rect 675114 372535 675170 372544
rect 675128 371566 675156 372535
rect 675128 371538 675418 371566
rect 703694 359380 703722 359516
rect 704154 359380 704182 359516
rect 704614 359380 704642 359516
rect 705074 359380 705102 359516
rect 705534 359380 705562 359516
rect 705994 359380 706022 359516
rect 706454 359380 706482 359516
rect 706914 359380 706942 359516
rect 707374 359380 707402 359516
rect 707834 359380 707862 359516
rect 708294 359380 708322 359516
rect 708754 359380 708782 359516
rect 709214 359380 709242 359516
rect 675298 358728 675354 358737
rect 675298 358663 675354 358672
rect 675114 358320 675170 358329
rect 675114 358255 675170 358264
rect 674654 357504 674710 357513
rect 675128 357474 675156 358255
rect 675312 357610 675340 358663
rect 675482 357912 675538 357921
rect 675482 357847 675538 357856
rect 675496 357746 675524 357847
rect 675484 357740 675536 357746
rect 675484 357682 675536 357688
rect 675300 357604 675352 357610
rect 675300 357546 675352 357552
rect 674654 357439 674710 357448
rect 675116 357468 675168 357474
rect 675116 357410 675168 357416
rect 674748 357332 674800 357338
rect 674748 357274 674800 357280
rect 674760 356697 674788 357274
rect 675482 357096 675538 357105
rect 675482 357031 675484 357040
rect 675536 357031 675538 357040
rect 675484 357002 675536 357008
rect 674746 356688 674802 356697
rect 674746 356623 674802 356632
rect 674654 356280 674710 356289
rect 674654 356215 674710 356224
rect 674470 349752 674526 349761
rect 674470 349687 674526 349696
rect 674286 348528 674342 348537
rect 674286 348463 674342 348472
rect 674104 158364 674156 158370
rect 674104 158306 674156 158312
rect 674300 138446 674328 348463
rect 674484 336734 674512 349687
rect 674472 336728 674524 336734
rect 674472 336670 674524 336676
rect 674472 335640 674524 335646
rect 674472 335582 674524 335588
rect 674484 335170 674512 335582
rect 674472 335164 674524 335170
rect 674472 335106 674524 335112
rect 674668 311681 674696 356215
rect 675482 355872 675538 355881
rect 675482 355807 675538 355816
rect 675298 355464 675354 355473
rect 675298 355399 675354 355408
rect 675312 354754 675340 355399
rect 675496 355230 675524 355807
rect 675484 355224 675536 355230
rect 675484 355166 675536 355172
rect 675482 355056 675538 355065
rect 675482 354991 675538 355000
rect 675496 354890 675524 354991
rect 675484 354884 675536 354890
rect 675484 354826 675536 354832
rect 675300 354748 675352 354754
rect 675300 354690 675352 354696
rect 675114 354648 675170 354657
rect 675114 354583 675170 354592
rect 675128 353462 675156 354583
rect 675298 353832 675354 353841
rect 675298 353767 675354 353776
rect 675116 353456 675168 353462
rect 675116 353398 675168 353404
rect 675312 353326 675340 353767
rect 675484 353592 675536 353598
rect 675484 353534 675536 353540
rect 675496 353433 675524 353534
rect 675482 353424 675538 353433
rect 675482 353359 675538 353368
rect 675300 353320 675352 353326
rect 675300 353262 675352 353268
rect 675482 352608 675538 352617
rect 675482 352543 675538 352552
rect 675496 351966 675524 352543
rect 675484 351960 675536 351966
rect 675484 351902 675536 351908
rect 675298 351384 675354 351393
rect 675298 351319 675354 351328
rect 675312 350606 675340 351319
rect 675484 350736 675536 350742
rect 675484 350678 675536 350684
rect 675300 350600 675352 350606
rect 675496 350577 675524 350678
rect 675300 350542 675352 350548
rect 675482 350568 675538 350577
rect 675482 350503 675538 350512
rect 675482 349344 675538 349353
rect 675482 349279 675484 349288
rect 675536 349279 675538 349288
rect 675484 349250 675536 349256
rect 675482 348936 675538 348945
rect 675482 348871 675484 348880
rect 675536 348871 675538 348880
rect 675484 348842 675536 348848
rect 683118 347712 683174 347721
rect 683118 347647 683174 347656
rect 675482 347304 675538 347313
rect 675482 347239 675538 347248
rect 675496 345030 675524 347239
rect 683132 346458 683160 347647
rect 675852 346452 675904 346458
rect 675852 346394 675904 346400
rect 683120 346452 683172 346458
rect 683120 346394 683172 346400
rect 675484 345024 675536 345030
rect 675484 344966 675536 344972
rect 675864 342145 675892 346394
rect 675850 342136 675906 342145
rect 675850 342071 675906 342080
rect 675116 340740 675168 340746
rect 675116 340682 675168 340688
rect 675128 340558 675156 340682
rect 675128 340530 675340 340558
rect 675312 340490 675340 340530
rect 675404 340490 675432 340544
rect 675312 340462 675432 340490
rect 675758 340368 675814 340377
rect 675758 340303 675814 340312
rect 675772 339864 675800 340303
rect 675666 339416 675722 339425
rect 675666 339351 675722 339360
rect 675680 339252 675708 339351
rect 675116 338020 675168 338026
rect 675116 337962 675168 337968
rect 675128 336857 675156 337962
rect 675574 337784 675630 337793
rect 675574 337719 675630 337728
rect 675588 337416 675616 337719
rect 675128 336829 675418 336857
rect 675116 336728 675168 336734
rect 675116 336670 675168 336676
rect 675758 336696 675814 336705
rect 675128 335594 675156 336670
rect 675758 336631 675814 336640
rect 675772 336192 675800 336631
rect 675128 335566 675340 335594
rect 675116 335504 675168 335510
rect 675116 335446 675168 335452
rect 675312 335458 675340 335566
rect 675404 335458 675432 335580
rect 674840 335164 674892 335170
rect 674840 335106 674892 335112
rect 674852 330049 674880 335106
rect 675128 332534 675156 335446
rect 675312 335430 675432 335458
rect 675300 333940 675352 333946
rect 675300 333882 675352 333888
rect 675312 333078 675340 333882
rect 675312 333050 675418 333078
rect 675128 332506 675418 332534
rect 675116 332444 675168 332450
rect 675116 332386 675168 332392
rect 675128 331242 675156 332386
rect 675758 332344 675814 332353
rect 675758 332279 675814 332288
rect 675772 331875 675800 332279
rect 675128 331214 675418 331242
rect 674852 330021 675418 330049
rect 675312 328222 675432 328250
rect 675312 328182 675340 328222
rect 674944 328154 675340 328182
rect 675404 328168 675432 328222
rect 674944 325650 674972 328154
rect 675128 327542 675418 327570
rect 674932 325644 674984 325650
rect 674932 325586 674984 325592
rect 675128 325514 675156 327542
rect 675758 326904 675814 326913
rect 675758 326839 675814 326848
rect 675772 326332 675800 326839
rect 675116 325508 675168 325514
rect 675116 325450 675168 325456
rect 703694 314364 703722 314500
rect 704154 314364 704182 314500
rect 704614 314364 704642 314500
rect 705074 314364 705102 314500
rect 705534 314364 705562 314500
rect 705994 314364 706022 314500
rect 706454 314364 706482 314500
rect 706914 314364 706942 314500
rect 707374 314364 707402 314500
rect 707834 314364 707862 314500
rect 708294 314364 708322 314500
rect 708754 314364 708782 314500
rect 709214 314364 709242 314500
rect 675482 313712 675538 313721
rect 675482 313647 675538 313656
rect 675496 313478 675524 313647
rect 675484 313472 675536 313478
rect 675484 313414 675536 313420
rect 675484 313336 675536 313342
rect 675482 313304 675484 313313
rect 675536 313304 675538 313313
rect 675482 313239 675538 313248
rect 675298 312896 675354 312905
rect 675298 312831 675354 312840
rect 675312 312050 675340 312831
rect 675484 312520 675536 312526
rect 675482 312488 675484 312497
rect 675536 312488 675538 312497
rect 675482 312423 675538 312432
rect 675482 312080 675538 312089
rect 675300 312044 675352 312050
rect 675482 312015 675538 312024
rect 675300 311986 675352 311992
rect 675496 311914 675524 312015
rect 675484 311908 675536 311914
rect 675484 311850 675536 311856
rect 674654 311672 674710 311681
rect 674654 311607 674710 311616
rect 675482 311264 675538 311273
rect 675482 311199 675538 311208
rect 675300 310888 675352 310894
rect 675298 310856 675300 310865
rect 675352 310856 675354 310865
rect 675298 310791 675354 310800
rect 675496 310554 675524 311199
rect 675484 310548 675536 310554
rect 675484 310490 675536 310496
rect 675298 310448 675354 310457
rect 675298 310383 675354 310392
rect 675312 309194 675340 310383
rect 675484 310072 675536 310078
rect 675482 310040 675484 310049
rect 675536 310040 675538 310049
rect 675482 309975 675538 309984
rect 675482 309632 675538 309641
rect 675482 309567 675538 309576
rect 675496 309398 675524 309567
rect 675484 309392 675536 309398
rect 675484 309334 675536 309340
rect 675482 309224 675538 309233
rect 675300 309188 675352 309194
rect 675482 309159 675538 309168
rect 675300 309130 675352 309136
rect 675022 308000 675078 308009
rect 675022 307935 675078 307944
rect 675036 307754 675064 307935
rect 675036 307726 675248 307754
rect 675022 307592 675078 307601
rect 675022 307527 675078 307536
rect 674470 306368 674526 306377
rect 674470 306303 674526 306312
rect 674484 292330 674512 306303
rect 674654 304328 674710 304337
rect 674654 304263 674710 304272
rect 674472 292324 674524 292330
rect 674472 292266 674524 292272
rect 674668 287518 674696 304263
rect 675036 298518 675064 307527
rect 674794 298512 674846 298518
rect 674760 298460 674794 298466
rect 674760 298454 674846 298460
rect 675024 298512 675076 298518
rect 675024 298454 675076 298460
rect 674760 298438 674834 298454
rect 674760 289814 674788 298438
rect 675220 298194 675248 307726
rect 675496 305674 675524 309159
rect 676034 308408 676090 308417
rect 676090 308366 676260 308394
rect 676034 308343 676090 308352
rect 674944 298166 675248 298194
rect 675312 305646 675524 305674
rect 674944 298058 674972 298166
rect 674944 298030 675156 298058
rect 675128 297378 675156 298030
rect 675036 297350 675156 297378
rect 675036 292414 675064 297350
rect 675312 296834 675340 305646
rect 675482 305552 675538 305561
rect 675482 305487 675484 305496
rect 675536 305487 675538 305496
rect 675484 305458 675536 305464
rect 676034 304736 676090 304745
rect 676034 304671 676090 304680
rect 675482 303920 675538 303929
rect 675482 303855 675484 303864
rect 675536 303855 675538 303864
rect 675484 303826 675536 303832
rect 675482 303512 675538 303521
rect 675482 303447 675484 303456
rect 675536 303447 675538 303456
rect 675484 303418 675536 303424
rect 676048 302977 676076 304671
rect 676034 302968 676090 302977
rect 676034 302903 676090 302912
rect 675482 302288 675538 302297
rect 675482 302223 675538 302232
rect 675496 300830 675524 302223
rect 675484 300824 675536 300830
rect 675484 300766 675536 300772
rect 676232 300665 676260 308366
rect 678242 307184 678298 307193
rect 678242 307119 678298 307128
rect 676402 305960 676458 305969
rect 676402 305895 676458 305904
rect 676416 301617 676444 305895
rect 676402 301608 676458 301617
rect 676402 301543 676458 301552
rect 675482 300656 675538 300665
rect 675482 300591 675538 300600
rect 676218 300656 676274 300665
rect 676218 300591 676274 300600
rect 675128 296806 675340 296834
rect 675128 294250 675156 296806
rect 675496 296274 675524 300591
rect 678256 297401 678284 307119
rect 681002 306776 681058 306785
rect 681002 306711 681058 306720
rect 680360 302252 680412 302258
rect 680360 302194 680412 302200
rect 680372 299441 680400 302194
rect 680358 299432 680414 299441
rect 680358 299367 680414 299376
rect 678242 297392 678298 297401
rect 678242 297327 678298 297336
rect 681016 297226 681044 306711
rect 683118 302696 683174 302705
rect 683118 302631 683174 302640
rect 683132 302258 683160 302631
rect 683120 302252 683172 302258
rect 683120 302194 683172 302200
rect 675852 297220 675904 297226
rect 675852 297162 675904 297168
rect 681004 297220 681056 297226
rect 681004 297162 681056 297168
rect 675864 296585 675892 297162
rect 675850 296576 675906 296585
rect 675850 296511 675906 296520
rect 675484 296268 675536 296274
rect 675484 296210 675536 296216
rect 675484 295928 675536 295934
rect 675484 295870 675536 295876
rect 675496 295528 675524 295870
rect 675574 295352 675630 295361
rect 675574 295287 675630 295296
rect 675588 294879 675616 295287
rect 675128 294222 675418 294250
rect 675036 292386 675418 292414
rect 675116 292324 675168 292330
rect 675116 292266 675168 292272
rect 675128 291870 675156 292266
rect 675128 291842 675418 291870
rect 675758 291544 675814 291553
rect 675758 291479 675814 291488
rect 675772 291176 675800 291479
rect 675758 291000 675814 291009
rect 675758 290935 675814 290944
rect 675772 290564 675800 290935
rect 674760 289786 674880 289814
rect 674852 288062 674880 289786
rect 675312 288102 675432 288130
rect 675312 288062 675340 288102
rect 674852 288034 675340 288062
rect 675404 288048 675432 288102
rect 674668 287490 675418 287518
rect 675758 287056 675814 287065
rect 675758 286991 675814 287000
rect 675772 286892 675800 286991
rect 675390 286512 675446 286521
rect 675390 286447 675446 286456
rect 675404 286212 675432 286447
rect 675114 285560 675170 285569
rect 675114 285495 675170 285504
rect 675128 285070 675156 285495
rect 675128 285042 675340 285070
rect 675312 285002 675340 285042
rect 675404 285002 675432 285056
rect 675312 284974 675432 285002
rect 675758 283656 675814 283665
rect 675758 283591 675814 283600
rect 675772 283220 675800 283591
rect 675666 282840 675722 282849
rect 675666 282775 675722 282784
rect 675680 282540 675708 282775
rect 675666 281616 675722 281625
rect 675666 281551 675722 281560
rect 675680 281355 675708 281551
rect 703694 269348 703722 269484
rect 704154 269348 704182 269484
rect 704614 269348 704642 269484
rect 705074 269348 705102 269484
rect 705534 269348 705562 269484
rect 705994 269348 706022 269484
rect 706454 269348 706482 269484
rect 706914 269348 706942 269484
rect 707374 269348 707402 269484
rect 707834 269348 707862 269484
rect 708294 269348 708322 269484
rect 708754 269348 708782 269484
rect 709214 269348 709242 269484
rect 675482 268696 675538 268705
rect 675482 268631 675538 268640
rect 675496 268530 675524 268631
rect 675484 268524 675536 268530
rect 675484 268466 675536 268472
rect 675484 268320 675536 268326
rect 675482 268288 675484 268297
rect 675536 268288 675538 268297
rect 675482 268223 675538 268232
rect 675482 267880 675538 267889
rect 675482 267815 675484 267824
rect 675536 267815 675538 267824
rect 675484 267786 675536 267792
rect 675482 267472 675538 267481
rect 675482 267407 675538 267416
rect 675298 267064 675354 267073
rect 675298 266999 675354 267008
rect 675312 266422 675340 266999
rect 675496 266830 675524 267407
rect 675484 266824 675536 266830
rect 675484 266766 675536 266772
rect 675482 266656 675538 266665
rect 675482 266591 675484 266600
rect 675536 266591 675538 266600
rect 675484 266562 675536 266568
rect 675300 266416 675352 266422
rect 675300 266358 675352 266364
rect 675482 266248 675538 266257
rect 675482 266183 675538 266192
rect 675298 265840 675354 265849
rect 675298 265775 675354 265784
rect 675312 265266 675340 265775
rect 675496 265606 675524 266183
rect 675484 265600 675536 265606
rect 675484 265542 675536 265548
rect 675484 265464 675536 265470
rect 675482 265432 675484 265441
rect 675536 265432 675538 265441
rect 675482 265367 675538 265376
rect 675300 265260 675352 265266
rect 675300 265202 675352 265208
rect 675484 265056 675536 265062
rect 675482 265024 675484 265033
rect 675536 265024 675538 265033
rect 675482 264959 675538 264968
rect 675482 264616 675538 264625
rect 675482 264551 675538 264560
rect 675496 263634 675524 264551
rect 675484 263628 675536 263634
rect 675484 263570 675536 263576
rect 676218 263256 676274 263265
rect 676218 263191 676274 263200
rect 675482 262576 675538 262585
rect 675482 262511 675484 262520
rect 675536 262511 675538 262520
rect 675484 262482 675536 262488
rect 675482 262168 675538 262177
rect 675482 262103 675484 262112
rect 675536 262103 675538 262112
rect 675484 262074 675536 262080
rect 674470 261352 674526 261361
rect 674470 261287 674526 261296
rect 674484 247042 674512 261287
rect 674838 261080 674894 261089
rect 674838 261015 674894 261024
rect 675850 261080 675906 261089
rect 675850 261015 675852 261024
rect 674654 259312 674710 259321
rect 674654 259247 674710 259256
rect 674472 247036 674524 247042
rect 674472 246978 674524 246984
rect 674668 244274 674696 259247
rect 674852 247926 674880 261015
rect 675904 261015 675906 261024
rect 675852 260986 675904 260992
rect 675482 260536 675538 260545
rect 675482 260471 675484 260480
rect 675536 260471 675538 260480
rect 675484 260442 675536 260448
rect 675482 260128 675538 260137
rect 675482 260063 675538 260072
rect 675496 259894 675524 260063
rect 675484 259888 675536 259894
rect 675484 259830 675536 259836
rect 675482 259720 675538 259729
rect 675482 259655 675484 259664
rect 675536 259655 675538 259664
rect 675484 259626 675536 259632
rect 676232 259570 676260 263191
rect 676402 262848 676458 262857
rect 676402 262783 676458 262792
rect 676416 261050 676444 262783
rect 676404 261044 676456 261050
rect 676404 260986 676456 260992
rect 675312 259542 676260 259570
rect 675022 254008 675078 254017
rect 675022 253943 675078 253952
rect 674840 247920 674892 247926
rect 674840 247862 674892 247868
rect 675036 246378 675064 253943
rect 675312 250526 675340 259542
rect 675482 258904 675538 258913
rect 675482 258839 675484 258848
rect 675536 258839 675538 258848
rect 675484 258810 675536 258816
rect 675482 258496 675538 258505
rect 675482 258431 675484 258440
rect 675536 258431 675538 258440
rect 675484 258402 675536 258408
rect 683118 257544 683174 257553
rect 683118 257479 683174 257488
rect 675482 257272 675538 257281
rect 675482 257207 675538 257216
rect 675496 253230 675524 257207
rect 683132 256766 683160 257479
rect 675852 256760 675904 256766
rect 675852 256702 675904 256708
rect 683120 256760 683172 256766
rect 683120 256702 683172 256708
rect 675864 254017 675892 256702
rect 675850 254008 675906 254017
rect 675850 253943 675906 253952
rect 675484 253224 675536 253230
rect 675484 253166 675536 253172
rect 675312 250498 675418 250526
rect 675206 249792 675262 249801
rect 675206 249727 675262 249736
rect 674576 244246 674696 244274
rect 674760 246350 675064 246378
rect 674576 242729 674604 244246
rect 674562 242720 674618 242729
rect 674562 242655 674618 242664
rect 674760 241346 674788 246350
rect 675220 244274 675248 249727
rect 675404 249642 675432 249900
rect 675312 249614 675432 249642
rect 675312 248414 675340 249614
rect 675574 249520 675630 249529
rect 675574 249455 675630 249464
rect 675588 249220 675616 249455
rect 675312 248386 675432 248414
rect 675404 248305 675432 248386
rect 675390 248296 675446 248305
rect 675390 248231 675446 248240
rect 675392 247920 675444 247926
rect 675392 247862 675444 247868
rect 675404 247384 675432 247862
rect 675392 247036 675444 247042
rect 675392 246978 675444 246984
rect 675404 246840 675432 246978
rect 675758 246664 675814 246673
rect 675758 246599 675814 246608
rect 675772 246199 675800 246599
rect 675390 245712 675446 245721
rect 675390 245647 675446 245656
rect 675404 245548 675432 245647
rect 675220 244246 675340 244274
rect 675312 243273 675340 244246
rect 675298 243264 675354 243273
rect 675298 243199 675354 243208
rect 675220 243057 675418 243085
rect 675220 242026 675248 243057
rect 675482 242720 675538 242729
rect 675482 242655 675538 242664
rect 675496 242519 675524 242655
rect 674944 241998 675248 242026
rect 675482 242040 675538 242049
rect 674944 241466 674972 241998
rect 675482 241975 675538 241984
rect 675496 241876 675524 241975
rect 675114 241768 675170 241777
rect 675114 241703 675170 241712
rect 675300 241732 675352 241738
rect 674932 241460 674984 241466
rect 674932 241402 674984 241408
rect 674760 241318 674880 241346
rect 674852 238134 674880 241318
rect 674840 238128 674892 238134
rect 674840 238070 674892 238076
rect 675128 236382 675156 241703
rect 675300 241674 675352 241680
rect 675312 241482 675340 241674
rect 675312 241454 675524 241482
rect 675496 241231 675524 241454
rect 675300 241120 675352 241126
rect 675300 241062 675352 241068
rect 675312 240054 675340 241062
rect 675312 240026 675418 240054
rect 675390 238640 675446 238649
rect 675390 238575 675446 238584
rect 675404 238204 675432 238575
rect 675300 238128 675352 238134
rect 675300 238070 675352 238076
rect 675312 237810 675340 238070
rect 675312 237782 675432 237810
rect 675404 237524 675432 237782
rect 675128 236354 675418 236382
rect 703694 224196 703722 224264
rect 704154 224196 704182 224264
rect 704614 224196 704642 224264
rect 705074 224196 705102 224264
rect 705534 224196 705562 224264
rect 705994 224196 706022 224264
rect 706454 224196 706482 224264
rect 706914 224196 706942 224264
rect 707374 224196 707402 224264
rect 707834 224196 707862 224264
rect 708294 224196 708322 224264
rect 708754 224196 708782 224264
rect 709214 224196 709242 224264
rect 675666 223544 675722 223553
rect 675666 223479 675722 223488
rect 675114 223136 675170 223145
rect 675114 223071 675170 223080
rect 675128 222630 675156 223071
rect 675484 222896 675536 222902
rect 675484 222838 675536 222844
rect 675300 222760 675352 222766
rect 675496 222737 675524 222838
rect 675300 222702 675352 222708
rect 675482 222728 675538 222737
rect 675116 222624 675168 222630
rect 675116 222566 675168 222572
rect 675312 222329 675340 222702
rect 675482 222663 675538 222672
rect 675680 222442 675708 223479
rect 675496 222414 675708 222442
rect 675298 222320 675354 222329
rect 675298 222255 675354 222264
rect 675496 222222 675524 222414
rect 675484 222216 675536 222222
rect 675484 222158 675536 222164
rect 675298 221912 675354 221921
rect 675298 221847 675354 221856
rect 675312 220862 675340 221847
rect 675482 221504 675538 221513
rect 675482 221439 675538 221448
rect 675496 221270 675524 221439
rect 675484 221264 675536 221270
rect 675484 221206 675536 221212
rect 675482 221096 675538 221105
rect 675482 221031 675484 221040
rect 675536 221031 675538 221040
rect 675484 221002 675536 221008
rect 675300 220856 675352 220862
rect 675300 220798 675352 220804
rect 675298 220688 675354 220697
rect 675298 220623 675354 220632
rect 674654 220280 674710 220289
rect 674654 220215 674710 220224
rect 674470 215384 674526 215393
rect 674470 215319 674526 215328
rect 674484 194546 674512 215319
rect 674668 195974 674696 220215
rect 675312 219638 675340 220623
rect 675482 219872 675538 219881
rect 675482 219807 675484 219816
rect 675536 219807 675538 219816
rect 675484 219778 675536 219784
rect 675300 219632 675352 219638
rect 675300 219574 675352 219580
rect 675484 219496 675536 219502
rect 675482 219464 675484 219473
rect 675536 219464 675538 219473
rect 675482 219399 675538 219408
rect 675574 219056 675630 219065
rect 675574 218991 675630 219000
rect 675206 217832 675262 217841
rect 675206 217767 675262 217776
rect 674930 214160 674986 214169
rect 674930 214095 674986 214104
rect 674944 213874 674972 214095
rect 674760 213846 674972 213874
rect 674760 201362 674788 213846
rect 675220 210746 675248 217767
rect 675390 217016 675446 217025
rect 675390 216951 675392 216960
rect 675444 216951 675446 216960
rect 675392 216922 675444 216928
rect 675390 216200 675446 216209
rect 675390 216135 675392 216144
rect 675444 216135 675446 216144
rect 675392 216106 675444 216112
rect 675588 215294 675616 218991
rect 675758 218240 675814 218249
rect 675758 218175 675814 218184
rect 675588 215266 675708 215294
rect 675482 213752 675538 213761
rect 675482 213687 675484 213696
rect 675536 213687 675538 213696
rect 675484 213658 675536 213664
rect 675482 213344 675538 213353
rect 675482 213279 675484 213288
rect 675536 213279 675538 213288
rect 675484 213250 675536 213256
rect 675482 212120 675538 212129
rect 675482 212055 675484 212064
rect 675536 212055 675538 212064
rect 675484 212026 675536 212032
rect 674852 210718 675248 210746
rect 674852 202209 674880 210718
rect 675680 210610 675708 215266
rect 675036 210582 675708 210610
rect 675036 204049 675064 210582
rect 675772 210474 675800 218175
rect 676034 214976 676090 214985
rect 676034 214911 676090 214920
rect 676048 211449 676076 214911
rect 683118 212528 683174 212537
rect 683118 212463 683174 212472
rect 676034 211440 676090 211449
rect 676034 211375 676090 211384
rect 683132 211177 683160 212463
rect 683118 211168 683174 211177
rect 683118 211103 683174 211112
rect 675312 210446 675800 210474
rect 675312 205337 675340 210446
rect 675312 205309 675418 205337
rect 675758 205048 675814 205057
rect 675758 204983 675814 204992
rect 675772 204680 675800 204983
rect 675036 204021 675418 204049
rect 674852 202181 675418 202209
rect 675392 201884 675444 201890
rect 675392 201826 675444 201832
rect 675404 201620 675432 201826
rect 674760 201334 674880 201362
rect 674852 200938 674880 201334
rect 675208 201340 675260 201346
rect 675208 201282 675260 201288
rect 675220 201022 675248 201282
rect 675220 200994 675418 201022
rect 674840 200932 674892 200938
rect 674840 200874 674892 200880
rect 675300 200932 675352 200938
rect 675300 200874 675352 200880
rect 675024 200524 675076 200530
rect 675024 200466 675076 200472
rect 675036 196058 675064 200466
rect 675312 197282 675340 200874
rect 675772 200025 675800 200328
rect 675758 200016 675814 200025
rect 675758 199951 675814 199960
rect 675758 198384 675814 198393
rect 675758 198319 675814 198328
rect 675772 197880 675800 198319
rect 675404 197282 675432 197336
rect 675312 197254 675432 197282
rect 675758 197024 675814 197033
rect 675758 196959 675814 196968
rect 675772 196656 675800 196959
rect 675036 196030 675418 196058
rect 674668 195946 674788 195974
rect 674472 194540 674524 194546
rect 674472 194482 674524 194488
rect 674760 180794 674788 195946
rect 675128 194806 675418 194834
rect 675128 194546 675156 194806
rect 675116 194540 675168 194546
rect 675116 194482 675168 194488
rect 675114 193352 675170 193361
rect 675114 193287 675170 193296
rect 675128 191162 675156 193287
rect 675758 193216 675814 193225
rect 675758 193151 675814 193160
rect 675772 192984 675800 193151
rect 675666 192808 675722 192817
rect 675666 192743 675722 192752
rect 675680 192372 675708 192743
rect 675128 191134 675418 191162
rect 675850 190088 675906 190097
rect 675850 190023 675906 190032
rect 675864 189786 675892 190023
rect 675852 189780 675904 189786
rect 675852 189722 675904 189728
rect 683120 189780 683172 189786
rect 683120 189722 683172 189728
rect 674576 180766 674788 180794
rect 674576 175681 674604 180766
rect 675298 178528 675354 178537
rect 675298 178463 675354 178472
rect 675312 178090 675340 178463
rect 675484 178288 675536 178294
rect 675484 178230 675536 178236
rect 675496 178129 675524 178230
rect 675482 178120 675538 178129
rect 675300 178084 675352 178090
rect 675482 178055 675538 178064
rect 675300 178026 675352 178032
rect 683132 177721 683160 189722
rect 703694 179180 703722 179316
rect 704154 179180 704182 179316
rect 704614 179180 704642 179316
rect 705074 179180 705102 179316
rect 705534 179180 705562 179316
rect 705994 179180 706022 179316
rect 706454 179180 706482 179316
rect 706914 179180 706942 179316
rect 707374 179180 707402 179316
rect 707834 179180 707862 179316
rect 708294 179180 708322 179316
rect 708754 179180 708782 179316
rect 709214 179180 709242 179316
rect 683118 177712 683174 177721
rect 683118 177647 683174 177656
rect 675298 177304 675354 177313
rect 675298 177239 675354 177248
rect 675312 176866 675340 177239
rect 675482 176896 675538 176905
rect 675300 176860 675352 176866
rect 675482 176831 675538 176840
rect 675300 176802 675352 176808
rect 675496 176730 675524 176831
rect 675484 176724 675536 176730
rect 675484 176666 675536 176672
rect 674746 176080 674802 176089
rect 674746 176015 674802 176024
rect 674562 175672 674618 175681
rect 674562 175607 674618 175616
rect 674470 174448 674526 174457
rect 674470 174383 674526 174392
rect 674288 138440 674340 138446
rect 674288 138382 674340 138388
rect 673920 133000 673972 133006
rect 673920 132942 673972 132948
rect 673368 131300 673420 131306
rect 673368 131242 673420 131248
rect 674104 130892 674156 130898
rect 674104 130834 674156 130840
rect 673092 130280 673144 130286
rect 673092 130222 673144 130228
rect 673184 125996 673236 126002
rect 673184 125938 673236 125944
rect 672908 124160 672960 124166
rect 672908 124102 672960 124108
rect 673196 111790 673224 125938
rect 673920 124772 673972 124778
rect 673920 124714 673972 124720
rect 673368 123004 673420 123010
rect 673368 122946 673420 122952
rect 673184 111784 673236 111790
rect 673184 111726 673236 111732
rect 672724 111172 672776 111178
rect 672724 111114 672776 111120
rect 669228 107704 669280 107710
rect 669226 107672 669228 107681
rect 669280 107672 669282 107681
rect 669226 107607 669282 107616
rect 673380 106321 673408 122946
rect 673932 107030 673960 124714
rect 674116 107710 674144 130834
rect 674484 129713 674512 174383
rect 674760 157334 674788 176015
rect 675482 175264 675538 175273
rect 675482 175199 675484 175208
rect 675536 175199 675538 175208
rect 675484 175170 675536 175176
rect 675298 174040 675354 174049
rect 675298 173975 675354 173984
rect 675114 172816 675170 172825
rect 675114 172751 675170 172760
rect 675128 157334 675156 172751
rect 675312 166994 675340 173975
rect 675850 173224 675906 173233
rect 675850 173159 675906 173168
rect 675482 172000 675538 172009
rect 675482 171935 675484 171944
rect 675536 171935 675538 171944
rect 675484 171906 675536 171912
rect 675484 171216 675536 171222
rect 675482 171184 675484 171193
rect 675536 171184 675538 171193
rect 675482 171119 675538 171128
rect 675482 170368 675538 170377
rect 675482 170303 675484 170312
rect 675536 170303 675538 170312
rect 675484 170274 675536 170280
rect 675482 169144 675538 169153
rect 675482 169079 675484 169088
rect 675536 169079 675538 169088
rect 675484 169050 675536 169056
rect 675482 168736 675538 168745
rect 675482 168671 675484 168680
rect 675536 168671 675538 168680
rect 675484 168642 675536 168648
rect 675482 168328 675538 168337
rect 675482 168263 675484 168272
rect 675536 168263 675538 168272
rect 675484 168234 675536 168240
rect 675482 167920 675538 167929
rect 675482 167855 675484 167864
rect 675536 167855 675538 167864
rect 675484 167826 675536 167832
rect 675482 167104 675538 167113
rect 675482 167039 675538 167048
rect 675220 166966 675340 166994
rect 675220 159066 675248 166966
rect 675496 166954 675524 167039
rect 675864 166994 675892 173159
rect 678242 171592 678298 171601
rect 678242 171527 678298 171536
rect 676678 169960 676734 169969
rect 676678 169895 676734 169904
rect 675404 166938 675524 166954
rect 675392 166932 675524 166938
rect 675444 166926 675524 166932
rect 675588 166966 675892 166994
rect 675392 166874 675444 166880
rect 675588 163690 675616 166966
rect 676692 166433 676720 169895
rect 676678 166424 676734 166433
rect 676678 166359 676734 166368
rect 675312 163662 675616 163690
rect 675312 160290 675340 163662
rect 678256 162722 678284 171527
rect 675852 162716 675904 162722
rect 675852 162658 675904 162664
rect 678244 162716 678296 162722
rect 678244 162658 678296 162664
rect 675864 161401 675892 162658
rect 675850 161392 675906 161401
rect 675850 161327 675906 161336
rect 675404 160290 675432 160344
rect 675312 160262 675432 160290
rect 675574 160168 675630 160177
rect 675574 160103 675630 160112
rect 675588 159664 675616 160103
rect 675220 159038 675340 159066
rect 675312 158930 675340 159038
rect 675404 158930 675432 159052
rect 675312 158902 675432 158930
rect 674668 157306 674788 157334
rect 675036 157306 675156 157334
rect 674668 131345 674696 157306
rect 675036 157230 675064 157306
rect 675036 157202 675340 157230
rect 675312 157162 675340 157202
rect 675404 157162 675432 157216
rect 675312 157134 675432 157162
rect 675116 157004 675168 157010
rect 675116 156946 675168 156952
rect 675128 156657 675156 156946
rect 675128 156629 675418 156657
rect 675758 156496 675814 156505
rect 675758 156431 675814 156440
rect 675772 155992 675800 156431
rect 675758 155680 675814 155689
rect 675758 155615 675814 155624
rect 675772 155380 675800 155615
rect 675116 153196 675168 153202
rect 675116 153138 675168 153144
rect 675128 152334 675156 153138
rect 675666 153096 675722 153105
rect 675666 153031 675722 153040
rect 675680 152864 675708 153031
rect 675128 152306 675418 152334
rect 675116 151768 675168 151774
rect 675116 151710 675168 151716
rect 675128 151042 675156 151710
rect 675772 151473 675800 151675
rect 675758 151464 675814 151473
rect 675758 151399 675814 151408
rect 675128 151014 675418 151042
rect 675128 149821 675418 149849
rect 675128 147626 675156 149821
rect 675300 149048 675352 149054
rect 675300 148990 675352 148996
rect 675116 147620 675168 147626
rect 675116 147562 675168 147568
rect 675312 146690 675340 148990
rect 675758 148472 675814 148481
rect 675758 148407 675814 148416
rect 675772 147968 675800 148407
rect 675666 147656 675722 147665
rect 675666 147591 675722 147600
rect 675680 147356 675708 147591
rect 675312 146662 675432 146690
rect 675404 146132 675432 146662
rect 703694 133892 703722 134028
rect 704154 133892 704182 134028
rect 704614 133892 704642 134028
rect 705074 133892 705102 134028
rect 705534 133892 705562 134028
rect 705994 133892 706022 134028
rect 706454 133892 706482 134028
rect 706914 133892 706942 134028
rect 707374 133892 707402 134028
rect 707834 133892 707862 134028
rect 708294 133892 708322 134028
rect 708754 133892 708782 134028
rect 709214 133892 709242 134028
rect 675298 133376 675354 133385
rect 675298 133311 675354 133320
rect 675312 132530 675340 133311
rect 675484 133000 675536 133006
rect 675482 132968 675484 132977
rect 675536 132968 675538 132977
rect 675482 132903 675538 132912
rect 675484 132796 675536 132802
rect 675484 132738 675536 132744
rect 675496 132569 675524 132738
rect 675482 132560 675538 132569
rect 675300 132524 675352 132530
rect 675482 132495 675538 132504
rect 675300 132466 675352 132472
rect 675298 132152 675354 132161
rect 675298 132087 675354 132096
rect 674654 131336 674710 131345
rect 675312 131306 675340 132087
rect 675482 131744 675538 131753
rect 675482 131679 675538 131688
rect 674654 131271 674710 131280
rect 675300 131300 675352 131306
rect 675300 131242 675352 131248
rect 675496 131170 675524 131679
rect 675484 131164 675536 131170
rect 675484 131106 675536 131112
rect 675482 130928 675538 130937
rect 675482 130863 675484 130872
rect 675536 130863 675538 130872
rect 675484 130834 675536 130840
rect 675482 130520 675538 130529
rect 675482 130455 675538 130464
rect 675496 130286 675524 130455
rect 675484 130280 675536 130286
rect 675484 130222 675536 130228
rect 675482 130112 675538 130121
rect 675482 130047 675538 130056
rect 675496 129946 675524 130047
rect 675484 129940 675536 129946
rect 675484 129882 675536 129888
rect 674470 129704 674526 129713
rect 674470 129639 674526 129648
rect 675482 129296 675538 129305
rect 675482 129231 675538 129240
rect 675496 128382 675524 129231
rect 675484 128376 675536 128382
rect 675484 128318 675536 128324
rect 679622 127800 679678 127809
rect 679622 127735 679678 127744
rect 674838 127664 674894 127673
rect 674838 127599 674894 127608
rect 674378 125216 674434 125225
rect 674378 125151 674434 125160
rect 674104 107704 674156 107710
rect 674104 107646 674156 107652
rect 673920 107024 673972 107030
rect 673920 106966 673972 106972
rect 673366 106312 673422 106321
rect 673366 106247 673422 106256
rect 669056 106134 669176 106162
rect 668950 106040 669006 106049
rect 668950 105975 669006 105984
rect 669148 104553 669176 106134
rect 674392 104666 674420 125151
rect 674654 123584 674710 123593
rect 674654 123519 674710 123528
rect 674668 105822 674696 123519
rect 674852 112010 674880 127599
rect 675022 126440 675078 126449
rect 675022 126375 675078 126384
rect 675036 114493 675064 126375
rect 675482 126032 675538 126041
rect 675482 125967 675484 125976
rect 675536 125967 675538 125976
rect 675484 125938 675536 125944
rect 675484 125656 675536 125662
rect 675482 125624 675484 125633
rect 675536 125624 675538 125633
rect 675482 125559 675538 125568
rect 675482 124808 675538 124817
rect 675482 124743 675484 124752
rect 675536 124743 675538 124752
rect 675484 124714 675536 124720
rect 675298 123992 675354 124001
rect 675298 123927 675354 123936
rect 675312 123010 675340 123927
rect 675482 123176 675538 123185
rect 675482 123111 675538 123120
rect 675300 123004 675352 123010
rect 675300 122946 675352 122952
rect 675496 122874 675524 123111
rect 675484 122868 675536 122874
rect 675484 122810 675536 122816
rect 675298 122496 675354 122505
rect 675298 122431 675354 122440
rect 675312 121514 675340 122431
rect 677598 122088 677654 122097
rect 677598 122023 677654 122032
rect 675482 121952 675538 121961
rect 675482 121887 675538 121896
rect 675300 121508 675352 121514
rect 675300 121450 675352 121456
rect 675496 120766 675524 121887
rect 675484 120760 675536 120766
rect 675484 120702 675536 120708
rect 675852 117292 675904 117298
rect 675852 117234 675904 117240
rect 675864 117178 675892 117234
rect 675312 117150 675892 117178
rect 675312 115138 675340 117150
rect 677612 117065 677640 122023
rect 679636 117298 679664 127735
rect 683118 126576 683174 126585
rect 683118 126511 683174 126520
rect 683132 124545 683160 126511
rect 683118 124536 683174 124545
rect 683118 124471 683174 124480
rect 683118 124128 683174 124137
rect 683118 124063 683174 124072
rect 683132 117337 683160 124063
rect 683118 117328 683174 117337
rect 679624 117292 679676 117298
rect 683118 117263 683174 117272
rect 679624 117234 679676 117240
rect 677598 117056 677654 117065
rect 677598 116991 677654 117000
rect 675312 115110 675418 115138
rect 675036 114465 675418 114493
rect 675312 113818 675418 113846
rect 675312 113121 675340 113818
rect 675298 113112 675354 113121
rect 675298 113047 675354 113056
rect 674852 111982 675418 112010
rect 675116 111784 675168 111790
rect 675116 111726 675168 111732
rect 675128 111466 675156 111726
rect 675128 111438 675418 111466
rect 675392 111172 675444 111178
rect 675392 111114 675444 111120
rect 675404 110772 675432 111114
rect 675758 110392 675814 110401
rect 675758 110327 675814 110336
rect 675772 110160 675800 110327
rect 675666 108080 675722 108089
rect 675666 108015 675722 108024
rect 675680 107644 675708 108015
rect 675312 107222 675432 107250
rect 675312 107114 675340 107222
rect 675128 107086 675340 107114
rect 675404 107100 675432 107222
rect 675128 106321 675156 107086
rect 675300 107024 675352 107030
rect 675300 106966 675352 106972
rect 675312 106502 675340 106966
rect 675312 106474 675418 106502
rect 675114 106312 675170 106321
rect 675114 106247 675170 106256
rect 675312 105862 675432 105890
rect 675312 105822 675340 105862
rect 674668 105794 675340 105822
rect 675404 105808 675432 105862
rect 674392 104638 675340 104666
rect 669134 104544 669190 104553
rect 675312 104530 675340 104638
rect 675404 104530 675432 104652
rect 675312 104502 675432 104530
rect 669134 104479 669190 104488
rect 675758 103184 675814 103193
rect 675758 103119 675814 103128
rect 668582 102912 668638 102921
rect 668582 102847 668638 102856
rect 675772 102816 675800 103119
rect 675666 102640 675722 102649
rect 675666 102575 675722 102584
rect 675680 102136 675708 102575
rect 675758 101416 675814 101425
rect 675758 101351 675814 101360
rect 675772 100980 675800 101351
rect 595272 100014 595608 100042
rect 596192 100014 596344 100042
rect 596560 100014 597080 100042
rect 597572 100014 597816 100042
rect 598032 100014 598552 100042
rect 598952 100014 599288 100042
rect 599504 100014 600024 100042
rect 600424 100014 600760 100042
rect 600884 100014 601496 100042
rect 601896 100014 602232 100042
rect 602632 100014 602968 100042
rect 603092 100014 603704 100042
rect 594064 97980 594116 97986
rect 594064 97922 594116 97928
rect 592684 97844 592736 97850
rect 592684 97786 592736 97792
rect 591304 97300 591356 97306
rect 591304 97242 591356 97248
rect 590108 96076 590160 96082
rect 590108 96018 590160 96024
rect 589924 74520 589976 74526
rect 589924 74462 589976 74468
rect 588544 55208 588596 55214
rect 588544 55150 588596 55156
rect 591316 53145 591344 97242
rect 591302 53136 591358 53145
rect 584588 53100 584640 53106
rect 591302 53071 591358 53080
rect 584588 53042 584640 53048
rect 577504 52488 577556 52494
rect 577504 52430 577556 52436
rect 497554 50552 497610 50561
rect 445208 50516 445260 50522
rect 549258 50552 549314 50561
rect 497554 50487 497610 50496
rect 498108 50516 498160 50522
rect 445208 50458 445260 50464
rect 549258 50487 549314 50496
rect 498108 50458 498160 50464
rect 445024 50380 445076 50386
rect 445024 50322 445076 50328
rect 445036 45121 445064 50322
rect 498120 47326 498148 50458
rect 498108 47320 498160 47326
rect 498108 47262 498160 47268
rect 499580 47320 499632 47326
rect 499580 47262 499632 47268
rect 499592 47025 499620 47262
rect 499578 47016 499634 47025
rect 499578 46951 499634 46960
rect 592696 46481 592724 97786
rect 594076 47841 594104 97922
rect 595272 97714 595300 100014
rect 596192 97986 596220 100014
rect 596180 97980 596232 97986
rect 596180 97922 596232 97928
rect 595260 97708 595312 97714
rect 595260 97650 595312 97656
rect 595628 97708 595680 97714
rect 595628 97650 595680 97656
rect 595444 97572 595496 97578
rect 595444 97514 595496 97520
rect 595456 51746 595484 97514
rect 595640 80714 595668 97650
rect 596560 84194 596588 100014
rect 597572 97850 597600 100014
rect 597560 97844 597612 97850
rect 597560 97786 597612 97792
rect 598032 84194 598060 100014
rect 598952 97578 598980 100014
rect 598940 97572 598992 97578
rect 598940 97514 598992 97520
rect 599504 84194 599532 100014
rect 600424 97306 600452 100014
rect 600412 97300 600464 97306
rect 600412 97242 600464 97248
rect 600884 84194 600912 100014
rect 601700 96960 601752 96966
rect 601700 96902 601752 96908
rect 596192 84166 596588 84194
rect 597572 84166 598060 84194
rect 598952 84166 599532 84194
rect 600332 84166 600912 84194
rect 595628 80708 595680 80714
rect 595628 80650 595680 80656
rect 595444 51740 595496 51746
rect 595444 51682 595496 51688
rect 596192 48929 596220 84166
rect 596178 48920 596234 48929
rect 596178 48855 596234 48864
rect 594062 47832 594118 47841
rect 594062 47767 594118 47776
rect 592682 46472 592738 46481
rect 592682 46407 592738 46416
rect 597572 46209 597600 84166
rect 598952 48113 598980 84166
rect 600332 49201 600360 84166
rect 600318 49192 600374 49201
rect 600318 49127 600374 49136
rect 598938 48104 598994 48113
rect 598938 48039 598994 48048
rect 597558 46200 597614 46209
rect 597558 46135 597614 46144
rect 445022 45112 445078 45121
rect 445022 45047 445078 45056
rect 601712 44849 601740 96902
rect 601896 50289 601924 100014
rect 602632 96966 602660 100014
rect 602620 96960 602672 96966
rect 602620 96902 602672 96908
rect 603092 51785 603120 100014
rect 604426 99770 604454 100028
rect 605176 100014 605512 100042
rect 605912 100014 606248 100042
rect 606648 100014 607168 100042
rect 607384 100014 607720 100042
rect 608120 100014 608456 100042
rect 608856 100014 609192 100042
rect 609592 100014 609928 100042
rect 610328 100014 610664 100042
rect 611064 100014 611308 100042
rect 611800 100014 612136 100042
rect 612536 100014 612688 100042
rect 613272 100014 613608 100042
rect 604426 99742 604500 99770
rect 603078 51776 603134 51785
rect 603078 51711 603134 51720
rect 601882 50280 601938 50289
rect 601882 50215 601938 50224
rect 601698 44840 601754 44849
rect 601698 44775 601754 44784
rect 604472 43489 604500 99742
rect 605484 97306 605512 100014
rect 605472 97300 605524 97306
rect 605472 97242 605524 97248
rect 606220 96966 606248 100014
rect 606208 96960 606260 96966
rect 606208 96902 606260 96908
rect 606944 96960 606996 96966
rect 606944 96902 606996 96908
rect 606956 93854 606984 96902
rect 607140 96506 607168 100014
rect 607140 96478 607352 96506
rect 606956 93826 607168 93854
rect 607140 75206 607168 93826
rect 607324 88330 607352 96478
rect 607692 94518 607720 100014
rect 608428 95946 608456 100014
rect 609164 96898 609192 100014
rect 609152 96892 609204 96898
rect 609152 96834 609204 96840
rect 609704 96892 609756 96898
rect 609704 96834 609756 96840
rect 608416 95940 608468 95946
rect 608416 95882 608468 95888
rect 607680 94512 607732 94518
rect 607680 94454 607732 94460
rect 609716 93158 609744 96834
rect 609704 93152 609756 93158
rect 609704 93094 609756 93100
rect 607312 88324 607364 88330
rect 607312 88266 607364 88272
rect 609900 85542 609928 100014
rect 610636 96082 610664 100014
rect 610624 96076 610676 96082
rect 610624 96018 610676 96024
rect 611280 91050 611308 100014
rect 611912 97300 611964 97306
rect 611912 97242 611964 97248
rect 611924 93854 611952 97242
rect 612108 96898 612136 100014
rect 612660 97034 612688 100014
rect 612648 97028 612700 97034
rect 612648 96970 612700 96976
rect 613384 97028 613436 97034
rect 613384 96970 613436 96976
rect 612096 96892 612148 96898
rect 612096 96834 612148 96840
rect 612648 96892 612700 96898
rect 612648 96834 612700 96840
rect 611924 93826 612044 93854
rect 611268 91044 611320 91050
rect 611268 90986 611320 90992
rect 609888 85536 609940 85542
rect 609888 85478 609940 85484
rect 607128 75200 607180 75206
rect 607128 75142 607180 75148
rect 612016 57254 612044 93826
rect 612660 80850 612688 96834
rect 612648 80844 612700 80850
rect 612648 80786 612700 80792
rect 613396 76566 613424 96970
rect 613580 96830 613608 100014
rect 613994 99770 614022 100028
rect 614744 100014 615080 100042
rect 615480 100014 615816 100042
rect 616216 100014 616552 100042
rect 616952 100014 617288 100042
rect 617688 100014 618116 100042
rect 618424 100014 618760 100042
rect 619160 100014 619588 100042
rect 619896 100014 620232 100042
rect 620632 100014 620968 100042
rect 621368 100014 621704 100042
rect 622104 100014 622348 100042
rect 622840 100014 623176 100042
rect 623576 100014 623728 100042
rect 624312 100014 624648 100042
rect 613994 99742 614068 99770
rect 614040 96966 614068 99742
rect 614028 96960 614080 96966
rect 614028 96902 614080 96908
rect 614764 96960 614816 96966
rect 614764 96902 614816 96908
rect 613568 96824 613620 96830
rect 613568 96766 613620 96772
rect 614028 96824 614080 96830
rect 614028 96766 614080 96772
rect 614040 77994 614068 96766
rect 614028 77988 614080 77994
rect 614028 77930 614080 77936
rect 614776 76702 614804 96902
rect 615052 93854 615080 100014
rect 615788 96966 615816 100014
rect 615776 96960 615828 96966
rect 615776 96902 615828 96908
rect 616524 95198 616552 100014
rect 617260 96966 617288 100014
rect 616788 96960 616840 96966
rect 616788 96902 616840 96908
rect 617248 96960 617300 96966
rect 617248 96902 617300 96908
rect 617892 96960 617944 96966
rect 617892 96902 617944 96908
rect 616512 95192 616564 95198
rect 616512 95134 616564 95140
rect 615052 93826 615448 93854
rect 614764 76696 614816 76702
rect 614764 76638 614816 76644
rect 613384 76560 613436 76566
rect 613384 76502 613436 76508
rect 615420 75342 615448 93826
rect 616800 79354 616828 96902
rect 617904 91050 617932 96902
rect 618088 92478 618116 100014
rect 618732 96898 618760 100014
rect 618720 96892 618772 96898
rect 618720 96834 618772 96840
rect 619560 93838 619588 100014
rect 620204 97986 620232 100014
rect 620192 97980 620244 97986
rect 620192 97922 620244 97928
rect 620940 96286 620968 100014
rect 621676 98802 621704 100014
rect 621664 98796 621716 98802
rect 621664 98738 621716 98744
rect 622320 98666 622348 100014
rect 622308 98660 622360 98666
rect 622308 98602 622360 98608
rect 623148 97714 623176 100014
rect 623700 99074 623728 100014
rect 623688 99068 623740 99074
rect 623688 99010 623740 99016
rect 623136 97708 623188 97714
rect 623136 97650 623188 97656
rect 624620 97578 624648 100014
rect 625034 99770 625062 100028
rect 625784 100014 625936 100042
rect 626520 100014 626856 100042
rect 627256 100014 627592 100042
rect 627992 100014 628236 100042
rect 628728 100014 629064 100042
rect 629464 100014 629800 100042
rect 630200 100014 630536 100042
rect 630936 100014 631272 100042
rect 631672 100014 631916 100042
rect 632408 100014 632744 100042
rect 633144 100014 633388 100042
rect 633880 100014 634216 100042
rect 634616 100014 634768 100042
rect 635352 100014 635688 100042
rect 625034 99742 625108 99770
rect 625080 99210 625108 99742
rect 625068 99204 625120 99210
rect 625068 99146 625120 99152
rect 625908 97850 625936 100014
rect 626828 97986 626856 100014
rect 626080 97980 626132 97986
rect 626080 97922 626132 97928
rect 626816 97980 626868 97986
rect 626816 97922 626868 97928
rect 625896 97844 625948 97850
rect 625896 97786 625948 97792
rect 624608 97572 624660 97578
rect 624608 97514 624660 97520
rect 620928 96280 620980 96286
rect 620928 96222 620980 96228
rect 621664 96076 621716 96082
rect 621664 96018 621716 96024
rect 620284 95940 620336 95946
rect 620284 95882 620336 95888
rect 619548 93832 619600 93838
rect 619548 93774 619600 93780
rect 618904 93152 618956 93158
rect 618904 93094 618956 93100
rect 618076 92472 618128 92478
rect 618076 92414 618128 92420
rect 617340 91044 617392 91050
rect 617340 90986 617392 90992
rect 617892 91044 617944 91050
rect 617892 90986 617944 90992
rect 617352 88194 617380 90986
rect 617340 88188 617392 88194
rect 617340 88130 617392 88136
rect 618916 84046 618944 93094
rect 620296 84182 620324 95882
rect 621676 86290 621704 96018
rect 622676 95192 622728 95198
rect 622676 95134 622728 95140
rect 622688 89690 622716 95134
rect 624976 94512 625028 94518
rect 626092 94489 626120 97922
rect 627564 97442 627592 100014
rect 627552 97436 627604 97442
rect 627552 97378 627604 97384
rect 628208 97306 628236 100014
rect 629036 98802 629064 100014
rect 629772 98938 629800 100014
rect 629760 98932 629812 98938
rect 629760 98874 629812 98880
rect 628380 98796 628432 98802
rect 628380 98738 628432 98744
rect 629024 98796 629076 98802
rect 629024 98738 629076 98744
rect 628196 97300 628248 97306
rect 628196 97242 628248 97248
rect 626264 96892 626316 96898
rect 626264 96834 626316 96840
rect 624976 94454 625028 94460
rect 626078 94480 626134 94489
rect 622676 89684 622728 89690
rect 622676 89626 622728 89632
rect 624988 88641 625016 94454
rect 626078 94415 626134 94424
rect 626276 92585 626304 96834
rect 626448 96280 626500 96286
rect 626448 96222 626500 96228
rect 626460 95441 626488 96222
rect 628392 95826 628420 98738
rect 630508 98666 630536 100014
rect 629484 98660 629536 98666
rect 629484 98602 629536 98608
rect 630496 98660 630548 98666
rect 630496 98602 630548 98608
rect 629496 95826 629524 98602
rect 630680 97708 630732 97714
rect 630680 97650 630732 97656
rect 630692 95826 630720 97650
rect 631244 96354 631272 100014
rect 631232 96348 631284 96354
rect 631232 96290 631284 96296
rect 631888 96218 631916 100014
rect 632152 99068 632204 99074
rect 632152 99010 632204 99016
rect 631876 96212 631928 96218
rect 631876 96154 631928 96160
rect 632164 95826 632192 99010
rect 632716 97714 632744 100014
rect 633360 97714 633388 100014
rect 632704 97708 632756 97714
rect 632704 97650 632756 97656
rect 633348 97708 633400 97714
rect 633348 97650 633400 97656
rect 632980 97572 633032 97578
rect 632980 97514 633032 97520
rect 628392 95798 628728 95826
rect 629496 95798 629832 95826
rect 630692 95798 631028 95826
rect 632132 95798 632192 95826
rect 632992 95826 633020 97514
rect 634188 97170 634216 100014
rect 634452 99204 634504 99210
rect 634452 99146 634504 99152
rect 634176 97164 634228 97170
rect 634176 97106 634228 97112
rect 634464 95826 634492 99146
rect 632992 95798 633328 95826
rect 634432 95798 634492 95826
rect 634740 95674 634768 100014
rect 635280 97844 635332 97850
rect 635280 97786 635332 97792
rect 635292 95826 635320 97786
rect 635660 96626 635688 100014
rect 635936 100014 636088 100042
rect 636824 100014 637068 100042
rect 637560 100014 637896 100042
rect 638296 100014 638632 100042
rect 639032 100014 639368 100042
rect 639768 100014 640104 100042
rect 640504 100014 640840 100042
rect 641240 100014 641576 100042
rect 641976 100014 642312 100042
rect 642712 100014 643048 100042
rect 643448 100014 643784 100042
rect 644184 100014 644336 100042
rect 644920 100014 645256 100042
rect 635648 96620 635700 96626
rect 635648 96562 635700 96568
rect 635292 95798 635628 95826
rect 635936 95713 635964 100014
rect 636384 97980 636436 97986
rect 636384 97922 636436 97928
rect 636396 95826 636424 97922
rect 637040 96937 637068 100014
rect 637580 97436 637632 97442
rect 637580 97378 637632 97384
rect 637026 96928 637082 96937
rect 637026 96863 637082 96872
rect 637592 95826 637620 97378
rect 637868 96082 637896 100014
rect 638604 96490 638632 100014
rect 639340 97442 639368 100014
rect 639328 97436 639380 97442
rect 639328 97378 639380 97384
rect 639052 97300 639104 97306
rect 639052 97242 639104 97248
rect 638592 96484 638644 96490
rect 638592 96426 638644 96432
rect 637856 96076 637908 96082
rect 637856 96018 637908 96024
rect 639064 95826 639092 97242
rect 636396 95798 636732 95826
rect 637592 95798 637928 95826
rect 639032 95798 639092 95826
rect 640076 95810 640104 100014
rect 640248 98796 640300 98802
rect 640248 98738 640300 98744
rect 640260 95826 640288 98738
rect 640812 95946 640840 100014
rect 640984 98932 641036 98938
rect 640984 98874 641036 98880
rect 640800 95940 640852 95946
rect 640800 95882 640852 95888
rect 640064 95804 640116 95810
rect 640228 95798 640288 95826
rect 640996 95826 641024 98874
rect 641548 97306 641576 100014
rect 642088 98660 642140 98666
rect 642088 98602 642140 98608
rect 641536 97300 641588 97306
rect 641536 97242 641588 97248
rect 640996 95798 641332 95826
rect 640064 95746 640116 95752
rect 635922 95704 635978 95713
rect 634728 95668 634780 95674
rect 642100 95690 642128 98602
rect 642284 96626 642312 100014
rect 643020 97850 643048 100014
rect 643008 97844 643060 97850
rect 643008 97786 643060 97792
rect 643008 97300 643060 97306
rect 643008 97242 643060 97248
rect 642824 96756 642876 96762
rect 642824 96698 642876 96704
rect 642272 96620 642324 96626
rect 642272 96562 642324 96568
rect 642836 96354 642864 96698
rect 642640 96348 642692 96354
rect 642640 96290 642692 96296
rect 642824 96348 642876 96354
rect 642824 96290 642876 96296
rect 642100 95662 642528 95690
rect 635922 95639 635978 95648
rect 634728 95610 634780 95616
rect 626446 95432 626502 95441
rect 626446 95367 626502 95376
rect 642652 95169 642680 96290
rect 643020 95826 643048 97242
rect 643468 97164 643520 97170
rect 643468 97106 643520 97112
rect 643284 96620 643336 96626
rect 643284 96562 643336 96568
rect 642928 95798 643048 95826
rect 642638 95160 642694 95169
rect 642638 95095 642694 95104
rect 642928 94518 642956 95798
rect 643100 95668 643152 95674
rect 643100 95610 643152 95616
rect 642916 94512 642968 94518
rect 642916 94454 642968 94460
rect 626448 93832 626500 93838
rect 626448 93774 626500 93780
rect 626460 93537 626488 93774
rect 626446 93528 626502 93537
rect 626446 93463 626502 93472
rect 626262 92576 626318 92585
rect 626262 92511 626318 92520
rect 625436 92472 625488 92478
rect 625436 92414 625488 92420
rect 625448 91633 625476 92414
rect 625434 91624 625490 91633
rect 625434 91559 625490 91568
rect 626448 91044 626500 91050
rect 626448 90986 626500 90992
rect 626460 90681 626488 90986
rect 626446 90672 626502 90681
rect 626446 90607 626502 90616
rect 626446 89720 626502 89729
rect 626446 89655 626448 89664
rect 626500 89655 626502 89664
rect 626448 89626 626500 89632
rect 624974 88632 625030 88641
rect 624974 88567 625030 88576
rect 626448 88324 626500 88330
rect 626448 88266 626500 88272
rect 625620 88188 625672 88194
rect 625620 88130 625672 88136
rect 625632 87009 625660 88130
rect 626460 87961 626488 88266
rect 626446 87952 626502 87961
rect 626446 87887 626502 87896
rect 625618 87000 625674 87009
rect 625618 86935 625674 86944
rect 621664 86284 621716 86290
rect 621664 86226 621716 86232
rect 626448 86284 626500 86290
rect 626448 86226 626500 86232
rect 626460 86057 626488 86226
rect 626446 86048 626502 86057
rect 626446 85983 626502 85992
rect 626448 85536 626500 85542
rect 626448 85478 626500 85484
rect 626460 85105 626488 85478
rect 626446 85096 626502 85105
rect 626446 85031 626502 85040
rect 620284 84176 620336 84182
rect 620284 84118 620336 84124
rect 626264 84176 626316 84182
rect 626264 84118 626316 84124
rect 626446 84144 626502 84153
rect 618904 84040 618956 84046
rect 618904 83982 618956 83988
rect 626276 83201 626304 84118
rect 626446 84079 626502 84088
rect 626460 83978 626488 84079
rect 626448 83972 626500 83978
rect 626448 83914 626500 83920
rect 626262 83192 626318 83201
rect 626262 83127 626318 83136
rect 643112 82793 643140 95610
rect 643296 93838 643324 96562
rect 643284 93832 643336 93838
rect 643284 93774 643336 93780
rect 643480 84697 643508 97106
rect 643756 94654 643784 100014
rect 643928 97708 643980 97714
rect 643928 97650 643980 97656
rect 643744 94648 643796 94654
rect 643744 94590 643796 94596
rect 643940 87145 643968 97650
rect 644308 97306 644336 100014
rect 644756 97572 644808 97578
rect 644756 97514 644808 97520
rect 644296 97300 644348 97306
rect 644296 97242 644348 97248
rect 644480 96212 644532 96218
rect 644480 96154 644532 96160
rect 644492 92177 644520 96154
rect 644478 92168 644534 92177
rect 644478 92103 644534 92112
rect 644768 89729 644796 97514
rect 645228 96762 645256 100014
rect 645642 99770 645670 100028
rect 646392 100014 646728 100042
rect 645596 99742 645670 99770
rect 645216 96756 645268 96762
rect 645216 96698 645268 96704
rect 645596 95674 645624 99742
rect 646504 97436 646556 97442
rect 646504 97378 646556 97384
rect 645768 96756 645820 96762
rect 645768 96698 645820 96704
rect 645584 95668 645636 95674
rect 645584 95610 645636 95616
rect 644754 89720 644810 89729
rect 644754 89655 644810 89664
rect 645780 87174 645808 96698
rect 646516 91050 646544 97378
rect 646700 96966 646728 100014
rect 647114 99770 647142 100028
rect 647864 100014 648384 100042
rect 647114 99742 647188 99770
rect 647160 97850 647188 99742
rect 647148 97844 647200 97850
rect 647148 97786 647200 97792
rect 646688 96960 646740 96966
rect 646688 96902 646740 96908
rect 647148 96960 647200 96966
rect 647148 96902 647200 96908
rect 646504 91044 646556 91050
rect 646504 90986 646556 90992
rect 647160 89010 647188 96902
rect 647148 89004 647200 89010
rect 647148 88946 647200 88952
rect 645768 87168 645820 87174
rect 643926 87136 643982 87145
rect 645768 87110 645820 87116
rect 643926 87071 643982 87080
rect 648356 87038 648384 100014
rect 648586 99770 648614 100028
rect 649336 100014 649672 100042
rect 650072 100014 650408 100042
rect 650808 100014 651144 100042
rect 651544 100014 651880 100042
rect 652280 100014 652616 100042
rect 653016 100014 653352 100042
rect 653752 100014 653996 100042
rect 654488 100014 654824 100042
rect 655224 100014 655468 100042
rect 648586 99742 648660 99770
rect 648632 96218 648660 99742
rect 648804 96348 648856 96354
rect 648804 96290 648856 96296
rect 648620 96212 648672 96218
rect 648620 96154 648672 96160
rect 648344 87032 648396 87038
rect 648344 86974 648396 86980
rect 643466 84688 643522 84697
rect 643466 84623 643522 84632
rect 643098 82784 643154 82793
rect 643098 82719 643154 82728
rect 628562 81696 628618 81705
rect 628562 81631 628618 81640
rect 628576 80986 628604 81631
rect 628564 80980 628616 80986
rect 628564 80922 628616 80928
rect 631520 80974 631856 81002
rect 638972 80974 639308 81002
rect 642456 80980 642508 80986
rect 629206 80880 629262 80889
rect 629206 80815 629262 80824
rect 629220 79490 629248 80815
rect 629208 79484 629260 79490
rect 629208 79426 629260 79432
rect 616788 79348 616840 79354
rect 616788 79290 616840 79296
rect 631048 78124 631100 78130
rect 631048 78066 631100 78072
rect 631060 77722 631088 78066
rect 631048 77716 631100 77722
rect 631048 77658 631100 77664
rect 628288 77580 628340 77586
rect 628288 77522 628340 77528
rect 624424 77444 624476 77450
rect 624424 77386 624476 77392
rect 625804 77444 625856 77450
rect 625804 77386 625856 77392
rect 615408 75336 615460 75342
rect 615408 75278 615460 75284
rect 612004 57248 612056 57254
rect 612004 57190 612056 57196
rect 624436 47569 624464 77386
rect 625816 52358 625844 77386
rect 628300 75954 628328 77522
rect 628288 75948 628340 75954
rect 628288 75890 628340 75896
rect 628300 75290 628328 75890
rect 631060 75290 631088 77658
rect 631520 77586 631548 80974
rect 636108 80708 636160 80714
rect 636108 80650 636160 80656
rect 633898 77752 633954 77761
rect 633898 77687 633954 77696
rect 631508 77580 631560 77586
rect 631508 77522 631560 77528
rect 633912 77450 633940 77687
rect 633900 77444 633952 77450
rect 633900 77386 633952 77392
rect 633912 75290 633940 77386
rect 636120 77294 636148 80650
rect 637488 79484 637540 79490
rect 637488 79426 637540 79432
rect 637118 78568 637174 78577
rect 637118 78503 637174 78512
rect 637132 77314 637160 78503
rect 637500 78266 637528 79426
rect 637488 78260 637540 78266
rect 637488 78202 637540 78208
rect 638972 78130 639000 80974
rect 642456 80922 642508 80928
rect 638960 78124 639012 78130
rect 638960 78066 639012 78072
rect 637120 77308 637172 77314
rect 636120 77266 636332 77294
rect 628176 75262 628328 75290
rect 631028 75262 631088 75290
rect 633880 75262 633940 75290
rect 636304 75154 636332 77266
rect 637120 77250 637172 77256
rect 639604 77308 639656 77314
rect 639604 77250 639656 77256
rect 639616 75290 639644 77250
rect 642468 75290 642496 80922
rect 645860 80844 645912 80850
rect 645860 80786 645912 80792
rect 645308 78260 645360 78266
rect 645308 78202 645360 78208
rect 645320 75290 645348 78202
rect 639584 75262 639644 75290
rect 642436 75262 642496 75290
rect 645288 75262 645348 75290
rect 636304 75126 636732 75154
rect 645872 66042 645900 80786
rect 647424 79348 647476 79354
rect 647424 79290 647476 79296
rect 646320 76696 646372 76702
rect 646320 76638 646372 76644
rect 646136 75336 646188 75342
rect 646136 75278 646188 75284
rect 646148 71777 646176 75278
rect 646134 71768 646190 71777
rect 646134 71703 646190 71712
rect 646332 70417 646360 76638
rect 646872 75200 646924 75206
rect 646872 75142 646924 75148
rect 646884 74497 646912 75142
rect 646870 74488 646926 74497
rect 646870 74423 646926 74432
rect 647436 73001 647464 79290
rect 647608 77988 647660 77994
rect 647608 77930 647660 77936
rect 647422 72992 647478 73001
rect 647422 72927 647478 72936
rect 646318 70408 646374 70417
rect 646318 70343 646374 70352
rect 647620 68513 647648 77930
rect 647606 68504 647662 68513
rect 647606 68439 647662 68448
rect 646134 66056 646190 66065
rect 645872 66014 646134 66042
rect 646134 65991 646190 66000
rect 648816 64025 648844 96290
rect 649644 94042 649672 100014
rect 650380 96966 650408 100014
rect 650368 96960 650420 96966
rect 650368 96902 650420 96908
rect 651116 96694 651144 100014
rect 651852 96830 651880 100014
rect 651840 96824 651892 96830
rect 651840 96766 651892 96772
rect 651104 96688 651156 96694
rect 651104 96630 651156 96636
rect 650920 96620 650972 96626
rect 650920 96562 650972 96568
rect 649632 94036 649684 94042
rect 649632 93978 649684 93984
rect 650644 94036 650696 94042
rect 650644 93978 650696 93984
rect 650656 86494 650684 93978
rect 650932 92478 650960 96562
rect 652588 96354 652616 100014
rect 653324 96490 653352 100014
rect 653312 96484 653364 96490
rect 653312 96426 653364 96432
rect 652576 96348 652628 96354
rect 652576 96290 652628 96296
rect 652024 95804 652076 95810
rect 652024 95746 652076 95752
rect 650920 92472 650972 92478
rect 650920 92414 650972 92420
rect 652036 86630 652064 95746
rect 653404 94648 653456 94654
rect 653404 94590 653456 94596
rect 653416 86766 653444 94590
rect 653968 94217 653996 100014
rect 654796 97238 654824 100014
rect 655440 97714 655468 100014
rect 655808 100014 655960 100042
rect 656696 100014 656848 100042
rect 657432 100014 657768 100042
rect 655428 97708 655480 97714
rect 655428 97650 655480 97656
rect 654784 97232 654836 97238
rect 654784 97174 654836 97180
rect 655244 97232 655296 97238
rect 655244 97174 655296 97180
rect 654324 96688 654376 96694
rect 654324 96630 654376 96636
rect 653954 94208 654010 94217
rect 653954 94143 654010 94152
rect 654140 93764 654192 93770
rect 654140 93706 654192 93712
rect 654152 92585 654180 93706
rect 654336 93401 654364 96630
rect 654322 93392 654378 93401
rect 654322 93327 654378 93336
rect 654138 92576 654194 92585
rect 654138 92511 654194 92520
rect 654324 92472 654376 92478
rect 654324 92414 654376 92420
rect 654336 91497 654364 92414
rect 654322 91488 654378 91497
rect 654322 91423 654378 91432
rect 654140 91044 654192 91050
rect 654140 90986 654192 90992
rect 654152 90681 654180 90986
rect 654138 90672 654194 90681
rect 654138 90607 654194 90616
rect 655256 88330 655284 97174
rect 655808 89865 655836 100014
rect 656820 97306 656848 100014
rect 656808 97300 656860 97306
rect 656808 97242 656860 97248
rect 656716 97096 656768 97102
rect 656716 97038 656768 97044
rect 656164 95668 656216 95674
rect 656164 95610 656216 95616
rect 655794 89856 655850 89865
rect 655794 89791 655850 89800
rect 656176 88806 656204 95610
rect 656164 88800 656216 88806
rect 656164 88742 656216 88748
rect 655244 88324 655296 88330
rect 655244 88266 655296 88272
rect 656532 87304 656584 87310
rect 656532 87246 656584 87252
rect 656544 87038 656572 87246
rect 656532 87032 656584 87038
rect 656532 86974 656584 86980
rect 656728 86970 656756 97038
rect 657740 95132 657768 100014
rect 658154 99770 658182 100028
rect 658904 100014 659240 100042
rect 659640 100014 659976 100042
rect 658154 99742 658228 99770
rect 658200 97442 658228 99742
rect 658832 97572 658884 97578
rect 658832 97514 658884 97520
rect 658188 97436 658240 97442
rect 658188 97378 658240 97384
rect 658280 96960 658332 96966
rect 658280 96902 658332 96908
rect 658292 95132 658320 96902
rect 658844 95132 658872 97514
rect 659212 95674 659240 100014
rect 659948 97986 659976 100014
rect 660132 100014 660376 100042
rect 659752 97980 659804 97986
rect 659752 97922 659804 97928
rect 659936 97980 659988 97986
rect 659936 97922 659988 97928
rect 659568 96824 659620 96830
rect 659568 96766 659620 96772
rect 659200 95668 659252 95674
rect 659200 95610 659252 95616
rect 659580 95132 659608 96766
rect 659764 95146 659792 97922
rect 660132 96966 660160 100014
rect 665732 97980 665784 97986
rect 665732 97922 665784 97928
rect 661960 97844 662012 97850
rect 661960 97786 662012 97792
rect 661408 97300 661460 97306
rect 661408 97242 661460 97248
rect 660120 96960 660172 96966
rect 660120 96902 660172 96908
rect 660672 96076 660724 96082
rect 660672 96018 660724 96024
rect 659764 95118 660146 95146
rect 660684 95132 660712 96018
rect 661420 95132 661448 97242
rect 661972 95132 662000 97786
rect 662512 97708 662564 97714
rect 662512 97650 662564 97656
rect 662524 95132 662552 97650
rect 663064 97436 663116 97442
rect 663064 97378 663116 97384
rect 663076 95132 663104 97378
rect 663984 96484 664036 96490
rect 663984 96426 664036 96432
rect 663800 96212 663852 96218
rect 663800 96154 663852 96160
rect 663248 94512 663300 94518
rect 663248 94454 663300 94460
rect 663260 93129 663288 94454
rect 663246 93120 663302 93129
rect 663246 93055 663302 93064
rect 663812 90409 663840 96154
rect 663798 90400 663854 90409
rect 663798 90335 663854 90344
rect 663996 89049 664024 96426
rect 665364 96348 665416 96354
rect 665364 96290 665416 96296
rect 665180 95940 665232 95946
rect 665180 95882 665232 95888
rect 664168 95668 664220 95674
rect 664168 95610 664220 95616
rect 663982 89040 664038 89049
rect 656900 89004 656952 89010
rect 663982 88975 664038 88984
rect 656900 88946 656952 88952
rect 656912 88890 656940 88946
rect 656912 88862 657202 88890
rect 664180 88806 664208 95610
rect 665192 91769 665220 95882
rect 665178 91760 665234 91769
rect 665178 91695 665234 91704
rect 665376 90681 665404 96290
rect 665744 93401 665772 97922
rect 665730 93392 665786 93401
rect 665730 93327 665786 93336
rect 665362 90672 665418 90681
rect 665362 90607 665418 90616
rect 657452 88800 657504 88806
rect 662328 88800 662380 88806
rect 657504 88748 657754 88754
rect 657452 88742 657754 88748
rect 657464 88726 657754 88742
rect 661986 88748 662328 88754
rect 661986 88742 662380 88748
rect 664168 88800 664220 88806
rect 664168 88742 664220 88748
rect 661986 88726 662368 88742
rect 658306 88330 658504 88346
rect 658306 88324 658516 88330
rect 658306 88318 658464 88324
rect 658464 88266 658516 88272
rect 656716 86964 656768 86970
rect 656716 86906 656768 86912
rect 653404 86760 653456 86766
rect 653404 86702 653456 86708
rect 652024 86624 652076 86630
rect 652024 86566 652076 86572
rect 658844 86494 658872 88196
rect 659580 86970 659608 88196
rect 659568 86964 659620 86970
rect 659568 86906 659620 86912
rect 660132 86630 660160 88196
rect 660684 87174 660712 88196
rect 660672 87168 660724 87174
rect 660672 87110 660724 87116
rect 661420 86766 661448 88196
rect 662524 87310 662552 88196
rect 662512 87304 662564 87310
rect 662512 87246 662564 87252
rect 661408 86760 661460 86766
rect 661408 86702 661460 86708
rect 660120 86624 660172 86630
rect 660120 86566 660172 86572
rect 650644 86488 650696 86494
rect 650644 86430 650696 86436
rect 658832 86488 658884 86494
rect 658832 86430 658884 86436
rect 648988 76560 649040 76566
rect 648988 76502 649040 76508
rect 649000 67017 649028 76502
rect 648986 67008 649042 67017
rect 648986 66943 649042 66952
rect 648802 64016 648858 64025
rect 648802 63951 648858 63960
rect 662420 57248 662472 57254
rect 662420 57190 662472 57196
rect 625804 52352 625856 52358
rect 625804 52294 625856 52300
rect 624422 47560 624478 47569
rect 624422 47495 624478 47504
rect 662432 47433 662460 57190
rect 663798 48512 663854 48521
rect 663798 48447 663854 48456
rect 662602 47832 662658 47841
rect 662602 47767 662658 47776
rect 662418 47424 662474 47433
rect 662418 47359 662474 47368
rect 662616 44878 662644 47767
rect 662604 44872 662656 44878
rect 662604 44814 662656 44820
rect 474462 43480 474518 43489
rect 474462 43415 474518 43424
rect 604458 43480 604514 43489
rect 663812 43450 663840 48447
rect 604458 43415 604514 43424
rect 663800 43444 663852 43450
rect 409602 42800 409658 42809
rect 409602 42735 409658 42744
rect 411074 42800 411130 42809
rect 411074 42735 411130 42744
rect 416594 42800 416650 42809
rect 416594 42735 416650 42744
rect 464894 42800 464950 42809
rect 464894 42735 464950 42744
rect 409616 42398 409644 42735
rect 411088 42500 411116 42735
rect 409604 42392 409656 42398
rect 409604 42334 409656 42340
rect 405108 42078 405582 42106
rect 416608 42092 416636 42735
rect 464908 42386 464936 42735
rect 474476 42500 474504 43415
rect 663800 43386 663852 43392
rect 518622 42392 518678 42401
rect 464896 42380 464948 42386
rect 464896 42322 464948 42328
rect 518678 42350 518834 42378
rect 518622 42327 518678 42336
rect 460570 42120 460626 42129
rect 460368 42078 460570 42106
rect 365166 42055 365222 42064
rect 471610 42120 471666 42129
rect 471408 42078 471610 42106
rect 460570 42055 460626 42064
rect 471610 42055 471666 42064
rect 514942 42120 514998 42129
rect 520462 42120 520518 42129
rect 514998 42078 515154 42106
rect 514942 42055 514998 42064
rect 525982 42120 526038 42129
rect 520518 42078 520674 42106
rect 520462 42055 520518 42064
rect 529570 42120 529626 42129
rect 526038 42078 526194 42106
rect 529322 42078 529570 42106
rect 525982 42055 526038 42064
rect 529570 42055 529626 42064
rect 521658 41984 521714 41993
rect 521714 41942 521870 41970
rect 521658 41919 521714 41928
rect 141896 40310 142200 40338
rect 141896 40202 141924 40310
rect 141758 40174 141924 40202
rect 141758 39984 141786 40174
<< via2 >>
rect 504546 1007020 504548 1007040
rect 504548 1007020 504600 1007040
rect 504600 1007020 504602 1007040
rect 504546 1006984 504602 1007020
rect 151726 1006868 151782 1006904
rect 151726 1006848 151728 1006868
rect 151728 1006848 151780 1006868
rect 151780 1006848 151782 1006868
rect 428002 1006868 428058 1006904
rect 506202 1006884 506204 1006904
rect 506204 1006884 506256 1006904
rect 506256 1006884 506258 1006904
rect 428002 1006848 428004 1006868
rect 428004 1006848 428056 1006868
rect 428056 1006848 428058 1006868
rect 506202 1006848 506258 1006884
rect 101126 1006460 101182 1006496
rect 101126 1006440 101128 1006460
rect 101128 1006440 101180 1006460
rect 101180 1006440 101182 1006460
rect 82266 995696 82322 995752
rect 81070 995424 81126 995480
rect 80150 994744 80206 994800
rect 84474 995152 84530 995208
rect 86590 995424 86646 995480
rect 87786 994952 87842 995008
rect 85670 994472 85726 994528
rect 92662 997192 92718 997248
rect 93122 995424 93178 995480
rect 93674 995832 93730 995888
rect 93674 995016 93730 995072
rect 85026 994200 85082 994256
rect 100298 1006324 100354 1006360
rect 100298 1006304 100300 1006324
rect 100300 1006304 100352 1006324
rect 100352 1006304 100354 1006324
rect 99470 1006188 99526 1006224
rect 99470 1006168 99472 1006188
rect 99472 1006168 99524 1006188
rect 99524 1006168 99526 1006188
rect 103978 1006188 104034 1006224
rect 103978 1006168 103980 1006188
rect 103980 1006168 104032 1006188
rect 104032 1006168 104034 1006188
rect 106830 1006188 106886 1006224
rect 106830 1006168 106832 1006188
rect 106832 1006168 106884 1006188
rect 106884 1006168 106886 1006188
rect 98274 1006052 98330 1006088
rect 98274 1006032 98276 1006052
rect 98276 1006032 98328 1006052
rect 98328 1006032 98330 1006052
rect 94686 994472 94742 994528
rect 94502 994200 94558 994256
rect 41786 968768 41842 968824
rect 41970 967136 42026 967192
rect 41786 962104 41842 962160
rect 41786 959112 41842 959168
rect 41786 956528 41842 956584
rect 41786 955440 41842 955496
rect 35162 952856 35218 952912
rect 39302 952176 39358 952232
rect 37922 938406 37978 938462
rect 40038 951768 40094 951824
rect 39302 937352 39358 937408
rect 35162 936944 35218 937000
rect 41418 951632 41474 951688
rect 41234 941840 41290 941896
rect 41234 941024 41290 941080
rect 41234 940208 41290 940264
rect 41050 939392 41106 939448
rect 41234 938406 41290 938462
rect 40038 935720 40094 935776
rect 40682 881864 40738 881920
rect 40222 819032 40278 819088
rect 39578 818624 39634 818680
rect 35622 817944 35678 818000
rect 35806 817264 35862 817320
rect 35438 816856 35494 816912
rect 35806 816448 35862 816504
rect 39762 817944 39818 818000
rect 35806 816040 35862 816096
rect 35622 815632 35678 815688
rect 35622 815224 35678 815280
rect 35806 814816 35862 814872
rect 35806 814428 35862 814464
rect 35806 814408 35808 814428
rect 35808 814408 35860 814428
rect 35860 814408 35862 814428
rect 41050 814000 41106 814056
rect 42246 937760 42302 937816
rect 42798 935312 42854 935368
rect 43074 934904 43130 934960
rect 43534 943472 43590 943528
rect 43626 942248 43682 942304
rect 43442 941332 43444 941352
rect 43444 941332 43496 941352
rect 43496 941332 43498 941352
rect 43442 941296 43498 941332
rect 43442 939820 43498 939856
rect 43442 939800 43444 939820
rect 43444 939800 43496 939820
rect 43496 939800 43498 939820
rect 43258 934496 43314 934552
rect 44638 943064 44694 943120
rect 47582 942656 47638 942712
rect 46202 940616 46258 940672
rect 98274 1001972 98330 1002008
rect 98274 1001952 98276 1001972
rect 98276 1001952 98328 1001972
rect 98328 1001952 98330 1001972
rect 97446 995968 97502 996024
rect 100298 1002380 100354 1002416
rect 100298 1002360 100300 1002380
rect 100300 1002360 100352 1002380
rect 100352 1002360 100354 1002380
rect 101126 1002244 101182 1002280
rect 101126 1002224 101128 1002244
rect 101128 1002224 101180 1002244
rect 101180 1002224 101182 1002244
rect 99102 1002108 99158 1002144
rect 99102 1002088 99104 1002108
rect 99104 1002088 99156 1002108
rect 99156 1002088 99158 1002108
rect 100206 995288 100262 995344
rect 100022 995016 100078 995072
rect 102322 1002652 102378 1002688
rect 102322 1002632 102324 1002652
rect 102324 1002632 102376 1002652
rect 102376 1002632 102378 1002652
rect 101954 1002516 102010 1002552
rect 101954 1002496 101956 1002516
rect 101956 1002496 102008 1002516
rect 102008 1002496 102010 1002516
rect 101954 1001972 102010 1002008
rect 101954 1001952 101956 1001972
rect 101956 1001952 102008 1001972
rect 102008 1001952 102010 1001972
rect 104806 1006052 104862 1006088
rect 104806 1006032 104808 1006052
rect 104808 1006032 104860 1006052
rect 104860 1006032 104862 1006052
rect 107658 1006052 107714 1006088
rect 107658 1006032 107660 1006052
rect 107660 1006032 107712 1006052
rect 107712 1006032 107714 1006052
rect 103150 1004692 103206 1004728
rect 103150 1004672 103152 1004692
rect 103152 1004672 103204 1004692
rect 103204 1004672 103206 1004692
rect 108486 1004692 108542 1004728
rect 108486 1004672 108488 1004692
rect 108488 1004672 108540 1004692
rect 108540 1004672 108542 1004692
rect 106002 1002532 106004 1002552
rect 106004 1002532 106056 1002552
rect 106056 1002532 106058 1002552
rect 106002 1002496 106058 1002532
rect 105634 1002260 105636 1002280
rect 105636 1002260 105688 1002280
rect 105688 1002260 105690 1002280
rect 105634 1002224 105690 1002260
rect 103150 1002108 103206 1002144
rect 103150 1002088 103152 1002108
rect 103152 1002088 103204 1002108
rect 103204 1002088 103206 1002108
rect 104806 1002124 104808 1002144
rect 104808 1002124 104860 1002144
rect 104860 1002124 104862 1002144
rect 104806 1002088 104862 1002124
rect 103978 1001952 104034 1002008
rect 106002 1001988 106004 1002008
rect 106004 1001988 106056 1002008
rect 106056 1001988 106058 1002008
rect 106002 1001952 106058 1001988
rect 103518 994744 103574 994800
rect 108026 1002396 108028 1002416
rect 108028 1002396 108080 1002416
rect 108080 1002396 108082 1002416
rect 108026 1002360 108082 1002396
rect 108486 1002260 108488 1002280
rect 108488 1002260 108540 1002280
rect 108540 1002260 108542 1002280
rect 106830 1002124 106832 1002144
rect 106832 1002124 106884 1002144
rect 106884 1002124 106886 1002144
rect 106830 1002088 106886 1002124
rect 108486 1002224 108542 1002260
rect 108854 1001972 108910 1002008
rect 108854 1001952 108856 1001972
rect 108856 1001952 108908 1001972
rect 108908 1001952 108910 1001972
rect 109682 1002108 109738 1002144
rect 109682 1002088 109684 1002108
rect 109684 1002088 109736 1002108
rect 109736 1002088 109738 1002108
rect 133602 995696 133658 995752
rect 139122 995696 139178 995752
rect 140962 995696 141018 995752
rect 142894 995696 142950 995752
rect 131578 994744 131634 994800
rect 132774 994472 132830 994528
rect 137098 995016 137154 995072
rect 141790 995288 141846 995344
rect 144366 996648 144422 996704
rect 144826 996376 144882 996432
rect 136454 994200 136510 994256
rect 307758 1006732 307814 1006768
rect 307758 1006712 307760 1006732
rect 307760 1006712 307812 1006732
rect 307812 1006712 307814 1006732
rect 357714 1006732 357770 1006768
rect 357714 1006712 357716 1006732
rect 357716 1006712 357768 1006732
rect 357768 1006712 357770 1006732
rect 430854 1006732 430910 1006768
rect 430854 1006712 430856 1006732
rect 430856 1006712 430908 1006732
rect 430908 1006712 430910 1006732
rect 146942 1006032 146998 1006088
rect 145746 996920 145802 996976
rect 146758 995288 146814 995344
rect 145562 994200 145618 994256
rect 150898 1006324 150954 1006360
rect 150898 1006304 150900 1006324
rect 150900 1006304 150952 1006324
rect 150952 1006304 150954 1006324
rect 151266 1006188 151322 1006224
rect 255318 1006460 255374 1006496
rect 255318 1006440 255320 1006460
rect 255320 1006440 255372 1006460
rect 255372 1006440 255374 1006460
rect 152094 1006340 152096 1006360
rect 152096 1006340 152148 1006360
rect 152148 1006340 152150 1006360
rect 152094 1006304 152150 1006340
rect 158258 1006324 158314 1006360
rect 158258 1006304 158260 1006324
rect 158260 1006304 158312 1006324
rect 158312 1006304 158314 1006324
rect 210422 1006340 210424 1006360
rect 210424 1006340 210476 1006360
rect 210476 1006340 210478 1006360
rect 210422 1006304 210478 1006340
rect 151266 1006168 151268 1006188
rect 151268 1006168 151320 1006188
rect 151320 1006168 151322 1006188
rect 159454 1006188 159510 1006224
rect 159454 1006168 159456 1006188
rect 159456 1006168 159508 1006188
rect 159508 1006168 159510 1006188
rect 160282 1006188 160338 1006224
rect 208398 1006204 208400 1006224
rect 208400 1006204 208452 1006224
rect 208452 1006204 208454 1006224
rect 160282 1006168 160284 1006188
rect 160284 1006168 160336 1006188
rect 160336 1006168 160338 1006188
rect 208398 1006168 208454 1006204
rect 148874 1006052 148930 1006088
rect 148874 1006032 148876 1006052
rect 148876 1006032 148928 1006052
rect 148928 1006032 148930 1006052
rect 150070 1006052 150126 1006088
rect 150070 1006032 150072 1006052
rect 150072 1006032 150124 1006052
rect 150124 1006032 150126 1006052
rect 158626 1006052 158682 1006088
rect 158626 1006032 158628 1006052
rect 158628 1006032 158680 1006052
rect 158680 1006032 158682 1006052
rect 152922 1005236 152978 1005272
rect 152922 1005216 152924 1005236
rect 152924 1005216 152976 1005236
rect 152976 1005216 152978 1005236
rect 148322 995016 148378 995072
rect 149242 1001972 149298 1002008
rect 149242 1001952 149244 1001972
rect 149244 1001952 149296 1001972
rect 149296 1001952 149298 1001972
rect 153750 1005100 153806 1005136
rect 153750 1005080 153752 1005100
rect 153752 1005080 153804 1005100
rect 153804 1005080 153806 1005100
rect 150898 1002108 150954 1002144
rect 150898 1002088 150900 1002108
rect 150900 1002088 150952 1002108
rect 150952 1002088 150954 1002108
rect 152922 1004964 152978 1005000
rect 152922 1004944 152924 1004964
rect 152924 1004944 152976 1004964
rect 152976 1004944 152978 1004964
rect 160650 1004964 160706 1005000
rect 160650 1004944 160652 1004964
rect 160652 1004944 160704 1004964
rect 160704 1004944 160706 1004964
rect 154118 1004828 154174 1004864
rect 154118 1004808 154120 1004828
rect 154120 1004808 154172 1004828
rect 154172 1004808 154174 1004828
rect 151266 995696 151322 995752
rect 153750 1001988 153752 1002008
rect 153752 1001988 153804 1002008
rect 153804 1001988 153806 1002008
rect 153750 1001952 153806 1001988
rect 149702 994472 149758 994528
rect 159454 1004828 159510 1004864
rect 159454 1004808 159456 1004828
rect 159456 1004808 159508 1004828
rect 159508 1004808 159510 1004828
rect 160650 1004692 160706 1004728
rect 160650 1004672 160652 1004692
rect 160652 1004672 160704 1004692
rect 160704 1004672 160706 1004692
rect 157430 1002516 157486 1002552
rect 157430 1002496 157432 1002516
rect 157432 1002496 157484 1002516
rect 157484 1002496 157486 1002516
rect 158626 1002380 158682 1002416
rect 158626 1002360 158628 1002380
rect 158628 1002360 158680 1002380
rect 158680 1002360 158682 1002380
rect 155774 1002260 155776 1002280
rect 155776 1002260 155828 1002280
rect 155828 1002260 155830 1002280
rect 155774 1002224 155830 1002260
rect 156602 1002244 156658 1002280
rect 156602 1002224 156604 1002244
rect 156604 1002224 156656 1002244
rect 156656 1002224 156658 1002244
rect 154578 1002124 154580 1002144
rect 154580 1002124 154632 1002144
rect 154632 1002124 154634 1002144
rect 154578 1002088 154634 1002124
rect 154946 1002108 155002 1002144
rect 154946 1002088 154948 1002108
rect 154948 1002088 155000 1002108
rect 155000 1002088 155002 1002108
rect 155774 1001972 155830 1002008
rect 155774 1001952 155776 1001972
rect 155776 1001952 155828 1001972
rect 155828 1001952 155830 1001972
rect 156602 1001952 156658 1002008
rect 157798 1001972 157854 1002008
rect 157798 1001952 157800 1001972
rect 157800 1001952 157852 1001972
rect 157852 1001952 157854 1001972
rect 157338 994744 157394 994800
rect 201038 1006052 201094 1006088
rect 201038 1006032 201040 1006052
rect 201040 1006032 201092 1006052
rect 201092 1006032 201094 1006052
rect 195150 997600 195206 997656
rect 184478 995696 184534 995752
rect 187514 995696 187570 995752
rect 189538 995696 189594 995752
rect 190458 995696 190514 995752
rect 195334 995696 195390 995752
rect 177302 995016 177358 995072
rect 180614 994492 180670 994528
rect 183834 995424 183890 995480
rect 184478 994744 184534 994800
rect 180614 994472 180616 994492
rect 180616 994472 180668 994492
rect 180668 994472 180670 994492
rect 188802 994472 188858 994528
rect 188158 993928 188214 993984
rect 192482 995424 192538 995480
rect 192942 994744 192998 994800
rect 193126 994744 193182 994800
rect 192942 994200 192998 994256
rect 209226 1004964 209282 1005000
rect 209226 1004944 209228 1004964
rect 209228 1004944 209280 1004964
rect 209280 1004944 209282 1004964
rect 207202 1004828 207258 1004864
rect 207202 1004808 207204 1004828
rect 207204 1004808 207256 1004828
rect 207256 1004808 207258 1004828
rect 209226 1004692 209282 1004728
rect 209226 1004672 209228 1004692
rect 209228 1004672 209280 1004692
rect 209280 1004672 209282 1004692
rect 206374 1002516 206430 1002552
rect 206374 1002496 206376 1002516
rect 206376 1002496 206428 1002516
rect 206428 1002496 206430 1002516
rect 198002 994744 198058 994800
rect 196622 993928 196678 993984
rect 191746 993112 191802 993168
rect 202694 998572 202750 998608
rect 202694 998552 202696 998572
rect 202696 998552 202748 998572
rect 202748 998552 202750 998572
rect 200670 997908 200672 997928
rect 200672 997908 200724 997928
rect 200724 997908 200726 997928
rect 200670 997872 200726 997908
rect 199842 996376 199898 996432
rect 199382 994200 199438 994256
rect 201866 997772 201868 997792
rect 201868 997772 201920 997792
rect 201920 997772 201922 997792
rect 201866 997736 201922 997772
rect 200210 997228 200212 997248
rect 200212 997228 200264 997248
rect 200264 997228 200266 997248
rect 200210 997192 200266 997228
rect 202694 998044 202696 998064
rect 202696 998044 202748 998064
rect 202748 998044 202750 998064
rect 202694 998008 202750 998044
rect 206374 1002244 206430 1002280
rect 206374 1002224 206376 1002244
rect 206376 1002224 206428 1002244
rect 206428 1002224 206430 1002244
rect 203890 1001972 203946 1002008
rect 203890 1001952 203892 1001972
rect 203892 1001952 203944 1001972
rect 203944 1001952 203946 1001972
rect 203522 999132 203524 999152
rect 203524 999132 203576 999152
rect 203576 999132 203578 999152
rect 203522 999096 203578 999132
rect 204350 998708 204406 998744
rect 204350 998688 204352 998708
rect 204352 998688 204404 998708
rect 204404 998688 204406 998708
rect 203522 997908 203524 997928
rect 203524 997908 203576 997928
rect 203576 997908 203578 997928
rect 203522 997872 203578 997908
rect 204718 997772 204720 997792
rect 204720 997772 204772 997792
rect 204772 997772 204774 997792
rect 204718 997736 204774 997772
rect 205546 1001972 205602 1002008
rect 205546 1001952 205548 1001972
rect 205548 1001952 205600 1001972
rect 205600 1001952 205602 1001972
rect 207202 1002088 207258 1002144
rect 205546 998180 205548 998200
rect 205548 998180 205600 998200
rect 205600 998180 205602 998200
rect 205546 998144 205602 998180
rect 202326 995424 202382 995480
rect 207570 1001952 207626 1002008
rect 208398 1001952 208454 1002008
rect 210422 1001952 210478 1002008
rect 211250 1002380 211306 1002416
rect 211250 1002360 211252 1002380
rect 211252 1002360 211304 1002380
rect 211304 1002360 211306 1002380
rect 211250 1002108 211306 1002144
rect 211250 1002088 211252 1002108
rect 211252 1002088 211304 1002108
rect 211304 1002088 211306 1002108
rect 212538 1004692 212594 1004728
rect 212538 1004672 212540 1004692
rect 212540 1004672 212592 1004692
rect 212592 1004672 212594 1004692
rect 212078 1001972 212134 1002008
rect 212078 1001952 212080 1001972
rect 212080 1001952 212132 1001972
rect 212132 1001952 212134 1001972
rect 200762 994472 200818 994528
rect 246670 996376 246726 996432
rect 240874 995696 240930 995752
rect 245566 995696 245622 995752
rect 239586 994880 239642 994936
rect 238666 994472 238722 994528
rect 236550 994200 236606 994256
rect 243910 995424 243966 995480
rect 242944 995152 243000 995208
rect 244232 995152 244288 995208
rect 254122 1006324 254178 1006360
rect 254122 1006304 254124 1006324
rect 254124 1006304 254176 1006324
rect 254176 1006304 254178 1006324
rect 253662 1006188 253718 1006224
rect 253662 1006168 253664 1006188
rect 253664 1006168 253716 1006188
rect 253716 1006168 253718 1006188
rect 262678 1006188 262734 1006224
rect 262678 1006168 262680 1006188
rect 262680 1006168 262732 1006188
rect 262732 1006168 262734 1006188
rect 252466 1006052 252522 1006088
rect 252466 1006032 252468 1006052
rect 252468 1006032 252520 1006052
rect 252520 1006032 252522 1006052
rect 261850 1006052 261906 1006088
rect 261850 1006032 261852 1006052
rect 261852 1006032 261904 1006052
rect 261904 1006032 261906 1006052
rect 247866 996648 247922 996704
rect 249338 995152 249394 995208
rect 247682 994880 247738 994936
rect 240138 993928 240194 993984
rect 263046 1005252 263048 1005272
rect 263048 1005252 263100 1005272
rect 263100 1005252 263102 1005272
rect 263046 1005216 263102 1005252
rect 255318 1002516 255374 1002552
rect 255318 1002496 255320 1002516
rect 255320 1002496 255372 1002516
rect 255372 1002496 255374 1002516
rect 261022 1002516 261078 1002552
rect 261022 1002496 261024 1002516
rect 261024 1002496 261076 1002516
rect 261076 1002496 261078 1002516
rect 256146 1002380 256202 1002416
rect 256146 1002360 256148 1002380
rect 256148 1002360 256200 1002380
rect 256200 1002360 256202 1002380
rect 252466 1001972 252522 1002008
rect 252466 1001952 252468 1001972
rect 252468 1001952 252520 1001972
rect 252520 1001952 252522 1001972
rect 254490 1002244 254546 1002280
rect 254490 1002224 254492 1002244
rect 254492 1002224 254544 1002244
rect 254544 1002224 254546 1002244
rect 253294 1002108 253350 1002144
rect 253294 1002088 253296 1002108
rect 253296 1002088 253348 1002108
rect 253348 1002088 253350 1002108
rect 256146 1002108 256202 1002144
rect 256146 1002088 256148 1002108
rect 256148 1002088 256200 1002108
rect 256200 1002088 256202 1002108
rect 263506 1002108 263562 1002144
rect 263506 1002088 263508 1002108
rect 263508 1002088 263560 1002108
rect 263560 1002088 263562 1002108
rect 261022 1001972 261078 1002008
rect 261022 1001952 261024 1001972
rect 261024 1001952 261076 1001972
rect 261076 1001952 261078 1001972
rect 263874 1001972 263930 1002008
rect 263874 1001952 263876 1001972
rect 263876 1001952 263928 1001972
rect 263928 1001952 263930 1001972
rect 258170 998164 258226 998200
rect 258170 998144 258172 998164
rect 258172 998144 258224 998164
rect 258224 998144 258226 998164
rect 257342 998028 257398 998064
rect 257342 998008 257344 998028
rect 257344 998008 257396 998028
rect 257396 998008 257398 998028
rect 256974 997892 257030 997928
rect 256974 997872 256976 997892
rect 256976 997872 257028 997892
rect 257028 997872 257030 997892
rect 256514 997736 256570 997792
rect 254582 994472 254638 994528
rect 258170 997872 258226 997928
rect 258998 997736 259054 997792
rect 260194 998044 260196 998064
rect 260196 998044 260248 998064
rect 260248 998044 260250 998064
rect 260194 998008 260250 998044
rect 259826 997908 259828 997928
rect 259828 997908 259880 997928
rect 259880 997908 259882 997928
rect 259826 997872 259882 997908
rect 260194 997772 260196 997792
rect 260196 997772 260248 997792
rect 260248 997772 260250 997792
rect 260194 997736 260250 997772
rect 261850 997736 261906 997792
rect 252006 994200 252062 994256
rect 251822 993928 251878 993984
rect 251454 993112 251510 993168
rect 291750 995696 291806 995752
rect 293498 995696 293554 995752
rect 297270 995696 297326 995752
rect 298282 997736 298338 997792
rect 286690 995424 286746 995480
rect 287794 994472 287850 994528
rect 287518 994200 287574 994256
rect 292486 995424 292542 995480
rect 290830 994744 290886 994800
rect 296166 995424 296222 995480
rect 296442 995052 296444 995072
rect 296444 995052 296496 995072
rect 296496 995052 296498 995072
rect 296442 995016 296498 995052
rect 298282 995696 298338 995752
rect 299018 996784 299074 996840
rect 304078 1006460 304134 1006496
rect 304078 1006440 304080 1006460
rect 304080 1006440 304132 1006460
rect 304132 1006440 304134 1006460
rect 305274 1006324 305330 1006360
rect 305274 1006304 305276 1006324
rect 305276 1006304 305328 1006324
rect 305328 1006304 305330 1006324
rect 314658 1006460 314714 1006496
rect 314658 1006440 314660 1006460
rect 314660 1006440 314712 1006460
rect 314712 1006440 314714 1006460
rect 361394 1006460 361450 1006496
rect 361394 1006440 361396 1006460
rect 361396 1006440 361448 1006460
rect 361448 1006440 361450 1006460
rect 306930 1006324 306986 1006360
rect 306930 1006304 306932 1006324
rect 306932 1006304 306984 1006324
rect 306984 1006304 306986 1006324
rect 311806 1006188 311862 1006224
rect 311806 1006168 311808 1006188
rect 311808 1006168 311860 1006188
rect 311860 1006168 311862 1006188
rect 314658 1006188 314714 1006224
rect 314658 1006168 314660 1006188
rect 314660 1006168 314712 1006188
rect 314712 1006168 314714 1006188
rect 301502 1006032 301558 1006088
rect 303250 1006052 303306 1006088
rect 303250 1006032 303252 1006052
rect 303252 1006032 303304 1006052
rect 303304 1006032 303306 1006052
rect 300858 996376 300914 996432
rect 300306 995968 300362 996024
rect 300122 995696 300178 995752
rect 298834 995016 298890 995072
rect 297914 994744 297970 994800
rect 304078 1006052 304134 1006088
rect 304078 1006032 304080 1006052
rect 304080 1006032 304132 1006052
rect 304132 1006032 304134 1006052
rect 305274 1006052 305330 1006088
rect 305274 1006032 305276 1006052
rect 305276 1006032 305328 1006052
rect 305328 1006032 305330 1006052
rect 307298 1005236 307354 1005272
rect 307298 1005216 307300 1005236
rect 307300 1005216 307352 1005236
rect 307352 1005216 307354 1005236
rect 303250 997772 303252 997792
rect 303252 997772 303304 997792
rect 303304 997772 303306 997792
rect 303250 997736 303306 997772
rect 301502 995424 301558 995480
rect 301042 994472 301098 994528
rect 308954 1004964 309010 1005000
rect 308954 1004944 308956 1004964
rect 308956 1004944 309008 1004964
rect 309008 1004944 309010 1004964
rect 306930 1004828 306986 1004864
rect 306930 1004808 306932 1004828
rect 306932 1004808 306984 1004828
rect 306984 1004808 306986 1004828
rect 313830 1004828 313886 1004864
rect 313830 1004808 313832 1004828
rect 313832 1004808 313884 1004828
rect 313884 1004808 313886 1004828
rect 308126 1004692 308182 1004728
rect 308126 1004672 308128 1004692
rect 308128 1004672 308180 1004692
rect 308180 1004672 308182 1004692
rect 315486 1004692 315542 1004728
rect 315486 1004672 315488 1004692
rect 315488 1004672 315540 1004692
rect 315540 1004672 315542 1004692
rect 310150 1002380 310206 1002416
rect 310150 1002360 310152 1002380
rect 310152 1002360 310204 1002380
rect 310204 1002360 310206 1002380
rect 306102 1002244 306158 1002280
rect 306102 1002224 306104 1002244
rect 306104 1002224 306156 1002244
rect 306156 1002224 306158 1002244
rect 308954 1002108 309010 1002144
rect 308954 1002088 308956 1002108
rect 308956 1002088 309008 1002108
rect 309008 1002088 309010 1002108
rect 306102 1001972 306158 1002008
rect 306102 1001952 306104 1001972
rect 306104 1001952 306156 1001972
rect 306156 1001952 306158 1001972
rect 304262 994200 304318 994256
rect 310150 1002088 310206 1002144
rect 310610 1002088 310666 1002144
rect 310978 1002108 311034 1002144
rect 310978 1002088 310980 1002108
rect 310980 1002088 311032 1002108
rect 311032 1002088 311034 1002108
rect 309782 1001972 309838 1002008
rect 309782 1001952 309784 1001972
rect 309784 1001952 309836 1001972
rect 309836 1001952 309838 1001972
rect 312634 1001972 312690 1002008
rect 312634 1001952 312636 1001972
rect 312636 1001952 312688 1001972
rect 312688 1001952 312690 1001972
rect 290278 993928 290334 993984
rect 307022 993928 307078 993984
rect 316406 992840 316462 992896
rect 365074 1006188 365130 1006224
rect 365074 1006168 365076 1006188
rect 365076 1006168 365128 1006188
rect 365128 1006168 365130 1006188
rect 354862 1006052 354918 1006088
rect 354862 1006032 354864 1006052
rect 354864 1006032 354916 1006052
rect 354916 1006032 354918 1006052
rect 357346 1006052 357402 1006088
rect 357346 1006032 357348 1006052
rect 357348 1006032 357400 1006052
rect 357400 1006032 357402 1006052
rect 356518 1005388 356520 1005408
rect 356520 1005388 356572 1005408
rect 356572 1005388 356574 1005408
rect 356518 1005352 356574 1005388
rect 355690 1004964 355746 1005000
rect 355690 1004944 355692 1004964
rect 355692 1004944 355744 1004964
rect 355744 1004944 355746 1004964
rect 355690 1004692 355746 1004728
rect 355690 1004672 355692 1004692
rect 355692 1004672 355744 1004692
rect 355744 1004672 355746 1004692
rect 354034 1001972 354090 1002008
rect 354034 1001952 354036 1001972
rect 354036 1001952 354088 1001972
rect 354088 1001952 354090 1001972
rect 360566 1005660 360568 1005680
rect 360568 1005660 360620 1005680
rect 360620 1005660 360622 1005680
rect 360566 1005624 360622 1005660
rect 359738 1005524 359740 1005544
rect 359740 1005524 359792 1005544
rect 359792 1005524 359794 1005544
rect 359738 1005488 359794 1005524
rect 356886 1005252 356888 1005272
rect 356888 1005252 356940 1005272
rect 356940 1005252 356942 1005272
rect 356886 1005216 356942 1005252
rect 363418 1005100 363474 1005136
rect 363418 1005080 363420 1005100
rect 363420 1005080 363472 1005100
rect 363472 1005080 363474 1005100
rect 365074 1005100 365130 1005136
rect 365074 1005080 365076 1005100
rect 365076 1005080 365128 1005100
rect 365128 1005080 365130 1005100
rect 361394 1004964 361450 1005000
rect 361394 1004944 361396 1004964
rect 361396 1004944 361448 1004964
rect 361448 1004944 361450 1004964
rect 364246 1004828 364302 1004864
rect 364246 1004808 364248 1004828
rect 364248 1004808 364300 1004828
rect 364300 1004808 364302 1004828
rect 362590 1004692 362646 1004728
rect 362590 1004672 362592 1004692
rect 362592 1004672 362644 1004692
rect 362644 1004672 362646 1004692
rect 358542 1002380 358598 1002416
rect 358542 1002360 358544 1002380
rect 358544 1002360 358596 1002380
rect 358596 1002360 358598 1002380
rect 359370 1002244 359426 1002280
rect 359370 1002224 359372 1002244
rect 359372 1002224 359424 1002244
rect 359424 1002224 359426 1002244
rect 358542 1002088 358598 1002144
rect 357346 1001972 357402 1002008
rect 357346 1001952 357348 1001972
rect 357348 1001952 357400 1001972
rect 357400 1001952 357402 1001972
rect 360566 1002108 360622 1002144
rect 360566 1002088 360568 1002108
rect 360568 1002088 360620 1002108
rect 360620 1002088 360622 1002108
rect 360198 1001972 360254 1002008
rect 360198 1001952 360200 1001972
rect 360200 1001952 360252 1001972
rect 360252 1001952 360254 1001972
rect 365902 1001972 365958 1002008
rect 365902 1001952 365904 1001972
rect 365904 1001952 365956 1001972
rect 365956 1001952 365958 1001972
rect 372342 996648 372398 996704
rect 372526 996376 372582 996432
rect 373262 995016 373318 995072
rect 376298 994744 376354 994800
rect 383106 995696 383162 995752
rect 385682 995696 385738 995752
rect 387890 995696 387946 995752
rect 388166 995696 388222 995752
rect 396538 995696 396594 995752
rect 381542 995288 381598 995344
rect 389362 995288 389418 995344
rect 392122 995016 392178 995072
rect 393318 995152 393374 995208
rect 393226 995016 393282 995072
rect 381266 994472 381322 994528
rect 392306 994472 392362 994528
rect 378414 994200 378470 994256
rect 395158 994744 395214 994800
rect 427174 1006596 427230 1006632
rect 427174 1006576 427176 1006596
rect 427176 1006576 427228 1006596
rect 427228 1006576 427230 1006596
rect 423494 1006460 423550 1006496
rect 423494 1006440 423496 1006460
rect 423496 1006440 423548 1006460
rect 423548 1006440 423550 1006460
rect 424322 1006324 424378 1006360
rect 424322 1006304 424324 1006324
rect 424324 1006304 424376 1006324
rect 424376 1006304 424378 1006324
rect 422666 1006032 422722 1006088
rect 423494 1006052 423550 1006088
rect 423494 1006032 423496 1006052
rect 423496 1006032 423548 1006052
rect 423548 1006032 423550 1006052
rect 429198 1006052 429254 1006088
rect 429198 1006032 429200 1006052
rect 429200 1006032 429252 1006052
rect 429252 1006032 429254 1006052
rect 427542 1005660 427544 1005680
rect 427544 1005660 427596 1005680
rect 427596 1005660 427598 1005680
rect 427542 1005624 427598 1005660
rect 425518 1005372 425574 1005408
rect 425518 1005352 425520 1005372
rect 425520 1005352 425572 1005372
rect 425572 1005352 425574 1005372
rect 424690 1005100 424746 1005136
rect 424690 1005080 424692 1005100
rect 424692 1005080 424744 1005100
rect 424744 1005080 424746 1005100
rect 421470 1001972 421526 1002008
rect 421470 1001952 421472 1001972
rect 421472 1001952 421524 1001972
rect 421524 1001952 421526 1001972
rect 393226 994200 393282 994256
rect 421010 996412 421012 996432
rect 421012 996412 421064 996432
rect 421064 996412 421066 996432
rect 421010 996376 421066 996412
rect 422666 1004672 422722 1004728
rect 425518 1003892 425520 1003912
rect 425520 1003892 425572 1003912
rect 425572 1003892 425574 1003912
rect 425518 1003856 425574 1003892
rect 424690 1002668 424692 1002688
rect 424692 1002668 424744 1002688
rect 424744 1002668 424746 1002688
rect 424690 1002632 424746 1002668
rect 428370 1005796 428372 1005816
rect 428372 1005796 428424 1005816
rect 428424 1005796 428426 1005816
rect 428370 1005760 428426 1005796
rect 430854 1005524 430856 1005544
rect 430856 1005524 430908 1005544
rect 430908 1005524 430910 1005544
rect 430854 1005488 430910 1005524
rect 430026 1005236 430082 1005272
rect 430026 1005216 430028 1005236
rect 430028 1005216 430080 1005236
rect 430080 1005216 430082 1005236
rect 431682 1005100 431738 1005136
rect 431682 1005080 431684 1005100
rect 431684 1005080 431736 1005100
rect 431736 1005080 431738 1005100
rect 432050 1005216 432106 1005272
rect 429198 1004964 429254 1005000
rect 429198 1004944 429200 1004964
rect 429200 1004944 429252 1004964
rect 429252 1004944 429254 1004964
rect 430026 1004828 430082 1004864
rect 430026 1004808 430028 1004828
rect 430028 1004808 430080 1004828
rect 430080 1004808 430082 1004828
rect 431682 1004692 431738 1004728
rect 431682 1004672 431684 1004692
rect 431684 1004672 431736 1004692
rect 431736 1004672 431738 1004692
rect 426346 1002224 426402 1002280
rect 426346 1001972 426402 1002008
rect 426346 1001952 426348 1001972
rect 426348 1001952 426400 1001972
rect 426400 1001952 426402 1001972
rect 428370 1001972 428426 1002008
rect 428370 1001952 428372 1001972
rect 428372 1001952 428424 1001972
rect 428424 1001952 428426 1001972
rect 432878 1004028 432880 1004048
rect 432880 1004028 432932 1004048
rect 432932 1004028 432934 1004048
rect 432878 1003992 432934 1004028
rect 433338 1002108 433394 1002144
rect 433338 1002088 433340 1002108
rect 433340 1002088 433392 1002108
rect 433392 1002088 433394 1002108
rect 439686 996648 439742 996704
rect 439870 996376 439926 996432
rect 501694 1006460 501750 1006496
rect 501694 1006440 501696 1006460
rect 501696 1006440 501748 1006460
rect 501748 1006440 501750 1006460
rect 502154 1006324 502210 1006360
rect 502154 1006304 502156 1006324
rect 502156 1006304 502208 1006324
rect 502208 1006304 502210 1006324
rect 500498 1006188 500554 1006224
rect 500498 1006168 500500 1006188
rect 500500 1006168 500552 1006188
rect 500552 1006168 500554 1006188
rect 499670 1006052 499726 1006088
rect 499670 1006032 499672 1006052
rect 499672 1006032 499724 1006052
rect 499724 1006032 499726 1006052
rect 505374 1006052 505430 1006088
rect 505374 1006032 505376 1006052
rect 505376 1006032 505428 1006052
rect 505428 1006032 505430 1006052
rect 451738 995016 451794 995072
rect 445758 994744 445814 994800
rect 456798 996104 456854 996160
rect 443458 993928 443514 993984
rect 454682 994200 454738 994256
rect 500498 1005252 500500 1005272
rect 500500 1005252 500552 1005272
rect 500552 1005252 500554 1005272
rect 500498 1005216 500554 1005252
rect 499670 1004828 499726 1004864
rect 499670 1004808 499672 1004828
rect 499672 1004808 499724 1004828
rect 499724 1004808 499726 1004828
rect 472622 995696 472678 995752
rect 477038 995696 477094 995752
rect 478326 995696 478382 995752
rect 485594 995696 485650 995752
rect 471794 994472 471850 994528
rect 474094 995424 474150 995480
rect 474738 995424 474794 995480
rect 476762 995016 476818 995072
rect 480810 995424 480866 995480
rect 482282 994744 482338 994800
rect 481546 994472 481602 994528
rect 477958 993928 478014 993984
rect 501326 1004692 501382 1004728
rect 501326 1004672 501328 1004692
rect 501328 1004672 501380 1004692
rect 501380 1004672 501382 1004692
rect 498474 1001972 498530 1002008
rect 498474 1001952 498476 1001972
rect 498476 1001952 498528 1001972
rect 498528 1001952 498530 1001972
rect 502522 1002532 502524 1002552
rect 502524 1002532 502576 1002552
rect 502576 1002532 502578 1002552
rect 502522 1002496 502578 1002532
rect 502522 1001972 502578 1002008
rect 502522 1001952 502524 1001972
rect 502524 1001952 502576 1001972
rect 502576 1001952 502578 1001972
rect 505006 1005524 505008 1005544
rect 505008 1005524 505060 1005544
rect 505060 1005524 505062 1005544
rect 505006 1005488 505062 1005524
rect 505374 1003892 505376 1003912
rect 505376 1003892 505428 1003912
rect 505428 1003892 505430 1003912
rect 505374 1003856 505430 1003892
rect 503350 1002244 503406 1002280
rect 503350 1002224 503352 1002244
rect 503352 1002224 503404 1002244
rect 503404 1002224 503406 1002244
rect 504178 1002108 504234 1002144
rect 504178 1002088 504180 1002108
rect 504180 1002088 504232 1002108
rect 504232 1002088 504234 1002108
rect 503350 1001972 503406 1002008
rect 503350 1001952 503352 1001972
rect 503352 1001952 503404 1001972
rect 503404 1001952 503406 1001972
rect 509054 1005796 509056 1005816
rect 509056 1005796 509108 1005816
rect 509108 1005796 509110 1005816
rect 509054 1005760 509110 1005796
rect 508226 1005388 508228 1005408
rect 508228 1005388 508280 1005408
rect 508280 1005388 508282 1005408
rect 508226 1005352 508282 1005388
rect 507030 1005116 507032 1005136
rect 507032 1005116 507084 1005136
rect 507084 1005116 507086 1005136
rect 507030 1005080 507086 1005116
rect 508226 1004980 508228 1005000
rect 508228 1004980 508280 1005000
rect 508280 1004980 508282 1005000
rect 508226 1004944 508282 1004980
rect 507858 1004844 507860 1004864
rect 507860 1004844 507912 1004864
rect 507912 1004844 507914 1004864
rect 507858 1004808 507914 1004844
rect 509054 1004692 509110 1004728
rect 509054 1004672 509056 1004692
rect 509056 1004672 509108 1004692
rect 509108 1004672 509110 1004692
rect 506202 1001972 506258 1002008
rect 506202 1001952 506204 1001972
rect 506204 1001952 506256 1001972
rect 506256 1001952 506258 1001972
rect 507030 1001952 507086 1002008
rect 509882 1002108 509938 1002144
rect 509882 1002088 509884 1002108
rect 509884 1002088 509936 1002108
rect 509936 1002088 509938 1002108
rect 510342 1004692 510398 1004728
rect 510342 1004672 510344 1004692
rect 510344 1004672 510396 1004692
rect 510396 1004672 510398 1004692
rect 511078 995832 511134 995888
rect 559654 1007004 559710 1007040
rect 559654 1006984 559656 1007004
rect 559656 1006984 559708 1007004
rect 559708 1006984 559710 1007004
rect 552294 1006460 552350 1006496
rect 552294 1006440 552296 1006460
rect 552296 1006440 552348 1006460
rect 552348 1006440 552350 1006460
rect 516874 996784 516930 996840
rect 516690 996376 516746 996432
rect 517058 995016 517114 995072
rect 519542 996240 519598 996296
rect 520186 995696 520242 995752
rect 551466 1006188 551522 1006224
rect 551466 1006168 551468 1006188
rect 551468 1006168 551520 1006188
rect 551520 1006168 551522 1006188
rect 551098 1006032 551154 1006088
rect 553122 1006052 553178 1006088
rect 553122 1006032 553124 1006052
rect 553124 1006032 553176 1006052
rect 553176 1006032 553178 1006052
rect 520922 994472 520978 994528
rect 518162 994200 518218 994256
rect 551098 997908 551100 997928
rect 551100 997908 551152 997928
rect 551152 997908 551154 997928
rect 526074 995696 526130 995752
rect 528006 995696 528062 995752
rect 528558 995696 528614 995752
rect 532790 995696 532846 995752
rect 536562 995696 536618 995752
rect 532514 995016 532570 995072
rect 535550 994472 535606 994528
rect 533710 994200 533766 994256
rect 551098 997872 551154 997908
rect 550270 997772 550272 997792
rect 550272 997772 550324 997792
rect 550324 997772 550326 997792
rect 550270 997736 550326 997772
rect 553950 1001988 553952 1002008
rect 553952 1001988 554004 1002008
rect 554004 1001988 554006 1002008
rect 553950 1001952 554006 1001988
rect 553122 998436 553178 998472
rect 553122 998416 553124 998436
rect 553124 998416 553176 998436
rect 553176 998416 553178 998436
rect 552294 997772 552296 997792
rect 552296 997772 552348 997792
rect 552348 997772 552350 997792
rect 552294 997736 552350 997772
rect 555146 1006868 555202 1006904
rect 555146 1006848 555148 1006868
rect 555148 1006848 555200 1006868
rect 555200 1006848 555202 1006868
rect 557170 1006732 557226 1006768
rect 557170 1006712 557172 1006732
rect 557172 1006712 557224 1006732
rect 557224 1006712 557226 1006732
rect 556802 1006460 556858 1006496
rect 556802 1006440 556804 1006460
rect 556804 1006440 556856 1006460
rect 556856 1006440 556858 1006460
rect 554318 1006324 554374 1006360
rect 554318 1006304 554320 1006324
rect 554320 1006304 554372 1006324
rect 554372 1006304 554374 1006324
rect 560850 1006188 560906 1006224
rect 560850 1006168 560852 1006188
rect 560852 1006168 560904 1006188
rect 560904 1006168 560906 1006188
rect 555146 1005388 555148 1005408
rect 555148 1005388 555200 1005408
rect 555200 1005388 555202 1005408
rect 555146 1005352 555202 1005388
rect 554318 1002260 554320 1002280
rect 554320 1002260 554372 1002280
rect 554372 1002260 554374 1002280
rect 554318 1002224 554374 1002260
rect 555974 1005660 555976 1005680
rect 555976 1005660 556028 1005680
rect 556028 1005660 556030 1005680
rect 555974 1005624 556030 1005660
rect 555974 1004828 556030 1004864
rect 555974 1004808 555976 1004828
rect 555976 1004808 556028 1004828
rect 556028 1004808 556030 1004828
rect 557630 1004692 557686 1004728
rect 557630 1004672 557632 1004692
rect 557632 1004672 557684 1004692
rect 557684 1004672 557686 1004692
rect 557998 1002652 558054 1002688
rect 557998 1002632 558000 1002652
rect 558000 1002632 558052 1002652
rect 558052 1002632 558054 1002652
rect 557998 1002396 558000 1002416
rect 558000 1002396 558052 1002416
rect 558052 1002396 558054 1002416
rect 557998 1002360 558054 1002396
rect 561678 1004692 561734 1004728
rect 561678 1004672 561680 1004692
rect 561680 1004672 561732 1004692
rect 561732 1004672 561734 1004692
rect 558826 1002788 558882 1002824
rect 558826 1002768 558828 1002788
rect 558828 1002768 558880 1002788
rect 558880 1002768 558882 1002788
rect 558826 1001972 558882 1002008
rect 558826 1001952 558828 1001972
rect 558828 1001952 558880 1001972
rect 558880 1001952 558882 1001972
rect 522946 993928 523002 993984
rect 536746 993928 536802 993984
rect 560022 1002124 560024 1002144
rect 560024 1002124 560076 1002144
rect 560076 1002124 560078 1002144
rect 560022 1002088 560078 1002124
rect 560482 1002260 560484 1002280
rect 560484 1002260 560536 1002280
rect 560536 1002260 560538 1002280
rect 560482 1002224 560538 1002260
rect 560850 1001988 560852 1002008
rect 560852 1001988 560904 1002008
rect 560904 1001988 560906 1002008
rect 560850 1001952 560906 1001988
rect 563702 995560 563758 995616
rect 570234 994744 570290 994800
rect 590566 996648 590622 996704
rect 590566 996376 590622 996432
rect 625250 995968 625306 996024
rect 625618 995696 625674 995752
rect 627182 995696 627238 995752
rect 627918 995696 627974 995752
rect 629758 995696 629814 995752
rect 630310 995424 630366 995480
rect 625618 995152 625674 995208
rect 634726 995152 634782 995208
rect 638866 994880 638922 994936
rect 637026 994744 637082 994800
rect 640798 994880 640854 994936
rect 62118 975976 62174 976032
rect 62118 962920 62174 962976
rect 62118 949864 62174 949920
rect 62118 936980 62120 937000
rect 62120 936980 62172 937000
rect 62172 936980 62174 937000
rect 62118 936944 62174 936980
rect 44822 936128 44878 936184
rect 44454 934088 44510 934144
rect 44178 933680 44234 933736
rect 42982 933272 43038 933328
rect 42430 932864 42486 932920
rect 42798 932048 42854 932104
rect 42430 881864 42486 881920
rect 42062 818624 42118 818680
rect 41878 817944 41934 818000
rect 41786 814000 41842 814056
rect 40774 812776 40830 812832
rect 35162 812368 35218 812424
rect 32402 811144 32458 811200
rect 31666 809920 31722 809976
rect 33782 809512 33838 809568
rect 40958 811960 41014 812016
rect 41326 811552 41382 811608
rect 41786 809240 41842 809296
rect 36542 809104 36598 809160
rect 35162 803800 35218 803856
rect 41326 807472 41382 807528
rect 41786 808288 41842 808344
rect 42062 806656 42118 806712
rect 41510 805024 41566 805080
rect 39762 802032 39818 802088
rect 40314 800672 40370 800728
rect 40590 800672 40646 800728
rect 41786 800264 41842 800320
rect 41786 799856 41842 799912
rect 42706 802032 42762 802088
rect 42062 797272 42118 797328
rect 41786 796184 41842 796240
rect 41786 794416 41842 794472
rect 41786 793464 41842 793520
rect 43258 813592 43314 813648
rect 43074 808696 43130 808752
rect 42062 790608 42118 790664
rect 42430 791560 42486 791616
rect 42246 789928 42302 789984
rect 42614 790200 42670 790256
rect 42246 788160 42302 788216
rect 42522 787888 42578 787944
rect 40038 774968 40094 775024
rect 35806 774324 35808 774344
rect 35808 774324 35860 774344
rect 35860 774324 35862 774344
rect 35806 774288 35862 774324
rect 35806 773880 35862 773936
rect 35346 773472 35402 773528
rect 35530 773064 35586 773120
rect 35806 773100 35808 773120
rect 35808 773100 35860 773120
rect 35860 773100 35862 773120
rect 35806 773064 35862 773100
rect 40866 773064 40922 773120
rect 42982 790608 43038 790664
rect 43074 773064 43130 773120
rect 35346 772248 35402 772304
rect 39762 772248 39818 772304
rect 42798 772248 42854 772304
rect 35530 771876 35532 771896
rect 35532 771876 35584 771896
rect 35584 771876 35586 771896
rect 35530 771840 35586 771876
rect 35714 771432 35770 771488
rect 39118 771452 39174 771488
rect 39118 771432 39120 771452
rect 39120 771432 39172 771452
rect 39172 771432 39174 771452
rect 35438 771024 35494 771080
rect 39854 771024 39910 771080
rect 42890 771024 42946 771080
rect 35622 770616 35678 770672
rect 35806 770208 35862 770264
rect 41418 770208 41474 770264
rect 35346 769392 35402 769448
rect 35530 768984 35586 769040
rect 35806 769004 35862 769040
rect 35806 768984 35808 769004
rect 35808 768984 35860 769004
rect 35860 768984 35862 769004
rect 35806 767760 35862 767816
rect 32402 767352 32458 767408
rect 35162 766944 35218 767000
rect 32402 759600 32458 759656
rect 35806 766536 35862 766592
rect 35806 766128 35862 766184
rect 35806 764496 35862 764552
rect 35622 764088 35678 764144
rect 35806 763700 35862 763736
rect 35806 763680 35808 763700
rect 35808 763680 35860 763700
rect 35860 763680 35862 763700
rect 35806 762864 35862 762920
rect 39854 768576 39910 768632
rect 42706 768576 42762 768632
rect 42246 768304 42302 768360
rect 40406 766164 40408 766184
rect 40408 766164 40460 766184
rect 40460 766164 40462 766184
rect 40406 766128 40462 766164
rect 40406 764496 40462 764552
rect 41510 763292 41566 763328
rect 41510 763272 41512 763292
rect 41512 763272 41564 763292
rect 41564 763272 41566 763292
rect 40498 760280 40554 760336
rect 40406 758276 40408 758296
rect 40408 758276 40460 758296
rect 40460 758276 40462 758296
rect 40406 758240 40462 758276
rect 39302 757696 39358 757752
rect 42430 758240 42486 758296
rect 41418 757288 41474 757344
rect 41786 756608 41842 756664
rect 42062 754024 42118 754080
rect 42062 752936 42118 752992
rect 42246 751576 42302 751632
rect 41786 751032 41842 751088
rect 41786 750352 41842 750408
rect 42614 750488 42670 750544
rect 42430 749400 42486 749456
rect 42246 745592 42302 745648
rect 41786 743688 41842 743744
rect 42430 745048 42486 745104
rect 42430 730904 42486 730960
rect 41142 730496 41198 730552
rect 43258 766128 43314 766184
rect 43626 797272 43682 797328
rect 44454 814000 44510 814056
rect 44638 807880 44694 807936
rect 46202 819032 46258 819088
rect 46202 806248 46258 806304
rect 44822 774968 44878 775024
rect 44178 771432 44234 771488
rect 44270 770208 44326 770264
rect 43442 754024 43498 754080
rect 43074 730088 43130 730144
rect 42890 729272 42946 729328
rect 40866 728626 40922 728682
rect 43074 728048 43130 728104
rect 41050 727402 41106 727458
rect 41326 727456 41382 727458
rect 41326 727404 41328 727456
rect 41328 727404 41380 727456
rect 41380 727404 41382 727456
rect 41326 727402 41382 727404
rect 41142 726824 41198 726880
rect 40958 726178 41014 726234
rect 37922 725192 37978 725248
rect 35162 724784 35218 724840
rect 33046 724376 33102 724432
rect 31758 720316 31814 720352
rect 31758 720296 31760 720316
rect 31760 720296 31812 720316
rect 31812 720296 31814 720316
rect 33782 723730 33838 723786
rect 33046 716760 33102 716816
rect 40682 723152 40738 723208
rect 39210 715128 39266 715184
rect 41326 726232 41382 726234
rect 41326 726180 41328 726232
rect 41328 726180 41380 726232
rect 41380 726180 41382 726232
rect 41326 726178 41382 726180
rect 41786 725736 41842 725792
rect 41326 725600 41382 725656
rect 41142 721712 41198 721768
rect 41786 722336 41842 722392
rect 41786 718528 41842 718584
rect 41326 714448 41382 714504
rect 40038 714176 40094 714232
rect 41510 714176 41566 714232
rect 42338 715128 42394 715184
rect 42522 715128 42578 715184
rect 41786 713904 41842 713960
rect 42522 714448 42578 714504
rect 41786 712136 41842 712192
rect 42154 711592 42210 711648
rect 42246 710368 42302 710424
rect 42246 709144 42302 709200
rect 41786 708464 41842 708520
rect 42062 707784 42118 707840
rect 42430 707240 42486 707296
rect 42062 706560 42118 706616
rect 42614 702480 42670 702536
rect 42430 701392 42486 701448
rect 42246 701120 42302 701176
rect 40958 688336 41014 688392
rect 42522 687248 42578 687304
rect 41142 686840 41198 686896
rect 40866 685854 40922 685910
rect 41326 685854 41382 685910
rect 41142 685208 41198 685264
rect 40774 684630 40830 684686
rect 41142 683984 41198 684040
rect 40958 683576 41014 683632
rect 34426 682352 34482 682408
rect 41326 683168 41382 683224
rect 41326 682760 41382 682816
rect 41786 682352 41842 682408
rect 32402 681128 32458 681184
rect 31022 680720 31078 680776
rect 40682 681944 40738 682000
rect 36542 681536 36598 681592
rect 32402 672696 32458 672752
rect 41786 680312 41842 680368
rect 41142 677048 41198 677104
rect 40682 675552 40738 675608
rect 42062 676640 42118 676696
rect 42062 675588 42064 675608
rect 42064 675588 42116 675608
rect 42116 675588 42118 675608
rect 42062 675552 42118 675588
rect 41142 672424 41198 672480
rect 42338 672424 42394 672480
rect 40406 671200 40462 671256
rect 39762 670928 39818 670984
rect 43258 723560 43314 723616
rect 43442 719888 43498 719944
rect 43442 687656 43498 687712
rect 43074 684528 43130 684584
rect 42614 667936 42670 667992
rect 42154 667664 42210 667720
rect 42430 667392 42486 667448
rect 42154 666304 42210 666360
rect 41970 663992 42026 664048
rect 42062 662768 42118 662824
rect 42706 659640 42762 659696
rect 42430 658552 42486 658608
rect 42154 658280 42210 658336
rect 38842 646040 38898 646096
rect 41234 645632 41290 645688
rect 35530 644680 35586 644736
rect 35806 644716 35808 644736
rect 35808 644716 35860 644736
rect 35860 644716 35862 644736
rect 35806 644680 35862 644716
rect 39670 644680 39726 644736
rect 35346 643864 35402 643920
rect 35530 643456 35586 643512
rect 35806 643492 35808 643512
rect 35808 643492 35860 643512
rect 35860 643492 35862 643512
rect 35806 643456 35862 643492
rect 35438 642640 35494 642696
rect 35622 642232 35678 642288
rect 39026 642252 39082 642288
rect 39026 642232 39028 642252
rect 39028 642232 39080 642252
rect 39080 642232 39082 642252
rect 35806 641824 35862 641880
rect 35346 641416 35402 641472
rect 39762 641416 39818 641472
rect 35530 641008 35586 641064
rect 35806 641008 35862 641064
rect 40314 641008 40370 641064
rect 43258 680584 43314 680640
rect 43442 678272 43498 678328
rect 43810 752936 43866 752992
rect 44822 760280 44878 760336
rect 44362 722744 44418 722800
rect 44362 707784 44418 707840
rect 43626 667664 43682 667720
rect 43074 642232 43130 642288
rect 39854 640192 39910 640248
rect 42890 640192 42946 640248
rect 34426 639784 34482 639840
rect 33782 638560 33838 638616
rect 32402 638152 32458 638208
rect 35530 639376 35586 639432
rect 35806 639376 35862 639432
rect 35530 637744 35586 637800
rect 35806 637764 35862 637800
rect 35806 637744 35808 637764
rect 35808 637744 35860 637764
rect 35860 637744 35862 637764
rect 40038 637336 40094 637392
rect 35806 636520 35862 636576
rect 41510 637764 41566 637800
rect 41510 637744 41512 637764
rect 41512 637744 41564 637764
rect 41564 637744 41566 637764
rect 41326 636112 41382 636168
rect 35622 635296 35678 635352
rect 40222 635296 40278 635352
rect 35806 634888 35862 634944
rect 39762 634888 39818 634944
rect 35622 634480 35678 634536
rect 35806 633684 35862 633720
rect 35806 633664 35808 633684
rect 35808 633664 35860 633684
rect 35860 633664 35862 633684
rect 42338 633800 42394 633856
rect 39302 631352 39358 631408
rect 42706 626728 42762 626784
rect 42154 623328 42210 623384
rect 41970 621424 42026 621480
rect 41970 620200 42026 620256
rect 42246 619792 42302 619848
rect 42430 618976 42486 619032
rect 42706 618704 42762 618760
rect 42246 615984 42302 616040
rect 41786 612720 41842 612776
rect 35806 601724 35862 601760
rect 35806 601704 35808 601724
rect 35808 601704 35860 601724
rect 35860 601704 35862 601724
rect 42614 600888 42670 600944
rect 41326 599256 41382 599312
rect 40866 598440 40922 598496
rect 41050 597794 41106 597850
rect 41326 597848 41382 597850
rect 41326 597796 41328 597848
rect 41328 597796 41380 597848
rect 41380 597796 41382 597848
rect 41326 597794 41382 597796
rect 41142 597216 41198 597272
rect 41326 596808 41382 596864
rect 41326 595992 41382 596048
rect 41786 595992 41842 596048
rect 33046 595584 33102 595640
rect 31022 594360 31078 594416
rect 35162 595176 35218 595232
rect 34426 594768 34482 594824
rect 34426 587152 34482 587208
rect 36542 593544 36598 593600
rect 41786 593952 41842 594008
rect 39946 590688 40002 590744
rect 41786 592864 41842 592920
rect 41786 592320 41842 592376
rect 40774 589600 40830 589656
rect 41786 589464 41842 589520
rect 40590 589328 40646 589384
rect 43166 598848 43222 598904
rect 40130 584840 40186 584896
rect 41418 584840 41474 584896
rect 39394 584568 39450 584624
rect 41602 584568 41658 584624
rect 41786 584296 41842 584352
rect 41786 583888 41842 583944
rect 41970 582528 42026 582584
rect 42154 581168 42210 581224
rect 41786 580216 41842 580272
rect 42246 579944 42302 580000
rect 42614 580488 42670 580544
rect 42062 578176 42118 578232
rect 42338 576544 42394 576600
rect 42062 575592 42118 575648
rect 41786 574640 41842 574696
rect 42706 573960 42762 574016
rect 42246 572192 42302 572248
rect 42430 571920 42486 571976
rect 43258 593136 43314 593192
rect 44270 686432 44326 686488
rect 43810 645632 43866 645688
rect 44638 679904 44694 679960
rect 44638 666304 44694 666360
rect 44454 644680 44510 644736
rect 44270 641416 44326 641472
rect 43994 636112 44050 636168
rect 43810 634888 43866 634944
rect 43994 623328 44050 623384
rect 43442 581168 43498 581224
rect 43258 578176 43314 578232
rect 41326 557676 41328 557696
rect 41328 557676 41380 557696
rect 41380 557676 41382 557696
rect 41326 557640 41382 557676
rect 40590 556008 40646 556064
rect 41142 555600 41198 555656
rect 42798 555192 42854 555248
rect 41050 555022 41106 555078
rect 40038 553352 40094 553408
rect 40958 553352 41014 553408
rect 29642 551928 29698 551984
rect 43442 558048 43498 558104
rect 43166 554376 43222 554432
rect 41878 549888 41934 549944
rect 31758 547460 31814 547496
rect 31758 547440 31760 547460
rect 31760 547440 31812 547460
rect 31812 547440 31814 547460
rect 41326 546352 41382 546408
rect 42062 549480 42118 549536
rect 41878 545536 41934 545592
rect 42338 548256 42394 548312
rect 42062 545264 42118 545320
rect 42706 549072 42762 549128
rect 42246 538192 42302 538248
rect 42062 537920 42118 537976
rect 42430 536968 42486 537024
rect 42246 533296 42302 533352
rect 42430 532616 42486 532672
rect 42614 529760 42670 529816
rect 41786 527584 41842 527640
rect 40682 522688 40738 522744
rect 42522 522688 42578 522744
rect 40682 431160 40738 431216
rect 41326 430480 41382 430536
rect 41142 430072 41198 430128
rect 42890 431160 42946 431216
rect 40958 429426 41014 429482
rect 41326 429426 41382 429482
rect 42982 428168 43038 428224
rect 41142 427624 41198 427680
rect 41142 425992 41198 426048
rect 40774 425176 40830 425232
rect 40774 418376 40830 418432
rect 41970 424360 42026 424416
rect 41142 417968 41198 418024
rect 42798 423136 42854 423192
rect 42246 419872 42302 419928
rect 42614 419464 42670 419520
rect 42430 417968 42486 418024
rect 41786 407496 41842 407552
rect 41786 403824 41842 403880
rect 43442 547032 43498 547088
rect 44086 600072 44142 600128
rect 44638 641008 44694 641064
rect 44454 637744 44510 637800
rect 44638 600480 44694 600536
rect 44270 599664 44326 599720
rect 43810 591504 43866 591560
rect 43810 558456 43866 558512
rect 44178 557232 44234 557288
rect 44638 591912 44694 591968
rect 44638 556824 44694 556880
rect 44454 556416 44510 556472
rect 43810 551520 43866 551576
rect 43626 537920 43682 537976
rect 43994 550704 44050 550760
rect 43166 427216 43222 427272
rect 43350 423544 43406 423600
rect 43166 422728 43222 422784
rect 41786 401920 41842 401976
rect 41786 400016 41842 400072
rect 41786 398792 41842 398848
rect 35346 387504 35402 387560
rect 39946 387524 40002 387560
rect 39946 387504 39948 387524
rect 39948 387504 40000 387524
rect 40000 387504 40002 387524
rect 35530 387096 35586 387152
rect 35806 387096 35862 387152
rect 40130 387096 40186 387152
rect 40314 386688 40370 386744
rect 35806 386280 35862 386336
rect 35346 385872 35402 385928
rect 35530 385464 35586 385520
rect 35806 385484 35862 385520
rect 35806 385464 35808 385484
rect 35808 385464 35860 385484
rect 35860 385464 35862 385484
rect 43626 387504 43682 387560
rect 39578 385056 39634 385112
rect 43074 385056 43130 385112
rect 35622 384648 35678 384704
rect 35806 384240 35862 384296
rect 35806 383832 35862 383888
rect 39670 383832 39726 383888
rect 35346 383424 35402 383480
rect 35530 383016 35586 383072
rect 35806 383016 35862 383072
rect 35806 382200 35862 382256
rect 40038 382200 40094 382256
rect 35622 381792 35678 381848
rect 32402 381384 32458 381440
rect 28814 376488 28870 376544
rect 35806 381384 35862 381440
rect 35622 380568 35678 380624
rect 39854 380568 39910 380624
rect 35438 380160 35494 380216
rect 35806 380160 35862 380216
rect 40038 380160 40094 380216
rect 35806 378936 35862 378992
rect 35622 377712 35678 377768
rect 41418 381792 41474 381848
rect 41050 379752 41106 379808
rect 42798 380568 42854 380624
rect 40222 378936 40278 378992
rect 41510 378120 41566 378176
rect 39762 377712 39818 377768
rect 35806 377304 35862 377360
rect 39578 377304 39634 377360
rect 41510 376932 41512 376952
rect 41512 376932 41564 376952
rect 41564 376932 41566 376952
rect 41510 376896 41566 376932
rect 35806 376080 35862 376136
rect 42062 369688 42118 369744
rect 41786 365608 41842 365664
rect 42062 364928 42118 364984
rect 41786 363704 41842 363760
rect 42798 369688 42854 369744
rect 41786 360576 41842 360632
rect 41878 358672 41934 358728
rect 41786 356904 41842 356960
rect 41970 355680 42026 355736
rect 40406 345752 40462 345808
rect 39762 344936 39818 344992
rect 39578 344664 39634 344720
rect 35346 344256 35402 344312
rect 35622 344256 35678 344312
rect 35806 343848 35862 343904
rect 39578 343440 39634 343496
rect 35346 343032 35402 343088
rect 35530 342624 35586 342680
rect 35806 342660 35808 342680
rect 35808 342660 35860 342680
rect 35860 342660 35862 342680
rect 35806 342624 35862 342660
rect 35622 341808 35678 341864
rect 43442 377712 43498 377768
rect 43626 377304 43682 377360
rect 44270 428848 44326 428904
rect 44178 426808 44234 426864
rect 43994 387096 44050 387152
rect 43994 383832 44050 383888
rect 44362 421232 44418 421288
rect 44178 381792 44234 381848
rect 43994 344936 44050 344992
rect 43810 344664 43866 344720
rect 43258 343440 43314 343496
rect 39946 343032 40002 343088
rect 42982 343032 43038 343088
rect 40314 342252 40316 342272
rect 40316 342252 40368 342272
rect 40368 342252 40370 342272
rect 40314 342216 40370 342252
rect 43258 342216 43314 342272
rect 35806 341436 35808 341456
rect 35808 341436 35860 341456
rect 35860 341436 35862 341456
rect 35806 341400 35862 341436
rect 35622 341028 35624 341048
rect 35624 341028 35676 341048
rect 35676 341028 35678 341048
rect 35622 340992 35678 341028
rect 40314 340992 40370 341048
rect 42890 340992 42946 341048
rect 35806 340584 35862 340640
rect 35622 340176 35678 340232
rect 35622 338952 35678 339008
rect 39578 338952 39634 339008
rect 35806 338544 35862 338600
rect 41510 338136 41566 338192
rect 35806 337728 35862 337784
rect 35530 336932 35586 336968
rect 35530 336912 35532 336932
rect 35532 336912 35584 336932
rect 35584 336912 35586 336932
rect 35806 336912 35862 336968
rect 40038 336912 40094 336968
rect 35622 336096 35678 336152
rect 35806 335688 35862 335744
rect 39670 335316 39672 335336
rect 39672 335316 39724 335336
rect 39724 335316 39726 335336
rect 39670 335280 39726 335316
rect 35438 334872 35494 334928
rect 35806 334872 35862 334928
rect 40314 334872 40370 334928
rect 35622 334464 35678 334520
rect 39578 334092 39580 334112
rect 39580 334092 39632 334112
rect 39632 334092 39634 334112
rect 39578 334056 39634 334092
rect 40314 333648 40370 333704
rect 35622 333240 35678 333296
rect 35806 332832 35862 332888
rect 39578 330520 39634 330576
rect 41786 324808 41842 324864
rect 41786 322768 41842 322824
rect 41786 315560 41842 315616
rect 41786 313656 41842 313712
rect 41786 312976 41842 313032
rect 41142 299240 41198 299296
rect 40958 298424 41014 298480
rect 42706 298832 42762 298888
rect 40958 298016 41014 298072
rect 42062 295568 42118 295624
rect 41786 295160 41842 295216
rect 41786 294888 41842 294944
rect 35162 294752 35218 294808
rect 41786 293528 41842 293584
rect 40498 292544 40500 292588
rect 40500 292544 40552 292588
rect 40552 292544 40554 292588
rect 40498 292532 40554 292544
rect 42062 292304 42118 292360
rect 41142 290672 41198 290728
rect 40958 290264 41014 290320
rect 41786 289992 41842 290048
rect 41326 289772 41382 289828
rect 44546 378120 44602 378176
rect 44362 376896 44418 376952
rect 44362 364928 44418 364984
rect 44178 338952 44234 339008
rect 43442 336912 43498 336968
rect 43626 334872 43682 334928
rect 43258 300056 43314 300112
rect 43258 297200 43314 297256
rect 43074 293936 43130 293992
rect 42890 291080 42946 291136
rect 41970 281424 42026 281480
rect 42246 277888 42302 277944
rect 41786 277344 41842 277400
rect 42062 277072 42118 277128
rect 42062 276528 42118 276584
rect 41786 273400 41842 273456
rect 41786 272312 41842 272368
rect 41786 270408 41842 270464
rect 40038 259392 40094 259448
rect 40406 258848 40462 258904
rect 35806 258032 35862 258088
rect 39578 257896 39634 257952
rect 35622 257488 35678 257544
rect 39946 257488 40002 257544
rect 35806 257116 35808 257136
rect 35808 257116 35860 257136
rect 35860 257116 35862 257136
rect 35806 257080 35862 257116
rect 35806 256672 35862 256728
rect 35806 256264 35862 256320
rect 35622 255856 35678 255912
rect 35806 255448 35862 255504
rect 35346 255040 35402 255096
rect 35162 254632 35218 254688
rect 35530 254224 35586 254280
rect 35806 254260 35808 254280
rect 35808 254260 35860 254280
rect 35860 254260 35862 254280
rect 35806 254224 35862 254260
rect 35806 253408 35862 253464
rect 35622 253000 35678 253056
rect 40314 256672 40370 256728
rect 43258 257488 43314 257544
rect 41418 255040 41474 255096
rect 39302 253000 39358 253056
rect 42890 253000 42946 253056
rect 35806 252612 35862 252648
rect 35806 252592 35808 252612
rect 35808 252592 35860 252612
rect 35860 252592 35862 252612
rect 41510 252612 41566 252648
rect 41510 252592 41512 252612
rect 41512 252592 41564 252612
rect 41564 252592 41566 252612
rect 35806 252184 35862 252240
rect 40590 252184 40646 252240
rect 35622 251776 35678 251832
rect 41326 251776 41382 251832
rect 35806 251388 35862 251424
rect 35806 251368 35808 251388
rect 35808 251368 35860 251388
rect 35860 251368 35862 251388
rect 41510 251368 41566 251424
rect 35438 250960 35494 251016
rect 35622 250552 35678 250608
rect 35806 250180 35808 250200
rect 35808 250180 35860 250200
rect 35860 250180 35862 250200
rect 35806 250144 35862 250180
rect 39394 250180 39396 250200
rect 39396 250180 39448 250200
rect 39448 250180 39450 250200
rect 39394 250144 39450 250180
rect 35530 248920 35586 248976
rect 35806 248920 35862 248976
rect 35622 248104 35678 248160
rect 35438 247696 35494 247752
rect 35806 247288 35862 247344
rect 35622 246880 35678 246936
rect 40130 248920 40186 248976
rect 39946 248512 40002 248568
rect 40130 248104 40186 248160
rect 41510 247696 41566 247752
rect 40130 247324 40132 247344
rect 40132 247324 40184 247344
rect 40184 247324 40186 247344
rect 40130 247288 40186 247324
rect 41510 246880 41566 246936
rect 41050 246064 41106 246120
rect 39578 245520 39634 245576
rect 42522 252184 42578 252240
rect 42154 247696 42210 247752
rect 42062 246880 42118 246936
rect 42246 238448 42302 238504
rect 41786 236544 41842 236600
rect 41786 234504 41842 234560
rect 42706 237360 42762 237416
rect 42062 227296 42118 227352
rect 41694 223624 41750 223680
rect 40682 222536 40738 222592
rect 28538 222264 28594 222320
rect 39762 218320 39818 218376
rect 40222 218048 40278 218104
rect 35346 214648 35402 214704
rect 35530 214240 35586 214296
rect 35806 214276 35808 214296
rect 35808 214276 35860 214296
rect 35860 214276 35862 214296
rect 35806 214240 35862 214276
rect 39762 214240 39818 214296
rect 35806 213424 35862 213480
rect 35622 213016 35678 213072
rect 28538 212608 28594 212664
rect 39302 213036 39358 213072
rect 39302 213016 39304 213036
rect 39304 213016 39356 213036
rect 39356 213016 39358 213036
rect 35806 212644 35808 212664
rect 35808 212644 35860 212664
rect 35860 212644 35862 212664
rect 35806 212608 35862 212644
rect 41234 212628 41290 212664
rect 41234 212608 41236 212628
rect 41236 212608 41288 212628
rect 41288 212608 41290 212628
rect 41050 212200 41106 212256
rect 35806 211792 35862 211848
rect 35622 211384 35678 211440
rect 39670 211404 39726 211440
rect 39670 211384 39672 211404
rect 39672 211384 39724 211404
rect 39724 211384 39726 211404
rect 41234 211792 41290 211848
rect 35806 210976 35862 211032
rect 35622 210568 35678 210624
rect 35806 210160 35862 210216
rect 42614 222536 42670 222592
rect 42154 212644 42156 212664
rect 42156 212644 42208 212664
rect 42208 212644 42210 212664
rect 42154 212608 42210 212644
rect 43074 250144 43130 250200
rect 43258 248920 43314 248976
rect 43994 335280 44050 335336
rect 43810 301552 43866 301608
rect 44638 334056 44694 334112
rect 44454 333648 44510 333704
rect 44546 299648 44602 299704
rect 44178 297608 44234 297664
rect 43994 293120 44050 293176
rect 43810 289992 43866 290048
rect 44178 291760 44234 291816
rect 44362 291488 44418 291544
rect 44178 277072 44234 277128
rect 44546 258848 44602 258904
rect 43626 257896 43682 257952
rect 44178 255040 44234 255096
rect 43626 248512 43682 248568
rect 43626 224984 43682 225040
rect 43442 218320 43498 218376
rect 43626 212200 43682 212256
rect 44546 248104 44602 248160
rect 44362 247288 44418 247344
rect 45190 764496 45246 764552
rect 45006 729680 45062 729736
rect 45190 728864 45246 728920
rect 45190 679496 45246 679552
rect 45006 677864 45062 677920
rect 45190 631352 45246 631408
rect 45558 552336 45614 552392
rect 45190 551112 45246 551168
rect 45374 548664 45430 548720
rect 45558 424768 45614 424824
rect 45374 421504 45430 421560
rect 45190 420688 45246 420744
rect 45374 379752 45430 379808
rect 45190 345752 45246 345808
rect 45558 330520 45614 330576
rect 45374 300872 45430 300928
rect 45558 295976 45614 296032
rect 45742 294888 45798 294944
rect 45926 294344 45982 294400
rect 45742 276528 45798 276584
rect 45190 256672 45246 256728
rect 45190 251776 45246 251832
rect 45006 229744 45062 229800
rect 45834 251368 45890 251424
rect 46018 246064 46074 246120
rect 46018 238448 46074 238504
rect 47582 763272 47638 763328
rect 46386 721112 46442 721168
rect 46938 423952 46994 424008
rect 47030 338136 47086 338192
rect 46754 259392 46810 259448
rect 46938 252592 46994 252648
rect 46386 227432 46442 227488
rect 47122 245520 47178 245576
rect 47766 731312 47822 731368
rect 47766 646040 47822 646096
rect 47766 601296 47822 601352
rect 47766 590280 47822 590336
rect 47950 386688 48006 386744
rect 48134 300464 48190 300520
rect 47766 226888 47822 226944
rect 47582 221584 47638 221640
rect 45558 214240 45614 214296
rect 44178 213016 44234 213072
rect 43810 211792 43866 211848
rect 42890 211384 42946 211440
rect 35622 209344 35678 209400
rect 30286 208936 30342 208992
rect 35806 208936 35862 208992
rect 39670 208564 39672 208584
rect 39672 208564 39724 208584
rect 39724 208564 39726 208584
rect 39670 208528 39726 208564
rect 35530 207304 35586 207360
rect 35806 207324 35862 207360
rect 35806 207304 35808 207324
rect 35808 207304 35860 207324
rect 35860 207304 35862 207324
rect 35622 206488 35678 206544
rect 35806 206080 35862 206136
rect 35622 205264 35678 205320
rect 35806 204876 35862 204912
rect 35806 204856 35808 204876
rect 35808 204856 35860 204876
rect 35860 204856 35862 204876
rect 39762 206896 39818 206952
rect 43074 208528 43130 208584
rect 40038 205672 40094 205728
rect 39578 205264 39634 205320
rect 42890 206896 42946 206952
rect 40314 204856 40370 204912
rect 35530 204468 35586 204504
rect 35530 204448 35532 204468
rect 35532 204448 35584 204468
rect 35584 204448 35586 204468
rect 35806 204448 35862 204504
rect 39394 204448 39450 204504
rect 39946 204040 40002 204096
rect 35622 203632 35678 203688
rect 41142 203632 41198 203688
rect 35806 203224 35862 203280
rect 41234 203244 41290 203280
rect 41234 203224 41236 203244
rect 41236 203224 41288 203244
rect 41288 203224 41290 203244
rect 30286 200640 30342 200696
rect 41786 197104 41842 197160
rect 44178 205264 44234 205320
rect 43258 204856 43314 204912
rect 41786 195200 41842 195256
rect 41786 191528 41842 191584
rect 43442 204448 43498 204504
rect 43626 203632 43682 203688
rect 43810 203224 43866 203280
rect 41786 185816 41842 185872
rect 41786 184048 41842 184104
rect 48962 278024 49018 278080
rect 50342 228520 50398 228576
rect 50526 228248 50582 228304
rect 53470 276664 53526 276720
rect 62118 923752 62174 923808
rect 62118 910696 62174 910752
rect 62118 897776 62174 897832
rect 62118 884740 62174 884776
rect 62118 884720 62120 884740
rect 62120 884720 62172 884740
rect 62172 884720 62174 884740
rect 62118 871664 62174 871720
rect 62118 858608 62174 858664
rect 62118 845552 62174 845608
rect 62118 832496 62174 832552
rect 62118 819440 62174 819496
rect 62118 806520 62174 806576
rect 62118 793620 62174 793656
rect 62118 793600 62120 793620
rect 62120 793600 62172 793620
rect 62172 793600 62174 793620
rect 62118 780408 62174 780464
rect 54850 265512 54906 265568
rect 54666 230016 54722 230072
rect 52090 227160 52146 227216
rect 62118 767372 62174 767408
rect 62118 767352 62120 767372
rect 62120 767352 62172 767372
rect 62172 767352 62174 767372
rect 62118 754296 62174 754352
rect 62118 741240 62174 741296
rect 62118 728184 62174 728240
rect 62118 715264 62174 715320
rect 62118 702208 62174 702264
rect 62118 689152 62174 689208
rect 62118 676096 62174 676152
rect 62118 663040 62174 663096
rect 62118 649984 62174 650040
rect 62118 637064 62174 637120
rect 62118 624008 62174 624064
rect 62118 610952 62174 611008
rect 62118 597896 62174 597952
rect 62118 584840 62174 584896
rect 62118 571784 62174 571840
rect 62118 558728 62174 558784
rect 62118 545808 62174 545864
rect 62762 532752 62818 532808
rect 62118 519696 62174 519752
rect 62118 506640 62174 506696
rect 62118 493584 62174 493640
rect 62118 480528 62174 480584
rect 62118 467472 62174 467528
rect 62762 454552 62818 454608
rect 62118 441496 62174 441552
rect 62118 428440 62174 428496
rect 62118 415420 62120 415440
rect 62120 415420 62172 415440
rect 62172 415420 62174 415440
rect 62118 415384 62174 415420
rect 62118 402328 62174 402384
rect 62118 389292 62174 389328
rect 62118 389272 62120 389292
rect 62120 389272 62172 389292
rect 62172 389272 62174 389292
rect 62118 376216 62174 376272
rect 62946 363296 63002 363352
rect 62762 350240 62818 350296
rect 62118 337184 62174 337240
rect 62118 324128 62174 324184
rect 62118 311072 62174 311128
rect 62118 298172 62174 298208
rect 62118 298152 62120 298172
rect 62120 298152 62172 298172
rect 62172 298152 62174 298172
rect 62762 285096 62818 285152
rect 56046 276936 56102 276992
rect 55862 226616 55918 226672
rect 50342 223896 50398 223952
rect 47950 218048 48006 218104
rect 44546 204040 44602 204096
rect 50986 219952 51042 220008
rect 54206 219700 54262 219736
rect 54206 219680 54208 219700
rect 54208 219680 54260 219700
rect 54260 219680 54262 219700
rect 58990 225528 59046 225584
rect 364154 267688 364210 267744
rect 366362 267688 366418 267744
rect 377678 267416 377734 267472
rect 379518 267416 379574 267472
rect 382186 269592 382242 269648
rect 384946 270272 385002 270328
rect 386602 270308 386604 270328
rect 386604 270308 386656 270328
rect 386656 270308 386658 270328
rect 386602 270272 386658 270308
rect 384486 269628 384488 269648
rect 384488 269628 384540 269648
rect 384540 269628 384542 269648
rect 384486 269592 384542 269628
rect 383658 267008 383714 267064
rect 384670 267028 384726 267064
rect 384670 267008 384672 267028
rect 384672 267008 384724 267028
rect 384724 267008 384726 267028
rect 388994 267008 389050 267064
rect 393410 269184 393466 269240
rect 393318 267028 393374 267064
rect 393318 267008 393320 267028
rect 393320 267008 393372 267028
rect 393372 267008 393374 267028
rect 400126 269728 400182 269784
rect 401138 267144 401194 267200
rect 402426 269184 402482 269240
rect 402610 267144 402666 267200
rect 403990 270580 403992 270600
rect 403992 270580 404044 270600
rect 404044 270580 404046 270600
rect 403990 270544 404046 270580
rect 408498 270544 408554 270600
rect 409510 270408 409566 270464
rect 412086 270716 412088 270736
rect 412088 270716 412140 270736
rect 412140 270716 412142 270736
rect 412086 270680 412142 270716
rect 412638 271088 412694 271144
rect 412730 270680 412786 270736
rect 412454 270408 412510 270464
rect 412454 270000 412510 270056
rect 412730 270000 412786 270056
rect 411994 267572 412050 267608
rect 411994 267552 411996 267572
rect 411996 267552 412048 267572
rect 412048 267552 412050 267572
rect 412730 267572 412786 267608
rect 412730 267552 412732 267572
rect 412732 267552 412784 267572
rect 412784 267552 412786 267572
rect 412638 267280 412694 267336
rect 415490 267824 415546 267880
rect 415122 267552 415178 267608
rect 417238 270544 417294 270600
rect 416318 267280 416374 267336
rect 417054 268096 417110 268152
rect 418986 271088 419042 271144
rect 418894 270680 418950 270736
rect 418250 270544 418306 270600
rect 418066 268096 418122 268152
rect 417790 267844 417846 267880
rect 417790 267824 417792 267844
rect 417792 267824 417844 267844
rect 417844 267824 417846 267844
rect 418342 267708 418398 267744
rect 418342 267688 418344 267708
rect 418344 267688 418396 267708
rect 418396 267688 418398 267708
rect 419262 267280 419318 267336
rect 420734 269456 420790 269512
rect 421102 267552 421158 267608
rect 423310 270716 423312 270736
rect 423312 270716 423364 270736
rect 423364 270716 423366 270736
rect 423310 270680 423366 270716
rect 424230 267552 424286 267608
rect 424966 267572 425022 267608
rect 424966 267552 424968 267572
rect 424968 267552 425020 267572
rect 425020 267552 425022 267572
rect 427818 272312 427874 272368
rect 427082 271940 427084 271960
rect 427084 271940 427136 271960
rect 427136 271940 427138 271960
rect 427082 271904 427138 271940
rect 427910 271904 427966 271960
rect 428186 271668 428188 271688
rect 428188 271668 428240 271688
rect 428240 271668 428242 271688
rect 428186 271632 428242 271668
rect 427818 270000 427874 270056
rect 427450 269456 427506 269512
rect 427634 269184 427690 269240
rect 428002 269184 428058 269240
rect 427634 268096 427690 268152
rect 427818 268096 427874 268152
rect 427910 267572 427966 267608
rect 427910 267552 427912 267572
rect 427912 267552 427964 267572
rect 427964 267552 427966 267572
rect 429382 271668 429384 271688
rect 429384 271668 429436 271688
rect 429436 271668 429438 271688
rect 429382 271632 429438 271668
rect 429106 271360 429162 271416
rect 428554 266872 428610 266928
rect 430946 272312 431002 272368
rect 431774 271632 431830 271688
rect 431406 270952 431462 271008
rect 429566 269456 429622 269512
rect 433154 272720 433210 272776
rect 432970 270988 432972 271008
rect 432972 270988 433024 271008
rect 433024 270988 433026 271008
rect 432970 270952 433026 270988
rect 434442 273944 434498 274000
rect 433522 271360 433578 271416
rect 433246 267688 433302 267744
rect 435362 273964 435418 274000
rect 435362 273944 435364 273964
rect 435364 273944 435416 273964
rect 435416 273944 435418 273964
rect 436926 273028 436928 273048
rect 436928 273028 436980 273048
rect 436980 273028 436982 273048
rect 436926 272992 436982 273028
rect 434810 270000 434866 270056
rect 436926 268368 436982 268424
rect 436558 267960 436614 268016
rect 435086 266192 435142 266248
rect 436742 266464 436798 266520
rect 438214 272992 438270 273048
rect 437294 272720 437350 272776
rect 437294 268660 437350 268696
rect 437294 268640 437296 268660
rect 437296 268640 437348 268660
rect 437348 268640 437350 268660
rect 437294 267688 437350 267744
rect 437294 266872 437350 266928
rect 437938 266464 437994 266520
rect 437754 266192 437810 266248
rect 441526 272040 441582 272096
rect 441158 271360 441214 271416
rect 439502 271088 439558 271144
rect 438858 268640 438914 268696
rect 441710 266348 441766 266384
rect 441710 266328 441712 266348
rect 441712 266328 441764 266348
rect 441764 266328 441766 266348
rect 442722 271360 442778 271416
rect 442998 267960 443054 268016
rect 442906 266348 442962 266384
rect 442906 266328 442908 266348
rect 442908 266328 442960 266348
rect 442960 266328 442962 266348
rect 443366 272076 443368 272096
rect 443368 272076 443420 272096
rect 443420 272076 443422 272096
rect 443366 272040 443422 272076
rect 445482 275440 445538 275496
rect 445390 272992 445446 273048
rect 444746 271088 444802 271144
rect 446770 272348 446772 272368
rect 446772 272348 446824 272368
rect 446824 272348 446826 272368
rect 446770 272312 446826 272348
rect 446126 271088 446182 271144
rect 446770 268640 446826 268696
rect 446770 267552 446826 267608
rect 446770 267028 446826 267064
rect 446770 267008 446772 267028
rect 446772 267008 446824 267028
rect 446824 267008 446826 267028
rect 446586 266736 446642 266792
rect 448150 273944 448206 274000
rect 447230 272992 447286 273048
rect 447414 272312 447470 272368
rect 447598 272312 447654 272368
rect 447414 267552 447470 267608
rect 447230 267008 447286 267064
rect 449714 273128 449770 273184
rect 448702 270136 448758 270192
rect 448518 268640 448574 268696
rect 451370 273964 451426 274000
rect 451370 273944 451372 273964
rect 451372 273944 451424 273964
rect 451424 273944 451426 273964
rect 450910 267008 450966 267064
rect 454590 274080 454646 274136
rect 454406 272348 454408 272368
rect 454408 272348 454460 272368
rect 454460 272348 454462 272368
rect 454406 272312 454462 272348
rect 456614 272720 456670 272776
rect 454774 266756 454830 266792
rect 454774 266736 454776 266756
rect 454776 266736 454828 266756
rect 454828 266736 454830 266756
rect 456614 271224 456670 271280
rect 456614 270544 456670 270600
rect 456614 270136 456670 270192
rect 456430 268912 456486 268968
rect 456614 267960 456670 268016
rect 457442 272756 457444 272776
rect 457444 272756 457496 272776
rect 457496 272756 457498 272776
rect 457442 272720 457498 272756
rect 458638 271904 458694 271960
rect 457442 270952 457498 271008
rect 457258 267008 457314 267064
rect 457166 266736 457222 266792
rect 460754 273672 460810 273728
rect 459926 270544 459982 270600
rect 459006 270272 459062 270328
rect 460938 273164 460940 273184
rect 460940 273164 460992 273184
rect 460992 273164 460994 273184
rect 460938 273128 460994 273164
rect 461582 275168 461638 275224
rect 461858 271224 461914 271280
rect 461030 268640 461086 268696
rect 461582 267960 461638 268016
rect 462778 271360 462834 271416
rect 462318 268912 462374 268968
rect 462502 268640 462558 268696
rect 461398 265784 461454 265840
rect 462778 266736 462834 266792
rect 463606 266736 463662 266792
rect 462686 266056 462742 266112
rect 462134 265784 462190 265840
rect 464894 272176 464950 272232
rect 466550 275188 466606 275224
rect 466550 275168 466552 275188
rect 466552 275168 466604 275188
rect 466604 275168 466606 275188
rect 466458 274896 466514 274952
rect 466412 274508 466468 274544
rect 466412 274488 466414 274508
rect 466414 274488 466466 274508
rect 466466 274488 466468 274508
rect 466550 273672 466606 273728
rect 466274 272448 466330 272504
rect 466274 271904 466330 271960
rect 466550 271396 466552 271416
rect 466552 271396 466604 271416
rect 466604 271396 466606 271416
rect 466550 271360 466606 271396
rect 466734 271360 466790 271416
rect 466274 269184 466330 269240
rect 466458 269184 466514 269240
rect 466734 268640 466790 268696
rect 466274 267008 466330 267064
rect 466734 267008 466790 267064
rect 466550 266736 466606 266792
rect 466550 266328 466606 266384
rect 469954 275984 470010 276040
rect 469770 274896 469826 274952
rect 469678 269184 469734 269240
rect 470506 275712 470562 275768
rect 471426 275712 471482 275768
rect 472162 274488 472218 274544
rect 472254 270680 472310 270736
rect 471426 268640 471482 268696
rect 473910 276004 473966 276040
rect 473910 275984 473912 276004
rect 473912 275984 473964 276004
rect 473964 275984 473966 276004
rect 473910 275712 473966 275768
rect 475750 277480 475806 277536
rect 475566 277208 475622 277264
rect 475750 276392 475806 276448
rect 475382 274488 475438 274544
rect 474094 268096 474150 268152
rect 473910 266328 473966 266384
rect 474646 267008 474702 267064
rect 476670 277480 476726 277536
rect 476394 277208 476450 277264
rect 476762 272720 476818 272776
rect 476762 272176 476818 272232
rect 475750 270036 475752 270056
rect 475752 270036 475804 270056
rect 475804 270036 475806 270056
rect 475750 270000 475806 270036
rect 476486 269184 476542 269240
rect 476670 269184 476726 269240
rect 476210 268096 476266 268152
rect 475750 267844 475806 267880
rect 475750 267824 475752 267844
rect 475752 267824 475804 267844
rect 475804 267824 475806 267844
rect 475750 267572 475806 267608
rect 475750 267552 475752 267572
rect 475752 267552 475804 267572
rect 475804 267552 475806 267572
rect 476118 267572 476174 267608
rect 476118 267552 476120 267572
rect 476120 267552 476172 267572
rect 476172 267552 476174 267572
rect 476302 267552 476358 267608
rect 476210 267008 476266 267064
rect 480994 275868 481050 275904
rect 480994 275848 480996 275868
rect 480996 275848 481048 275868
rect 481048 275848 481050 275868
rect 481270 275168 481326 275224
rect 480350 274508 480406 274544
rect 480350 274488 480352 274508
rect 480352 274488 480404 274508
rect 480404 274488 480406 274508
rect 477866 270000 477922 270056
rect 479982 270000 480038 270056
rect 479246 265240 479302 265296
rect 481454 274352 481510 274408
rect 644662 278024 644718 278080
rect 484122 275848 484178 275904
rect 484306 274896 484362 274952
rect 484122 269184 484178 269240
rect 482282 267552 482338 267608
rect 481822 265784 481878 265840
rect 483294 266464 483350 266520
rect 485870 276392 485926 276448
rect 486054 275984 486110 276040
rect 485870 275868 485926 275904
rect 485870 275848 485872 275868
rect 485872 275848 485924 275868
rect 485924 275848 485926 275868
rect 487342 275712 487398 275768
rect 486698 274896 486754 274952
rect 486698 274624 486754 274680
rect 486422 274352 486478 274408
rect 484858 270000 484914 270056
rect 484674 268912 484730 268968
rect 484858 268640 484914 268696
rect 485042 268096 485098 268152
rect 486882 274352 486938 274408
rect 487066 273808 487122 273864
rect 485870 272212 485872 272232
rect 485872 272212 485924 272232
rect 485924 272212 485926 272232
rect 485870 272176 485926 272212
rect 486054 272176 486110 272232
rect 485778 271904 485834 271960
rect 485870 271360 485926 271416
rect 485502 270952 485558 271008
rect 486882 270680 486938 270736
rect 486606 269184 486662 269240
rect 486422 268912 486478 268968
rect 486238 268640 486294 268696
rect 485686 267824 485742 267880
rect 486054 267960 486110 268016
rect 485870 267688 485926 267744
rect 485594 267008 485650 267064
rect 485594 265240 485650 265296
rect 488354 270000 488410 270056
rect 490746 275712 490802 275768
rect 492218 275984 492274 276040
rect 492586 275848 492642 275904
rect 488722 273828 488778 273864
rect 488722 273808 488724 273828
rect 488724 273808 488776 273828
rect 488776 273808 488778 273828
rect 489366 273808 489422 273864
rect 488538 269728 488594 269784
rect 491022 272720 491078 272776
rect 490194 268640 490250 268696
rect 491574 269184 491630 269240
rect 490010 267008 490066 267064
rect 490194 266872 490250 266928
rect 491574 267960 491630 268016
rect 491206 266892 491262 266928
rect 491206 266872 491208 266892
rect 491208 266872 491260 266892
rect 491260 266872 491262 266892
rect 493138 276392 493194 276448
rect 492954 271904 493010 271960
rect 494150 274896 494206 274952
rect 493966 270816 494022 270872
rect 493230 269184 493286 269240
rect 493046 268640 493102 268696
rect 492770 267708 492826 267744
rect 492770 267688 492772 267708
rect 492772 267688 492824 267708
rect 492824 267688 492826 267708
rect 492126 266736 492182 266792
rect 494978 274624 495034 274680
rect 495254 274644 495310 274680
rect 495254 274624 495256 274644
rect 495256 274624 495308 274644
rect 495308 274624 495310 274644
rect 495254 274352 495310 274408
rect 494886 273264 494942 273320
rect 495898 272992 495954 273048
rect 495898 272176 495954 272232
rect 499394 277208 499450 277264
rect 499394 275848 499450 275904
rect 498934 274896 498990 274952
rect 499394 274896 499450 274952
rect 499670 274896 499726 274952
rect 497186 274644 497242 274680
rect 497186 274624 497188 274644
rect 497188 274624 497240 274644
rect 497240 274624 497242 274644
rect 497462 273536 497518 273592
rect 495806 271088 495862 271144
rect 496358 271088 496414 271144
rect 495438 270580 495440 270600
rect 495440 270580 495492 270600
rect 495492 270580 495494 270600
rect 495438 270544 495494 270580
rect 496726 271088 496782 271144
rect 496542 270816 496598 270872
rect 494702 269728 494758 269784
rect 494518 268096 494574 268152
rect 495530 269184 495586 269240
rect 495070 268640 495126 268696
rect 495530 268640 495586 268696
rect 502522 277208 502578 277264
rect 500866 273264 500922 273320
rect 505282 273536 505338 273592
rect 504178 270544 504234 270600
rect 509422 277208 509478 277264
rect 508870 276392 508926 276448
rect 509054 276392 509110 276448
rect 509238 276392 509294 276448
rect 512182 277208 512238 277264
rect 507858 272992 507914 273048
rect 511354 272720 511410 272776
rect 504914 268640 504970 268696
rect 506478 268640 506534 268696
rect 504914 268096 504970 268152
rect 502154 267824 502210 267880
rect 499946 267552 500002 267608
rect 498014 267008 498070 267064
rect 504822 267008 504878 267064
rect 499946 266736 500002 266792
rect 504730 266464 504786 266520
rect 507122 266464 507178 266520
rect 518898 267280 518954 267336
rect 535458 269456 535514 269512
rect 541070 275440 541126 275496
rect 539874 271632 539930 271688
rect 547878 268368 547934 268424
rect 569498 274080 569554 274136
rect 582746 270272 582802 270328
rect 578882 267552 578938 267608
rect 585782 267008 585838 267064
rect 589278 266056 589334 266112
rect 593142 272448 593198 272504
rect 619086 275168 619142 275224
rect 626170 271360 626226 271416
rect 632150 273808 632206 273864
rect 630678 270000 630734 270056
rect 642730 271088 642786 271144
rect 640614 269728 640670 269784
rect 619638 265784 619694 265840
rect 511538 262656 511594 262712
rect 510986 260208 511042 260264
rect 510802 257760 510858 257816
rect 511538 255312 511594 255368
rect 511906 252864 511962 252920
rect 510802 250416 510858 250472
rect 79322 230288 79378 230344
rect 68742 222808 68798 222864
rect 71410 223080 71466 223136
rect 73066 220088 73122 220144
rect 77206 218592 77262 218648
rect 126426 219156 126482 219192
rect 126426 219136 126428 219156
rect 126428 219136 126480 219156
rect 126480 219136 126482 219156
rect 510986 247968 511042 248024
rect 131762 245656 131818 245712
rect 129002 221720 129058 221776
rect 128634 219156 128690 219192
rect 128634 219136 128636 219156
rect 128636 219136 128688 219156
rect 128688 219136 128690 219156
rect 130198 218864 130254 218920
rect 511262 245520 511318 245576
rect 511906 243072 511962 243128
rect 511078 240624 511134 240680
rect 510894 235728 510950 235784
rect 511262 238176 511318 238232
rect 507490 233008 507546 233064
rect 147126 231240 147182 231296
rect 144274 230832 144330 230888
rect 132866 230560 132922 230616
rect 140778 230288 140834 230344
rect 140778 229472 140834 229528
rect 131762 221992 131818 222048
rect 137926 219136 137982 219192
rect 138478 219136 138534 219192
rect 143446 226344 143502 226400
rect 141606 225936 141662 225992
rect 140686 224168 140742 224224
rect 142158 224440 142214 224496
rect 142250 224204 142252 224224
rect 142252 224204 142304 224224
rect 142304 224204 142306 224224
rect 142250 224168 142306 224204
rect 142250 219136 142306 219192
rect 143446 218048 143502 218104
rect 147310 230832 147366 230888
rect 147310 230560 147366 230616
rect 147034 230308 147090 230344
rect 147034 230288 147036 230308
rect 147036 230288 147088 230308
rect 147088 230288 147090 230308
rect 147494 229084 147550 229120
rect 147494 229064 147496 229084
rect 147496 229064 147548 229084
rect 147548 229064 147550 229084
rect 147310 228792 147366 228848
rect 148690 231240 148746 231296
rect 148874 231240 148930 231296
rect 148690 230560 148746 230616
rect 145930 222536 145986 222592
rect 144734 220360 144790 220416
rect 144734 219136 144790 219192
rect 147954 227840 148010 227896
rect 147678 226344 147734 226400
rect 147770 225392 147826 225448
rect 146666 224168 146722 224224
rect 147126 222572 147128 222592
rect 147128 222572 147180 222592
rect 147180 222572 147182 222592
rect 147126 222536 147182 222572
rect 147034 221176 147090 221232
rect 148506 225936 148562 225992
rect 149426 230968 149482 231024
rect 149978 229064 150034 229120
rect 149058 224440 149114 224496
rect 148322 221176 148378 221232
rect 149518 227704 149574 227760
rect 149242 220360 149298 220416
rect 150990 228792 151046 228848
rect 151358 228792 151414 228848
rect 151082 226344 151138 226400
rect 150806 224168 150862 224224
rect 150714 221176 150770 221232
rect 150070 218320 150126 218376
rect 151726 230288 151782 230344
rect 151910 229472 151966 229528
rect 151542 225664 151598 225720
rect 151910 222536 151966 222592
rect 153014 231240 153070 231296
rect 153290 230288 153346 230344
rect 154118 229472 154174 229528
rect 152922 228792 152978 228848
rect 152278 224168 152334 224224
rect 152278 221176 152334 221232
rect 151450 218048 151506 218104
rect 153934 220360 153990 220416
rect 151910 218320 151966 218376
rect 154762 227976 154818 228032
rect 156326 229064 156382 229120
rect 157614 231104 157670 231160
rect 155498 227704 155554 227760
rect 155222 222808 155278 222864
rect 152554 218184 152610 218240
rect 156510 225936 156566 225992
rect 157614 229472 157670 229528
rect 156878 226344 156934 226400
rect 157430 225936 157486 225992
rect 157292 225616 157348 225618
rect 157292 225564 157294 225616
rect 157294 225564 157346 225616
rect 157346 225564 157348 225616
rect 157292 225562 157348 225564
rect 157154 225392 157210 225448
rect 158166 229064 158222 229120
rect 156418 222808 156474 222864
rect 156234 220360 156290 220416
rect 157430 223216 157486 223272
rect 156602 219136 156658 219192
rect 156602 218592 156658 218648
rect 159822 230696 159878 230752
rect 159546 230560 159602 230616
rect 159270 224168 159326 224224
rect 158810 220088 158866 220144
rect 160466 223352 160522 223408
rect 162306 225528 162362 225584
rect 162674 225392 162730 225448
rect 161110 222808 161166 222864
rect 160926 222536 160982 222592
rect 161570 222536 161626 222592
rect 161386 221176 161442 221232
rect 161570 221176 161626 221232
rect 161294 218476 161350 218512
rect 161294 218456 161296 218476
rect 161296 218456 161348 218476
rect 161348 218456 161350 218476
rect 161754 218456 161810 218512
rect 161294 218184 161350 218240
rect 161478 218204 161534 218240
rect 161478 218184 161480 218204
rect 161480 218184 161532 218204
rect 161532 218184 161534 218204
rect 163778 223352 163834 223408
rect 164790 228928 164846 228984
rect 164606 222536 164662 222592
rect 163226 219136 163282 219192
rect 164422 219952 164478 220008
rect 166354 229200 166410 229256
rect 167182 230324 167184 230344
rect 167184 230324 167236 230344
rect 167236 230324 167238 230344
rect 167182 230288 167238 230324
rect 166998 228928 167054 228984
rect 167182 228792 167238 228848
rect 167826 230696 167882 230752
rect 167550 218184 167606 218240
rect 169298 231104 169354 231160
rect 169206 229472 169262 229528
rect 169022 225392 169078 225448
rect 168562 219952 168618 220008
rect 172334 229200 172390 229256
rect 172242 224304 172298 224360
rect 174910 228792 174966 228848
rect 176014 230732 176016 230752
rect 176016 230732 176068 230752
rect 176068 230732 176070 230752
rect 176014 230696 176070 230732
rect 176842 230968 176898 231024
rect 176382 230288 176438 230344
rect 176566 229472 176622 229528
rect 176382 224304 176438 224360
rect 177578 230696 177634 230752
rect 178314 230968 178370 231024
rect 179050 228792 179106 228848
rect 181258 225936 181314 225992
rect 181994 225972 181996 225992
rect 181996 225972 182048 225992
rect 182048 225972 182050 225992
rect 181994 225936 182050 225972
rect 183282 228812 183338 228848
rect 183282 228792 183284 228812
rect 183284 228792 183336 228812
rect 183336 228792 183338 228812
rect 183190 219136 183246 219192
rect 183558 218476 183614 218512
rect 183558 218456 183560 218476
rect 183560 218456 183612 218476
rect 183612 218456 183614 218476
rect 184846 229472 184902 229528
rect 186134 230288 186190 230344
rect 186134 229472 186190 229528
rect 186134 225392 186190 225448
rect 184202 218864 184258 218920
rect 185306 218456 185362 218512
rect 189170 230288 189226 230344
rect 190182 225664 190238 225720
rect 190274 225392 190330 225448
rect 190734 225664 190790 225720
rect 189906 219136 189962 219192
rect 193034 230288 193090 230344
rect 192666 228792 192722 228848
rect 191930 218612 191986 218648
rect 191930 218592 191932 218612
rect 191932 218592 191984 218612
rect 191984 218592 191986 218612
rect 194598 230288 194654 230344
rect 195702 228792 195758 228848
rect 196622 218592 196678 218648
rect 199290 225972 199292 225992
rect 199292 225972 199344 225992
rect 199344 225972 199346 225992
rect 199290 225936 199346 225972
rect 200118 229356 200174 229392
rect 200118 229336 200126 229356
rect 200126 229336 200174 229356
rect 199842 225936 199898 225992
rect 201406 229336 201462 229392
rect 203890 224712 203946 224768
rect 204994 224712 205050 224768
rect 202878 218748 202934 218784
rect 202878 218728 202880 218748
rect 202880 218728 202932 218748
rect 202932 218728 202934 218748
rect 205500 218748 205556 218784
rect 205500 218728 205502 218748
rect 205502 218728 205554 218748
rect 205554 218728 205556 218748
rect 205454 218476 205510 218512
rect 205454 218456 205456 218476
rect 205456 218456 205508 218476
rect 205508 218456 205510 218476
rect 205638 218456 205694 218512
rect 215206 218204 215262 218240
rect 215206 218184 215208 218204
rect 215208 218184 215260 218204
rect 215260 218184 215262 218204
rect 217322 218184 217378 218240
rect 435362 218592 435418 218648
rect 440974 225528 441030 225584
rect 442446 218864 442502 218920
rect 449530 222808 449586 222864
rect 455878 229356 455934 229392
rect 455878 229336 455880 229356
rect 455880 229336 455932 229356
rect 455932 229336 455934 229356
rect 458822 229356 458878 229392
rect 458822 229336 458824 229356
rect 458824 229336 458876 229356
rect 458876 229336 458878 229356
rect 480166 229356 480222 229392
rect 480166 229336 480168 229356
rect 480168 229336 480220 229356
rect 480220 229336 480222 229356
rect 480534 229356 480590 229392
rect 480534 229336 480536 229356
rect 480536 229336 480588 229356
rect 480588 229336 480590 229356
rect 481822 224168 481878 224224
rect 482650 224168 482706 224224
rect 483018 223032 483074 223034
rect 483018 222980 483020 223032
rect 483020 222980 483072 223032
rect 483072 222980 483074 223032
rect 483018 222978 483074 222980
rect 483662 226208 483718 226264
rect 484306 225936 484362 225992
rect 483662 224748 483664 224768
rect 483664 224748 483716 224768
rect 483716 224748 483718 224768
rect 483662 224712 483718 224748
rect 483294 220088 483350 220144
rect 485318 227704 485374 227760
rect 486238 224748 486240 224768
rect 486240 224748 486292 224768
rect 486292 224748 486294 224768
rect 486238 224712 486294 224748
rect 484858 224476 484860 224496
rect 484860 224476 484912 224496
rect 484912 224476 484914 224496
rect 484858 224440 484914 224476
rect 485870 224440 485926 224496
rect 484674 222536 484730 222592
rect 478786 218320 478842 218376
rect 482190 218340 482246 218376
rect 482190 218320 482192 218340
rect 482192 218320 482244 218340
rect 482244 218320 482246 218340
rect 486238 222536 486294 222592
rect 485870 220108 485926 220144
rect 485870 220088 485872 220108
rect 485872 220088 485924 220108
rect 485924 220088 485926 220108
rect 487342 229336 487398 229392
rect 486790 223352 486846 223408
rect 487066 223080 487122 223136
rect 484582 218592 484638 218648
rect 484582 218048 484638 218104
rect 495438 230288 495494 230344
rect 499854 230288 499910 230344
rect 490194 229472 490250 229528
rect 495622 229472 495678 229528
rect 499670 229492 499726 229528
rect 499670 229472 499672 229492
rect 499672 229472 499724 229492
rect 499724 229472 499726 229492
rect 495898 229200 495954 229256
rect 490194 229064 490250 229120
rect 489918 228792 489974 228848
rect 495806 228792 495862 228848
rect 495438 227840 495494 227896
rect 490746 227704 490802 227760
rect 488078 225936 488134 225992
rect 487894 218748 487950 218784
rect 487894 218728 487896 218748
rect 487896 218728 487948 218748
rect 487948 218728 487950 218748
rect 487618 218456 487674 218512
rect 489872 225972 489874 225992
rect 489874 225972 489926 225992
rect 489926 225972 489928 225992
rect 489872 225936 489928 225972
rect 491942 226208 491998 226264
rect 493874 225256 493930 225312
rect 489550 219136 489606 219192
rect 489826 218048 489882 218104
rect 490562 218204 490618 218240
rect 491114 218456 491170 218512
rect 490562 218184 490564 218204
rect 490564 218184 490616 218204
rect 490616 218184 490618 218204
rect 490378 218048 490434 218104
rect 491298 218184 491354 218240
rect 491114 217232 491170 217288
rect 491390 217116 491446 217152
rect 491390 217096 491392 217116
rect 491392 217096 491444 217116
rect 491444 217096 491446 217116
rect 494426 219136 494482 219192
rect 493690 217912 493746 217968
rect 495254 217232 495310 217288
rect 498198 223352 498254 223408
rect 502522 223080 502578 223136
rect 499578 219000 499634 219056
rect 500222 219000 500278 219056
rect 501234 217504 501290 217560
rect 503534 219952 503590 220008
rect 503350 217504 503406 217560
rect 505098 228792 505154 228848
rect 504914 227840 504970 227896
rect 505098 226344 505154 226400
rect 504914 225936 504970 225992
rect 504730 225564 504732 225584
rect 504732 225564 504784 225584
rect 504784 225564 504786 225584
rect 504730 225528 504786 225564
rect 505190 225564 505192 225584
rect 505192 225564 505244 225584
rect 505244 225564 505246 225584
rect 505190 225528 505246 225564
rect 505742 218592 505798 218648
rect 510158 226380 510160 226400
rect 510160 226380 510212 226400
rect 510212 226380 510214 226400
rect 510158 226344 510214 226380
rect 510158 222808 510214 222864
rect 508318 218592 508374 218648
rect 507122 218048 507178 218104
rect 507674 218048 507730 218104
rect 508318 218048 508374 218104
rect 510158 218592 510214 218648
rect 513562 228792 513618 228848
rect 514574 225972 514576 225992
rect 514576 225972 514628 225992
rect 514628 225972 514630 225992
rect 514574 225936 514630 225972
rect 512734 218864 512790 218920
rect 516782 225936 516838 225992
rect 518898 222536 518954 222592
rect 524326 220224 524382 220280
rect 525982 221176 526038 221232
rect 525062 220904 525118 220960
rect 529754 221176 529810 221232
rect 533526 221176 533582 221232
rect 533986 220904 534042 220960
rect 536654 221176 536710 221232
rect 538402 220768 538458 220824
rect 543554 221040 543610 221096
rect 543370 220496 543426 220552
rect 545210 220768 545266 220824
rect 545762 220496 545818 220552
rect 548706 222808 548762 222864
rect 550822 221040 550878 221096
rect 555422 223352 555478 223408
rect 553490 221176 553546 221232
rect 553306 221040 553362 221096
rect 553122 220652 553178 220688
rect 553122 220632 553124 220652
rect 553124 220632 553176 220652
rect 553176 220632 553178 220652
rect 553490 220496 553546 220552
rect 553674 220496 553730 220552
rect 554870 221176 554926 221232
rect 556342 222808 556398 222864
rect 557354 224440 557410 224496
rect 557998 222808 558054 222864
rect 558550 224440 558606 224496
rect 558550 223352 558606 223408
rect 559838 222808 559894 222864
rect 560666 220496 560722 220552
rect 562782 220904 562838 220960
rect 562966 220668 562968 220688
rect 562968 220668 563020 220688
rect 563020 220668 563022 220688
rect 562966 220632 563022 220668
rect 564622 220496 564678 220552
rect 565358 220496 565414 220552
rect 564806 217776 564862 217832
rect 567290 220768 567346 220824
rect 567474 219156 567530 219192
rect 567474 219136 567476 219156
rect 567476 219136 567528 219156
rect 567528 219136 567530 219156
rect 567290 217776 567346 217832
rect 572534 220496 572590 220552
rect 572534 219136 572590 219192
rect 574190 219136 574246 219192
rect 574282 217776 574338 217832
rect 574374 216416 574430 216472
rect 574926 220496 574982 220552
rect 575110 219136 575166 219192
rect 574926 216044 574928 216064
rect 574928 216044 574980 216064
rect 574980 216044 574982 216064
rect 574926 216008 574982 216044
rect 575478 216688 575534 216744
rect 41786 183368 41842 183424
rect 613290 225256 613346 225312
rect 592038 221176 592094 221232
rect 578882 215328 578938 215384
rect 578330 212880 578386 212936
rect 579526 210296 579582 210352
rect 579526 208528 579582 208584
rect 579526 205828 579582 205864
rect 579526 205808 579528 205828
rect 579528 205808 579580 205828
rect 579580 205808 579582 205828
rect 594154 221212 594156 221232
rect 594156 221212 594208 221232
rect 594208 221212 594210 221232
rect 594154 221176 594210 221212
rect 596270 220224 596326 220280
rect 595166 217504 595222 217560
rect 595718 217232 595774 217288
rect 596822 216960 596878 217016
rect 611634 224168 611690 224224
rect 598018 219952 598074 220008
rect 601514 217540 601516 217560
rect 601516 217540 601568 217560
rect 601568 217540 601570 217560
rect 601514 217504 601570 217540
rect 601330 217232 601386 217288
rect 603446 217504 603502 217560
rect 603078 217232 603134 217288
rect 609610 218320 609666 218376
rect 612830 216688 612886 216744
rect 614394 223080 614450 223136
rect 616878 218864 616934 218920
rect 616142 218592 616198 218648
rect 615038 218048 615094 218104
rect 618534 222536 618590 222592
rect 648618 229744 648674 229800
rect 647238 228520 647294 228576
rect 646410 226616 646466 226672
rect 647514 227432 647570 227488
rect 650550 228248 650606 228304
rect 651654 975840 651710 975896
rect 651654 962512 651710 962568
rect 651654 949320 651710 949376
rect 651654 936128 651710 936184
rect 651654 922664 651710 922720
rect 651654 909492 651710 909528
rect 651654 909472 651656 909492
rect 651656 909472 651708 909492
rect 651708 909472 651710 909492
rect 651654 896144 651710 896200
rect 651654 882816 651710 882872
rect 651654 869624 651710 869680
rect 651654 856296 651710 856352
rect 651654 842968 651710 843024
rect 651654 829776 651710 829832
rect 651654 816448 651710 816504
rect 651654 803276 651710 803312
rect 651654 803256 651656 803276
rect 651656 803256 651708 803276
rect 651708 803256 651710 803276
rect 651654 789928 651710 789984
rect 651654 776600 651710 776656
rect 651654 763292 651710 763328
rect 651654 763272 651656 763292
rect 651656 763272 651708 763292
rect 651708 763272 651710 763292
rect 651654 736752 651710 736808
rect 651654 723424 651710 723480
rect 651654 710232 651710 710288
rect 651654 696940 651656 696960
rect 651656 696940 651708 696960
rect 651708 696940 651710 696960
rect 651654 696904 651710 696940
rect 651654 683576 651710 683632
rect 651654 670384 651710 670440
rect 651654 657056 651710 657112
rect 651654 643728 651710 643784
rect 651654 617208 651710 617264
rect 651654 590708 651710 590744
rect 651654 590688 651656 590708
rect 651656 590688 651708 590708
rect 651708 590688 651710 590708
rect 651654 577360 651710 577416
rect 651654 564032 651710 564088
rect 651654 550840 651710 550896
rect 651654 524184 651710 524240
rect 651654 510992 651710 511048
rect 651654 497664 651710 497720
rect 651654 484492 651710 484528
rect 651654 484472 651656 484492
rect 651656 484472 651708 484492
rect 651708 484472 651710 484492
rect 651654 471144 651710 471200
rect 651654 457816 651710 457872
rect 651654 444508 651710 444544
rect 651654 444488 651656 444508
rect 651656 444488 651708 444508
rect 651708 444488 651710 444508
rect 651654 417968 651710 418024
rect 651654 404640 651710 404696
rect 651654 391448 651710 391504
rect 651654 378156 651656 378176
rect 651656 378156 651708 378176
rect 651708 378156 651710 378176
rect 651654 378120 651710 378156
rect 651654 364792 651710 364848
rect 651654 351600 651710 351656
rect 651654 338272 651710 338328
rect 651654 324944 651710 325000
rect 651654 285232 651710 285288
rect 651654 226888 651710 226944
rect 652022 750080 652078 750136
rect 652022 630536 652078 630592
rect 652022 603880 652078 603936
rect 652022 537512 652078 537568
rect 652022 431296 652078 431352
rect 652022 311752 652078 311808
rect 652206 298424 652262 298480
rect 653034 276936 653090 276992
rect 656898 276664 656954 276720
rect 654322 230016 654378 230072
rect 656346 227160 656402 227216
rect 658462 265512 658518 265568
rect 661498 221992 661554 222048
rect 662418 223896 662474 223952
rect 662602 221720 662658 221776
rect 663798 221448 663854 221504
rect 663982 219680 664038 219736
rect 665822 211112 665878 211168
rect 664442 210840 664498 210896
rect 578330 203224 578386 203280
rect 579158 200640 579214 200696
rect 589462 208276 589518 208312
rect 589462 208256 589464 208276
rect 589464 208256 589516 208276
rect 589516 208256 589518 208276
rect 589554 206932 589556 206952
rect 589556 206932 589608 206952
rect 589608 206932 589610 206952
rect 589554 206896 589610 206932
rect 589462 205128 589518 205184
rect 589462 203632 589518 203688
rect 589462 202136 589518 202192
rect 589462 199824 589518 199880
rect 590566 198600 590622 198656
rect 578882 198056 578938 198112
rect 589462 196968 589518 197024
rect 579526 196036 579582 196072
rect 579526 196016 579528 196036
rect 579528 196016 579580 196036
rect 579580 196016 579582 196036
rect 589554 195472 589610 195528
rect 579526 193860 579582 193896
rect 579526 193840 579528 193860
rect 579528 193840 579580 193860
rect 579580 193840 579582 193860
rect 589554 193568 589610 193624
rect 589462 191664 589518 191720
rect 579526 191140 579582 191176
rect 579526 191120 579528 191140
rect 579528 191120 579580 191140
rect 579580 191120 579582 191140
rect 589462 190032 589518 190088
rect 579526 188980 579528 189000
rect 579528 188980 579580 189000
rect 579580 188980 579582 189000
rect 579526 188944 579582 188980
rect 589646 188400 589702 188456
rect 589462 186768 589518 186824
rect 579526 186632 579582 186688
rect 589462 185136 589518 185192
rect 578514 184320 578570 184376
rect 589462 183504 589518 183560
rect 579434 182008 579490 182064
rect 589462 181872 589518 181928
rect 578330 179152 578386 179208
rect 579526 176432 579582 176488
rect 578698 174664 578754 174720
rect 579526 172080 579582 172136
rect 589462 180240 589518 180296
rect 589462 178608 589518 178664
rect 589462 176976 589518 177032
rect 589278 175364 589334 175400
rect 589278 175344 589280 175364
rect 589280 175344 589332 175364
rect 589332 175344 589334 175364
rect 579250 169532 579252 169552
rect 579252 169532 579304 169552
rect 579304 169532 579306 169552
rect 579250 169496 579306 169532
rect 578882 166912 578938 166968
rect 589738 173712 589794 173768
rect 589462 172080 589518 172136
rect 588542 170448 588598 170504
rect 579526 164464 579582 164520
rect 579526 162424 579582 162480
rect 579526 159704 579582 159760
rect 579250 157120 579306 157176
rect 578698 155080 578754 155136
rect 578330 152632 578386 152688
rect 579526 150048 579582 150104
rect 578422 147600 578478 147656
rect 578790 144608 578846 144664
rect 578330 137672 578386 137728
rect 578330 133048 578386 133104
rect 579250 142840 579306 142896
rect 579526 140256 579582 140312
rect 579342 135124 579344 135144
rect 579344 135124 579396 135144
rect 579396 135124 579398 135144
rect 579342 135088 579398 135124
rect 579066 130600 579122 130656
rect 578882 125296 578938 125352
rect 578882 122612 578884 122632
rect 578884 122612 578936 122632
rect 578936 122612 578938 122632
rect 578882 122576 578938 122612
rect 578422 120808 578478 120864
rect 578514 118260 578516 118280
rect 578516 118260 578568 118280
rect 578568 118260 578570 118280
rect 578514 118224 578570 118260
rect 578330 105848 578386 105904
rect 578606 96192 578662 96248
rect 578514 88984 578570 89040
rect 78586 50224 78642 50280
rect 131026 49680 131082 49736
rect 151910 47232 151966 47288
rect 151910 45872 151966 45928
rect 187514 42064 187570 42120
rect 306976 42336 307032 42392
rect 310104 42336 310160 42392
rect 361946 42064 362002 42120
rect 365166 42064 365222 42120
rect 579526 127880 579582 127936
rect 579250 115640 579306 115696
rect 579526 113092 579528 113112
rect 579528 113092 579580 113112
rect 579580 113092 579582 113112
rect 579526 113056 579582 113092
rect 579526 111016 579582 111072
rect 579250 108432 579306 108488
rect 579526 103420 579582 103456
rect 579526 103400 579528 103420
rect 579528 103400 579580 103420
rect 579580 103400 579582 103420
rect 579250 100544 579306 100600
rect 579526 98776 579582 98832
rect 579526 93608 579582 93664
rect 579526 91044 579582 91080
rect 579526 91024 579528 91044
rect 579528 91024 579580 91044
rect 579580 91024 579582 91044
rect 579526 86400 579582 86456
rect 579342 83816 579398 83872
rect 579526 81388 579582 81424
rect 579526 81368 579528 81388
rect 579528 81368 579580 81388
rect 579580 81368 579582 81388
rect 579066 79192 579122 79248
rect 578882 76744 578938 76800
rect 578514 68720 578570 68776
rect 579526 74160 579582 74216
rect 579526 71476 579528 71496
rect 579528 71476 579580 71496
rect 579580 71476 579582 71496
rect 579526 71440 579582 71476
rect 579526 66952 579582 67008
rect 579250 64504 579306 64560
rect 578514 61784 578570 61840
rect 579526 58964 579528 58984
rect 579528 58964 579580 58984
rect 579580 58964 579582 58984
rect 579526 58928 579582 58964
rect 589462 168816 589518 168872
rect 589462 167184 589518 167240
rect 589462 165552 589518 165608
rect 589738 163920 589794 163976
rect 590106 162288 590162 162344
rect 589462 160656 589518 160712
rect 588726 159024 588782 159080
rect 579066 57160 579122 57216
rect 578514 54712 578570 54768
rect 588542 144336 588598 144392
rect 589462 157412 589518 157448
rect 589462 157392 589464 157412
rect 589464 157392 589516 157412
rect 589516 157392 589518 157412
rect 589370 155760 589426 155816
rect 589462 154128 589518 154184
rect 589738 152496 589794 152552
rect 589922 150864 589978 150920
rect 589278 149232 589334 149288
rect 589462 147600 589518 147656
rect 589462 145968 589518 146024
rect 589462 141072 589518 141128
rect 589462 139440 589518 139496
rect 590290 142704 590346 142760
rect 589922 137808 589978 137864
rect 589462 136176 589518 136232
rect 589462 134544 589518 134600
rect 589462 132912 589518 132968
rect 588910 131280 588966 131336
rect 588726 124752 588782 124808
rect 589462 129648 589518 129704
rect 589278 126384 589334 126440
rect 589462 121508 589518 121544
rect 589462 121488 589464 121508
rect 589464 121488 589516 121508
rect 589516 121488 589518 121508
rect 590106 128016 590162 128072
rect 589462 119856 589518 119912
rect 589462 118224 589518 118280
rect 589462 116592 589518 116648
rect 589922 114960 589978 115016
rect 589462 113328 589518 113384
rect 589646 111696 589702 111752
rect 589462 110064 589518 110120
rect 589462 108432 589518 108488
rect 589462 106800 589518 106856
rect 589462 105168 589518 105224
rect 589462 103556 589518 103592
rect 589462 103536 589464 103556
rect 589464 103536 589516 103556
rect 589516 103536 589518 103556
rect 589370 101904 589426 101960
rect 590290 123120 590346 123176
rect 666742 245928 666798 245984
rect 666926 245656 666982 245712
rect 666742 222264 666798 222320
rect 666558 184728 666614 184784
rect 666926 192616 666982 192672
rect 667386 246064 667442 246120
rect 668122 245928 668178 245984
rect 675390 966456 675446 966512
rect 672906 959112 672962 959168
rect 668582 728728 668638 728784
rect 669410 774968 669466 775024
rect 668766 688608 668822 688664
rect 669042 685072 669098 685128
rect 669594 735120 669650 735176
rect 669410 710640 669466 710696
rect 669042 617208 669098 617264
rect 668306 245656 668362 245712
rect 668398 219408 668454 219464
rect 666926 159976 666982 160032
rect 668122 187720 668178 187776
rect 667938 177948 667994 177984
rect 667938 177928 667940 177948
rect 667940 177928 667992 177948
rect 667992 177928 667994 177948
rect 667938 174700 667940 174720
rect 667940 174700 667992 174720
rect 667992 174700 667994 174720
rect 667938 174664 667994 174700
rect 667938 169668 667940 169688
rect 667940 169668 667992 169688
rect 667992 169668 667994 169688
rect 667938 169632 667994 169668
rect 668030 164908 668032 164928
rect 668032 164908 668084 164928
rect 668084 164908 668086 164928
rect 668030 164872 668086 164908
rect 667938 130600 667994 130656
rect 667938 125704 667994 125760
rect 669042 593544 669098 593600
rect 669594 642096 669650 642152
rect 668582 168136 668638 168192
rect 668582 165688 668638 165744
rect 668582 163240 668638 163296
rect 669226 342080 669282 342136
rect 669134 241984 669190 242040
rect 669134 224984 669190 225040
rect 668950 223624 669006 223680
rect 668766 158344 668822 158400
rect 668766 150220 668768 150240
rect 668768 150220 668820 150240
rect 668820 150220 668822 150240
rect 668766 150184 668822 150220
rect 668766 145288 668822 145344
rect 668582 143656 668638 143712
rect 668674 140428 668676 140448
rect 668676 140428 668728 140448
rect 668728 140428 668730 140448
rect 668674 140392 668730 140428
rect 668766 138624 668822 138680
rect 668766 135496 668822 135552
rect 668214 120808 668270 120864
rect 667938 117544 667994 117600
rect 668398 115812 668400 115832
rect 668400 115812 668452 115832
rect 668452 115812 668454 115832
rect 668398 115776 668454 115812
rect 668398 114316 668400 114336
rect 668400 114316 668452 114336
rect 668452 114316 668454 114336
rect 668398 114280 668454 114316
rect 668030 112648 668086 112704
rect 666742 109316 666798 109372
rect 669226 182860 669228 182880
rect 669228 182860 669280 182880
rect 669280 182860 669282 182880
rect 669226 182824 669282 182860
rect 669134 176568 669190 176624
rect 669226 129004 669228 129024
rect 669228 129004 669280 129024
rect 669280 129004 669282 129024
rect 669226 128968 669282 129004
rect 670422 734440 670478 734496
rect 669226 124108 669228 124128
rect 669228 124108 669280 124128
rect 669280 124108 669282 124128
rect 669226 124072 669282 124108
rect 669134 119212 669136 119232
rect 669136 119212 669188 119232
rect 669188 119212 669190 119232
rect 669134 119176 669190 119212
rect 671250 734168 671306 734224
rect 672354 867992 672410 868048
rect 670790 647400 670846 647456
rect 675758 965096 675814 965152
rect 675206 963328 675262 963384
rect 674470 952176 674526 952232
rect 674470 933408 674526 933464
rect 675758 961968 675814 962024
rect 674930 959384 674986 959440
rect 675114 959112 675170 959168
rect 675758 958296 675814 958352
rect 675758 956392 675814 956448
rect 674930 948912 674986 948968
rect 675666 953944 675722 954000
rect 675390 952176 675446 952232
rect 677506 951496 677562 951552
rect 675942 949184 675998 949240
rect 674930 941840 674986 941896
rect 674930 938304 674986 938360
rect 675850 941840 675906 941896
rect 675482 939936 675538 939992
rect 675666 939528 675722 939584
rect 675298 939120 675354 939176
rect 675482 938712 675538 938768
rect 675298 937896 675354 937952
rect 675482 937524 675484 937544
rect 675484 937524 675536 937544
rect 675536 937524 675538 937544
rect 675482 937488 675538 937524
rect 675482 937080 675538 937136
rect 675666 936672 675722 936728
rect 675482 936264 675538 936320
rect 675298 935856 675354 935912
rect 675850 934632 675906 934688
rect 675114 934088 675170 934144
rect 675298 933816 675354 933872
rect 675482 933036 675484 933056
rect 675484 933036 675536 933056
rect 675536 933036 675538 933056
rect 675482 933000 675538 933036
rect 674654 932592 674710 932648
rect 674286 932184 674342 932240
rect 675482 931404 675484 931424
rect 675484 931404 675536 931424
rect 675536 931404 675538 931424
rect 675482 931368 675538 931404
rect 683302 950000 683358 950056
rect 677506 931096 677562 931152
rect 675482 930164 675538 930200
rect 675482 930144 675484 930164
rect 675484 930144 675536 930164
rect 675536 930144 675538 930164
rect 683302 935584 683358 935640
rect 682382 935176 682438 935232
rect 675482 929736 675538 929792
rect 683118 929464 683174 929520
rect 672998 864184 673054 864240
rect 675482 928512 675538 928568
rect 675758 877104 675814 877160
rect 675298 876424 675354 876480
rect 675390 873976 675446 874032
rect 673274 773608 673330 773664
rect 672998 752256 673054 752312
rect 675758 872752 675814 872808
rect 675390 872208 675446 872264
rect 674470 854256 674526 854312
rect 672814 730088 672870 730144
rect 671802 667800 671858 667856
rect 670606 217912 670662 217968
rect 671894 616800 671950 616856
rect 671526 608640 671582 608696
rect 670974 344936 671030 344992
rect 670974 278704 671030 278760
rect 670974 216552 671030 216608
rect 670790 211112 670846 211168
rect 670790 210840 670846 210896
rect 670790 201456 670846 201512
rect 670606 193296 670662 193352
rect 668766 111016 668822 111072
rect 671802 345208 671858 345264
rect 671894 245656 671950 245712
rect 671894 216144 671950 216200
rect 672906 663448 672962 663504
rect 672814 553968 672870 554024
rect 672538 377984 672594 378040
rect 673458 734848 673514 734904
rect 673826 732672 673882 732728
rect 673642 725872 673698 725928
rect 673642 683032 673698 683088
rect 673458 682760 673514 682816
rect 674838 869624 674894 869680
rect 675666 869624 675722 869680
rect 675482 867992 675538 868048
rect 674838 863776 674894 863832
rect 675482 864184 675538 864240
rect 675482 863776 675538 863832
rect 675390 784216 675446 784272
rect 674930 780272 674986 780328
rect 675482 779864 675538 779920
rect 674746 775376 674802 775432
rect 674562 772656 674618 772712
rect 675390 774968 675446 775024
rect 675390 773608 675446 773664
rect 675390 773336 675446 773392
rect 675114 771704 675170 771760
rect 675850 772656 675906 772712
rect 679622 772656 679678 772712
rect 675850 771704 675906 771760
rect 675482 761540 675484 761560
rect 675484 761540 675536 761560
rect 675536 761540 675538 761560
rect 675482 761504 675538 761540
rect 675298 761096 675354 761152
rect 675482 760688 675538 760744
rect 675482 760300 675538 760336
rect 675482 760280 675484 760300
rect 675484 760280 675536 760300
rect 675536 760280 675538 760300
rect 675482 759892 675538 759928
rect 675482 759872 675484 759892
rect 675484 759872 675536 759892
rect 675536 759872 675538 759892
rect 675482 759500 675484 759520
rect 675484 759500 675536 759520
rect 675536 759500 675538 759520
rect 675482 759464 675538 759500
rect 675482 759076 675538 759112
rect 675482 759056 675484 759076
rect 675484 759056 675536 759076
rect 675536 759056 675538 759076
rect 675482 758684 675484 758704
rect 675484 758684 675536 758704
rect 675536 758684 675538 758704
rect 675482 758648 675538 758684
rect 675482 758260 675538 758296
rect 675482 758240 675484 758260
rect 675484 758240 675536 758260
rect 675536 758240 675538 758260
rect 675298 757832 675354 757888
rect 675482 757444 675538 757480
rect 675482 757424 675484 757444
rect 675484 757424 675536 757444
rect 675536 757424 675538 757444
rect 676954 761776 677010 761832
rect 676954 757016 677010 757072
rect 683394 772384 683450 772440
rect 682382 771296 682438 771352
rect 681002 756608 681058 756664
rect 679622 756200 679678 756256
rect 675850 755792 675906 755848
rect 682382 755384 682438 755440
rect 675482 755012 675484 755032
rect 675484 755012 675536 755032
rect 675536 755012 675538 755032
rect 675482 754976 675538 755012
rect 675482 754604 675484 754624
rect 675484 754604 675536 754624
rect 675536 754604 675538 754624
rect 675482 754568 675538 754604
rect 675482 753380 675484 753400
rect 675484 753380 675536 753400
rect 675536 753380 675538 753400
rect 675482 753344 675538 753380
rect 675482 752972 675484 752992
rect 675484 752972 675536 752992
rect 675536 752972 675538 752992
rect 675482 752936 675538 752972
rect 675850 752256 675906 752312
rect 675482 751748 675484 751768
rect 675484 751748 675536 751768
rect 675536 751748 675538 751768
rect 675482 751712 675538 751748
rect 675482 751324 675538 751360
rect 675482 751304 675484 751324
rect 675484 751304 675536 751324
rect 675536 751304 675538 751324
rect 684038 771976 684094 772032
rect 684038 754160 684094 754216
rect 683394 752528 683450 752584
rect 683210 752120 683266 752176
rect 674930 751032 674986 751088
rect 683118 750692 683174 750748
rect 675482 750100 675538 750136
rect 675482 750080 675484 750100
rect 675484 750080 675536 750100
rect 675536 750080 675538 750100
rect 675574 743008 675630 743064
rect 675390 738656 675446 738712
rect 675114 738112 675170 738168
rect 675482 734848 675538 734904
rect 675482 734440 675538 734496
rect 675482 734168 675538 734224
rect 675298 733624 675354 733680
rect 675390 732672 675446 732728
rect 675390 730088 675446 730144
rect 674562 728048 674618 728104
rect 674286 723152 674342 723208
rect 674838 715300 674840 715320
rect 674840 715300 674892 715320
rect 674892 715300 674894 715320
rect 674838 715264 674894 715300
rect 674470 707104 674526 707160
rect 675390 728728 675446 728784
rect 676034 728048 676090 728104
rect 675850 723152 675906 723208
rect 675206 721520 675262 721576
rect 675482 716488 675538 716544
rect 675298 716080 675354 716136
rect 675482 715672 675538 715728
rect 675482 714876 675538 714912
rect 675482 714856 675484 714876
rect 675484 714856 675536 714876
rect 675536 714856 675538 714876
rect 675482 714484 675484 714504
rect 675484 714484 675536 714504
rect 675536 714484 675538 714504
rect 675482 714448 675538 714484
rect 675482 714060 675538 714096
rect 675482 714040 675484 714060
rect 675484 714040 675536 714060
rect 675536 714040 675538 714060
rect 675482 713668 675484 713688
rect 675484 713668 675536 713688
rect 675536 713668 675538 713688
rect 675482 713632 675538 713668
rect 677690 713448 677746 713488
rect 677690 713432 677692 713448
rect 677692 713432 677744 713448
rect 677744 713432 677746 713448
rect 675482 713244 675538 713280
rect 675482 713224 675484 713244
rect 675484 713224 675536 713244
rect 675536 713224 675538 713244
rect 675482 712852 675484 712872
rect 675484 712852 675536 712872
rect 675536 712852 675538 712872
rect 675482 712816 675538 712852
rect 675482 712428 675538 712464
rect 675482 712408 675484 712428
rect 675484 712408 675536 712428
rect 675536 712408 675538 712428
rect 675482 712036 675484 712056
rect 675484 712036 675536 712056
rect 675536 712036 675538 712056
rect 675482 712000 675538 712036
rect 676034 711592 676090 711648
rect 675482 711220 675484 711240
rect 675484 711220 675536 711240
rect 675536 711220 675538 711240
rect 675482 711184 675538 711220
rect 683118 710776 683174 710832
rect 675850 710640 675906 710696
rect 675482 710368 675538 710424
rect 675298 709996 675300 710016
rect 675300 709996 675352 710016
rect 675352 709996 675354 710016
rect 675298 709960 675354 709996
rect 675482 709588 675484 709608
rect 675484 709588 675536 709608
rect 675536 709588 675538 709608
rect 675482 709552 675538 709588
rect 675482 708772 675484 708792
rect 675484 708772 675536 708792
rect 675536 708772 675538 708792
rect 675482 708736 675538 708772
rect 675482 708364 675484 708384
rect 675484 708364 675536 708384
rect 675536 708364 675538 708384
rect 675482 708328 675538 708364
rect 675482 707548 675484 707568
rect 675484 707548 675536 707568
rect 675536 707548 675538 707568
rect 675482 707512 675538 707548
rect 675482 706308 675538 706344
rect 675482 706288 675484 706308
rect 675484 706288 675536 706308
rect 675536 706288 675538 706308
rect 683486 707920 683542 707976
rect 683302 706696 683358 706752
rect 683118 705472 683174 705528
rect 675482 705084 675538 705120
rect 675482 705064 675484 705084
rect 675484 705064 675536 705084
rect 675536 705064 675538 705084
rect 674010 668888 674066 668944
rect 674010 644680 674066 644736
rect 673734 644272 673790 644328
rect 673550 599800 673606 599856
rect 673918 643456 673974 643512
rect 675390 696768 675446 696824
rect 675114 694592 675170 694648
rect 674930 694048 674986 694104
rect 675114 692960 675170 693016
rect 674470 618568 674526 618624
rect 674286 617752 674342 617808
rect 675114 688608 675170 688664
rect 674838 684256 674894 684312
rect 674838 669704 674894 669760
rect 674838 664028 674840 664048
rect 674840 664028 674892 664048
rect 674892 664028 674894 664048
rect 674838 663992 674894 664028
rect 675298 685616 675354 685672
rect 675482 685072 675538 685128
rect 675482 684256 675538 684312
rect 675850 683032 675906 683088
rect 676034 682760 676090 682816
rect 681002 681808 681058 681864
rect 675482 671336 675538 671392
rect 675482 670928 675538 670984
rect 675482 670520 675538 670576
rect 675482 670112 675538 670168
rect 675482 669296 675538 669352
rect 675482 668516 675484 668536
rect 675484 668516 675536 668536
rect 675536 668516 675538 668536
rect 675482 668480 675538 668516
rect 675482 667700 675484 667720
rect 675484 667700 675536 667720
rect 675536 667700 675538 667720
rect 675482 667664 675538 667700
rect 675482 667276 675538 667312
rect 675482 667256 675484 667276
rect 675484 667256 675536 667276
rect 675536 667256 675538 667276
rect 681002 666984 681058 667040
rect 675482 666068 675484 666088
rect 675484 666068 675536 666088
rect 675536 666068 675538 666088
rect 675482 666032 675538 666068
rect 675482 665624 675538 665680
rect 675666 664808 675722 664864
rect 675482 664400 675538 664456
rect 675850 663448 675906 663504
rect 675482 663212 675484 663232
rect 675484 663212 675536 663232
rect 675536 663212 675538 663232
rect 675482 663176 675538 663212
rect 675482 662804 675484 662824
rect 675484 662804 675536 662824
rect 675536 662804 675538 662824
rect 675482 662768 675538 662804
rect 675482 661580 675484 661600
rect 675484 661580 675536 661600
rect 675536 661580 675538 661600
rect 675482 661544 675538 661580
rect 675482 661156 675538 661192
rect 675482 661136 675484 661156
rect 675484 661136 675536 661156
rect 675536 661136 675538 661156
rect 675482 659932 675538 659968
rect 675482 659912 675484 659932
rect 675484 659912 675536 659932
rect 675536 659912 675538 659932
rect 683210 662496 683266 662552
rect 684038 674056 684094 674112
rect 684038 663720 684094 663776
rect 683394 662088 683450 662144
rect 683118 660048 683174 660104
rect 675574 652840 675630 652896
rect 675206 650120 675262 650176
rect 674930 643864 674986 643920
rect 675390 648896 675446 648952
rect 675390 647944 675446 648000
rect 675666 647400 675722 647456
rect 675390 644680 675446 644736
rect 675390 644272 675446 644328
rect 675390 643456 675446 643512
rect 675390 642096 675446 642152
rect 675666 640328 675722 640384
rect 675482 638152 675538 638208
rect 675298 637880 675354 637936
rect 675206 637608 675262 637664
rect 675850 637880 675906 637936
rect 675482 636520 675538 636576
rect 675206 631352 675262 631408
rect 675390 631352 675446 631408
rect 675298 626320 675354 626376
rect 675114 625912 675170 625968
rect 675482 625504 675538 625560
rect 675298 625096 675354 625152
rect 675114 624688 675170 624744
rect 675482 624300 675538 624336
rect 675482 624280 675484 624300
rect 675484 624280 675536 624300
rect 675536 624280 675538 624300
rect 675482 623908 675484 623928
rect 675484 623908 675536 623928
rect 675536 623908 675538 623928
rect 675482 623872 675538 623908
rect 675298 623600 675354 623656
rect 676402 623600 676458 623656
rect 675482 623464 675538 623520
rect 675298 623056 675354 623112
rect 675482 622648 675538 622704
rect 675298 622240 675354 622296
rect 683394 636792 683450 636848
rect 683210 636520 683266 636576
rect 679622 621968 679678 622024
rect 682382 621560 682438 621616
rect 675482 621016 675538 621072
rect 683394 623600 683450 623656
rect 683210 620744 683266 620800
rect 675482 620200 675538 620256
rect 675298 619828 675300 619848
rect 675300 619828 675352 619848
rect 675352 619828 675354 619848
rect 675298 619792 675354 619828
rect 675482 619420 675484 619440
rect 675484 619420 675536 619440
rect 675536 619420 675538 619440
rect 675482 619384 675538 619420
rect 675482 618196 675484 618216
rect 675484 618196 675536 618216
rect 675536 618196 675538 618216
rect 675482 618160 675538 618196
rect 683578 619112 683634 619168
rect 683394 617480 683450 617536
rect 675850 617208 675906 617264
rect 674654 616936 674710 616992
rect 675482 616528 675538 616584
rect 675298 616140 675354 616176
rect 675298 616120 675300 616140
rect 675300 616120 675352 616140
rect 675352 616120 675354 616140
rect 683118 615440 683174 615496
rect 675482 614896 675538 614952
rect 674102 592864 674158 592920
rect 673642 574504 673698 574560
rect 673550 547032 673606 547088
rect 675114 604424 675170 604480
rect 675114 602928 675170 602984
rect 675482 599800 675538 599856
rect 674838 586200 674894 586256
rect 674746 579808 674802 579864
rect 674930 571512 674986 571568
rect 675390 593544 675446 593600
rect 675850 592864 675906 592920
rect 678242 592864 678298 592920
rect 676034 592592 676090 592648
rect 675482 581052 675538 581088
rect 675482 581032 675484 581052
rect 675484 581032 675536 581052
rect 675536 581032 675538 581052
rect 675298 580624 675354 580680
rect 675482 580216 675538 580272
rect 675482 579420 675538 579456
rect 675482 579400 675484 579420
rect 675484 579400 675536 579420
rect 675536 579400 675538 579420
rect 675482 579028 675484 579048
rect 675484 579028 675536 579048
rect 675536 579028 675538 579048
rect 675482 578992 675538 579028
rect 675482 578604 675538 578640
rect 675482 578584 675484 578604
rect 675484 578584 675536 578604
rect 675536 578584 675538 578604
rect 675298 578176 675354 578232
rect 675298 577788 675354 577824
rect 675298 577768 675300 577788
rect 675300 577768 675352 577788
rect 675352 577768 675354 577788
rect 675298 577396 675300 577416
rect 675300 577396 675352 577416
rect 675352 577396 675354 577416
rect 675298 577360 675354 577396
rect 675298 576972 675354 577008
rect 675298 576952 675300 576972
rect 675300 576952 675352 576972
rect 675352 576952 675354 576972
rect 675482 576544 675538 576600
rect 676034 575728 676090 575784
rect 678242 575592 678298 575648
rect 675298 574912 675354 574968
rect 675482 574096 675538 574152
rect 675482 573724 675484 573744
rect 675484 573724 675536 573744
rect 675536 573724 675538 573744
rect 675482 573688 675538 573724
rect 675482 572908 675484 572928
rect 675484 572908 675536 572928
rect 675536 572908 675538 572928
rect 675482 572872 675538 572908
rect 675482 572500 675484 572520
rect 675484 572500 675536 572520
rect 675536 572500 675538 572520
rect 675482 572464 675538 572500
rect 675482 572056 675538 572112
rect 683210 571920 683266 571976
rect 683394 571104 683450 571160
rect 675482 570852 675538 570888
rect 675482 570832 675484 570852
rect 675484 570832 675536 570852
rect 675536 570832 675538 570852
rect 683118 570288 683174 570344
rect 675482 569628 675538 569664
rect 675482 569608 675484 569628
rect 675484 569608 675536 569628
rect 675536 569608 675538 569628
rect 674102 483112 674158 483168
rect 675390 561856 675446 561912
rect 675482 559408 675538 559464
rect 675758 559000 675814 559056
rect 675482 553968 675538 554024
rect 675390 550296 675446 550352
rect 675022 549752 675078 549808
rect 675482 549208 675538 549264
rect 674746 547304 674802 547360
rect 674562 546760 674618 546816
rect 674562 535064 674618 535120
rect 674746 534112 674802 534168
rect 674562 533568 674618 533624
rect 674746 531936 674802 531992
rect 674746 492088 674802 492144
rect 674562 490048 674618 490104
rect 674746 485152 674802 485208
rect 674378 482704 674434 482760
rect 673274 394576 673330 394632
rect 673274 340448 673330 340504
rect 673366 286456 673422 286512
rect 673090 285504 673146 285560
rect 672538 278704 672594 278760
rect 671986 215464 672042 215520
rect 672538 212608 672594 212664
rect 672354 210432 672410 210488
rect 672354 209208 672410 209264
rect 672354 183504 672410 183560
rect 672170 168272 672226 168328
rect 672906 241712 672962 241768
rect 675482 547848 675538 547904
rect 675206 545808 675262 545864
rect 675758 547576 675814 547632
rect 675114 508816 675170 508872
rect 675114 491680 675170 491736
rect 675482 536016 675538 536072
rect 675482 535492 675538 535528
rect 675482 535472 675484 535492
rect 675484 535472 675536 535492
rect 675536 535472 675538 535492
rect 675482 534792 675538 534848
rect 675482 534384 675538 534440
rect 675482 533160 675538 533216
rect 675482 532344 675538 532400
rect 675482 531564 675484 531584
rect 675484 531564 675536 531584
rect 675536 531564 675538 531584
rect 675482 531528 675538 531564
rect 675482 530712 675538 530768
rect 675482 529932 675484 529952
rect 675484 529932 675536 529952
rect 675536 529932 675538 529952
rect 675482 529896 675538 529932
rect 675482 529372 675538 529408
rect 675482 529352 675484 529372
rect 675484 529352 675536 529372
rect 675536 529352 675538 529372
rect 675482 529080 675538 529136
rect 675482 528300 675484 528320
rect 675484 528300 675536 528320
rect 675536 528300 675538 528320
rect 675482 528264 675538 528300
rect 675482 527620 675484 527640
rect 675484 527620 675536 527640
rect 675536 527620 675538 527640
rect 675482 527584 675538 527620
rect 675482 526088 675538 526144
rect 675482 524592 675538 524648
rect 675482 491272 675538 491328
rect 675482 490864 675538 490920
rect 675482 488416 675538 488472
rect 675942 547324 675998 547360
rect 675942 547304 675944 547324
rect 675944 547304 675996 547324
rect 675996 547304 675998 547324
rect 675942 547032 675998 547088
rect 676126 546760 676182 546816
rect 675942 532820 675998 532876
rect 682382 545128 682438 545184
rect 682382 530576 682438 530632
rect 683394 528128 683450 528184
rect 683210 526904 683266 526960
rect 683118 525716 683120 525736
rect 683120 525716 683172 525736
rect 683172 525716 683174 525736
rect 683118 525680 683174 525716
rect 676126 508816 676182 508872
rect 677414 490456 677470 490512
rect 677230 489640 677286 489696
rect 675942 489232 675998 489288
rect 676034 488824 676090 488880
rect 675942 488008 675998 488064
rect 675758 487600 675814 487656
rect 675298 486784 675354 486840
rect 675482 486376 675538 486432
rect 675482 485988 675538 486024
rect 675482 485968 675484 485988
rect 675484 485968 675536 485988
rect 675536 485968 675538 485988
rect 675482 485560 675538 485616
rect 675482 484336 675538 484392
rect 675298 483964 675300 483984
rect 675300 483964 675352 483984
rect 675352 483964 675354 483984
rect 675298 483928 675354 483964
rect 675298 483556 675300 483576
rect 675300 483556 675352 483576
rect 675352 483556 675354 483576
rect 675298 483520 675354 483556
rect 675482 482332 675484 482352
rect 675484 482332 675536 482352
rect 675536 482332 675538 482352
rect 675482 482296 675538 482332
rect 675482 481908 675538 481944
rect 675482 481888 675484 481908
rect 675484 481888 675536 481908
rect 675536 481888 675538 481908
rect 674930 481480 674986 481536
rect 675482 480684 675538 480720
rect 675482 480664 675484 480684
rect 675484 480664 675536 480684
rect 675536 480664 675538 480684
rect 675298 403824 675354 403880
rect 675482 403416 675538 403472
rect 675482 403028 675538 403064
rect 675482 403008 675484 403028
rect 675484 403008 675536 403028
rect 675536 403008 675538 403028
rect 674654 402192 674710 402248
rect 674286 396072 674342 396128
rect 674102 393624 674158 393680
rect 673918 249736 673974 249792
rect 673918 213968 673974 214024
rect 673734 210432 673790 210488
rect 673550 190032 673606 190088
rect 673182 183504 673238 183560
rect 674470 395664 674526 395720
rect 675482 401396 675538 401432
rect 675482 401376 675484 401396
rect 675484 401376 675536 401396
rect 675536 401376 675538 401396
rect 675482 400580 675538 400616
rect 675482 400560 675484 400580
rect 675484 400560 675536 400580
rect 675536 400560 675538 400580
rect 683302 500928 683358 500984
rect 679622 487192 679678 487248
rect 683302 484744 683358 484800
rect 677414 402872 677470 402928
rect 677230 402056 677286 402112
rect 676034 400968 676090 401024
rect 675850 400152 675906 400208
rect 675482 399764 675538 399800
rect 675482 399744 675484 399764
rect 675484 399744 675536 399764
rect 675536 399744 675538 399764
rect 675666 399336 675722 399392
rect 675114 398112 675170 398168
rect 675298 397296 675354 397352
rect 675482 396480 675538 396536
rect 676218 398384 676274 398440
rect 681002 397568 681058 397624
rect 675482 394440 675538 394496
rect 675482 394032 675538 394088
rect 675482 392400 675538 392456
rect 683026 392672 683082 392728
rect 683026 389816 683082 389872
rect 681002 388456 681058 388512
rect 675758 384920 675814 384976
rect 675758 380568 675814 380624
rect 675758 378664 675814 378720
rect 675758 377304 675814 377360
rect 675298 374992 675354 375048
rect 675666 372952 675722 373008
rect 675114 372544 675170 372600
rect 675298 358672 675354 358728
rect 675114 358264 675170 358320
rect 674654 357448 674710 357504
rect 675482 357856 675538 357912
rect 675482 357060 675538 357096
rect 675482 357040 675484 357060
rect 675484 357040 675536 357060
rect 675536 357040 675538 357060
rect 674746 356632 674802 356688
rect 674654 356224 674710 356280
rect 674470 349696 674526 349752
rect 674286 348472 674342 348528
rect 675482 355816 675538 355872
rect 675298 355408 675354 355464
rect 675482 355000 675538 355056
rect 675114 354592 675170 354648
rect 675298 353776 675354 353832
rect 675482 353368 675538 353424
rect 675482 352552 675538 352608
rect 675298 351328 675354 351384
rect 675482 350512 675538 350568
rect 675482 349308 675538 349344
rect 675482 349288 675484 349308
rect 675484 349288 675536 349308
rect 675536 349288 675538 349308
rect 675482 348900 675538 348936
rect 675482 348880 675484 348900
rect 675484 348880 675536 348900
rect 675536 348880 675538 348900
rect 683118 347656 683174 347712
rect 675482 347248 675538 347304
rect 675850 342080 675906 342136
rect 675758 340312 675814 340368
rect 675666 339360 675722 339416
rect 675574 337728 675630 337784
rect 675758 336640 675814 336696
rect 675758 332288 675814 332344
rect 675758 326848 675814 326904
rect 675482 313656 675538 313712
rect 675482 313284 675484 313304
rect 675484 313284 675536 313304
rect 675536 313284 675538 313304
rect 675482 313248 675538 313284
rect 675298 312840 675354 312896
rect 675482 312468 675484 312488
rect 675484 312468 675536 312488
rect 675536 312468 675538 312488
rect 675482 312432 675538 312468
rect 675482 312024 675538 312080
rect 674654 311616 674710 311672
rect 675482 311208 675538 311264
rect 675298 310836 675300 310856
rect 675300 310836 675352 310856
rect 675352 310836 675354 310856
rect 675298 310800 675354 310836
rect 675298 310392 675354 310448
rect 675482 310020 675484 310040
rect 675484 310020 675536 310040
rect 675536 310020 675538 310040
rect 675482 309984 675538 310020
rect 675482 309576 675538 309632
rect 675482 309168 675538 309224
rect 675022 307944 675078 308000
rect 675022 307536 675078 307592
rect 674470 306312 674526 306368
rect 674654 304272 674710 304328
rect 676034 308352 676090 308408
rect 675482 305516 675538 305552
rect 675482 305496 675484 305516
rect 675484 305496 675536 305516
rect 675536 305496 675538 305516
rect 676034 304680 676090 304736
rect 675482 303884 675538 303920
rect 675482 303864 675484 303884
rect 675484 303864 675536 303884
rect 675536 303864 675538 303884
rect 675482 303476 675538 303512
rect 675482 303456 675484 303476
rect 675484 303456 675536 303476
rect 675536 303456 675538 303476
rect 676034 302912 676090 302968
rect 675482 302232 675538 302288
rect 678242 307128 678298 307184
rect 676402 305904 676458 305960
rect 676402 301552 676458 301608
rect 675482 300600 675538 300656
rect 676218 300600 676274 300656
rect 681002 306720 681058 306776
rect 680358 299376 680414 299432
rect 678242 297336 678298 297392
rect 683118 302640 683174 302696
rect 675850 296520 675906 296576
rect 675574 295296 675630 295352
rect 675758 291488 675814 291544
rect 675758 290944 675814 291000
rect 675758 287000 675814 287056
rect 675390 286456 675446 286512
rect 675114 285504 675170 285560
rect 675758 283600 675814 283656
rect 675666 282784 675722 282840
rect 675666 281560 675722 281616
rect 675482 268640 675538 268696
rect 675482 268268 675484 268288
rect 675484 268268 675536 268288
rect 675536 268268 675538 268288
rect 675482 268232 675538 268268
rect 675482 267844 675538 267880
rect 675482 267824 675484 267844
rect 675484 267824 675536 267844
rect 675536 267824 675538 267844
rect 675482 267416 675538 267472
rect 675298 267008 675354 267064
rect 675482 266620 675538 266656
rect 675482 266600 675484 266620
rect 675484 266600 675536 266620
rect 675536 266600 675538 266620
rect 675482 266192 675538 266248
rect 675298 265784 675354 265840
rect 675482 265412 675484 265432
rect 675484 265412 675536 265432
rect 675536 265412 675538 265432
rect 675482 265376 675538 265412
rect 675482 265004 675484 265024
rect 675484 265004 675536 265024
rect 675536 265004 675538 265024
rect 675482 264968 675538 265004
rect 675482 264560 675538 264616
rect 676218 263200 676274 263256
rect 675482 262540 675538 262576
rect 675482 262520 675484 262540
rect 675484 262520 675536 262540
rect 675536 262520 675538 262540
rect 675482 262132 675538 262168
rect 675482 262112 675484 262132
rect 675484 262112 675536 262132
rect 675536 262112 675538 262132
rect 674470 261296 674526 261352
rect 674838 261024 674894 261080
rect 675850 261044 675906 261080
rect 675850 261024 675852 261044
rect 675852 261024 675904 261044
rect 675904 261024 675906 261044
rect 674654 259256 674710 259312
rect 675482 260500 675538 260536
rect 675482 260480 675484 260500
rect 675484 260480 675536 260500
rect 675536 260480 675538 260500
rect 675482 260072 675538 260128
rect 675482 259684 675538 259720
rect 675482 259664 675484 259684
rect 675484 259664 675536 259684
rect 675536 259664 675538 259684
rect 676402 262792 676458 262848
rect 675022 253952 675078 254008
rect 675482 258868 675538 258904
rect 675482 258848 675484 258868
rect 675484 258848 675536 258868
rect 675536 258848 675538 258868
rect 675482 258460 675538 258496
rect 675482 258440 675484 258460
rect 675484 258440 675536 258460
rect 675536 258440 675538 258460
rect 683118 257488 683174 257544
rect 675482 257216 675538 257272
rect 675850 253952 675906 254008
rect 675206 249736 675262 249792
rect 674562 242664 674618 242720
rect 675574 249464 675630 249520
rect 675390 248240 675446 248296
rect 675758 246608 675814 246664
rect 675390 245656 675446 245712
rect 675298 243208 675354 243264
rect 675482 242664 675538 242720
rect 675482 241984 675538 242040
rect 675114 241712 675170 241768
rect 675390 238584 675446 238640
rect 675666 223488 675722 223544
rect 675114 223080 675170 223136
rect 675482 222672 675538 222728
rect 675298 222264 675354 222320
rect 675298 221856 675354 221912
rect 675482 221448 675538 221504
rect 675482 221060 675538 221096
rect 675482 221040 675484 221060
rect 675484 221040 675536 221060
rect 675536 221040 675538 221060
rect 675298 220632 675354 220688
rect 674654 220224 674710 220280
rect 674470 215328 674526 215384
rect 675482 219836 675538 219872
rect 675482 219816 675484 219836
rect 675484 219816 675536 219836
rect 675536 219816 675538 219836
rect 675482 219444 675484 219464
rect 675484 219444 675536 219464
rect 675536 219444 675538 219464
rect 675482 219408 675538 219444
rect 675574 219000 675630 219056
rect 675206 217776 675262 217832
rect 674930 214104 674986 214160
rect 675390 216980 675446 217016
rect 675390 216960 675392 216980
rect 675392 216960 675444 216980
rect 675444 216960 675446 216980
rect 675390 216164 675446 216200
rect 675390 216144 675392 216164
rect 675392 216144 675444 216164
rect 675444 216144 675446 216164
rect 675758 218184 675814 218240
rect 675482 213716 675538 213752
rect 675482 213696 675484 213716
rect 675484 213696 675536 213716
rect 675536 213696 675538 213716
rect 675482 213308 675538 213344
rect 675482 213288 675484 213308
rect 675484 213288 675536 213308
rect 675536 213288 675538 213308
rect 675482 212084 675538 212120
rect 675482 212064 675484 212084
rect 675484 212064 675536 212084
rect 675536 212064 675538 212084
rect 676034 214920 676090 214976
rect 683118 212472 683174 212528
rect 676034 211384 676090 211440
rect 683118 211112 683174 211168
rect 675758 204992 675814 205048
rect 675758 199960 675814 200016
rect 675758 198328 675814 198384
rect 675758 196968 675814 197024
rect 675114 193296 675170 193352
rect 675758 193160 675814 193216
rect 675666 192752 675722 192808
rect 675850 190032 675906 190088
rect 675298 178472 675354 178528
rect 675482 178064 675538 178120
rect 683118 177656 683174 177712
rect 675298 177248 675354 177304
rect 675482 176840 675538 176896
rect 674746 176024 674802 176080
rect 674562 175616 674618 175672
rect 674470 174392 674526 174448
rect 669226 107652 669228 107672
rect 669228 107652 669280 107672
rect 669280 107652 669282 107672
rect 669226 107616 669282 107652
rect 675482 175228 675538 175264
rect 675482 175208 675484 175228
rect 675484 175208 675536 175228
rect 675536 175208 675538 175228
rect 675298 173984 675354 174040
rect 675114 172760 675170 172816
rect 675850 173168 675906 173224
rect 675482 171964 675538 172000
rect 675482 171944 675484 171964
rect 675484 171944 675536 171964
rect 675536 171944 675538 171964
rect 675482 171164 675484 171184
rect 675484 171164 675536 171184
rect 675536 171164 675538 171184
rect 675482 171128 675538 171164
rect 675482 170332 675538 170368
rect 675482 170312 675484 170332
rect 675484 170312 675536 170332
rect 675536 170312 675538 170332
rect 675482 169108 675538 169144
rect 675482 169088 675484 169108
rect 675484 169088 675536 169108
rect 675536 169088 675538 169108
rect 675482 168700 675538 168736
rect 675482 168680 675484 168700
rect 675484 168680 675536 168700
rect 675536 168680 675538 168700
rect 675482 168292 675538 168328
rect 675482 168272 675484 168292
rect 675484 168272 675536 168292
rect 675536 168272 675538 168292
rect 675482 167884 675538 167920
rect 675482 167864 675484 167884
rect 675484 167864 675536 167884
rect 675536 167864 675538 167884
rect 675482 167048 675538 167104
rect 678242 171536 678298 171592
rect 676678 169904 676734 169960
rect 676678 166368 676734 166424
rect 675850 161336 675906 161392
rect 675574 160112 675630 160168
rect 675758 156440 675814 156496
rect 675758 155624 675814 155680
rect 675666 153040 675722 153096
rect 675758 151408 675814 151464
rect 675758 148416 675814 148472
rect 675666 147600 675722 147656
rect 675298 133320 675354 133376
rect 675482 132948 675484 132968
rect 675484 132948 675536 132968
rect 675536 132948 675538 132968
rect 675482 132912 675538 132948
rect 675482 132504 675538 132560
rect 675298 132096 675354 132152
rect 674654 131280 674710 131336
rect 675482 131688 675538 131744
rect 675482 130892 675538 130928
rect 675482 130872 675484 130892
rect 675484 130872 675536 130892
rect 675536 130872 675538 130892
rect 675482 130464 675538 130520
rect 675482 130056 675538 130112
rect 674470 129648 674526 129704
rect 675482 129240 675538 129296
rect 679622 127744 679678 127800
rect 674838 127608 674894 127664
rect 674378 125160 674434 125216
rect 673366 106256 673422 106312
rect 668950 105984 669006 106040
rect 674654 123528 674710 123584
rect 675022 126384 675078 126440
rect 675482 125996 675538 126032
rect 675482 125976 675484 125996
rect 675484 125976 675536 125996
rect 675536 125976 675538 125996
rect 675482 125604 675484 125624
rect 675484 125604 675536 125624
rect 675536 125604 675538 125624
rect 675482 125568 675538 125604
rect 675482 124772 675538 124808
rect 675482 124752 675484 124772
rect 675484 124752 675536 124772
rect 675536 124752 675538 124772
rect 675298 123936 675354 123992
rect 675482 123120 675538 123176
rect 675298 122440 675354 122496
rect 677598 122032 677654 122088
rect 675482 121896 675538 121952
rect 683118 126520 683174 126576
rect 683118 124480 683174 124536
rect 683118 124072 683174 124128
rect 683118 117272 683174 117328
rect 677598 117000 677654 117056
rect 675298 113056 675354 113112
rect 675758 110336 675814 110392
rect 675666 108024 675722 108080
rect 675114 106256 675170 106312
rect 669134 104488 669190 104544
rect 675758 103128 675814 103184
rect 668582 102856 668638 102912
rect 675666 102584 675722 102640
rect 675758 101360 675814 101416
rect 591302 53080 591358 53136
rect 497554 50496 497610 50552
rect 549258 50496 549314 50552
rect 499578 46960 499634 47016
rect 596178 48864 596234 48920
rect 594062 47776 594118 47832
rect 592682 46416 592738 46472
rect 600318 49136 600374 49192
rect 598938 48048 598994 48104
rect 597558 46144 597614 46200
rect 445022 45056 445078 45112
rect 603078 51720 603134 51776
rect 601882 50224 601938 50280
rect 601698 44784 601754 44840
rect 626078 94424 626134 94480
rect 637026 96872 637082 96928
rect 635922 95648 635978 95704
rect 626446 95376 626502 95432
rect 642638 95104 642694 95160
rect 626446 93472 626502 93528
rect 626262 92520 626318 92576
rect 625434 91568 625490 91624
rect 626446 90616 626502 90672
rect 626446 89684 626502 89720
rect 626446 89664 626448 89684
rect 626448 89664 626500 89684
rect 626500 89664 626502 89684
rect 624974 88576 625030 88632
rect 626446 87896 626502 87952
rect 625618 86944 625674 87000
rect 626446 85992 626502 86048
rect 626446 85040 626502 85096
rect 626446 84088 626502 84144
rect 626262 83136 626318 83192
rect 644478 92112 644534 92168
rect 644754 89664 644810 89720
rect 643926 87080 643982 87136
rect 643466 84632 643522 84688
rect 643098 82728 643154 82784
rect 628562 81640 628618 81696
rect 629206 80824 629262 80880
rect 633898 77696 633954 77752
rect 637118 78512 637174 78568
rect 646134 71712 646190 71768
rect 646870 74432 646926 74488
rect 647422 72936 647478 72992
rect 646318 70352 646374 70408
rect 647606 68448 647662 68504
rect 646134 66000 646190 66056
rect 653954 94152 654010 94208
rect 654322 93336 654378 93392
rect 654138 92520 654194 92576
rect 654322 91432 654378 91488
rect 654138 90616 654194 90672
rect 655794 89800 655850 89856
rect 663246 93064 663302 93120
rect 663798 90344 663854 90400
rect 663982 88984 664038 89040
rect 665178 91704 665234 91760
rect 665730 93336 665786 93392
rect 665362 90616 665418 90672
rect 648986 66952 649042 67008
rect 648802 63960 648858 64016
rect 624422 47504 624478 47560
rect 663798 48456 663854 48512
rect 662602 47776 662658 47832
rect 662418 47368 662474 47424
rect 474462 43424 474518 43480
rect 604458 43424 604514 43480
rect 409602 42744 409658 42800
rect 411074 42744 411130 42800
rect 416594 42744 416650 42800
rect 464894 42744 464950 42800
rect 518622 42336 518678 42392
rect 460570 42064 460626 42120
rect 471610 42064 471666 42120
rect 514942 42064 514998 42120
rect 520462 42064 520518 42120
rect 525982 42064 526038 42120
rect 529570 42064 529626 42120
rect 521658 41928 521714 41984
<< metal3 >>
rect 504541 1007042 504607 1007045
rect 559649 1007042 559715 1007045
rect 504436 1007040 504607 1007042
rect 504436 1006984 504546 1007040
rect 504602 1006984 504607 1007040
rect 504436 1006982 504607 1006984
rect 559452 1007040 559715 1007042
rect 559452 1006984 559654 1007040
rect 559710 1006984 559715 1007040
rect 559452 1006982 559715 1006984
rect 504541 1006979 504607 1006982
rect 559649 1006979 559715 1006982
rect 151721 1006906 151787 1006909
rect 427997 1006906 428063 1006909
rect 506197 1006906 506263 1006909
rect 151721 1006904 151892 1006906
rect 151721 1006848 151726 1006904
rect 151782 1006848 151892 1006904
rect 151721 1006846 151892 1006848
rect 427800 1006904 428063 1006906
rect 427800 1006848 428002 1006904
rect 428058 1006848 428063 1006904
rect 427800 1006846 428063 1006848
rect 506000 1006904 506263 1006906
rect 506000 1006848 506202 1006904
rect 506258 1006848 506263 1006904
rect 506000 1006846 506263 1006848
rect 151721 1006843 151787 1006846
rect 427997 1006843 428063 1006846
rect 506197 1006843 506263 1006846
rect 555141 1006906 555207 1006909
rect 555141 1006904 555404 1006906
rect 555141 1006848 555146 1006904
rect 555202 1006848 555404 1006904
rect 555141 1006846 555404 1006848
rect 555141 1006843 555207 1006846
rect 307753 1006770 307819 1006773
rect 357709 1006770 357775 1006773
rect 430849 1006770 430915 1006773
rect 557165 1006770 557231 1006773
rect 307753 1006768 307924 1006770
rect 307753 1006712 307758 1006768
rect 307814 1006712 307924 1006768
rect 307753 1006710 307924 1006712
rect 357709 1006768 357972 1006770
rect 357709 1006712 357714 1006768
rect 357770 1006712 357972 1006768
rect 357709 1006710 357972 1006712
rect 430849 1006768 431020 1006770
rect 430849 1006712 430854 1006768
rect 430910 1006712 431020 1006768
rect 430849 1006710 431020 1006712
rect 557060 1006768 557231 1006770
rect 557060 1006712 557170 1006768
rect 557226 1006712 557231 1006768
rect 557060 1006710 557231 1006712
rect 307753 1006707 307819 1006710
rect 357709 1006707 357775 1006710
rect 430849 1006707 430915 1006710
rect 557165 1006707 557231 1006710
rect 427169 1006634 427235 1006637
rect 426972 1006632 427235 1006634
rect 426972 1006576 427174 1006632
rect 427230 1006576 427235 1006632
rect 426972 1006574 427235 1006576
rect 427169 1006571 427235 1006574
rect 101121 1006498 101187 1006501
rect 100924 1006496 101187 1006498
rect 100924 1006440 101126 1006496
rect 101182 1006440 101187 1006496
rect 100924 1006438 101187 1006440
rect 101121 1006435 101187 1006438
rect 255313 1006498 255379 1006501
rect 304073 1006498 304139 1006501
rect 255313 1006496 255576 1006498
rect 255313 1006440 255318 1006496
rect 255374 1006440 255576 1006496
rect 255313 1006438 255576 1006440
rect 303876 1006496 304139 1006498
rect 303876 1006440 304078 1006496
rect 304134 1006440 304139 1006496
rect 303876 1006438 304139 1006440
rect 255313 1006435 255379 1006438
rect 304073 1006435 304139 1006438
rect 314653 1006498 314719 1006501
rect 361389 1006498 361455 1006501
rect 314653 1006496 314916 1006498
rect 314653 1006440 314658 1006496
rect 314714 1006440 314916 1006496
rect 314653 1006438 314916 1006440
rect 361192 1006496 361455 1006498
rect 361192 1006440 361394 1006496
rect 361450 1006440 361455 1006496
rect 361192 1006438 361455 1006440
rect 314653 1006435 314719 1006438
rect 361389 1006435 361455 1006438
rect 423489 1006498 423555 1006501
rect 501689 1006498 501755 1006501
rect 552289 1006498 552355 1006501
rect 556797 1006498 556863 1006501
rect 423489 1006496 423752 1006498
rect 423489 1006440 423494 1006496
rect 423550 1006440 423752 1006496
rect 423489 1006438 423752 1006440
rect 501492 1006496 501755 1006498
rect 501492 1006440 501694 1006496
rect 501750 1006440 501755 1006496
rect 501492 1006438 501755 1006440
rect 552092 1006496 552355 1006498
rect 552092 1006440 552294 1006496
rect 552350 1006440 552355 1006496
rect 552092 1006438 552355 1006440
rect 556600 1006496 556863 1006498
rect 556600 1006440 556802 1006496
rect 556858 1006440 556863 1006496
rect 556600 1006438 556863 1006440
rect 423489 1006435 423555 1006438
rect 501689 1006435 501755 1006438
rect 552289 1006435 552355 1006438
rect 556797 1006435 556863 1006438
rect 100293 1006362 100359 1006365
rect 100096 1006360 100359 1006362
rect 100096 1006304 100298 1006360
rect 100354 1006304 100359 1006360
rect 100096 1006302 100359 1006304
rect 100293 1006299 100359 1006302
rect 150893 1006362 150959 1006365
rect 152089 1006362 152155 1006365
rect 158253 1006362 158319 1006365
rect 210417 1006362 210483 1006365
rect 150893 1006360 151156 1006362
rect 150893 1006304 150898 1006360
rect 150954 1006304 151156 1006360
rect 150893 1006302 151156 1006304
rect 152089 1006360 152352 1006362
rect 152089 1006304 152094 1006360
rect 152150 1006304 152352 1006360
rect 152089 1006302 152352 1006304
rect 158056 1006360 158319 1006362
rect 158056 1006304 158258 1006360
rect 158314 1006304 158319 1006360
rect 158056 1006302 158319 1006304
rect 210220 1006360 210483 1006362
rect 210220 1006304 210422 1006360
rect 210478 1006304 210483 1006360
rect 210220 1006302 210483 1006304
rect 150893 1006299 150959 1006302
rect 152089 1006299 152155 1006302
rect 158253 1006299 158319 1006302
rect 210417 1006299 210483 1006302
rect 254117 1006362 254183 1006365
rect 305269 1006362 305335 1006365
rect 306925 1006362 306991 1006365
rect 424317 1006362 424383 1006365
rect 502149 1006362 502215 1006365
rect 554313 1006362 554379 1006365
rect 254117 1006360 254380 1006362
rect 254117 1006304 254122 1006360
rect 254178 1006304 254380 1006360
rect 254117 1006302 254380 1006304
rect 305269 1006360 305532 1006362
rect 305269 1006304 305274 1006360
rect 305330 1006304 305532 1006360
rect 305269 1006302 305532 1006304
rect 306728 1006360 306991 1006362
rect 306728 1006304 306930 1006360
rect 306986 1006304 306991 1006360
rect 306728 1006302 306991 1006304
rect 424120 1006360 424383 1006362
rect 424120 1006304 424322 1006360
rect 424378 1006304 424383 1006360
rect 424120 1006302 424383 1006304
rect 501952 1006360 502215 1006362
rect 501952 1006304 502154 1006360
rect 502210 1006304 502215 1006360
rect 501952 1006302 502215 1006304
rect 554116 1006360 554379 1006362
rect 554116 1006304 554318 1006360
rect 554374 1006304 554379 1006360
rect 554116 1006302 554379 1006304
rect 254117 1006299 254183 1006302
rect 305269 1006299 305335 1006302
rect 306925 1006299 306991 1006302
rect 424317 1006299 424383 1006302
rect 502149 1006299 502215 1006302
rect 554313 1006299 554379 1006302
rect 99465 1006226 99531 1006229
rect 103973 1006226 104039 1006229
rect 106825 1006226 106891 1006229
rect 99465 1006224 99728 1006226
rect 99465 1006168 99470 1006224
rect 99526 1006168 99728 1006224
rect 99465 1006166 99728 1006168
rect 103973 1006224 104236 1006226
rect 103973 1006168 103978 1006224
rect 104034 1006168 104236 1006224
rect 103973 1006166 104236 1006168
rect 106628 1006224 106891 1006226
rect 106628 1006168 106830 1006224
rect 106886 1006168 106891 1006224
rect 106628 1006166 106891 1006168
rect 99465 1006163 99531 1006166
rect 103973 1006163 104039 1006166
rect 106825 1006163 106891 1006166
rect 151261 1006226 151327 1006229
rect 159449 1006226 159515 1006229
rect 160277 1006226 160343 1006229
rect 151261 1006224 151524 1006226
rect 151261 1006168 151266 1006224
rect 151322 1006168 151524 1006224
rect 151261 1006166 151524 1006168
rect 159252 1006224 159515 1006226
rect 159252 1006168 159454 1006224
rect 159510 1006168 159515 1006224
rect 159252 1006166 159515 1006168
rect 160080 1006224 160343 1006226
rect 160080 1006168 160282 1006224
rect 160338 1006168 160343 1006224
rect 160080 1006166 160343 1006168
rect 151261 1006163 151327 1006166
rect 159449 1006163 159515 1006166
rect 160277 1006163 160343 1006166
rect 208393 1006226 208459 1006229
rect 253657 1006226 253723 1006229
rect 262673 1006226 262739 1006229
rect 208393 1006224 208656 1006226
rect 208393 1006168 208398 1006224
rect 208454 1006168 208656 1006224
rect 208393 1006166 208656 1006168
rect 253657 1006224 253920 1006226
rect 253657 1006168 253662 1006224
rect 253718 1006168 253920 1006224
rect 253657 1006166 253920 1006168
rect 262476 1006224 262739 1006226
rect 262476 1006168 262678 1006224
rect 262734 1006168 262739 1006224
rect 262476 1006166 262739 1006168
rect 208393 1006163 208459 1006166
rect 253657 1006163 253723 1006166
rect 262673 1006163 262739 1006166
rect 311801 1006226 311867 1006229
rect 314653 1006226 314719 1006229
rect 365069 1006226 365135 1006229
rect 500493 1006226 500559 1006229
rect 311801 1006224 312064 1006226
rect 311801 1006168 311806 1006224
rect 311862 1006168 312064 1006224
rect 311801 1006166 312064 1006168
rect 314548 1006224 314719 1006226
rect 314548 1006168 314658 1006224
rect 314714 1006168 314719 1006224
rect 314548 1006166 314719 1006168
rect 364872 1006224 365135 1006226
rect 364872 1006168 365074 1006224
rect 365130 1006168 365135 1006224
rect 364872 1006166 365135 1006168
rect 500296 1006224 500559 1006226
rect 500296 1006168 500498 1006224
rect 500554 1006168 500559 1006224
rect 500296 1006166 500559 1006168
rect 311801 1006163 311867 1006166
rect 314653 1006163 314719 1006166
rect 365069 1006163 365135 1006166
rect 500493 1006163 500559 1006166
rect 551461 1006226 551527 1006229
rect 560845 1006226 560911 1006229
rect 551461 1006224 551724 1006226
rect 551461 1006168 551466 1006224
rect 551522 1006168 551724 1006224
rect 551461 1006166 551724 1006168
rect 560740 1006224 560911 1006226
rect 560740 1006168 560850 1006224
rect 560906 1006168 560911 1006224
rect 560740 1006166 560911 1006168
rect 551461 1006163 551527 1006166
rect 560845 1006163 560911 1006166
rect 98269 1006090 98335 1006093
rect 104801 1006090 104867 1006093
rect 107653 1006090 107719 1006093
rect 98269 1006088 98900 1006090
rect 98269 1006032 98274 1006088
rect 98330 1006032 98900 1006088
rect 98269 1006030 98900 1006032
rect 104801 1006088 104972 1006090
rect 104801 1006032 104806 1006088
rect 104862 1006032 104972 1006088
rect 104801 1006030 104972 1006032
rect 107456 1006088 107719 1006090
rect 107456 1006032 107658 1006088
rect 107714 1006032 107719 1006088
rect 107456 1006030 107719 1006032
rect 98269 1006027 98335 1006030
rect 104801 1006027 104867 1006030
rect 107653 1006027 107719 1006030
rect 146937 1006090 147003 1006093
rect 148869 1006090 148935 1006093
rect 150065 1006090 150131 1006093
rect 158621 1006090 158687 1006093
rect 201033 1006090 201099 1006093
rect 252461 1006090 252527 1006093
rect 261845 1006090 261911 1006093
rect 146937 1006088 148935 1006090
rect 146937 1006032 146942 1006088
rect 146998 1006032 148874 1006088
rect 148930 1006032 148935 1006088
rect 146937 1006030 148935 1006032
rect 149868 1006088 150328 1006090
rect 149868 1006032 150070 1006088
rect 150126 1006032 150328 1006088
rect 149868 1006030 150328 1006032
rect 158621 1006088 158884 1006090
rect 158621 1006032 158626 1006088
rect 158682 1006032 158884 1006088
rect 158621 1006030 158884 1006032
rect 201033 1006088 201756 1006090
rect 201033 1006032 201038 1006088
rect 201094 1006032 201756 1006088
rect 201033 1006030 201756 1006032
rect 252461 1006088 253092 1006090
rect 252461 1006032 252466 1006088
rect 252522 1006032 253092 1006088
rect 252461 1006030 253092 1006032
rect 261648 1006088 261911 1006090
rect 261648 1006032 261850 1006088
rect 261906 1006032 261911 1006088
rect 261648 1006030 261911 1006032
rect 146937 1006027 147003 1006030
rect 148869 1006027 148935 1006030
rect 150065 1006027 150131 1006030
rect 158621 1006027 158687 1006030
rect 201033 1006027 201099 1006030
rect 252461 1006027 252527 1006030
rect 261845 1006027 261911 1006030
rect 301497 1006090 301563 1006093
rect 303245 1006090 303311 1006093
rect 301497 1006088 303311 1006090
rect 301497 1006032 301502 1006088
rect 301558 1006032 303250 1006088
rect 303306 1006032 303311 1006088
rect 301497 1006030 303311 1006032
rect 301497 1006027 301563 1006030
rect 303245 1006027 303311 1006030
rect 304073 1006090 304139 1006093
rect 305269 1006090 305335 1006093
rect 354857 1006090 354923 1006093
rect 357341 1006090 357407 1006093
rect 422661 1006090 422727 1006093
rect 423489 1006090 423555 1006093
rect 429193 1006090 429259 1006093
rect 499665 1006090 499731 1006093
rect 505369 1006090 505435 1006093
rect 551093 1006090 551159 1006093
rect 304073 1006088 304704 1006090
rect 304073 1006032 304078 1006088
rect 304134 1006032 304704 1006088
rect 304073 1006030 304704 1006032
rect 305164 1006088 305335 1006090
rect 305164 1006032 305274 1006088
rect 305330 1006032 305335 1006088
rect 305164 1006030 305335 1006032
rect 354660 1006088 355120 1006090
rect 354660 1006032 354862 1006088
rect 354918 1006032 355120 1006088
rect 354660 1006030 355120 1006032
rect 357144 1006088 357407 1006090
rect 357144 1006032 357346 1006088
rect 357402 1006032 357407 1006088
rect 357144 1006030 357407 1006032
rect 422096 1006088 422727 1006090
rect 422096 1006032 422666 1006088
rect 422722 1006032 422727 1006088
rect 422096 1006030 422727 1006032
rect 423292 1006088 423555 1006090
rect 423292 1006032 423494 1006088
rect 423550 1006032 423555 1006088
rect 423292 1006030 423555 1006032
rect 428996 1006088 429259 1006090
rect 428996 1006032 429198 1006088
rect 429254 1006032 429259 1006088
rect 428996 1006030 429259 1006032
rect 499100 1006088 499731 1006090
rect 499100 1006032 499670 1006088
rect 499726 1006032 499731 1006088
rect 499100 1006030 499731 1006032
rect 505172 1006088 505435 1006090
rect 505172 1006032 505374 1006088
rect 505430 1006032 505435 1006088
rect 505172 1006030 505435 1006032
rect 550436 1006088 551159 1006090
rect 550436 1006032 551098 1006088
rect 551154 1006032 551159 1006088
rect 550436 1006030 551159 1006032
rect 304073 1006027 304139 1006030
rect 305269 1006027 305335 1006030
rect 354857 1006027 354923 1006030
rect 357341 1006027 357407 1006030
rect 422661 1006027 422727 1006030
rect 423489 1006027 423555 1006030
rect 429193 1006027 429259 1006030
rect 499665 1006027 499731 1006030
rect 505369 1006027 505435 1006030
rect 551093 1006027 551159 1006030
rect 553117 1006090 553183 1006093
rect 553117 1006088 553380 1006090
rect 553117 1006032 553122 1006088
rect 553178 1006032 553380 1006088
rect 553117 1006030 553380 1006032
rect 553117 1006027 553183 1006030
rect 428365 1005818 428431 1005821
rect 428260 1005816 428431 1005818
rect 428260 1005760 428370 1005816
rect 428426 1005760 428431 1005816
rect 428260 1005758 428431 1005760
rect 428365 1005755 428431 1005758
rect 509049 1005818 509115 1005821
rect 509049 1005816 509312 1005818
rect 509049 1005760 509054 1005816
rect 509110 1005760 509312 1005816
rect 509049 1005758 509312 1005760
rect 509049 1005755 509115 1005758
rect 360561 1005682 360627 1005685
rect 427537 1005682 427603 1005685
rect 360364 1005680 360627 1005682
rect 360364 1005624 360566 1005680
rect 360622 1005624 360627 1005680
rect 360364 1005622 360627 1005624
rect 427340 1005680 427603 1005682
rect 427340 1005624 427542 1005680
rect 427598 1005624 427603 1005680
rect 427340 1005622 427603 1005624
rect 360561 1005619 360627 1005622
rect 427537 1005619 427603 1005622
rect 555969 1005682 556035 1005685
rect 555969 1005680 556232 1005682
rect 555969 1005624 555974 1005680
rect 556030 1005624 556232 1005680
rect 555969 1005622 556232 1005624
rect 555969 1005619 556035 1005622
rect 359733 1005546 359799 1005549
rect 430849 1005546 430915 1005549
rect 505001 1005546 505067 1005549
rect 359628 1005544 359799 1005546
rect 359628 1005488 359738 1005544
rect 359794 1005488 359799 1005544
rect 359628 1005486 359799 1005488
rect 430652 1005544 430915 1005546
rect 430652 1005488 430854 1005544
rect 430910 1005488 430915 1005544
rect 430652 1005486 430915 1005488
rect 504804 1005544 505067 1005546
rect 504804 1005488 505006 1005544
rect 505062 1005488 505067 1005544
rect 504804 1005486 505067 1005488
rect 359733 1005483 359799 1005486
rect 430849 1005483 430915 1005486
rect 505001 1005483 505067 1005486
rect 356513 1005410 356579 1005413
rect 425513 1005410 425579 1005413
rect 508221 1005410 508287 1005413
rect 555141 1005410 555207 1005413
rect 356316 1005408 356579 1005410
rect 356316 1005352 356518 1005408
rect 356574 1005352 356579 1005408
rect 356316 1005350 356579 1005352
rect 425316 1005408 425579 1005410
rect 425316 1005352 425518 1005408
rect 425574 1005352 425579 1005408
rect 425316 1005350 425579 1005352
rect 508116 1005408 508287 1005410
rect 508116 1005352 508226 1005408
rect 508282 1005352 508287 1005408
rect 508116 1005350 508287 1005352
rect 555036 1005408 555207 1005410
rect 555036 1005352 555146 1005408
rect 555202 1005352 555207 1005408
rect 555036 1005350 555207 1005352
rect 356513 1005347 356579 1005350
rect 425513 1005347 425579 1005350
rect 508221 1005347 508287 1005350
rect 555141 1005347 555207 1005350
rect 152917 1005274 152983 1005277
rect 263041 1005274 263107 1005277
rect 152917 1005272 153180 1005274
rect 152917 1005216 152922 1005272
rect 152978 1005216 153180 1005272
rect 152917 1005214 153180 1005216
rect 262844 1005272 263107 1005274
rect 262844 1005216 263046 1005272
rect 263102 1005216 263107 1005272
rect 262844 1005214 263107 1005216
rect 152917 1005211 152983 1005214
rect 263041 1005211 263107 1005214
rect 307293 1005274 307359 1005277
rect 356881 1005274 356947 1005277
rect 430021 1005274 430087 1005277
rect 307293 1005272 307556 1005274
rect 307293 1005216 307298 1005272
rect 307354 1005216 307556 1005272
rect 307293 1005214 307556 1005216
rect 356684 1005272 356947 1005274
rect 356684 1005216 356886 1005272
rect 356942 1005216 356947 1005272
rect 356684 1005214 356947 1005216
rect 429824 1005272 430087 1005274
rect 429824 1005216 430026 1005272
rect 430082 1005216 430087 1005272
rect 429824 1005214 430087 1005216
rect 307293 1005211 307359 1005214
rect 356881 1005211 356947 1005214
rect 430021 1005211 430087 1005214
rect 432045 1005274 432111 1005277
rect 500493 1005274 500559 1005277
rect 432045 1005272 432308 1005274
rect 432045 1005216 432050 1005272
rect 432106 1005216 432308 1005272
rect 432045 1005214 432308 1005216
rect 500493 1005272 500756 1005274
rect 500493 1005216 500498 1005272
rect 500554 1005216 500756 1005272
rect 500493 1005214 500756 1005216
rect 432045 1005211 432111 1005214
rect 500493 1005211 500559 1005214
rect 153745 1005138 153811 1005141
rect 363413 1005138 363479 1005141
rect 153745 1005136 153916 1005138
rect 153745 1005080 153750 1005136
rect 153806 1005080 153916 1005136
rect 153745 1005078 153916 1005080
rect 363308 1005136 363479 1005138
rect 363308 1005080 363418 1005136
rect 363474 1005080 363479 1005136
rect 363308 1005078 363479 1005080
rect 153745 1005075 153811 1005078
rect 363413 1005075 363479 1005078
rect 365069 1005138 365135 1005141
rect 424685 1005138 424751 1005141
rect 431677 1005138 431743 1005141
rect 507025 1005138 507091 1005141
rect 365069 1005136 365332 1005138
rect 365069 1005080 365074 1005136
rect 365130 1005080 365332 1005136
rect 365069 1005078 365332 1005080
rect 424580 1005136 424751 1005138
rect 424580 1005080 424690 1005136
rect 424746 1005080 424751 1005136
rect 424580 1005078 424751 1005080
rect 431480 1005136 431743 1005138
rect 431480 1005080 431682 1005136
rect 431738 1005080 431743 1005136
rect 431480 1005078 431743 1005080
rect 506828 1005136 507091 1005138
rect 506828 1005080 507030 1005136
rect 507086 1005080 507091 1005136
rect 506828 1005078 507091 1005080
rect 365069 1005075 365135 1005078
rect 424685 1005075 424751 1005078
rect 431677 1005075 431743 1005078
rect 507025 1005075 507091 1005078
rect 152917 1005002 152983 1005005
rect 152720 1005000 152983 1005002
rect 152720 1004944 152922 1005000
rect 152978 1004944 152983 1005000
rect 152720 1004942 152983 1004944
rect 152917 1004939 152983 1004942
rect 160645 1005002 160711 1005005
rect 209221 1005002 209287 1005005
rect 308949 1005002 309015 1005005
rect 160645 1005000 160908 1005002
rect 160645 1004944 160650 1005000
rect 160706 1004944 160908 1005000
rect 160645 1004942 160908 1004944
rect 209221 1005000 209484 1005002
rect 209221 1004944 209226 1005000
rect 209282 1004944 209484 1005000
rect 209221 1004942 209484 1004944
rect 308752 1005000 309015 1005002
rect 308752 1004944 308954 1005000
rect 309010 1004944 309015 1005000
rect 308752 1004942 309015 1004944
rect 160645 1004939 160711 1004942
rect 209221 1004939 209287 1004942
rect 308949 1004939 309015 1004942
rect 355685 1005002 355751 1005005
rect 361389 1005002 361455 1005005
rect 429193 1005002 429259 1005005
rect 508221 1005002 508287 1005005
rect 355685 1005000 355948 1005002
rect 355685 1004944 355690 1005000
rect 355746 1004944 355948 1005000
rect 355685 1004942 355948 1004944
rect 361389 1005000 361652 1005002
rect 361389 1004944 361394 1005000
rect 361450 1004944 361652 1005000
rect 361389 1004942 361652 1004944
rect 429193 1005000 429456 1005002
rect 429193 1004944 429198 1005000
rect 429254 1004944 429456 1005000
rect 429193 1004942 429456 1004944
rect 508221 1005000 508484 1005002
rect 508221 1004944 508226 1005000
rect 508282 1004944 508484 1005000
rect 508221 1004942 508484 1004944
rect 355685 1004939 355751 1004942
rect 361389 1004939 361455 1004942
rect 429193 1004939 429259 1004942
rect 508221 1004939 508287 1004942
rect 154113 1004866 154179 1004869
rect 159449 1004866 159515 1004869
rect 207197 1004866 207263 1004869
rect 154113 1004864 154376 1004866
rect 154113 1004808 154118 1004864
rect 154174 1004808 154376 1004864
rect 154113 1004806 154376 1004808
rect 159449 1004864 159712 1004866
rect 159449 1004808 159454 1004864
rect 159510 1004808 159712 1004864
rect 159449 1004806 159712 1004808
rect 207000 1004864 207263 1004866
rect 207000 1004808 207202 1004864
rect 207258 1004808 207263 1004864
rect 207000 1004806 207263 1004808
rect 154113 1004803 154179 1004806
rect 159449 1004803 159515 1004806
rect 207197 1004803 207263 1004806
rect 306925 1004866 306991 1004869
rect 313825 1004866 313891 1004869
rect 364241 1004866 364307 1004869
rect 306925 1004864 307188 1004866
rect 306925 1004808 306930 1004864
rect 306986 1004808 307188 1004864
rect 306925 1004806 307188 1004808
rect 313628 1004864 313891 1004866
rect 313628 1004808 313830 1004864
rect 313886 1004808 313891 1004864
rect 313628 1004806 313891 1004808
rect 364044 1004864 364307 1004866
rect 364044 1004808 364246 1004864
rect 364302 1004808 364307 1004864
rect 364044 1004806 364307 1004808
rect 306925 1004803 306991 1004806
rect 313825 1004803 313891 1004806
rect 364241 1004803 364307 1004806
rect 430021 1004866 430087 1004869
rect 499665 1004866 499731 1004869
rect 507853 1004866 507919 1004869
rect 555969 1004866 556035 1004869
rect 430021 1004864 430284 1004866
rect 430021 1004808 430026 1004864
rect 430082 1004808 430284 1004864
rect 430021 1004806 430284 1004808
rect 499665 1004864 499928 1004866
rect 499665 1004808 499670 1004864
rect 499726 1004808 499928 1004864
rect 499665 1004806 499928 1004808
rect 507656 1004864 507919 1004866
rect 507656 1004808 507858 1004864
rect 507914 1004808 507919 1004864
rect 507656 1004806 507919 1004808
rect 555772 1004864 556035 1004866
rect 555772 1004808 555974 1004864
rect 556030 1004808 556035 1004864
rect 555772 1004806 556035 1004808
rect 430021 1004803 430087 1004806
rect 499665 1004803 499731 1004806
rect 507853 1004803 507919 1004806
rect 555969 1004803 556035 1004806
rect 103145 1004730 103211 1004733
rect 102948 1004728 103211 1004730
rect 102948 1004672 103150 1004728
rect 103206 1004672 103211 1004728
rect 102948 1004670 103211 1004672
rect 103145 1004667 103211 1004670
rect 108481 1004730 108547 1004733
rect 160645 1004730 160711 1004733
rect 209221 1004730 209287 1004733
rect 212533 1004730 212599 1004733
rect 108481 1004728 108652 1004730
rect 108481 1004672 108486 1004728
rect 108542 1004672 108652 1004728
rect 108481 1004670 108652 1004672
rect 160540 1004728 160711 1004730
rect 160540 1004672 160650 1004728
rect 160706 1004672 160711 1004728
rect 160540 1004670 160711 1004672
rect 209024 1004728 209287 1004730
rect 209024 1004672 209226 1004728
rect 209282 1004672 209287 1004728
rect 209024 1004670 209287 1004672
rect 212336 1004728 212599 1004730
rect 212336 1004672 212538 1004728
rect 212594 1004672 212599 1004728
rect 212336 1004670 212599 1004672
rect 108481 1004667 108547 1004670
rect 160645 1004667 160711 1004670
rect 209221 1004667 209287 1004670
rect 212533 1004667 212599 1004670
rect 308121 1004730 308187 1004733
rect 315481 1004730 315547 1004733
rect 355685 1004730 355751 1004733
rect 362585 1004730 362651 1004733
rect 308121 1004728 308384 1004730
rect 308121 1004672 308126 1004728
rect 308182 1004672 308384 1004728
rect 308121 1004670 308384 1004672
rect 315284 1004728 315547 1004730
rect 315284 1004672 315486 1004728
rect 315542 1004672 315547 1004728
rect 315284 1004670 315547 1004672
rect 355488 1004728 355751 1004730
rect 355488 1004672 355690 1004728
rect 355746 1004672 355751 1004728
rect 355488 1004670 355751 1004672
rect 362388 1004728 362651 1004730
rect 362388 1004672 362590 1004728
rect 362646 1004672 362651 1004728
rect 362388 1004670 362651 1004672
rect 308121 1004667 308187 1004670
rect 315481 1004667 315547 1004670
rect 355685 1004667 355751 1004670
rect 362585 1004667 362651 1004670
rect 422661 1004730 422727 1004733
rect 431677 1004730 431743 1004733
rect 501321 1004730 501387 1004733
rect 509049 1004730 509115 1004733
rect 510337 1004730 510403 1004733
rect 557625 1004730 557691 1004733
rect 561673 1004730 561739 1004733
rect 422661 1004728 422924 1004730
rect 422661 1004672 422666 1004728
rect 422722 1004672 422924 1004728
rect 422661 1004670 422924 1004672
rect 431677 1004728 431940 1004730
rect 431677 1004672 431682 1004728
rect 431738 1004672 431940 1004728
rect 431677 1004670 431940 1004672
rect 501124 1004728 501387 1004730
rect 501124 1004672 501326 1004728
rect 501382 1004672 501387 1004728
rect 501124 1004670 501387 1004672
rect 508852 1004728 509115 1004730
rect 508852 1004672 509054 1004728
rect 509110 1004672 509115 1004728
rect 508852 1004670 509115 1004672
rect 510140 1004728 510403 1004730
rect 510140 1004672 510342 1004728
rect 510398 1004672 510403 1004728
rect 510140 1004670 510403 1004672
rect 557428 1004728 557691 1004730
rect 557428 1004672 557630 1004728
rect 557686 1004672 557691 1004728
rect 557428 1004670 557691 1004672
rect 561476 1004728 561739 1004730
rect 561476 1004672 561678 1004728
rect 561734 1004672 561739 1004728
rect 561476 1004670 561739 1004672
rect 422661 1004667 422727 1004670
rect 431677 1004667 431743 1004670
rect 501321 1004667 501387 1004670
rect 509049 1004667 509115 1004670
rect 510337 1004667 510403 1004670
rect 557625 1004667 557691 1004670
rect 561673 1004667 561739 1004670
rect 432873 1004050 432939 1004053
rect 432676 1004048 432939 1004050
rect 432676 1003992 432878 1004048
rect 432934 1003992 432939 1004048
rect 432676 1003990 432939 1003992
rect 432873 1003987 432939 1003990
rect 425513 1003914 425579 1003917
rect 505369 1003914 505435 1003917
rect 425513 1003912 425776 1003914
rect 425513 1003856 425518 1003912
rect 425574 1003856 425776 1003912
rect 425513 1003854 425776 1003856
rect 505369 1003912 505632 1003914
rect 505369 1003856 505374 1003912
rect 505430 1003856 505632 1003912
rect 505369 1003854 505632 1003856
rect 425513 1003851 425579 1003854
rect 505369 1003851 505435 1003854
rect 558821 1002826 558887 1002829
rect 558821 1002824 559084 1002826
rect 558821 1002768 558826 1002824
rect 558882 1002768 559084 1002824
rect 558821 1002766 559084 1002768
rect 558821 1002763 558887 1002766
rect 102317 1002690 102383 1002693
rect 424685 1002690 424751 1002693
rect 557993 1002690 558059 1002693
rect 102317 1002688 102580 1002690
rect 102317 1002632 102322 1002688
rect 102378 1002632 102580 1002688
rect 102317 1002630 102580 1002632
rect 424685 1002688 424948 1002690
rect 424685 1002632 424690 1002688
rect 424746 1002632 424948 1002688
rect 424685 1002630 424948 1002632
rect 557796 1002688 558059 1002690
rect 557796 1002632 557998 1002688
rect 558054 1002632 558059 1002688
rect 557796 1002630 558059 1002632
rect 102317 1002627 102383 1002630
rect 424685 1002627 424751 1002630
rect 557993 1002627 558059 1002630
rect 101949 1002554 102015 1002557
rect 105997 1002554 106063 1002557
rect 157425 1002554 157491 1002557
rect 206369 1002554 206435 1002557
rect 255313 1002554 255379 1002557
rect 261017 1002554 261083 1002557
rect 502517 1002554 502583 1002557
rect 101752 1002552 102015 1002554
rect 101752 1002496 101954 1002552
rect 102010 1002496 102015 1002552
rect 101752 1002494 102015 1002496
rect 105892 1002552 106063 1002554
rect 105892 1002496 106002 1002552
rect 106058 1002496 106063 1002552
rect 105892 1002494 106063 1002496
rect 157228 1002552 157491 1002554
rect 157228 1002496 157430 1002552
rect 157486 1002496 157491 1002552
rect 157228 1002494 157491 1002496
rect 206172 1002552 206435 1002554
rect 206172 1002496 206374 1002552
rect 206430 1002496 206435 1002552
rect 206172 1002494 206435 1002496
rect 255116 1002552 255379 1002554
rect 255116 1002496 255318 1002552
rect 255374 1002496 255379 1002552
rect 255116 1002494 255379 1002496
rect 260820 1002552 261083 1002554
rect 260820 1002496 261022 1002552
rect 261078 1002496 261083 1002552
rect 260820 1002494 261083 1002496
rect 502412 1002552 502583 1002554
rect 502412 1002496 502522 1002552
rect 502578 1002496 502583 1002552
rect 502412 1002494 502583 1002496
rect 101949 1002491 102015 1002494
rect 105997 1002491 106063 1002494
rect 157425 1002491 157491 1002494
rect 206369 1002491 206435 1002494
rect 255313 1002491 255379 1002494
rect 261017 1002491 261083 1002494
rect 502517 1002491 502583 1002494
rect 100293 1002418 100359 1002421
rect 108021 1002418 108087 1002421
rect 158621 1002418 158687 1002421
rect 100293 1002416 100556 1002418
rect 100293 1002360 100298 1002416
rect 100354 1002360 100556 1002416
rect 100293 1002358 100556 1002360
rect 107916 1002416 108087 1002418
rect 107916 1002360 108026 1002416
rect 108082 1002360 108087 1002416
rect 107916 1002358 108087 1002360
rect 158516 1002416 158687 1002418
rect 158516 1002360 158626 1002416
rect 158682 1002360 158687 1002416
rect 158516 1002358 158687 1002360
rect 100293 1002355 100359 1002358
rect 108021 1002355 108087 1002358
rect 158621 1002355 158687 1002358
rect 211245 1002418 211311 1002421
rect 256141 1002418 256207 1002421
rect 310145 1002418 310211 1002421
rect 211245 1002416 211508 1002418
rect 211245 1002360 211250 1002416
rect 211306 1002360 211508 1002416
rect 211245 1002358 211508 1002360
rect 256141 1002416 256404 1002418
rect 256141 1002360 256146 1002416
rect 256202 1002360 256404 1002416
rect 256141 1002358 256404 1002360
rect 309948 1002416 310211 1002418
rect 309948 1002360 310150 1002416
rect 310206 1002360 310211 1002416
rect 309948 1002358 310211 1002360
rect 211245 1002355 211311 1002358
rect 256141 1002355 256207 1002358
rect 310145 1002355 310211 1002358
rect 358537 1002418 358603 1002421
rect 557993 1002418 558059 1002421
rect 358537 1002416 358800 1002418
rect 358537 1002360 358542 1002416
rect 358598 1002360 358800 1002416
rect 358537 1002358 358800 1002360
rect 557993 1002416 558256 1002418
rect 557993 1002360 557998 1002416
rect 558054 1002360 558256 1002416
rect 557993 1002358 558256 1002360
rect 358537 1002355 358603 1002358
rect 557993 1002355 558059 1002358
rect 101121 1002282 101187 1002285
rect 105629 1002282 105695 1002285
rect 108481 1002282 108547 1002285
rect 101121 1002280 101292 1002282
rect 101121 1002224 101126 1002280
rect 101182 1002224 101292 1002280
rect 101121 1002222 101292 1002224
rect 105432 1002280 105695 1002282
rect 105432 1002224 105634 1002280
rect 105690 1002224 105695 1002280
rect 105432 1002222 105695 1002224
rect 108284 1002280 108547 1002282
rect 108284 1002224 108486 1002280
rect 108542 1002224 108547 1002280
rect 108284 1002222 108547 1002224
rect 101121 1002219 101187 1002222
rect 105629 1002219 105695 1002222
rect 108481 1002219 108547 1002222
rect 155769 1002282 155835 1002285
rect 156597 1002282 156663 1002285
rect 206369 1002282 206435 1002285
rect 254485 1002282 254551 1002285
rect 306097 1002282 306163 1002285
rect 359365 1002282 359431 1002285
rect 155769 1002280 156032 1002282
rect 155769 1002224 155774 1002280
rect 155830 1002224 156032 1002280
rect 155769 1002222 156032 1002224
rect 156597 1002280 156860 1002282
rect 156597 1002224 156602 1002280
rect 156658 1002224 156860 1002280
rect 156597 1002222 156860 1002224
rect 206369 1002280 206540 1002282
rect 206369 1002224 206374 1002280
rect 206430 1002224 206540 1002280
rect 206369 1002222 206540 1002224
rect 254485 1002280 254748 1002282
rect 254485 1002224 254490 1002280
rect 254546 1002224 254748 1002280
rect 254485 1002222 254748 1002224
rect 306097 1002280 306360 1002282
rect 306097 1002224 306102 1002280
rect 306158 1002224 306360 1002280
rect 306097 1002222 306360 1002224
rect 359168 1002280 359431 1002282
rect 359168 1002224 359370 1002280
rect 359426 1002224 359431 1002280
rect 359168 1002222 359431 1002224
rect 155769 1002219 155835 1002222
rect 156597 1002219 156663 1002222
rect 206369 1002219 206435 1002222
rect 254485 1002219 254551 1002222
rect 306097 1002219 306163 1002222
rect 359365 1002219 359431 1002222
rect 426341 1002282 426407 1002285
rect 503345 1002282 503411 1002285
rect 426341 1002280 426604 1002282
rect 426341 1002224 426346 1002280
rect 426402 1002224 426604 1002280
rect 426341 1002222 426604 1002224
rect 503148 1002280 503411 1002282
rect 503148 1002224 503350 1002280
rect 503406 1002224 503411 1002280
rect 503148 1002222 503411 1002224
rect 426341 1002219 426407 1002222
rect 503345 1002219 503411 1002222
rect 554313 1002282 554379 1002285
rect 560477 1002282 560543 1002285
rect 554313 1002280 554576 1002282
rect 554313 1002224 554318 1002280
rect 554374 1002224 554576 1002280
rect 554313 1002222 554576 1002224
rect 560280 1002280 560543 1002282
rect 560280 1002224 560482 1002280
rect 560538 1002224 560543 1002280
rect 560280 1002222 560543 1002224
rect 554313 1002219 554379 1002222
rect 560477 1002219 560543 1002222
rect 99097 1002146 99163 1002149
rect 103145 1002146 103211 1002149
rect 104801 1002146 104867 1002149
rect 99097 1002144 99268 1002146
rect 99097 1002088 99102 1002144
rect 99158 1002088 99268 1002144
rect 99097 1002086 99268 1002088
rect 103145 1002144 103408 1002146
rect 103145 1002088 103150 1002144
rect 103206 1002088 103408 1002144
rect 103145 1002086 103408 1002088
rect 104604 1002144 104867 1002146
rect 104604 1002088 104806 1002144
rect 104862 1002088 104867 1002144
rect 104604 1002086 104867 1002088
rect 99097 1002083 99163 1002086
rect 103145 1002083 103211 1002086
rect 104801 1002083 104867 1002086
rect 106825 1002146 106891 1002149
rect 109677 1002146 109743 1002149
rect 150893 1002146 150959 1002149
rect 106825 1002144 107088 1002146
rect 106825 1002088 106830 1002144
rect 106886 1002088 107088 1002144
rect 106825 1002086 107088 1002088
rect 109480 1002144 109743 1002146
rect 109480 1002088 109682 1002144
rect 109738 1002088 109743 1002144
rect 109480 1002086 109743 1002088
rect 150696 1002144 150959 1002146
rect 150696 1002088 150898 1002144
rect 150954 1002088 150959 1002144
rect 150696 1002086 150959 1002088
rect 106825 1002083 106891 1002086
rect 109677 1002083 109743 1002086
rect 150893 1002083 150959 1002086
rect 154573 1002146 154639 1002149
rect 154941 1002146 155007 1002149
rect 207197 1002146 207263 1002149
rect 211245 1002146 211311 1002149
rect 154573 1002144 154836 1002146
rect 154573 1002088 154578 1002144
rect 154634 1002088 154836 1002144
rect 154573 1002086 154836 1002088
rect 154941 1002144 155204 1002146
rect 154941 1002088 154946 1002144
rect 155002 1002088 155204 1002144
rect 154941 1002086 155204 1002088
rect 207197 1002144 207460 1002146
rect 207197 1002088 207202 1002144
rect 207258 1002088 207460 1002144
rect 207197 1002086 207460 1002088
rect 211140 1002144 211311 1002146
rect 211140 1002088 211250 1002144
rect 211306 1002088 211311 1002144
rect 211140 1002086 211311 1002088
rect 154573 1002083 154639 1002086
rect 154941 1002083 155007 1002086
rect 207197 1002083 207263 1002086
rect 211245 1002083 211311 1002086
rect 253289 1002146 253355 1002149
rect 256141 1002146 256207 1002149
rect 263501 1002146 263567 1002149
rect 253289 1002144 253460 1002146
rect 253289 1002088 253294 1002144
rect 253350 1002088 253460 1002144
rect 253289 1002086 253460 1002088
rect 255944 1002144 256207 1002146
rect 255944 1002088 256146 1002144
rect 256202 1002088 256207 1002144
rect 255944 1002086 256207 1002088
rect 263304 1002144 263567 1002146
rect 263304 1002088 263506 1002144
rect 263562 1002088 263567 1002144
rect 263304 1002086 263567 1002088
rect 253289 1002083 253355 1002086
rect 256141 1002083 256207 1002086
rect 263501 1002083 263567 1002086
rect 308949 1002146 309015 1002149
rect 310145 1002146 310211 1002149
rect 310605 1002146 310671 1002149
rect 310973 1002146 311039 1002149
rect 358537 1002146 358603 1002149
rect 308949 1002144 309212 1002146
rect 308949 1002088 308954 1002144
rect 309010 1002088 309212 1002144
rect 308949 1002086 309212 1002088
rect 310145 1002144 310408 1002146
rect 310145 1002088 310150 1002144
rect 310206 1002088 310408 1002144
rect 310145 1002086 310408 1002088
rect 310605 1002144 310868 1002146
rect 310605 1002088 310610 1002144
rect 310666 1002088 310868 1002144
rect 310605 1002086 310868 1002088
rect 310973 1002144 311236 1002146
rect 310973 1002088 310978 1002144
rect 311034 1002088 311236 1002144
rect 310973 1002086 311236 1002088
rect 358340 1002144 358603 1002146
rect 358340 1002088 358542 1002144
rect 358598 1002088 358603 1002144
rect 358340 1002086 358603 1002088
rect 308949 1002083 309015 1002086
rect 310145 1002083 310211 1002086
rect 310605 1002083 310671 1002086
rect 310973 1002083 311039 1002086
rect 358537 1002083 358603 1002086
rect 360561 1002146 360627 1002149
rect 433333 1002146 433399 1002149
rect 504173 1002146 504239 1002149
rect 509877 1002146 509943 1002149
rect 560017 1002146 560083 1002149
rect 360561 1002144 360824 1002146
rect 360561 1002088 360566 1002144
rect 360622 1002088 360824 1002144
rect 360561 1002086 360824 1002088
rect 433136 1002144 433399 1002146
rect 433136 1002088 433338 1002144
rect 433394 1002088 433399 1002144
rect 433136 1002086 433399 1002088
rect 503976 1002144 504239 1002146
rect 503976 1002088 504178 1002144
rect 504234 1002088 504239 1002144
rect 503976 1002086 504239 1002088
rect 509680 1002144 509943 1002146
rect 509680 1002088 509882 1002144
rect 509938 1002088 509943 1002144
rect 509680 1002086 509943 1002088
rect 559820 1002144 560083 1002146
rect 559820 1002088 560022 1002144
rect 560078 1002088 560083 1002144
rect 559820 1002086 560083 1002088
rect 360561 1002083 360627 1002086
rect 433333 1002083 433399 1002086
rect 504173 1002083 504239 1002086
rect 509877 1002083 509943 1002086
rect 560017 1002083 560083 1002086
rect 98269 1002010 98335 1002013
rect 98072 1002008 98335 1002010
rect 98072 1001952 98274 1002008
rect 98330 1001952 98335 1002008
rect 98072 1001950 98335 1001952
rect 98269 1001947 98335 1001950
rect 101949 1002010 102015 1002013
rect 103973 1002010 104039 1002013
rect 101949 1002008 102212 1002010
rect 101949 1001952 101954 1002008
rect 102010 1001952 102212 1002008
rect 101949 1001950 102212 1001952
rect 103776 1002008 104039 1002010
rect 103776 1001952 103978 1002008
rect 104034 1001952 104039 1002008
rect 103776 1001950 104039 1001952
rect 101949 1001947 102015 1001950
rect 103973 1001947 104039 1001950
rect 105997 1002010 106063 1002013
rect 108849 1002010 108915 1002013
rect 149237 1002010 149303 1002013
rect 153745 1002010 153811 1002013
rect 155769 1002010 155835 1002013
rect 156597 1002010 156663 1002013
rect 157793 1002010 157859 1002013
rect 105997 1002008 106260 1002010
rect 105997 1001952 106002 1002008
rect 106058 1001952 106260 1002008
rect 105997 1001950 106260 1001952
rect 108849 1002008 109112 1002010
rect 108849 1001952 108854 1002008
rect 108910 1001952 109112 1002008
rect 108849 1001950 109112 1001952
rect 149237 1002008 149500 1002010
rect 149237 1001952 149242 1002008
rect 149298 1001952 149500 1002008
rect 149237 1001950 149500 1001952
rect 153548 1002008 153811 1002010
rect 153548 1001952 153750 1002008
rect 153806 1001952 153811 1002008
rect 153548 1001950 153811 1001952
rect 155572 1002008 155835 1002010
rect 155572 1001952 155774 1002008
rect 155830 1001952 155835 1002008
rect 155572 1001950 155835 1001952
rect 156400 1002008 156663 1002010
rect 156400 1001952 156602 1002008
rect 156658 1001952 156663 1002008
rect 156400 1001950 156663 1001952
rect 157596 1002008 157859 1002010
rect 157596 1001952 157798 1002008
rect 157854 1001952 157859 1002008
rect 157596 1001950 157859 1001952
rect 105997 1001947 106063 1001950
rect 108849 1001947 108915 1001950
rect 149237 1001947 149303 1001950
rect 153745 1001947 153811 1001950
rect 155769 1001947 155835 1001950
rect 156597 1001947 156663 1001950
rect 157793 1001947 157859 1001950
rect 203885 1002010 203951 1002013
rect 205541 1002010 205607 1002013
rect 207565 1002010 207631 1002013
rect 208393 1002010 208459 1002013
rect 203885 1002008 204148 1002010
rect 203885 1001952 203890 1002008
rect 203946 1001952 204148 1002008
rect 203885 1001950 204148 1001952
rect 205541 1002008 205804 1002010
rect 205541 1001952 205546 1002008
rect 205602 1001952 205804 1002008
rect 205541 1001950 205804 1001952
rect 207565 1002008 207828 1002010
rect 207565 1001952 207570 1002008
rect 207626 1001952 207828 1002008
rect 207565 1001950 207828 1001952
rect 208196 1002008 208459 1002010
rect 208196 1001952 208398 1002008
rect 208454 1001952 208459 1002008
rect 208196 1001950 208459 1001952
rect 203885 1001947 203951 1001950
rect 205541 1001947 205607 1001950
rect 207565 1001947 207631 1001950
rect 208393 1001947 208459 1001950
rect 210417 1002010 210483 1002013
rect 212073 1002010 212139 1002013
rect 252461 1002010 252527 1002013
rect 210417 1002008 210680 1002010
rect 210417 1001952 210422 1002008
rect 210478 1001952 210680 1002008
rect 210417 1001950 210680 1001952
rect 211876 1002008 212139 1002010
rect 211876 1001952 212078 1002008
rect 212134 1001952 212139 1002008
rect 211876 1001950 212139 1001952
rect 252264 1002008 252527 1002010
rect 252264 1001952 252466 1002008
rect 252522 1001952 252527 1002008
rect 252264 1001950 252527 1001952
rect 210417 1001947 210483 1001950
rect 212073 1001947 212139 1001950
rect 252461 1001947 252527 1001950
rect 261017 1002010 261083 1002013
rect 263869 1002010 263935 1002013
rect 306097 1002010 306163 1002013
rect 309777 1002010 309843 1002013
rect 261017 1002008 261280 1002010
rect 261017 1001952 261022 1002008
rect 261078 1001952 261280 1002008
rect 261017 1001950 261280 1001952
rect 263764 1002008 263935 1002010
rect 263764 1001952 263874 1002008
rect 263930 1001952 263935 1002008
rect 263764 1001950 263935 1001952
rect 305900 1002008 306163 1002010
rect 305900 1001952 306102 1002008
rect 306158 1001952 306163 1002008
rect 305900 1001950 306163 1001952
rect 309580 1002008 309843 1002010
rect 309580 1001952 309782 1002008
rect 309838 1001952 309843 1002008
rect 309580 1001950 309843 1001952
rect 261017 1001947 261083 1001950
rect 263869 1001947 263935 1001950
rect 306097 1001947 306163 1001950
rect 309777 1001947 309843 1001950
rect 312629 1002010 312695 1002013
rect 354029 1002010 354095 1002013
rect 357341 1002010 357407 1002013
rect 360193 1002010 360259 1002013
rect 365897 1002010 365963 1002013
rect 312629 1002008 312892 1002010
rect 312629 1001952 312634 1002008
rect 312690 1001952 312892 1002008
rect 312629 1001950 312892 1001952
rect 354029 1002008 354292 1002010
rect 354029 1001952 354034 1002008
rect 354090 1001952 354292 1002008
rect 354029 1001950 354292 1001952
rect 357341 1002008 357604 1002010
rect 357341 1001952 357346 1002008
rect 357402 1001952 357604 1002008
rect 357341 1001950 357604 1001952
rect 359996 1002008 360259 1002010
rect 359996 1001952 360198 1002008
rect 360254 1001952 360259 1002008
rect 359996 1001950 360259 1001952
rect 365700 1002008 365963 1002010
rect 365700 1001952 365902 1002008
rect 365958 1001952 365963 1002008
rect 365700 1001950 365963 1001952
rect 312629 1001947 312695 1001950
rect 354029 1001947 354095 1001950
rect 357341 1001947 357407 1001950
rect 360193 1001947 360259 1001950
rect 365897 1001947 365963 1001950
rect 421465 1002010 421531 1002013
rect 426341 1002010 426407 1002013
rect 421465 1002008 421636 1002010
rect 421465 1001952 421470 1002008
rect 421526 1001952 421636 1002008
rect 421465 1001950 421636 1001952
rect 426144 1002008 426407 1002010
rect 426144 1001952 426346 1002008
rect 426402 1001952 426407 1002008
rect 426144 1001950 426407 1001952
rect 421465 1001947 421531 1001950
rect 426341 1001947 426407 1001950
rect 428365 1002010 428431 1002013
rect 498469 1002010 498535 1002013
rect 502517 1002010 502583 1002013
rect 503345 1002010 503411 1002013
rect 506197 1002010 506263 1002013
rect 507025 1002010 507091 1002013
rect 553945 1002010 554011 1002013
rect 558821 1002010 558887 1002013
rect 428365 1002008 428628 1002010
rect 428365 1001952 428370 1002008
rect 428426 1001952 428628 1002008
rect 428365 1001950 428628 1001952
rect 498469 1002008 498732 1002010
rect 498469 1001952 498474 1002008
rect 498530 1001952 498732 1002008
rect 498469 1001950 498732 1001952
rect 502517 1002008 502780 1002010
rect 502517 1001952 502522 1002008
rect 502578 1001952 502780 1002008
rect 502517 1001950 502780 1001952
rect 503345 1002008 503608 1002010
rect 503345 1001952 503350 1002008
rect 503406 1001952 503608 1002008
rect 503345 1001950 503608 1001952
rect 506197 1002008 506460 1002010
rect 506197 1001952 506202 1002008
rect 506258 1001952 506460 1002008
rect 506197 1001950 506460 1001952
rect 507025 1002008 507196 1002010
rect 507025 1001952 507030 1002008
rect 507086 1001952 507196 1002008
rect 507025 1001950 507196 1001952
rect 553748 1002008 554011 1002010
rect 553748 1001952 553950 1002008
rect 554006 1001952 554011 1002008
rect 553748 1001950 554011 1001952
rect 558624 1002008 558887 1002010
rect 558624 1001952 558826 1002008
rect 558882 1001952 558887 1002008
rect 558624 1001950 558887 1001952
rect 428365 1001947 428431 1001950
rect 498469 1001947 498535 1001950
rect 502517 1001947 502583 1001950
rect 503345 1001947 503411 1001950
rect 506197 1001947 506263 1001950
rect 507025 1001947 507091 1001950
rect 553945 1001947 554011 1001950
rect 558821 1001947 558887 1001950
rect 560845 1002010 560911 1002013
rect 560845 1002008 561108 1002010
rect 560845 1001952 560850 1002008
rect 560906 1001952 561108 1002008
rect 560845 1001950 561108 1001952
rect 560845 1001947 560911 1001950
rect 203517 999154 203583 999157
rect 203320 999152 203583 999154
rect 203320 999096 203522 999152
rect 203578 999096 203583 999152
rect 203320 999094 203583 999096
rect 203517 999091 203583 999094
rect 204345 998746 204411 998749
rect 204345 998744 204516 998746
rect 204345 998688 204350 998744
rect 204406 998688 204516 998744
rect 204345 998686 204516 998688
rect 204345 998683 204411 998686
rect 202689 998610 202755 998613
rect 202689 998608 202952 998610
rect 202689 998552 202694 998608
rect 202750 998552 202952 998608
rect 202689 998550 202952 998552
rect 202689 998547 202755 998550
rect 553117 998474 553183 998477
rect 552920 998472 553183 998474
rect 552920 998416 553122 998472
rect 553178 998416 553183 998472
rect 552920 998414 553183 998416
rect 553117 998411 553183 998414
rect 205541 998202 205607 998205
rect 258165 998202 258231 998205
rect 205344 998200 205607 998202
rect 205344 998144 205546 998200
rect 205602 998144 205607 998200
rect 205344 998142 205607 998144
rect 257968 998200 258231 998202
rect 257968 998144 258170 998200
rect 258226 998144 258231 998200
rect 257968 998142 258231 998144
rect 205541 998139 205607 998142
rect 258165 998139 258231 998142
rect 202689 998066 202755 998069
rect 202492 998064 202755 998066
rect 202492 998008 202694 998064
rect 202750 998008 202755 998064
rect 202492 998006 202755 998008
rect 202689 998003 202755 998006
rect 257337 998066 257403 998069
rect 260189 998066 260255 998069
rect 257337 998064 257600 998066
rect 257337 998008 257342 998064
rect 257398 998008 257600 998064
rect 257337 998006 257600 998008
rect 260084 998064 260255 998066
rect 260084 998008 260194 998064
rect 260250 998008 260255 998064
rect 260084 998006 260255 998008
rect 257337 998003 257403 998006
rect 260189 998003 260255 998006
rect 200665 997930 200731 997933
rect 203517 997930 203583 997933
rect 256969 997930 257035 997933
rect 258165 997930 258231 997933
rect 259821 997930 259887 997933
rect 200665 997928 200836 997930
rect 200665 997872 200670 997928
rect 200726 997872 200836 997928
rect 200665 997870 200836 997872
rect 203517 997928 203780 997930
rect 203517 997872 203522 997928
rect 203578 997872 203780 997928
rect 203517 997870 203780 997872
rect 256969 997928 257140 997930
rect 256969 997872 256974 997928
rect 257030 997872 257140 997928
rect 256969 997870 257140 997872
rect 258165 997928 258428 997930
rect 258165 997872 258170 997928
rect 258226 997872 258428 997928
rect 258165 997870 258428 997872
rect 259624 997928 259887 997930
rect 259624 997872 259826 997928
rect 259882 997872 259887 997928
rect 259624 997870 259887 997872
rect 200665 997867 200731 997870
rect 203517 997867 203583 997870
rect 256969 997867 257035 997870
rect 258165 997867 258231 997870
rect 259821 997867 259887 997870
rect 551093 997930 551159 997933
rect 551093 997928 551356 997930
rect 551093 997872 551098 997928
rect 551154 997872 551356 997928
rect 551093 997870 551356 997872
rect 551093 997867 551159 997870
rect 201861 997794 201927 997797
rect 204713 997794 204779 997797
rect 256509 997794 256575 997797
rect 258993 997794 259059 997797
rect 260189 997794 260255 997797
rect 261845 997794 261911 997797
rect 298277 997794 298343 997797
rect 303245 997794 303311 997797
rect 550265 997794 550331 997797
rect 201861 997792 202124 997794
rect 201861 997736 201866 997792
rect 201922 997736 202124 997792
rect 201861 997734 202124 997736
rect 204713 997792 204976 997794
rect 204713 997736 204718 997792
rect 204774 997736 204976 997792
rect 204713 997734 204976 997736
rect 256509 997792 256772 997794
rect 256509 997736 256514 997792
rect 256570 997736 256772 997792
rect 256509 997734 256772 997736
rect 258993 997792 259164 997794
rect 258993 997736 258998 997792
rect 259054 997736 259164 997792
rect 258993 997734 259164 997736
rect 260189 997792 260452 997794
rect 260189 997736 260194 997792
rect 260250 997736 260452 997792
rect 260189 997734 260452 997736
rect 261845 997792 262108 997794
rect 261845 997736 261850 997792
rect 261906 997736 262108 997792
rect 261845 997734 262108 997736
rect 298277 997792 303311 997794
rect 298277 997736 298282 997792
rect 298338 997736 303250 997792
rect 303306 997736 303311 997792
rect 298277 997734 303311 997736
rect 550068 997792 550331 997794
rect 550068 997736 550270 997792
rect 550326 997736 550331 997792
rect 550068 997734 550331 997736
rect 201861 997731 201927 997734
rect 204713 997731 204779 997734
rect 256509 997731 256575 997734
rect 258993 997731 259059 997734
rect 260189 997731 260255 997734
rect 261845 997731 261911 997734
rect 298277 997731 298343 997734
rect 303245 997731 303311 997734
rect 550265 997731 550331 997734
rect 552289 997794 552355 997797
rect 552289 997792 552552 997794
rect 552289 997736 552294 997792
rect 552350 997736 552552 997792
rect 552289 997734 552552 997736
rect 552289 997731 552355 997734
rect 195145 997660 195211 997661
rect 195094 997596 195100 997660
rect 195164 997658 195211 997660
rect 195164 997656 195256 997658
rect 195206 997600 195256 997656
rect 195164 997598 195256 997600
rect 195164 997596 195211 997598
rect 195145 997595 195211 997596
rect 87822 997188 87828 997252
rect 87892 997250 87898 997252
rect 92657 997250 92723 997253
rect 87892 997248 92723 997250
rect 87892 997192 92662 997248
rect 92718 997192 92723 997248
rect 87892 997190 92723 997192
rect 87892 997188 87898 997190
rect 92657 997187 92723 997190
rect 180558 997188 180564 997252
rect 180628 997250 180634 997252
rect 183870 997250 183876 997252
rect 180628 997190 183876 997250
rect 180628 997188 180634 997190
rect 183870 997188 183876 997190
rect 183940 997188 183946 997252
rect 200205 997250 200271 997253
rect 190410 997248 200271 997250
rect 190410 997192 200210 997248
rect 200266 997192 200271 997248
rect 190410 997190 200271 997192
rect 145741 996978 145807 996981
rect 133646 996976 145807 996978
rect 133646 996920 145746 996976
rect 145802 996920 145807 996976
rect 133646 996918 145807 996920
rect 82310 996374 85682 996434
rect 82310 995757 82370 996374
rect 85622 996298 85682 996374
rect 85622 996238 93870 996298
rect 93810 996026 93870 996238
rect 97441 996026 97507 996029
rect 93810 996024 97507 996026
rect 93810 995968 97446 996024
rect 97502 995968 97507 996024
rect 93810 995966 97507 995968
rect 97441 995963 97507 995966
rect 93669 995890 93735 995893
rect 82261 995752 82370 995757
rect 82261 995696 82266 995752
rect 82322 995696 82370 995752
rect 82261 995694 82370 995696
rect 82494 995888 93735 995890
rect 82494 995832 93674 995888
rect 93730 995832 93735 995888
rect 82494 995830 93735 995832
rect 82261 995691 82327 995694
rect 81065 995482 81131 995485
rect 82494 995482 82554 995830
rect 93669 995827 93735 995830
rect 133646 995757 133706 996918
rect 145741 996915 145807 996918
rect 144361 996706 144427 996709
rect 139166 996704 144427 996706
rect 139166 996648 144366 996704
rect 144422 996648 144427 996704
rect 139166 996646 144427 996648
rect 139166 995757 139226 996646
rect 144361 996643 144427 996646
rect 144821 996434 144887 996437
rect 190410 996434 190470 997190
rect 200205 997187 200271 997190
rect 292798 996780 292804 996844
rect 292868 996842 292874 996844
rect 299013 996842 299079 996845
rect 292868 996840 299079 996842
rect 292868 996784 299018 996840
rect 299074 996784 299079 996840
rect 292868 996782 299079 996784
rect 292868 996780 292874 996782
rect 299013 996779 299079 996782
rect 516869 996842 516935 996845
rect 527950 996842 527956 996844
rect 516869 996840 527956 996842
rect 516869 996784 516874 996840
rect 516930 996784 527956 996840
rect 516869 996782 527956 996784
rect 516869 996779 516935 996782
rect 527950 996780 527956 996782
rect 528020 996780 528026 996844
rect 247861 996706 247927 996709
rect 240918 996704 247927 996706
rect 240918 996648 247866 996704
rect 247922 996648 247927 996704
rect 240918 996646 247927 996648
rect 141006 996432 144887 996434
rect 141006 996376 144826 996432
rect 144882 996376 144887 996432
rect 141006 996374 144887 996376
rect 141006 995757 141066 996374
rect 144821 996371 144887 996374
rect 187558 996374 190470 996434
rect 187558 995757 187618 996374
rect 192518 996372 192524 996436
rect 192588 996434 192594 996436
rect 199837 996434 199903 996437
rect 192588 996432 199903 996434
rect 192588 996376 199842 996432
rect 199898 996376 199903 996432
rect 192588 996374 199903 996376
rect 192588 996372 192594 996374
rect 199837 996371 199903 996374
rect 133597 995752 133706 995757
rect 133597 995696 133602 995752
rect 133658 995696 133706 995752
rect 133597 995694 133706 995696
rect 139117 995752 139226 995757
rect 139117 995696 139122 995752
rect 139178 995696 139226 995752
rect 139117 995694 139226 995696
rect 140957 995752 141066 995757
rect 140957 995696 140962 995752
rect 141018 995696 141066 995752
rect 140957 995694 141066 995696
rect 142889 995754 142955 995757
rect 151261 995754 151327 995757
rect 142889 995752 151327 995754
rect 142889 995696 142894 995752
rect 142950 995696 151266 995752
rect 151322 995696 151327 995752
rect 142889 995694 151327 995696
rect 133597 995691 133663 995694
rect 139117 995691 139183 995694
rect 140957 995691 141023 995694
rect 142889 995691 142955 995694
rect 151261 995691 151327 995694
rect 183870 995692 183876 995756
rect 183940 995754 183946 995756
rect 184473 995754 184539 995757
rect 183940 995752 184539 995754
rect 183940 995696 184478 995752
rect 184534 995696 184539 995752
rect 183940 995694 184539 995696
rect 183940 995692 183946 995694
rect 184473 995691 184539 995694
rect 187509 995752 187618 995757
rect 189533 995756 189599 995757
rect 189533 995754 189580 995756
rect 187509 995696 187514 995752
rect 187570 995696 187618 995752
rect 187509 995694 187618 995696
rect 189488 995752 189580 995754
rect 189488 995696 189538 995752
rect 189488 995694 189580 995696
rect 187509 995691 187575 995694
rect 189533 995692 189580 995694
rect 189644 995692 189650 995756
rect 190453 995754 190519 995757
rect 195329 995754 195395 995757
rect 190453 995752 195395 995754
rect 190453 995696 190458 995752
rect 190514 995696 195334 995752
rect 195390 995696 195395 995752
rect 190453 995694 195395 995696
rect 189533 995691 189599 995692
rect 190453 995691 190519 995694
rect 195329 995691 195395 995694
rect 81065 995480 82554 995482
rect 81065 995424 81070 995480
rect 81126 995424 82554 995480
rect 81065 995422 82554 995424
rect 86585 995482 86651 995485
rect 93117 995482 93183 995485
rect 86585 995480 93183 995482
rect 86585 995424 86590 995480
rect 86646 995424 93122 995480
rect 93178 995424 93183 995480
rect 86585 995422 93183 995424
rect 81065 995419 81131 995422
rect 86585 995419 86651 995422
rect 93117 995419 93183 995422
rect 183829 995482 183895 995485
rect 192477 995484 192543 995485
rect 186262 995482 186268 995484
rect 183829 995480 186268 995482
rect 183829 995424 183834 995480
rect 183890 995424 186268 995480
rect 183829 995422 186268 995424
rect 183829 995419 183895 995422
rect 186262 995420 186268 995422
rect 186332 995420 186338 995484
rect 192477 995482 192524 995484
rect 192432 995480 192524 995482
rect 192432 995424 192482 995480
rect 192432 995422 192524 995424
rect 192477 995420 192524 995422
rect 192588 995420 192594 995484
rect 194542 995420 194548 995484
rect 194612 995482 194618 995484
rect 202321 995482 202387 995485
rect 194612 995480 202387 995482
rect 194612 995424 202326 995480
rect 202382 995424 202387 995480
rect 194612 995422 202387 995424
rect 194612 995420 194618 995422
rect 192477 995419 192543 995420
rect 202321 995419 202387 995422
rect 100201 995346 100267 995349
rect 93534 995344 100267 995346
rect 93534 995288 100206 995344
rect 100262 995288 100267 995344
rect 93534 995286 100267 995288
rect 84469 995210 84535 995213
rect 93534 995210 93594 995286
rect 100201 995283 100267 995286
rect 141785 995346 141851 995349
rect 146753 995346 146819 995349
rect 141785 995344 146819 995346
rect 141785 995288 141790 995344
rect 141846 995288 146758 995344
rect 146814 995288 146819 995344
rect 141785 995286 146819 995288
rect 141785 995283 141851 995286
rect 146753 995283 146819 995286
rect 84469 995208 93594 995210
rect 84469 995152 84474 995208
rect 84530 995152 93594 995208
rect 84469 995150 93594 995152
rect 84469 995147 84535 995150
rect 93669 995074 93735 995077
rect 100017 995074 100083 995077
rect 93669 995072 100083 995074
rect 93669 995016 93674 995072
rect 93730 995016 100022 995072
rect 100078 995016 100083 995072
rect 93669 995014 100083 995016
rect 87781 995012 87847 995013
rect 87781 995010 87828 995012
rect 87736 995008 87828 995010
rect 87736 994952 87786 995008
rect 87736 994950 87828 994952
rect 87781 994948 87828 994950
rect 87892 994948 87898 995012
rect 93669 995011 93735 995014
rect 100017 995011 100083 995014
rect 137093 995074 137159 995077
rect 148317 995074 148383 995077
rect 137093 995072 148383 995074
rect 137093 995016 137098 995072
rect 137154 995016 148322 995072
rect 148378 995016 148383 995072
rect 137093 995014 148383 995016
rect 137093 995011 137159 995014
rect 148317 995011 148383 995014
rect 177297 995074 177363 995077
rect 209822 995074 209882 996132
rect 240918 995757 240978 996646
rect 247861 996643 247927 996646
rect 372337 996706 372403 996709
rect 439681 996706 439747 996709
rect 474038 996706 474044 996708
rect 372337 996704 388178 996706
rect 372337 996648 372342 996704
rect 372398 996648 388178 996704
rect 372337 996646 388178 996648
rect 372337 996643 372403 996646
rect 246665 996434 246731 996437
rect 240869 995752 240978 995757
rect 240869 995696 240874 995752
rect 240930 995696 240978 995752
rect 240869 995694 240978 995696
rect 245518 996432 246731 996434
rect 245518 996376 246670 996432
rect 246726 996376 246731 996432
rect 245518 996374 246731 996376
rect 245518 995757 245578 996374
rect 246665 996371 246731 996374
rect 293534 996372 293540 996436
rect 293604 996434 293610 996436
rect 300853 996434 300919 996437
rect 293604 996432 300919 996434
rect 293604 996376 300858 996432
rect 300914 996376 300919 996432
rect 293604 996374 300919 996376
rect 293604 996372 293610 996374
rect 300853 996371 300919 996374
rect 372521 996434 372587 996437
rect 372521 996432 387994 996434
rect 372521 996376 372526 996432
rect 372582 996376 387994 996432
rect 372521 996374 387994 996376
rect 372521 996371 372587 996374
rect 245518 995752 245627 995757
rect 245518 995696 245566 995752
rect 245622 995696 245627 995752
rect 245518 995694 245627 995696
rect 240869 995691 240935 995694
rect 245561 995691 245627 995694
rect 243905 995482 243971 995485
rect 258766 995482 258826 996132
rect 300301 996026 300367 996029
rect 292530 996024 300367 996026
rect 292530 995968 300306 996024
rect 300362 995968 300367 996024
rect 292530 995966 300367 995968
rect 291745 995754 291811 995757
rect 292530 995754 292590 995966
rect 300301 995963 300367 995966
rect 387934 995757 387994 996374
rect 293493 995756 293559 995757
rect 293493 995754 293540 995756
rect 291745 995752 292590 995754
rect 291745 995696 291750 995752
rect 291806 995696 292590 995752
rect 291745 995694 292590 995696
rect 293448 995752 293540 995754
rect 293448 995696 293498 995752
rect 293448 995694 293540 995696
rect 291745 995691 291811 995694
rect 293493 995692 293540 995694
rect 293604 995692 293610 995756
rect 297265 995754 297331 995757
rect 298277 995754 298343 995757
rect 297265 995752 298343 995754
rect 297265 995696 297270 995752
rect 297326 995696 298282 995752
rect 298338 995696 298343 995752
rect 297265 995694 298343 995696
rect 293493 995691 293559 995692
rect 297265 995691 297331 995694
rect 298277 995691 298343 995694
rect 298502 995692 298508 995756
rect 298572 995754 298578 995756
rect 300117 995754 300183 995757
rect 298572 995752 300183 995754
rect 298572 995696 300122 995752
rect 300178 995696 300183 995752
rect 298572 995694 300183 995696
rect 298572 995692 298578 995694
rect 300117 995691 300183 995694
rect 383101 995754 383167 995757
rect 385677 995754 385743 995757
rect 383101 995752 385743 995754
rect 383101 995696 383106 995752
rect 383162 995696 385682 995752
rect 385738 995696 385743 995752
rect 383101 995694 385743 995696
rect 383101 995691 383167 995694
rect 385677 995691 385743 995694
rect 387885 995752 387994 995757
rect 387885 995696 387890 995752
rect 387946 995696 387994 995752
rect 387885 995694 387994 995696
rect 388118 995757 388178 996646
rect 439681 996704 474044 996706
rect 439681 996648 439686 996704
rect 439742 996648 474044 996704
rect 439681 996646 474044 996648
rect 439681 996643 439747 996646
rect 474038 996644 474044 996646
rect 474108 996644 474114 996708
rect 590561 996706 590627 996709
rect 627862 996706 627868 996708
rect 590561 996704 627868 996706
rect 590561 996648 590566 996704
rect 590622 996648 627868 996704
rect 590561 996646 627868 996648
rect 590561 996643 590627 996646
rect 627862 996644 627868 996646
rect 627932 996644 627938 996708
rect 528318 996570 528324 996572
rect 518942 996510 528324 996570
rect 421005 996434 421071 996437
rect 396582 996432 421071 996434
rect 396582 996376 421010 996432
rect 421066 996376 421071 996432
rect 396582 996374 421071 996376
rect 396582 995757 396642 996374
rect 421005 996371 421071 996374
rect 439865 996434 439931 996437
rect 474774 996434 474780 996436
rect 439865 996432 474780 996434
rect 439865 996376 439870 996432
rect 439926 996376 474780 996432
rect 439865 996374 474780 996376
rect 439865 996371 439931 996374
rect 474774 996372 474780 996374
rect 474844 996372 474850 996436
rect 516685 996434 516751 996437
rect 518942 996434 519002 996510
rect 528318 996508 528324 996510
rect 528388 996508 528394 996572
rect 590561 996434 590627 996437
rect 475886 996374 478338 996434
rect 456793 996162 456859 996165
rect 475886 996162 475946 996374
rect 456793 996160 475946 996162
rect 456793 996104 456798 996160
rect 456854 996104 475946 996160
rect 456793 996102 475946 996104
rect 456793 996099 456859 996102
rect 478278 995757 478338 996374
rect 516685 996432 519002 996434
rect 516685 996376 516690 996432
rect 516746 996376 519002 996432
rect 516685 996374 519002 996376
rect 528510 996374 532802 996434
rect 516685 996371 516751 996374
rect 519537 996298 519603 996301
rect 528510 996298 528570 996374
rect 519537 996296 528570 996298
rect 519537 996240 519542 996296
rect 519598 996240 528570 996296
rect 519537 996238 528570 996240
rect 519537 996235 519603 996238
rect 506422 995828 506428 995892
rect 506492 995890 506498 995892
rect 511073 995890 511139 995893
rect 506492 995888 511139 995890
rect 506492 995832 511078 995888
rect 511134 995832 511139 995888
rect 506492 995830 511139 995832
rect 506492 995828 506498 995830
rect 511073 995827 511139 995830
rect 532742 995757 532802 996374
rect 590561 996432 629770 996434
rect 590561 996376 590566 996432
rect 590622 996376 629770 996432
rect 590561 996374 629770 996376
rect 590561 996371 590627 996374
rect 625245 996026 625311 996029
rect 625245 996024 625354 996026
rect 625245 995968 625250 996024
rect 625306 995968 625354 996024
rect 625245 995963 625354 995968
rect 388118 995752 388227 995757
rect 388118 995696 388166 995752
rect 388222 995696 388227 995752
rect 388118 995694 388227 995696
rect 387885 995691 387951 995694
rect 388161 995691 388227 995694
rect 396533 995752 396642 995757
rect 396533 995696 396538 995752
rect 396594 995696 396642 995752
rect 396533 995694 396642 995696
rect 472617 995754 472683 995757
rect 477033 995754 477099 995757
rect 472617 995752 477099 995754
rect 472617 995696 472622 995752
rect 472678 995696 477038 995752
rect 477094 995696 477099 995752
rect 472617 995694 477099 995696
rect 478278 995752 478387 995757
rect 485589 995756 485655 995757
rect 485589 995754 485636 995756
rect 478278 995696 478326 995752
rect 478382 995696 478387 995752
rect 478278 995694 478387 995696
rect 485544 995752 485636 995754
rect 485544 995696 485594 995752
rect 485544 995694 485636 995696
rect 396533 995691 396599 995694
rect 472617 995691 472683 995694
rect 477033 995691 477099 995694
rect 478321 995691 478387 995694
rect 485589 995692 485636 995694
rect 485700 995692 485706 995756
rect 520181 995754 520247 995757
rect 526069 995754 526135 995757
rect 528001 995756 528067 995757
rect 520181 995752 526135 995754
rect 520181 995696 520186 995752
rect 520242 995696 526074 995752
rect 526130 995696 526135 995752
rect 520181 995694 526135 995696
rect 485589 995691 485655 995692
rect 520181 995691 520247 995694
rect 526069 995691 526135 995694
rect 527950 995692 527956 995756
rect 528020 995754 528067 995756
rect 528020 995752 528112 995754
rect 528062 995696 528112 995752
rect 528020 995694 528112 995696
rect 528020 995692 528067 995694
rect 528318 995692 528324 995756
rect 528388 995754 528394 995756
rect 528553 995754 528619 995757
rect 528388 995752 528619 995754
rect 528388 995696 528558 995752
rect 528614 995696 528619 995752
rect 528388 995694 528619 995696
rect 532742 995752 532851 995757
rect 536557 995756 536623 995757
rect 536557 995754 536604 995756
rect 532742 995696 532790 995752
rect 532846 995696 532851 995752
rect 532742 995694 532851 995696
rect 536512 995752 536604 995754
rect 536512 995696 536562 995752
rect 536512 995694 536604 995696
rect 528388 995692 528394 995694
rect 528001 995691 528067 995692
rect 528553 995691 528619 995694
rect 532785 995691 532851 995694
rect 536557 995692 536604 995694
rect 536668 995692 536674 995756
rect 536557 995691 536623 995692
rect 556102 995556 556108 995620
rect 556172 995618 556178 995620
rect 563697 995618 563763 995621
rect 556172 995616 563763 995618
rect 556172 995560 563702 995616
rect 563758 995560 563763 995616
rect 556172 995558 563763 995560
rect 556172 995556 556178 995558
rect 563697 995555 563763 995558
rect 243905 995480 258826 995482
rect 243905 995424 243910 995480
rect 243966 995424 258826 995480
rect 243905 995422 258826 995424
rect 286685 995484 286751 995485
rect 286685 995480 286732 995484
rect 286796 995482 286802 995484
rect 292481 995482 292547 995485
rect 292798 995482 292804 995484
rect 286685 995424 286690 995480
rect 243905 995419 243971 995422
rect 286685 995420 286732 995424
rect 286796 995422 286842 995482
rect 292481 995480 292804 995482
rect 292481 995424 292486 995480
rect 292542 995424 292804 995480
rect 292481 995422 292804 995424
rect 286796 995420 286802 995422
rect 286685 995419 286751 995420
rect 292481 995419 292547 995422
rect 292798 995420 292804 995422
rect 292868 995420 292874 995484
rect 296161 995482 296227 995485
rect 301497 995482 301563 995485
rect 474089 995484 474155 995485
rect 296161 995480 301563 995482
rect 296161 995424 296166 995480
rect 296222 995424 301502 995480
rect 301558 995424 301563 995480
rect 296161 995422 301563 995424
rect 296161 995419 296227 995422
rect 301497 995419 301563 995422
rect 474038 995420 474044 995484
rect 474108 995482 474155 995484
rect 474733 995484 474799 995485
rect 474733 995482 474780 995484
rect 474108 995480 474200 995482
rect 474150 995424 474200 995480
rect 474108 995422 474200 995424
rect 474688 995480 474780 995482
rect 474688 995424 474738 995480
rect 474688 995422 474780 995424
rect 474108 995420 474155 995422
rect 474089 995419 474155 995420
rect 474733 995420 474780 995422
rect 474844 995420 474850 995484
rect 480110 995420 480116 995484
rect 480180 995482 480186 995484
rect 480805 995482 480871 995485
rect 480180 995480 480871 995482
rect 480180 995424 480810 995480
rect 480866 995424 480871 995480
rect 480180 995422 480871 995424
rect 625294 995482 625354 995963
rect 629710 995757 629770 996374
rect 625613 995754 625679 995757
rect 627177 995754 627243 995757
rect 627913 995756 627979 995757
rect 625613 995752 627243 995754
rect 625613 995696 625618 995752
rect 625674 995696 627182 995752
rect 627238 995696 627243 995752
rect 625613 995694 627243 995696
rect 625613 995691 625679 995694
rect 627177 995691 627243 995694
rect 627862 995692 627868 995756
rect 627932 995754 627979 995756
rect 627932 995752 628024 995754
rect 627974 995696 628024 995752
rect 627932 995694 628024 995696
rect 629710 995752 629819 995757
rect 629710 995696 629758 995752
rect 629814 995696 629819 995752
rect 629710 995694 629819 995696
rect 627932 995692 627979 995694
rect 627913 995691 627979 995692
rect 629753 995691 629819 995694
rect 630305 995482 630371 995485
rect 625294 995480 630371 995482
rect 625294 995424 630310 995480
rect 630366 995424 630371 995480
rect 625294 995422 630371 995424
rect 480180 995420 480186 995422
rect 474733 995419 474799 995420
rect 480805 995419 480871 995422
rect 630305 995419 630371 995422
rect 381537 995346 381603 995349
rect 389357 995346 389423 995349
rect 381537 995344 389423 995346
rect 381537 995288 381542 995344
rect 381598 995288 389362 995344
rect 389418 995288 389423 995344
rect 381537 995286 389423 995288
rect 381537 995283 381603 995286
rect 389357 995283 389423 995286
rect 242939 995212 243005 995213
rect 242934 995210 242940 995212
rect 242848 995150 242940 995210
rect 242934 995148 242940 995150
rect 243004 995148 243010 995212
rect 244227 995210 244293 995213
rect 249333 995210 249399 995213
rect 393313 995210 393379 995213
rect 244227 995208 249399 995210
rect 244227 995152 244232 995208
rect 244288 995152 249338 995208
rect 249394 995152 249399 995208
rect 244227 995150 249399 995152
rect 242939 995147 243005 995148
rect 244227 995147 244293 995150
rect 249333 995147 249399 995150
rect 393270 995208 393379 995210
rect 393270 995152 393318 995208
rect 393374 995152 393379 995208
rect 393270 995147 393379 995152
rect 625613 995210 625679 995213
rect 634721 995210 634787 995213
rect 625613 995208 634787 995210
rect 625613 995152 625618 995208
rect 625674 995152 634726 995208
rect 634782 995152 634787 995208
rect 625613 995150 634787 995152
rect 625613 995147 625679 995150
rect 634721 995147 634787 995150
rect 393270 995077 393330 995147
rect 177297 995072 209882 995074
rect 177297 995016 177302 995072
rect 177358 995016 209882 995072
rect 177297 995014 209882 995016
rect 296437 995074 296503 995077
rect 298829 995074 298895 995077
rect 296437 995072 298895 995074
rect 296437 995016 296442 995072
rect 296498 995016 298834 995072
rect 298890 995016 298895 995072
rect 296437 995014 298895 995016
rect 177297 995011 177363 995014
rect 296437 995011 296503 995014
rect 298829 995011 298895 995014
rect 373257 995074 373323 995077
rect 392117 995074 392183 995077
rect 373257 995072 392183 995074
rect 373257 995016 373262 995072
rect 373318 995016 392122 995072
rect 392178 995016 392183 995072
rect 373257 995014 392183 995016
rect 373257 995011 373323 995014
rect 392117 995011 392183 995014
rect 393221 995072 393330 995077
rect 393221 995016 393226 995072
rect 393282 995016 393330 995072
rect 393221 995014 393330 995016
rect 451733 995074 451799 995077
rect 476757 995074 476823 995077
rect 451733 995072 476823 995074
rect 451733 995016 451738 995072
rect 451794 995016 476762 995072
rect 476818 995016 476823 995072
rect 451733 995014 476823 995016
rect 393221 995011 393287 995014
rect 451733 995011 451799 995014
rect 476757 995011 476823 995014
rect 517053 995074 517119 995077
rect 532509 995074 532575 995077
rect 517053 995072 532575 995074
rect 517053 995016 517058 995072
rect 517114 995016 532514 995072
rect 532570 995016 532575 995072
rect 517053 995014 532575 995016
rect 517053 995011 517119 995014
rect 532509 995011 532575 995014
rect 87781 994947 87847 994948
rect 239581 994938 239647 994941
rect 247677 994938 247743 994941
rect 239581 994936 247743 994938
rect 239581 994880 239586 994936
rect 239642 994880 247682 994936
rect 247738 994880 247743 994936
rect 239581 994878 247743 994880
rect 239581 994875 239647 994878
rect 247677 994875 247743 994878
rect 638861 994938 638927 994941
rect 640793 994938 640859 994941
rect 638861 994936 640859 994938
rect 638861 994880 638866 994936
rect 638922 994880 640798 994936
rect 640854 994880 640859 994936
rect 638861 994878 640859 994880
rect 638861 994875 638927 994878
rect 640793 994875 640859 994878
rect 80145 994802 80211 994805
rect 103513 994802 103579 994805
rect 80145 994800 103579 994802
rect 80145 994744 80150 994800
rect 80206 994744 103518 994800
rect 103574 994744 103579 994800
rect 80145 994742 103579 994744
rect 80145 994739 80211 994742
rect 103513 994739 103579 994742
rect 131573 994802 131639 994805
rect 157333 994802 157399 994805
rect 131573 994800 157399 994802
rect 131573 994744 131578 994800
rect 131634 994744 157338 994800
rect 157394 994744 157399 994800
rect 131573 994742 157399 994744
rect 131573 994739 131639 994742
rect 157333 994739 157399 994742
rect 184473 994802 184539 994805
rect 192937 994802 193003 994805
rect 184473 994800 193003 994802
rect 184473 994744 184478 994800
rect 184534 994744 192942 994800
rect 192998 994744 193003 994800
rect 184473 994742 193003 994744
rect 184473 994739 184539 994742
rect 192937 994739 193003 994742
rect 193121 994802 193187 994805
rect 197997 994802 198063 994805
rect 193121 994800 198063 994802
rect 193121 994744 193126 994800
rect 193182 994744 198002 994800
rect 198058 994744 198063 994800
rect 193121 994742 198063 994744
rect 193121 994739 193187 994742
rect 197997 994739 198063 994742
rect 290825 994802 290891 994805
rect 297909 994802 297975 994805
rect 290825 994800 297975 994802
rect 290825 994744 290830 994800
rect 290886 994744 297914 994800
rect 297970 994744 297975 994800
rect 290825 994742 297975 994744
rect 290825 994739 290891 994742
rect 297909 994739 297975 994742
rect 376293 994802 376359 994805
rect 395153 994802 395219 994805
rect 376293 994800 395219 994802
rect 376293 994744 376298 994800
rect 376354 994744 395158 994800
rect 395214 994744 395219 994800
rect 376293 994742 395219 994744
rect 376293 994739 376359 994742
rect 395153 994739 395219 994742
rect 445753 994802 445819 994805
rect 482277 994802 482343 994805
rect 445753 994800 482343 994802
rect 445753 994744 445758 994800
rect 445814 994744 482282 994800
rect 482338 994744 482343 994800
rect 445753 994742 482343 994744
rect 445753 994739 445819 994742
rect 482277 994739 482343 994742
rect 570229 994802 570295 994805
rect 637021 994802 637087 994805
rect 570229 994800 637087 994802
rect 570229 994744 570234 994800
rect 570290 994744 637026 994800
rect 637082 994744 637087 994800
rect 570229 994742 637087 994744
rect 570229 994739 570295 994742
rect 637021 994739 637087 994742
rect 85665 994530 85731 994533
rect 94681 994530 94747 994533
rect 85665 994528 94747 994530
rect 85665 994472 85670 994528
rect 85726 994472 94686 994528
rect 94742 994472 94747 994528
rect 85665 994470 94747 994472
rect 85665 994467 85731 994470
rect 94681 994467 94747 994470
rect 132769 994530 132835 994533
rect 149697 994530 149763 994533
rect 180609 994532 180675 994533
rect 132769 994528 149763 994530
rect 132769 994472 132774 994528
rect 132830 994472 149702 994528
rect 149758 994472 149763 994528
rect 132769 994470 149763 994472
rect 132769 994467 132835 994470
rect 149697 994467 149763 994470
rect 180558 994468 180564 994532
rect 180628 994530 180675 994532
rect 188797 994530 188863 994533
rect 200757 994530 200823 994533
rect 180628 994528 180720 994530
rect 180670 994472 180720 994528
rect 180628 994470 180720 994472
rect 188797 994528 200823 994530
rect 188797 994472 188802 994528
rect 188858 994472 200762 994528
rect 200818 994472 200823 994528
rect 188797 994470 200823 994472
rect 180628 994468 180675 994470
rect 180609 994467 180675 994468
rect 188797 994467 188863 994470
rect 200757 994467 200823 994470
rect 238661 994530 238727 994533
rect 254577 994530 254643 994533
rect 238661 994528 254643 994530
rect 238661 994472 238666 994528
rect 238722 994472 254582 994528
rect 254638 994472 254643 994528
rect 238661 994470 254643 994472
rect 238661 994467 238727 994470
rect 254577 994467 254643 994470
rect 287789 994530 287855 994533
rect 301037 994530 301103 994533
rect 287789 994528 301103 994530
rect 287789 994472 287794 994528
rect 287850 994472 301042 994528
rect 301098 994472 301103 994528
rect 287789 994470 301103 994472
rect 287789 994467 287855 994470
rect 301037 994467 301103 994470
rect 381261 994530 381327 994533
rect 392301 994530 392367 994533
rect 381261 994528 392367 994530
rect 381261 994472 381266 994528
rect 381322 994472 392306 994528
rect 392362 994472 392367 994528
rect 381261 994470 392367 994472
rect 381261 994467 381327 994470
rect 392301 994467 392367 994470
rect 471789 994530 471855 994533
rect 481541 994530 481607 994533
rect 471789 994528 481607 994530
rect 471789 994472 471794 994528
rect 471850 994472 481546 994528
rect 481602 994472 481607 994528
rect 471789 994470 481607 994472
rect 471789 994467 471855 994470
rect 481541 994467 481607 994470
rect 520917 994530 520983 994533
rect 535545 994530 535611 994533
rect 520917 994528 535611 994530
rect 520917 994472 520922 994528
rect 520978 994472 535550 994528
rect 535606 994472 535611 994528
rect 520917 994470 535611 994472
rect 520917 994467 520983 994470
rect 535545 994467 535611 994470
rect 85021 994258 85087 994261
rect 94497 994258 94563 994261
rect 85021 994256 94563 994258
rect 85021 994200 85026 994256
rect 85082 994200 94502 994256
rect 94558 994200 94563 994256
rect 85021 994198 94563 994200
rect 85021 994195 85087 994198
rect 94497 994195 94563 994198
rect 136449 994258 136515 994261
rect 145557 994258 145623 994261
rect 136449 994256 145623 994258
rect 136449 994200 136454 994256
rect 136510 994200 145562 994256
rect 145618 994200 145623 994256
rect 136449 994198 145623 994200
rect 136449 994195 136515 994198
rect 145557 994195 145623 994198
rect 192937 994258 193003 994261
rect 199377 994258 199443 994261
rect 192937 994256 199443 994258
rect 192937 994200 192942 994256
rect 192998 994200 199382 994256
rect 199438 994200 199443 994256
rect 192937 994198 199443 994200
rect 192937 994195 193003 994198
rect 199377 994195 199443 994198
rect 236545 994258 236611 994261
rect 252001 994258 252067 994261
rect 236545 994256 252067 994258
rect 236545 994200 236550 994256
rect 236606 994200 252006 994256
rect 252062 994200 252067 994256
rect 236545 994198 252067 994200
rect 236545 994195 236611 994198
rect 252001 994195 252067 994198
rect 287513 994258 287579 994261
rect 304257 994258 304323 994261
rect 287513 994256 304323 994258
rect 287513 994200 287518 994256
rect 287574 994200 304262 994256
rect 304318 994200 304323 994256
rect 287513 994198 304323 994200
rect 287513 994195 287579 994198
rect 304257 994195 304323 994198
rect 378409 994258 378475 994261
rect 393221 994258 393287 994261
rect 378409 994256 393287 994258
rect 378409 994200 378414 994256
rect 378470 994200 393226 994256
rect 393282 994200 393287 994256
rect 378409 994198 393287 994200
rect 378409 994195 378475 994198
rect 393221 994195 393287 994198
rect 454677 994258 454743 994261
rect 480110 994258 480116 994260
rect 454677 994256 480116 994258
rect 454677 994200 454682 994256
rect 454738 994200 480116 994256
rect 454677 994198 480116 994200
rect 454677 994195 454743 994198
rect 480110 994196 480116 994198
rect 480180 994196 480186 994260
rect 518157 994258 518223 994261
rect 533705 994258 533771 994261
rect 518157 994256 533771 994258
rect 518157 994200 518162 994256
rect 518218 994200 533710 994256
rect 533766 994200 533771 994256
rect 518157 994198 533771 994200
rect 518157 994195 518223 994198
rect 533705 994195 533771 994198
rect 188153 993986 188219 993989
rect 196617 993986 196683 993989
rect 188153 993984 196683 993986
rect 188153 993928 188158 993984
rect 188214 993928 196622 993984
rect 196678 993928 196683 993984
rect 188153 993926 196683 993928
rect 188153 993923 188219 993926
rect 196617 993923 196683 993926
rect 240133 993986 240199 993989
rect 251817 993986 251883 993989
rect 240133 993984 251883 993986
rect 240133 993928 240138 993984
rect 240194 993928 251822 993984
rect 251878 993928 251883 993984
rect 240133 993926 251883 993928
rect 240133 993923 240199 993926
rect 251817 993923 251883 993926
rect 290273 993986 290339 993989
rect 307017 993986 307083 993989
rect 290273 993984 307083 993986
rect 290273 993928 290278 993984
rect 290334 993928 307022 993984
rect 307078 993928 307083 993984
rect 290273 993926 307083 993928
rect 290273 993923 290339 993926
rect 307017 993923 307083 993926
rect 443453 993986 443519 993989
rect 477953 993986 478019 993989
rect 443453 993984 478019 993986
rect 443453 993928 443458 993984
rect 443514 993928 477958 993984
rect 478014 993928 478019 993984
rect 443453 993926 478019 993928
rect 443453 993923 443519 993926
rect 477953 993923 478019 993926
rect 522941 993986 523007 993989
rect 536741 993986 536807 993989
rect 522941 993984 536807 993986
rect 522941 993928 522946 993984
rect 523002 993928 536746 993984
rect 536802 993928 536807 993984
rect 522941 993926 536807 993928
rect 522941 993923 523007 993926
rect 536741 993923 536807 993926
rect 191741 993170 191807 993173
rect 251449 993170 251515 993173
rect 191741 993168 251515 993170
rect 191741 993112 191746 993168
rect 191802 993112 251454 993168
rect 251510 993112 251515 993168
rect 191741 993110 251515 993112
rect 191741 993107 191807 993110
rect 251449 993107 251515 993110
rect 242934 992836 242940 992900
rect 243004 992898 243010 992900
rect 316401 992898 316467 992901
rect 243004 992896 316467 992898
rect 243004 992840 316406 992896
rect 316462 992840 316467 992896
rect 243004 992838 316467 992840
rect 243004 992836 243010 992838
rect 316401 992835 316467 992838
rect 62113 976034 62179 976037
rect 62113 976032 64492 976034
rect 62113 975976 62118 976032
rect 62174 975976 64492 976032
rect 62113 975974 64492 975976
rect 62113 975971 62179 975974
rect 651649 975898 651715 975901
rect 650164 975896 651715 975898
rect 650164 975840 651654 975896
rect 651710 975840 651715 975896
rect 650164 975838 651715 975840
rect 651649 975835 651715 975838
rect 41454 968764 41460 968828
rect 41524 968826 41530 968828
rect 41781 968826 41847 968829
rect 41524 968824 41847 968826
rect 41524 968768 41786 968824
rect 41842 968768 41847 968824
rect 41524 968766 41847 968768
rect 41524 968764 41530 968766
rect 41781 968763 41847 968766
rect 41965 967196 42031 967197
rect 41965 967192 42012 967196
rect 42076 967194 42082 967196
rect 41965 967136 41970 967192
rect 41965 967132 42012 967136
rect 42076 967134 42122 967194
rect 42076 967132 42082 967134
rect 41965 967131 42031 967132
rect 675385 966516 675451 966517
rect 675334 966514 675340 966516
rect 675294 966454 675340 966514
rect 675404 966512 675451 966516
rect 675446 966456 675451 966512
rect 675334 966452 675340 966454
rect 675404 966452 675451 966456
rect 675385 966451 675451 966452
rect 675753 965154 675819 965157
rect 676070 965154 676076 965156
rect 675753 965152 676076 965154
rect 675753 965096 675758 965152
rect 675814 965096 676076 965152
rect 675753 965094 676076 965096
rect 675753 965091 675819 965094
rect 676070 965092 676076 965094
rect 676140 965092 676146 965156
rect 675201 963388 675267 963389
rect 675150 963386 675156 963388
rect 675110 963326 675156 963386
rect 675220 963384 675267 963388
rect 675262 963328 675267 963384
rect 675150 963324 675156 963326
rect 675220 963324 675267 963328
rect 675201 963323 675267 963324
rect 62113 962978 62179 962981
rect 62113 962976 64492 962978
rect 62113 962920 62118 962976
rect 62174 962920 64492 962976
rect 62113 962918 64492 962920
rect 62113 962915 62179 962918
rect 651649 962570 651715 962573
rect 650164 962568 651715 962570
rect 650164 962512 651654 962568
rect 651710 962512 651715 962568
rect 650164 962510 651715 962512
rect 651649 962507 651715 962510
rect 41781 962164 41847 962165
rect 41781 962160 41828 962164
rect 41892 962162 41898 962164
rect 41781 962104 41786 962160
rect 41781 962100 41828 962104
rect 41892 962102 41938 962162
rect 41892 962100 41898 962102
rect 41781 962099 41847 962100
rect 675753 962026 675819 962029
rect 676622 962026 676628 962028
rect 675753 962024 676628 962026
rect 675753 961968 675758 962024
rect 675814 961968 676628 962024
rect 675753 961966 676628 961968
rect 675753 961963 675819 961966
rect 676622 961964 676628 961966
rect 676692 961964 676698 962028
rect 674925 959442 674991 959445
rect 675150 959442 675156 959444
rect 674925 959440 675156 959442
rect 674925 959384 674930 959440
rect 674986 959384 675156 959440
rect 674925 959382 675156 959384
rect 674925 959379 674991 959382
rect 675150 959380 675156 959382
rect 675220 959380 675226 959444
rect 41270 959108 41276 959172
rect 41340 959170 41346 959172
rect 41781 959170 41847 959173
rect 41340 959168 41847 959170
rect 41340 959112 41786 959168
rect 41842 959112 41847 959168
rect 41340 959110 41847 959112
rect 41340 959108 41346 959110
rect 41781 959107 41847 959110
rect 672901 959170 672967 959173
rect 675109 959170 675175 959173
rect 672901 959168 675175 959170
rect 672901 959112 672906 959168
rect 672962 959112 675114 959168
rect 675170 959112 675175 959168
rect 672901 959110 675175 959112
rect 672901 959107 672967 959110
rect 675109 959107 675175 959110
rect 675753 958354 675819 958357
rect 676806 958354 676812 958356
rect 675753 958352 676812 958354
rect 675753 958296 675758 958352
rect 675814 958296 676812 958352
rect 675753 958294 676812 958296
rect 675753 958291 675819 958294
rect 676806 958292 676812 958294
rect 676876 958292 676882 958356
rect 40718 956524 40724 956588
rect 40788 956586 40794 956588
rect 41781 956586 41847 956589
rect 40788 956584 41847 956586
rect 40788 956528 41786 956584
rect 41842 956528 41847 956584
rect 40788 956526 41847 956528
rect 40788 956524 40794 956526
rect 41781 956523 41847 956526
rect 675753 956450 675819 956453
rect 676990 956450 676996 956452
rect 675753 956448 676996 956450
rect 675753 956392 675758 956448
rect 675814 956392 676996 956448
rect 675753 956390 676996 956392
rect 675753 956387 675819 956390
rect 676990 956388 676996 956390
rect 677060 956388 677066 956452
rect 40534 955436 40540 955500
rect 40604 955498 40610 955500
rect 41781 955498 41847 955501
rect 40604 955496 41847 955498
rect 40604 955440 41786 955496
rect 41842 955440 41847 955496
rect 40604 955438 41847 955440
rect 40604 955436 40610 955438
rect 41781 955435 41847 955438
rect 675661 954002 675727 954005
rect 675886 954002 675892 954004
rect 675661 954000 675892 954002
rect 675661 953944 675666 954000
rect 675722 953944 675892 954000
rect 675661 953942 675892 953944
rect 675661 953939 675727 953942
rect 675886 953940 675892 953942
rect 675956 953940 675962 954004
rect 35157 952914 35223 952917
rect 41454 952914 41460 952916
rect 35157 952912 41460 952914
rect 35157 952856 35162 952912
rect 35218 952856 41460 952912
rect 35157 952854 41460 952856
rect 35157 952851 35223 952854
rect 41454 952852 41460 952854
rect 41524 952852 41530 952916
rect 39297 952234 39363 952237
rect 41638 952234 41644 952236
rect 39297 952232 41644 952234
rect 39297 952176 39302 952232
rect 39358 952176 41644 952232
rect 39297 952174 41644 952176
rect 39297 952171 39363 952174
rect 41638 952172 41644 952174
rect 41708 952172 41714 952236
rect 674465 952234 674531 952237
rect 675385 952234 675451 952237
rect 674465 952232 675451 952234
rect 674465 952176 674470 952232
rect 674526 952176 675390 952232
rect 675446 952176 675451 952232
rect 674465 952174 675451 952176
rect 674465 952171 674531 952174
rect 675385 952171 675451 952174
rect 40033 951826 40099 951829
rect 41270 951826 41276 951828
rect 40033 951824 41276 951826
rect 40033 951768 40038 951824
rect 40094 951768 41276 951824
rect 40033 951766 41276 951768
rect 40033 951763 40099 951766
rect 41270 951764 41276 951766
rect 41340 951764 41346 951828
rect 41413 951690 41479 951693
rect 42006 951690 42012 951692
rect 41413 951688 42012 951690
rect 41413 951632 41418 951688
rect 41474 951632 42012 951688
rect 41413 951630 42012 951632
rect 41413 951627 41479 951630
rect 42006 951628 42012 951630
rect 42076 951628 42082 951692
rect 676622 951492 676628 951556
rect 676692 951554 676698 951556
rect 677501 951554 677567 951557
rect 676692 951552 677567 951554
rect 676692 951496 677506 951552
rect 677562 951496 677567 951552
rect 676692 951494 677567 951496
rect 676692 951492 676698 951494
rect 677501 951491 677567 951494
rect 676070 949996 676076 950060
rect 676140 950058 676146 950060
rect 683297 950058 683363 950061
rect 676140 950056 683363 950058
rect 676140 950000 683302 950056
rect 683358 950000 683363 950056
rect 676140 949998 683363 950000
rect 676140 949996 676146 949998
rect 683297 949995 683363 949998
rect 62113 949922 62179 949925
rect 62113 949920 64492 949922
rect 62113 949864 62118 949920
rect 62174 949864 64492 949920
rect 62113 949862 64492 949864
rect 62113 949859 62179 949862
rect 651649 949378 651715 949381
rect 650164 949376 651715 949378
rect 650164 949320 651654 949376
rect 651710 949320 651715 949376
rect 650164 949318 651715 949320
rect 651649 949315 651715 949318
rect 675937 949244 676003 949245
rect 675886 949242 675892 949244
rect 675846 949182 675892 949242
rect 675956 949240 676003 949244
rect 675998 949184 676003 949240
rect 675886 949180 675892 949182
rect 675956 949180 676003 949184
rect 675937 949179 676003 949180
rect 674925 948970 674991 948973
rect 675334 948970 675340 948972
rect 674925 948968 675340 948970
rect 674925 948912 674930 948968
rect 674986 948912 675340 948968
rect 674925 948910 675340 948912
rect 674925 948907 674991 948910
rect 675334 948908 675340 948910
rect 675404 948908 675410 948972
rect 43529 943530 43595 943533
rect 41492 943528 43595 943530
rect 41492 943472 43534 943528
rect 43590 943472 43595 943528
rect 41492 943470 43595 943472
rect 43529 943467 43595 943470
rect 44633 943122 44699 943125
rect 41492 943120 44699 943122
rect 41492 943064 44638 943120
rect 44694 943064 44699 943120
rect 41492 943062 44699 943064
rect 44633 943059 44699 943062
rect 47577 942714 47643 942717
rect 41492 942712 47643 942714
rect 41492 942656 47582 942712
rect 47638 942656 47643 942712
rect 41492 942654 47643 942656
rect 47577 942651 47643 942654
rect 43621 942306 43687 942309
rect 41492 942304 43687 942306
rect 41492 942248 43626 942304
rect 43682 942248 43687 942304
rect 41492 942246 43687 942248
rect 43621 942243 43687 942246
rect 41229 941898 41295 941901
rect 674925 941898 674991 941901
rect 675845 941898 675911 941901
rect 41229 941896 41308 941898
rect 41229 941840 41234 941896
rect 41290 941840 41308 941896
rect 41229 941838 41308 941840
rect 674925 941896 675911 941898
rect 674925 941840 674930 941896
rect 674986 941840 675850 941896
rect 675906 941840 675911 941896
rect 674925 941838 675911 941840
rect 41229 941835 41295 941838
rect 674925 941835 674991 941838
rect 675845 941835 675911 941838
rect 41492 941430 41890 941490
rect 41830 941354 41890 941430
rect 43437 941354 43503 941357
rect 41830 941352 43503 941354
rect 41830 941296 43442 941352
rect 43498 941296 43503 941352
rect 41830 941294 43503 941296
rect 43437 941291 43503 941294
rect 41229 941082 41295 941085
rect 41229 941080 41308 941082
rect 41229 941024 41234 941080
rect 41290 941024 41308 941080
rect 41229 941022 41308 941024
rect 41229 941019 41295 941022
rect 46197 940674 46263 940677
rect 41492 940672 46263 940674
rect 41492 940616 46202 940672
rect 46258 940616 46263 940672
rect 41492 940614 46263 940616
rect 46197 940611 46263 940614
rect 41229 940266 41295 940269
rect 41229 940264 41308 940266
rect 41229 940208 41234 940264
rect 41290 940208 41308 940264
rect 41229 940206 41308 940208
rect 41229 940203 41295 940206
rect 675477 939994 675543 939997
rect 675477 939992 676292 939994
rect 675477 939936 675482 939992
rect 675538 939936 676292 939992
rect 675477 939934 676292 939936
rect 675477 939931 675543 939934
rect 43437 939858 43503 939861
rect 41492 939856 43503 939858
rect 41492 939800 43442 939856
rect 43498 939800 43503 939856
rect 41492 939798 43503 939800
rect 43437 939795 43503 939798
rect 675661 939586 675727 939589
rect 675661 939584 676292 939586
rect 675661 939528 675666 939584
rect 675722 939528 676292 939584
rect 675661 939526 676292 939528
rect 675661 939523 675727 939526
rect 41045 939450 41111 939453
rect 41045 939448 41124 939450
rect 41045 939392 41050 939448
rect 41106 939392 41124 939448
rect 41045 939390 41124 939392
rect 41045 939387 41111 939390
rect 675293 939178 675359 939181
rect 675293 939176 676292 939178
rect 675293 939120 675298 939176
rect 675354 939120 676292 939176
rect 675293 939118 676292 939120
rect 675293 939115 675359 939118
rect 41822 939042 41828 939044
rect 41492 938982 41828 939042
rect 41822 938980 41828 938982
rect 41892 938980 41898 939044
rect 675477 938770 675543 938773
rect 675477 938768 676292 938770
rect 675477 938712 675482 938768
rect 675538 938712 676292 938768
rect 675477 938710 676292 938712
rect 675477 938707 675543 938710
rect 41278 938467 41338 938604
rect 37917 938464 37983 938467
rect 37917 938462 38026 938464
rect 37917 938406 37922 938462
rect 37978 938406 38026 938462
rect 37917 938401 38026 938406
rect 41229 938462 41338 938467
rect 41229 938406 41234 938462
rect 41290 938406 41338 938462
rect 41229 938404 41338 938406
rect 41229 938401 41295 938404
rect 37966 938196 38026 938401
rect 674925 938362 674991 938365
rect 674925 938360 676292 938362
rect 674925 938304 674930 938360
rect 674986 938304 676292 938360
rect 674925 938302 676292 938304
rect 674925 938299 674991 938302
rect 675293 937954 675359 937957
rect 675293 937952 676292 937954
rect 675293 937896 675298 937952
rect 675354 937896 676292 937952
rect 675293 937894 676292 937896
rect 675293 937891 675359 937894
rect 42241 937818 42307 937821
rect 41492 937816 42307 937818
rect 41492 937760 42246 937816
rect 42302 937760 42307 937816
rect 41492 937758 42307 937760
rect 42241 937755 42307 937758
rect 675477 937546 675543 937549
rect 675477 937544 676292 937546
rect 675477 937488 675482 937544
rect 675538 937488 676292 937544
rect 675477 937486 676292 937488
rect 675477 937483 675543 937486
rect 39297 937410 39363 937413
rect 39284 937408 39363 937410
rect 39284 937352 39302 937408
rect 39358 937352 39363 937408
rect 39284 937350 39363 937352
rect 39297 937347 39363 937350
rect 675477 937138 675543 937141
rect 675477 937136 676292 937138
rect 675477 937080 675482 937136
rect 675538 937080 676292 937136
rect 675477 937078 676292 937080
rect 675477 937075 675543 937078
rect 35157 937002 35223 937005
rect 62113 937002 62179 937005
rect 35157 937000 35236 937002
rect 35157 936944 35162 937000
rect 35218 936944 35236 937000
rect 35157 936942 35236 936944
rect 62113 937000 64492 937002
rect 62113 936944 62118 937000
rect 62174 936944 64492 937000
rect 62113 936942 64492 936944
rect 35157 936939 35223 936942
rect 62113 936939 62179 936942
rect 675661 936730 675727 936733
rect 675661 936728 676292 936730
rect 675661 936672 675666 936728
rect 675722 936672 676292 936728
rect 675661 936670 676292 936672
rect 675661 936667 675727 936670
rect 41822 936594 41828 936596
rect 41492 936534 41828 936594
rect 41822 936532 41828 936534
rect 41892 936532 41898 936596
rect 675477 936322 675543 936325
rect 675477 936320 676292 936322
rect 675477 936264 675482 936320
rect 675538 936264 676292 936320
rect 675477 936262 676292 936264
rect 675477 936259 675543 936262
rect 44817 936186 44883 936189
rect 651649 936186 651715 936189
rect 41492 936184 44883 936186
rect 41492 936128 44822 936184
rect 44878 936128 44883 936184
rect 41492 936126 44883 936128
rect 650164 936184 651715 936186
rect 650164 936128 651654 936184
rect 651710 936128 651715 936184
rect 650164 936126 651715 936128
rect 44817 936123 44883 936126
rect 651649 936123 651715 936126
rect 675293 935914 675359 935917
rect 675293 935912 676292 935914
rect 675293 935856 675298 935912
rect 675354 935856 676292 935912
rect 675293 935854 676292 935856
rect 675293 935851 675359 935854
rect 40033 935778 40099 935781
rect 40020 935776 40099 935778
rect 40020 935720 40038 935776
rect 40094 935720 40099 935776
rect 40020 935718 40099 935720
rect 40033 935715 40099 935718
rect 683297 935642 683363 935645
rect 683254 935640 683363 935642
rect 683254 935584 683302 935640
rect 683358 935584 683363 935640
rect 683254 935579 683363 935584
rect 683254 935476 683314 935579
rect 42793 935370 42859 935373
rect 41492 935368 42859 935370
rect 41492 935312 42798 935368
rect 42854 935312 42859 935368
rect 41492 935310 42859 935312
rect 42793 935307 42859 935310
rect 682377 935234 682443 935237
rect 682334 935232 682443 935234
rect 682334 935176 682382 935232
rect 682438 935176 682443 935232
rect 682334 935171 682443 935176
rect 682334 935068 682394 935171
rect 43069 934962 43135 934965
rect 41492 934960 43135 934962
rect 41492 934904 43074 934960
rect 43130 934904 43135 934960
rect 41492 934902 43135 934904
rect 43069 934899 43135 934902
rect 675845 934690 675911 934693
rect 675845 934688 676292 934690
rect 675845 934632 675850 934688
rect 675906 934632 676292 934688
rect 675845 934630 676292 934632
rect 675845 934627 675911 934630
rect 43253 934554 43319 934557
rect 41492 934552 43319 934554
rect 41492 934496 43258 934552
rect 43314 934496 43319 934552
rect 41492 934494 43319 934496
rect 43253 934491 43319 934494
rect 44449 934146 44515 934149
rect 41492 934144 44515 934146
rect 41492 934088 44454 934144
rect 44510 934088 44515 934144
rect 41492 934086 44515 934088
rect 44449 934083 44515 934086
rect 675109 934146 675175 934149
rect 676262 934146 676322 934252
rect 675109 934144 676322 934146
rect 675109 934088 675114 934144
rect 675170 934088 676322 934144
rect 675109 934086 676322 934088
rect 675109 934083 675175 934086
rect 675293 933874 675359 933877
rect 675293 933872 676292 933874
rect 675293 933816 675298 933872
rect 675354 933816 676292 933872
rect 675293 933814 676292 933816
rect 675293 933811 675359 933814
rect 44173 933738 44239 933741
rect 41492 933736 44239 933738
rect 41492 933680 44178 933736
rect 44234 933680 44239 933736
rect 41492 933678 44239 933680
rect 44173 933675 44239 933678
rect 674465 933466 674531 933469
rect 674465 933464 676292 933466
rect 674465 933408 674470 933464
rect 674526 933408 676292 933464
rect 674465 933406 676292 933408
rect 674465 933403 674531 933406
rect 42977 933330 43043 933333
rect 41492 933328 43043 933330
rect 41492 933272 42982 933328
rect 43038 933272 43043 933328
rect 41492 933270 43043 933272
rect 42977 933267 43043 933270
rect 675477 933058 675543 933061
rect 675477 933056 676292 933058
rect 675477 933000 675482 933056
rect 675538 933000 676292 933056
rect 675477 932998 676292 933000
rect 675477 932995 675543 932998
rect 42425 932922 42491 932925
rect 41492 932920 42491 932922
rect 27662 932484 27722 932892
rect 41492 932864 42430 932920
rect 42486 932864 42491 932920
rect 41492 932862 42491 932864
rect 42425 932859 42491 932862
rect 674649 932650 674715 932653
rect 674649 932648 676292 932650
rect 674649 932592 674654 932648
rect 674710 932592 676292 932648
rect 674649 932590 676292 932592
rect 674649 932587 674715 932590
rect 674281 932242 674347 932245
rect 674281 932240 676292 932242
rect 674281 932184 674286 932240
rect 674342 932184 676292 932240
rect 674281 932182 676292 932184
rect 674281 932179 674347 932182
rect 42793 932106 42859 932109
rect 41492 932104 42859 932106
rect 41492 932048 42798 932104
rect 42854 932048 42859 932104
rect 41492 932046 42859 932048
rect 42793 932043 42859 932046
rect 676990 931908 676996 931972
rect 677060 931908 677066 931972
rect 676998 931804 677058 931908
rect 675477 931426 675543 931429
rect 675477 931424 676292 931426
rect 675477 931368 675482 931424
rect 675538 931368 676292 931424
rect 675477 931366 676292 931368
rect 675477 931363 675543 931366
rect 677501 931154 677567 931157
rect 677501 931152 677610 931154
rect 677501 931096 677506 931152
rect 677562 931096 677610 931152
rect 677501 931091 677610 931096
rect 677550 930988 677610 931091
rect 676806 930684 676812 930748
rect 676876 930684 676882 930748
rect 676814 930580 676874 930684
rect 675477 930202 675543 930205
rect 675477 930200 676292 930202
rect 675477 930144 675482 930200
rect 675538 930144 676292 930200
rect 675477 930142 676292 930144
rect 675477 930139 675543 930142
rect 675477 929794 675543 929797
rect 675477 929792 676292 929794
rect 675477 929736 675482 929792
rect 675538 929736 676292 929792
rect 675477 929734 676292 929736
rect 675477 929731 675543 929734
rect 683113 929522 683179 929525
rect 683070 929520 683179 929522
rect 683070 929464 683118 929520
rect 683174 929464 683179 929520
rect 683070 929459 683179 929464
rect 683070 928948 683130 929459
rect 675477 928570 675543 928573
rect 675477 928568 676292 928570
rect 675477 928512 675482 928568
rect 675538 928512 676292 928568
rect 675477 928510 676292 928512
rect 675477 928507 675543 928510
rect 62113 923810 62179 923813
rect 62113 923808 64492 923810
rect 62113 923752 62118 923808
rect 62174 923752 64492 923808
rect 62113 923750 64492 923752
rect 62113 923747 62179 923750
rect 651649 922722 651715 922725
rect 650164 922720 651715 922722
rect 650164 922664 651654 922720
rect 651710 922664 651715 922720
rect 650164 922662 651715 922664
rect 651649 922659 651715 922662
rect 62113 910754 62179 910757
rect 62113 910752 64492 910754
rect 62113 910696 62118 910752
rect 62174 910696 64492 910752
rect 62113 910694 64492 910696
rect 62113 910691 62179 910694
rect 651649 909530 651715 909533
rect 650164 909528 651715 909530
rect 650164 909472 651654 909528
rect 651710 909472 651715 909528
rect 650164 909470 651715 909472
rect 651649 909467 651715 909470
rect 62113 897834 62179 897837
rect 62113 897832 64492 897834
rect 62113 897776 62118 897832
rect 62174 897776 64492 897832
rect 62113 897774 64492 897776
rect 62113 897771 62179 897774
rect 651649 896202 651715 896205
rect 650164 896200 651715 896202
rect 650164 896144 651654 896200
rect 651710 896144 651715 896200
rect 650164 896142 651715 896144
rect 651649 896139 651715 896142
rect 62113 884778 62179 884781
rect 62113 884776 64492 884778
rect 62113 884720 62118 884776
rect 62174 884720 64492 884776
rect 62113 884718 64492 884720
rect 62113 884715 62179 884718
rect 651649 882874 651715 882877
rect 650164 882872 651715 882874
rect 650164 882816 651654 882872
rect 651710 882816 651715 882872
rect 650164 882814 651715 882816
rect 651649 882811 651715 882814
rect 40677 881922 40743 881925
rect 42425 881922 42491 881925
rect 40677 881920 42491 881922
rect 40677 881864 40682 881920
rect 40738 881864 42430 881920
rect 42486 881864 42491 881920
rect 40677 881862 42491 881864
rect 40677 881859 40743 881862
rect 42425 881859 42491 881862
rect 675753 877162 675819 877165
rect 676070 877162 676076 877164
rect 675753 877160 676076 877162
rect 675753 877104 675758 877160
rect 675814 877104 676076 877160
rect 675753 877102 676076 877104
rect 675753 877099 675819 877102
rect 676070 877100 676076 877102
rect 676140 877100 676146 877164
rect 675293 876482 675359 876485
rect 676990 876482 676996 876484
rect 675293 876480 676996 876482
rect 675293 876424 675298 876480
rect 675354 876424 676996 876480
rect 675293 876422 676996 876424
rect 675293 876419 675359 876422
rect 676990 876420 676996 876422
rect 677060 876420 677066 876484
rect 675385 874036 675451 874037
rect 675334 874034 675340 874036
rect 675294 873974 675340 874034
rect 675404 874032 675451 874036
rect 675446 873976 675451 874032
rect 675334 873972 675340 873974
rect 675404 873972 675451 873976
rect 675385 873971 675451 873972
rect 675753 872810 675819 872813
rect 676806 872810 676812 872812
rect 675753 872808 676812 872810
rect 675753 872752 675758 872808
rect 675814 872752 676812 872808
rect 675753 872750 676812 872752
rect 675753 872747 675819 872750
rect 676806 872748 676812 872750
rect 676876 872748 676882 872812
rect 673862 872204 673868 872268
rect 673932 872266 673938 872268
rect 675385 872266 675451 872269
rect 673932 872264 675451 872266
rect 673932 872208 675390 872264
rect 675446 872208 675451 872264
rect 673932 872206 675451 872208
rect 673932 872204 673938 872206
rect 675385 872203 675451 872206
rect 62113 871722 62179 871725
rect 62113 871720 64492 871722
rect 62113 871664 62118 871720
rect 62174 871664 64492 871720
rect 62113 871662 64492 871664
rect 62113 871659 62179 871662
rect 651649 869682 651715 869685
rect 650164 869680 651715 869682
rect 650164 869624 651654 869680
rect 651710 869624 651715 869680
rect 650164 869622 651715 869624
rect 651649 869619 651715 869622
rect 674833 869682 674899 869685
rect 675334 869682 675340 869684
rect 674833 869680 675340 869682
rect 674833 869624 674838 869680
rect 674894 869624 675340 869680
rect 674833 869622 675340 869624
rect 674833 869619 674899 869622
rect 675334 869620 675340 869622
rect 675404 869620 675410 869684
rect 675661 869682 675727 869685
rect 675886 869682 675892 869684
rect 675661 869680 675892 869682
rect 675661 869624 675666 869680
rect 675722 869624 675892 869680
rect 675661 869622 675892 869624
rect 675661 869619 675727 869622
rect 675886 869620 675892 869622
rect 675956 869620 675962 869684
rect 672349 868050 672415 868053
rect 675477 868050 675543 868053
rect 672349 868048 675543 868050
rect 672349 867992 672354 868048
rect 672410 867992 675482 868048
rect 675538 867992 675543 868048
rect 672349 867990 675543 867992
rect 672349 867987 672415 867990
rect 675477 867987 675543 867990
rect 672993 864242 673059 864245
rect 675477 864242 675543 864245
rect 672993 864240 675543 864242
rect 672993 864184 672998 864240
rect 673054 864184 675482 864240
rect 675538 864184 675543 864240
rect 672993 864182 675543 864184
rect 672993 864179 673059 864182
rect 675477 864179 675543 864182
rect 674833 863834 674899 863837
rect 675477 863834 675543 863837
rect 674833 863832 675543 863834
rect 674833 863776 674838 863832
rect 674894 863776 675482 863832
rect 675538 863776 675543 863832
rect 674833 863774 675543 863776
rect 674833 863771 674899 863774
rect 675477 863771 675543 863774
rect 62113 858666 62179 858669
rect 62113 858664 64492 858666
rect 62113 858608 62118 858664
rect 62174 858608 64492 858664
rect 62113 858606 64492 858608
rect 62113 858603 62179 858606
rect 651649 856354 651715 856357
rect 650164 856352 651715 856354
rect 650164 856296 651654 856352
rect 651710 856296 651715 856352
rect 650164 856294 651715 856296
rect 651649 856291 651715 856294
rect 674465 854316 674531 854317
rect 674414 854314 674420 854316
rect 674374 854254 674420 854314
rect 674484 854312 674531 854316
rect 674526 854256 674531 854312
rect 674414 854252 674420 854254
rect 674484 854252 674531 854256
rect 674465 854251 674531 854252
rect 62113 845610 62179 845613
rect 62113 845608 64492 845610
rect 62113 845552 62118 845608
rect 62174 845552 64492 845608
rect 62113 845550 64492 845552
rect 62113 845547 62179 845550
rect 651649 843026 651715 843029
rect 650164 843024 651715 843026
rect 650164 842968 651654 843024
rect 651710 842968 651715 843024
rect 650164 842966 651715 842968
rect 651649 842963 651715 842966
rect 62113 832554 62179 832557
rect 62113 832552 64492 832554
rect 62113 832496 62118 832552
rect 62174 832496 64492 832552
rect 62113 832494 64492 832496
rect 62113 832491 62179 832494
rect 651649 829834 651715 829837
rect 650164 829832 651715 829834
rect 650164 829776 651654 829832
rect 651710 829776 651715 829832
rect 650164 829774 651715 829776
rect 651649 829771 651715 829774
rect 62113 819498 62179 819501
rect 62113 819496 64492 819498
rect 62113 819440 62118 819496
rect 62174 819440 64492 819496
rect 62113 819438 64492 819440
rect 62113 819435 62179 819438
rect 40217 819090 40283 819093
rect 46197 819090 46263 819093
rect 40217 819088 46263 819090
rect 40217 819032 40222 819088
rect 40278 819032 46202 819088
rect 46258 819032 46263 819088
rect 40217 819030 46263 819032
rect 40217 819027 40283 819030
rect 46197 819027 46263 819030
rect 39573 818682 39639 818685
rect 42057 818682 42123 818685
rect 39573 818680 42123 818682
rect 39573 818624 39578 818680
rect 39634 818624 42062 818680
rect 42118 818624 42123 818680
rect 39573 818622 42123 818624
rect 39573 818619 39639 818622
rect 42057 818619 42123 818622
rect 35617 818002 35683 818005
rect 35574 818000 35683 818002
rect 35574 817944 35622 818000
rect 35678 817944 35683 818000
rect 35574 817939 35683 817944
rect 39757 818002 39823 818005
rect 41873 818002 41939 818005
rect 39757 818000 41939 818002
rect 39757 817944 39762 818000
rect 39818 817944 41878 818000
rect 41934 817944 41939 818000
rect 39757 817942 41939 817944
rect 39757 817939 39823 817942
rect 41873 817939 41939 817942
rect 35574 817700 35634 817939
rect 35801 817322 35867 817325
rect 35788 817320 35867 817322
rect 35788 817264 35806 817320
rect 35862 817264 35867 817320
rect 35788 817262 35867 817264
rect 35801 817259 35867 817262
rect 35433 816914 35499 816917
rect 35420 816912 35499 816914
rect 35420 816856 35438 816912
rect 35494 816856 35499 816912
rect 35420 816854 35499 816856
rect 35433 816851 35499 816854
rect 35801 816506 35867 816509
rect 651649 816506 651715 816509
rect 35788 816504 35867 816506
rect 35788 816448 35806 816504
rect 35862 816448 35867 816504
rect 35788 816446 35867 816448
rect 650164 816504 651715 816506
rect 650164 816448 651654 816504
rect 651710 816448 651715 816504
rect 650164 816446 651715 816448
rect 35801 816443 35867 816446
rect 651649 816443 651715 816446
rect 35801 816098 35867 816101
rect 35788 816096 35867 816098
rect 35788 816040 35806 816096
rect 35862 816040 35867 816096
rect 35788 816038 35867 816040
rect 35801 816035 35867 816038
rect 35617 815690 35683 815693
rect 35604 815688 35683 815690
rect 35604 815632 35622 815688
rect 35678 815632 35683 815688
rect 35604 815630 35683 815632
rect 35617 815627 35683 815630
rect 35617 815282 35683 815285
rect 35604 815280 35683 815282
rect 35604 815224 35622 815280
rect 35678 815224 35683 815280
rect 35604 815222 35683 815224
rect 35617 815219 35683 815222
rect 35801 814874 35867 814877
rect 35788 814872 35867 814874
rect 35788 814816 35806 814872
rect 35862 814816 35867 814872
rect 35788 814814 35867 814816
rect 35801 814811 35867 814814
rect 35801 814466 35867 814469
rect 35788 814464 35867 814466
rect 35788 814408 35806 814464
rect 35862 814408 35867 814464
rect 35788 814406 35867 814408
rect 35801 814403 35867 814406
rect 41045 814058 41111 814061
rect 41781 814058 41847 814061
rect 44449 814058 44515 814061
rect 41045 814056 41124 814058
rect 41045 814000 41050 814056
rect 41106 814000 41124 814056
rect 41045 813998 41124 814000
rect 41781 814056 44515 814058
rect 41781 814000 41786 814056
rect 41842 814000 44454 814056
rect 44510 814000 44515 814056
rect 41781 813998 44515 814000
rect 41045 813995 41111 813998
rect 41781 813995 41847 813998
rect 44449 813995 44515 813998
rect 43253 813650 43319 813653
rect 41492 813648 43319 813650
rect 41492 813592 43258 813648
rect 43314 813592 43319 813648
rect 41492 813590 43319 813592
rect 43253 813587 43319 813590
rect 42006 813242 42012 813244
rect 41492 813182 42012 813242
rect 42006 813180 42012 813182
rect 42076 813180 42082 813244
rect 40769 812834 40835 812837
rect 40756 812832 40835 812834
rect 40756 812776 40774 812832
rect 40830 812776 40835 812832
rect 40756 812774 40835 812776
rect 40769 812771 40835 812774
rect 35157 812426 35223 812429
rect 35157 812424 35236 812426
rect 35157 812368 35162 812424
rect 35218 812368 35236 812424
rect 35157 812366 35236 812368
rect 35157 812363 35223 812366
rect 40953 812018 41019 812021
rect 40940 812016 41019 812018
rect 40940 811960 40958 812016
rect 41014 811960 41019 812016
rect 40940 811958 41019 811960
rect 40953 811955 41019 811958
rect 41321 811610 41387 811613
rect 41308 811608 41387 811610
rect 41308 811552 41326 811608
rect 41382 811552 41387 811608
rect 41308 811550 41387 811552
rect 41321 811547 41387 811550
rect 32397 811202 32463 811205
rect 32397 811200 32476 811202
rect 32397 811144 32402 811200
rect 32458 811144 32476 811200
rect 32397 811142 32476 811144
rect 32397 811139 32463 811142
rect 40542 810762 40602 810764
rect 40534 810698 40540 810762
rect 40604 810698 40610 810762
rect 40718 810562 40724 810626
rect 40788 810562 40794 810626
rect 40726 810356 40786 810562
rect 31661 809978 31727 809981
rect 31661 809976 31740 809978
rect 31661 809920 31666 809976
rect 31722 809920 31740 809976
rect 31661 809918 31740 809920
rect 31661 809915 31727 809918
rect 33777 809570 33843 809573
rect 33764 809568 33843 809570
rect 33764 809512 33782 809568
rect 33838 809512 33843 809568
rect 33764 809510 33843 809512
rect 33777 809507 33843 809510
rect 41781 809300 41847 809301
rect 41781 809296 41828 809300
rect 41892 809298 41898 809300
rect 41781 809240 41786 809296
rect 41781 809236 41828 809240
rect 41892 809238 41938 809298
rect 41892 809236 41898 809238
rect 41781 809235 41847 809236
rect 36537 809162 36603 809165
rect 36524 809160 36603 809162
rect 36524 809104 36542 809160
rect 36598 809104 36603 809160
rect 36524 809102 36603 809104
rect 36537 809099 36603 809102
rect 43069 808754 43135 808757
rect 41492 808752 43135 808754
rect 41492 808696 43074 808752
rect 43130 808696 43135 808752
rect 41492 808694 43135 808696
rect 43069 808691 43135 808694
rect 41781 808346 41847 808349
rect 41492 808344 41847 808346
rect 41492 808288 41786 808344
rect 41842 808288 41847 808344
rect 41492 808286 41847 808288
rect 41781 808283 41847 808286
rect 44633 807938 44699 807941
rect 41492 807936 44699 807938
rect 41492 807880 44638 807936
rect 44694 807880 44699 807936
rect 41492 807878 44699 807880
rect 44633 807875 44699 807878
rect 41321 807530 41387 807533
rect 41308 807528 41387 807530
rect 41308 807472 41326 807528
rect 41382 807472 41387 807528
rect 41308 807470 41387 807472
rect 41321 807467 41387 807470
rect 41462 806714 41522 807092
rect 42057 806714 42123 806717
rect 41462 806712 42123 806714
rect 41462 806684 42062 806712
rect 41492 806656 42062 806684
rect 42118 806656 42123 806712
rect 41492 806654 42123 806656
rect 42057 806651 42123 806654
rect 62113 806578 62179 806581
rect 62113 806576 64492 806578
rect 62113 806520 62118 806576
rect 62174 806520 64492 806576
rect 62113 806518 64492 806520
rect 62113 806515 62179 806518
rect 46197 806306 46263 806309
rect 41492 806304 46263 806306
rect 41492 806248 46202 806304
rect 46258 806248 46263 806304
rect 41492 806246 46263 806248
rect 46197 806243 46263 806246
rect 40902 805020 40908 805084
rect 40972 805082 40978 805084
rect 41505 805082 41571 805085
rect 40972 805080 41571 805082
rect 40972 805024 41510 805080
rect 41566 805024 41571 805080
rect 40972 805022 41571 805024
rect 40972 805020 40978 805022
rect 41505 805019 41571 805022
rect 35157 803858 35223 803861
rect 41822 803858 41828 803860
rect 35157 803856 41828 803858
rect 35157 803800 35162 803856
rect 35218 803800 41828 803856
rect 35157 803798 41828 803800
rect 35157 803795 35223 803798
rect 41822 803796 41828 803798
rect 41892 803796 41898 803860
rect 651649 803314 651715 803317
rect 650164 803312 651715 803314
rect 650164 803256 651654 803312
rect 651710 803256 651715 803312
rect 650164 803254 651715 803256
rect 651649 803251 651715 803254
rect 39757 802090 39823 802093
rect 42701 802090 42767 802093
rect 39757 802088 42767 802090
rect 39757 802032 39762 802088
rect 39818 802032 42706 802088
rect 42762 802032 42767 802088
rect 39757 802030 42767 802032
rect 39757 802027 39823 802030
rect 42701 802027 42767 802030
rect 40309 800732 40375 800733
rect 40309 800730 40356 800732
rect 40264 800728 40356 800730
rect 40264 800672 40314 800728
rect 40264 800670 40356 800672
rect 40309 800668 40356 800670
rect 40420 800668 40426 800732
rect 40585 800730 40651 800733
rect 41086 800730 41092 800732
rect 40585 800728 41092 800730
rect 40585 800672 40590 800728
rect 40646 800672 41092 800728
rect 40585 800670 41092 800672
rect 40309 800667 40375 800668
rect 40585 800667 40651 800670
rect 41086 800668 41092 800670
rect 41156 800668 41162 800732
rect 41781 800320 41847 800325
rect 41781 800264 41786 800320
rect 41842 800264 41847 800320
rect 41781 800259 41847 800264
rect 41784 799917 41844 800259
rect 41781 799912 41847 799917
rect 41781 799856 41786 799912
rect 41842 799856 41847 799912
rect 41781 799851 41847 799856
rect 42057 797330 42123 797333
rect 43621 797330 43687 797333
rect 42057 797328 43687 797330
rect 42057 797272 42062 797328
rect 42118 797272 43626 797328
rect 43682 797272 43687 797328
rect 42057 797270 43687 797272
rect 42057 797267 42123 797270
rect 43621 797267 43687 797270
rect 41086 796180 41092 796244
rect 41156 796242 41162 796244
rect 41781 796242 41847 796245
rect 41156 796240 41847 796242
rect 41156 796184 41786 796240
rect 41842 796184 41847 796240
rect 41156 796182 41847 796184
rect 41156 796180 41162 796182
rect 41781 796179 41847 796182
rect 40350 794412 40356 794476
rect 40420 794474 40426 794476
rect 41781 794474 41847 794477
rect 40420 794472 41847 794474
rect 40420 794416 41786 794472
rect 41842 794416 41847 794472
rect 40420 794414 41847 794416
rect 40420 794412 40426 794414
rect 41781 794411 41847 794414
rect 62113 793658 62179 793661
rect 62113 793656 64492 793658
rect 62113 793600 62118 793656
rect 62174 793600 64492 793656
rect 62113 793598 64492 793600
rect 62113 793595 62179 793598
rect 40902 793460 40908 793524
rect 40972 793522 40978 793524
rect 41781 793522 41847 793525
rect 40972 793520 41847 793522
rect 40972 793464 41786 793520
rect 41842 793464 41847 793520
rect 40972 793462 41847 793464
rect 40972 793460 40978 793462
rect 41781 793459 41847 793462
rect 41638 791556 41644 791620
rect 41708 791618 41714 791620
rect 42425 791618 42491 791621
rect 41708 791616 42491 791618
rect 41708 791560 42430 791616
rect 42486 791560 42491 791616
rect 41708 791558 42491 791560
rect 41708 791556 41714 791558
rect 42425 791555 42491 791558
rect 42057 790666 42123 790669
rect 42977 790666 43043 790669
rect 42057 790664 43043 790666
rect 42057 790608 42062 790664
rect 42118 790608 42982 790664
rect 43038 790608 43043 790664
rect 42057 790606 43043 790608
rect 42057 790603 42123 790606
rect 42977 790603 43043 790606
rect 40534 790196 40540 790260
rect 40604 790258 40610 790260
rect 42609 790258 42675 790261
rect 40604 790256 42675 790258
rect 40604 790200 42614 790256
rect 42670 790200 42675 790256
rect 40604 790198 42675 790200
rect 40604 790196 40610 790198
rect 42609 790195 42675 790198
rect 40718 789924 40724 789988
rect 40788 789986 40794 789988
rect 42241 789986 42307 789989
rect 651649 789986 651715 789989
rect 40788 789984 42307 789986
rect 40788 789928 42246 789984
rect 42302 789928 42307 789984
rect 40788 789926 42307 789928
rect 650164 789984 651715 789986
rect 650164 789928 651654 789984
rect 651710 789928 651715 789984
rect 650164 789926 651715 789928
rect 40788 789924 40794 789926
rect 42241 789923 42307 789926
rect 651649 789923 651715 789926
rect 41454 788156 41460 788220
rect 41524 788218 41530 788220
rect 42241 788218 42307 788221
rect 41524 788216 42307 788218
rect 41524 788160 42246 788216
rect 42302 788160 42307 788216
rect 41524 788158 42307 788160
rect 41524 788156 41530 788158
rect 42241 788155 42307 788158
rect 41822 787884 41828 787948
rect 41892 787946 41898 787948
rect 42517 787946 42583 787949
rect 41892 787944 42583 787946
rect 41892 787888 42522 787944
rect 42578 787888 42583 787944
rect 41892 787886 42583 787888
rect 41892 787884 41898 787886
rect 42517 787883 42583 787886
rect 674230 784212 674236 784276
rect 674300 784274 674306 784276
rect 675385 784274 675451 784277
rect 674300 784272 675451 784274
rect 674300 784216 675390 784272
rect 675446 784216 675451 784272
rect 674300 784214 675451 784216
rect 674300 784212 674306 784214
rect 675385 784211 675451 784214
rect 62113 780466 62179 780469
rect 62113 780464 64492 780466
rect 62113 780408 62118 780464
rect 62174 780408 64492 780464
rect 62113 780406 64492 780408
rect 62113 780403 62179 780406
rect 674925 780332 674991 780333
rect 674925 780330 674972 780332
rect 674880 780328 674972 780330
rect 674880 780272 674930 780328
rect 674880 780270 674972 780272
rect 674925 780268 674972 780270
rect 675036 780268 675042 780332
rect 674925 780267 674991 780268
rect 675150 779860 675156 779924
rect 675220 779922 675226 779924
rect 675477 779922 675543 779925
rect 675220 779920 675543 779922
rect 675220 779864 675482 779920
rect 675538 779864 675543 779920
rect 675220 779862 675543 779864
rect 675220 779860 675226 779862
rect 675477 779859 675543 779862
rect 651649 776658 651715 776661
rect 650164 776656 651715 776658
rect 650164 776600 651654 776656
rect 651710 776600 651715 776656
rect 650164 776598 651715 776600
rect 651649 776595 651715 776598
rect 674741 775434 674807 775437
rect 675150 775434 675156 775436
rect 674741 775432 675156 775434
rect 674741 775376 674746 775432
rect 674802 775376 675156 775432
rect 674741 775374 675156 775376
rect 674741 775371 674807 775374
rect 675150 775372 675156 775374
rect 675220 775372 675226 775436
rect 40033 775026 40099 775029
rect 44817 775026 44883 775029
rect 40033 775024 44883 775026
rect 40033 774968 40038 775024
rect 40094 774968 44822 775024
rect 44878 774968 44883 775024
rect 40033 774966 44883 774968
rect 40033 774963 40099 774966
rect 44817 774963 44883 774966
rect 669405 775026 669471 775029
rect 675385 775026 675451 775029
rect 669405 775024 675451 775026
rect 669405 774968 669410 775024
rect 669466 774968 675390 775024
rect 675446 774968 675451 775024
rect 669405 774966 675451 774968
rect 669405 774963 669471 774966
rect 675385 774963 675451 774966
rect 35758 774349 35818 774452
rect 35758 774344 35867 774349
rect 35758 774288 35806 774344
rect 35862 774288 35867 774344
rect 35758 774286 35867 774288
rect 35801 774283 35867 774286
rect 35758 773941 35818 774044
rect 35758 773936 35867 773941
rect 35758 773880 35806 773936
rect 35862 773880 35867 773936
rect 35758 773878 35867 773880
rect 35801 773875 35867 773878
rect 673269 773666 673335 773669
rect 675385 773666 675451 773669
rect 673269 773664 675451 773666
rect 35390 773533 35450 773636
rect 673269 773608 673274 773664
rect 673330 773608 675390 773664
rect 675446 773608 675451 773664
rect 673269 773606 675451 773608
rect 673269 773603 673335 773606
rect 675385 773603 675451 773606
rect 35341 773528 35450 773533
rect 35341 773472 35346 773528
rect 35402 773472 35450 773528
rect 35341 773470 35450 773472
rect 35341 773467 35407 773470
rect 674966 773332 674972 773396
rect 675036 773394 675042 773396
rect 675385 773394 675451 773397
rect 675036 773392 675451 773394
rect 675036 773336 675390 773392
rect 675446 773336 675451 773392
rect 675036 773334 675451 773336
rect 675036 773332 675042 773334
rect 675385 773331 675451 773334
rect 35758 773125 35818 773228
rect 35525 773122 35591 773125
rect 35525 773120 35634 773122
rect 35525 773064 35530 773120
rect 35586 773064 35634 773120
rect 35525 773059 35634 773064
rect 35758 773120 35867 773125
rect 35758 773064 35806 773120
rect 35862 773064 35867 773120
rect 35758 773062 35867 773064
rect 35801 773059 35867 773062
rect 40861 773122 40927 773125
rect 43069 773122 43135 773125
rect 40861 773120 43135 773122
rect 40861 773064 40866 773120
rect 40922 773064 43074 773120
rect 43130 773064 43135 773120
rect 40861 773062 43135 773064
rect 40861 773059 40927 773062
rect 43069 773059 43135 773062
rect 35574 772820 35634 773059
rect 674557 772714 674623 772717
rect 675845 772714 675911 772717
rect 674557 772712 675911 772714
rect 674557 772656 674562 772712
rect 674618 772656 675850 772712
rect 675906 772656 675911 772712
rect 674557 772654 675911 772656
rect 674557 772651 674623 772654
rect 675845 772651 675911 772654
rect 676070 772652 676076 772716
rect 676140 772714 676146 772716
rect 679617 772714 679683 772717
rect 676140 772712 679683 772714
rect 676140 772656 679622 772712
rect 679678 772656 679683 772712
rect 676140 772654 679683 772656
rect 676140 772652 676146 772654
rect 679617 772651 679683 772654
rect 35390 772309 35450 772412
rect 673862 772380 673868 772444
rect 673932 772442 673938 772444
rect 683389 772442 683455 772445
rect 673932 772440 683455 772442
rect 673932 772384 683394 772440
rect 683450 772384 683455 772440
rect 673932 772382 683455 772384
rect 673932 772380 673938 772382
rect 683389 772379 683455 772382
rect 35341 772304 35450 772309
rect 35341 772248 35346 772304
rect 35402 772248 35450 772304
rect 35341 772246 35450 772248
rect 39757 772306 39823 772309
rect 42793 772306 42859 772309
rect 39757 772304 42859 772306
rect 39757 772248 39762 772304
rect 39818 772248 42798 772304
rect 42854 772248 42859 772304
rect 39757 772246 42859 772248
rect 35341 772243 35407 772246
rect 39757 772243 39823 772246
rect 42793 772243 42859 772246
rect 35574 771901 35634 772004
rect 674414 771972 674420 772036
rect 674484 772034 674490 772036
rect 684033 772034 684099 772037
rect 674484 772032 684099 772034
rect 674484 771976 684038 772032
rect 684094 771976 684099 772032
rect 674484 771974 684099 771976
rect 674484 771972 674490 771974
rect 684033 771971 684099 771974
rect 35525 771896 35634 771901
rect 35525 771840 35530 771896
rect 35586 771840 35634 771896
rect 35525 771838 35634 771840
rect 35525 771835 35591 771838
rect 675109 771762 675175 771765
rect 675845 771762 675911 771765
rect 675109 771760 675911 771762
rect 675109 771704 675114 771760
rect 675170 771704 675850 771760
rect 675906 771704 675911 771760
rect 675109 771702 675911 771704
rect 675109 771699 675175 771702
rect 675845 771699 675911 771702
rect 35758 771493 35818 771596
rect 35709 771488 35818 771493
rect 35709 771432 35714 771488
rect 35770 771432 35818 771488
rect 35709 771430 35818 771432
rect 39113 771490 39179 771493
rect 44173 771490 44239 771493
rect 39113 771488 44239 771490
rect 39113 771432 39118 771488
rect 39174 771432 44178 771488
rect 44234 771432 44239 771488
rect 39113 771430 44239 771432
rect 35709 771427 35775 771430
rect 39113 771427 39179 771430
rect 44173 771427 44239 771430
rect 675886 771292 675892 771356
rect 675956 771354 675962 771356
rect 682377 771354 682443 771357
rect 675956 771352 682443 771354
rect 675956 771296 682382 771352
rect 682438 771296 682443 771352
rect 675956 771294 682443 771296
rect 675956 771292 675962 771294
rect 682377 771291 682443 771294
rect 35390 771085 35450 771188
rect 35390 771080 35499 771085
rect 35390 771024 35438 771080
rect 35494 771024 35499 771080
rect 35390 771022 35499 771024
rect 35433 771019 35499 771022
rect 39849 771082 39915 771085
rect 42885 771082 42951 771085
rect 39849 771080 42951 771082
rect 39849 771024 39854 771080
rect 39910 771024 42890 771080
rect 42946 771024 42951 771080
rect 39849 771022 42951 771024
rect 39849 771019 39915 771022
rect 42885 771019 42951 771022
rect 35574 770677 35634 770780
rect 35574 770672 35683 770677
rect 35574 770616 35622 770672
rect 35678 770616 35683 770672
rect 35574 770614 35683 770616
rect 35617 770611 35683 770614
rect 35758 770269 35818 770372
rect 35758 770264 35867 770269
rect 35758 770208 35806 770264
rect 35862 770208 35867 770264
rect 35758 770206 35867 770208
rect 35801 770203 35867 770206
rect 41413 770266 41479 770269
rect 44265 770266 44331 770269
rect 41413 770264 44331 770266
rect 41413 770208 41418 770264
rect 41474 770208 44270 770264
rect 44326 770208 44331 770264
rect 41413 770206 44331 770208
rect 41413 770203 41479 770206
rect 44265 770203 44331 770206
rect 41462 769860 41522 769964
rect 41454 769796 41460 769860
rect 41524 769796 41530 769860
rect 35390 769453 35450 769556
rect 35341 769448 35450 769453
rect 35341 769392 35346 769448
rect 35402 769392 35450 769448
rect 35341 769390 35450 769392
rect 35341 769387 35407 769390
rect 35574 769045 35634 769148
rect 35525 769040 35634 769045
rect 35801 769042 35867 769045
rect 35525 768984 35530 769040
rect 35586 768984 35634 769040
rect 35525 768982 35634 768984
rect 35758 769040 35867 769042
rect 35758 768984 35806 769040
rect 35862 768984 35867 769040
rect 35525 768979 35591 768982
rect 35758 768979 35867 768984
rect 35758 768740 35818 768979
rect 39849 768634 39915 768637
rect 42701 768634 42767 768637
rect 39849 768632 42767 768634
rect 39849 768576 39854 768632
rect 39910 768576 42706 768632
rect 42762 768576 42767 768632
rect 39849 768574 42767 768576
rect 39849 768571 39915 768574
rect 42701 768571 42767 768574
rect 42241 768362 42307 768365
rect 41492 768360 42307 768362
rect 41492 768304 42246 768360
rect 42302 768304 42307 768360
rect 41492 768302 42307 768304
rect 42241 768299 42307 768302
rect 35758 767821 35818 767924
rect 35758 767816 35867 767821
rect 35758 767760 35806 767816
rect 35862 767760 35867 767816
rect 35758 767758 35867 767760
rect 35801 767755 35867 767758
rect 32446 767413 32506 767516
rect 32397 767408 32506 767413
rect 32397 767352 32402 767408
rect 32458 767352 32506 767408
rect 32397 767350 32506 767352
rect 62113 767410 62179 767413
rect 62113 767408 64492 767410
rect 62113 767352 62118 767408
rect 62174 767352 64492 767408
rect 62113 767350 64492 767352
rect 32397 767347 32463 767350
rect 62113 767347 62179 767350
rect 35206 767005 35266 767108
rect 35157 767000 35266 767005
rect 35157 766944 35162 767000
rect 35218 766944 35266 767000
rect 35157 766942 35266 766944
rect 35157 766939 35223 766942
rect 35758 766597 35818 766700
rect 35758 766592 35867 766597
rect 35758 766536 35806 766592
rect 35862 766536 35867 766592
rect 35758 766534 35867 766536
rect 35801 766531 35867 766534
rect 35758 766189 35818 766292
rect 35758 766184 35867 766189
rect 35758 766128 35806 766184
rect 35862 766128 35867 766184
rect 35758 766126 35867 766128
rect 35801 766123 35867 766126
rect 40401 766186 40467 766189
rect 43253 766186 43319 766189
rect 40401 766184 43319 766186
rect 40401 766128 40406 766184
rect 40462 766128 43258 766184
rect 43314 766128 43319 766184
rect 40401 766126 43319 766128
rect 40401 766123 40467 766126
rect 43253 766123 43319 766126
rect 40910 765780 40970 765884
rect 40902 765716 40908 765780
rect 40972 765716 40978 765780
rect 40542 765372 40602 765476
rect 40534 765308 40540 765372
rect 40604 765308 40610 765372
rect 40726 764964 40786 765068
rect 40718 764900 40724 764964
rect 40788 764900 40794 764964
rect 35758 764557 35818 764660
rect 35758 764552 35867 764557
rect 35758 764496 35806 764552
rect 35862 764496 35867 764552
rect 35758 764494 35867 764496
rect 35801 764491 35867 764494
rect 40401 764554 40467 764557
rect 45185 764554 45251 764557
rect 40401 764552 45251 764554
rect 40401 764496 40406 764552
rect 40462 764496 45190 764552
rect 45246 764496 45251 764552
rect 40401 764494 45251 764496
rect 40401 764491 40467 764494
rect 45185 764491 45251 764494
rect 35574 764149 35634 764252
rect 35574 764144 35683 764149
rect 35574 764088 35622 764144
rect 35678 764088 35683 764144
rect 35574 764086 35683 764088
rect 35617 764083 35683 764086
rect 35758 763741 35818 763844
rect 35758 763736 35867 763741
rect 35758 763680 35806 763736
rect 35862 763680 35867 763736
rect 35758 763675 35867 763680
rect 35758 763436 35818 763675
rect 41505 763330 41571 763333
rect 47577 763330 47643 763333
rect 651649 763330 651715 763333
rect 41505 763328 47643 763330
rect 41505 763272 41510 763328
rect 41566 763272 47582 763328
rect 47638 763272 47643 763328
rect 41505 763270 47643 763272
rect 650164 763328 651715 763330
rect 650164 763272 651654 763328
rect 651710 763272 651715 763328
rect 650164 763270 651715 763272
rect 41505 763267 41571 763270
rect 47577 763267 47643 763270
rect 651649 763267 651715 763270
rect 35758 762925 35818 763028
rect 35758 762920 35867 762925
rect 35758 762864 35806 762920
rect 35862 762864 35867 762920
rect 35758 762862 35867 762864
rect 35801 762859 35867 762862
rect 676949 761836 677015 761837
rect 676949 761832 676996 761836
rect 677060 761834 677066 761836
rect 676949 761776 676954 761832
rect 676949 761772 676996 761776
rect 677060 761774 677106 761834
rect 677060 761772 677066 761774
rect 676949 761771 677015 761772
rect 675477 761562 675543 761565
rect 675477 761560 676292 761562
rect 675477 761504 675482 761560
rect 675538 761504 676292 761560
rect 675477 761502 676292 761504
rect 675477 761499 675543 761502
rect 675293 761154 675359 761157
rect 675293 761152 676292 761154
rect 675293 761096 675298 761152
rect 675354 761096 676292 761152
rect 675293 761094 676292 761096
rect 675293 761091 675359 761094
rect 675477 760746 675543 760749
rect 675477 760744 676292 760746
rect 675477 760688 675482 760744
rect 675538 760688 676292 760744
rect 675477 760686 676292 760688
rect 675477 760683 675543 760686
rect 40493 760338 40559 760341
rect 44817 760338 44883 760341
rect 40493 760336 44883 760338
rect 40493 760280 40498 760336
rect 40554 760280 44822 760336
rect 44878 760280 44883 760336
rect 40493 760278 44883 760280
rect 40493 760275 40559 760278
rect 44817 760275 44883 760278
rect 675477 760338 675543 760341
rect 675477 760336 676292 760338
rect 675477 760280 675482 760336
rect 675538 760280 676292 760336
rect 675477 760278 676292 760280
rect 675477 760275 675543 760278
rect 675477 759930 675543 759933
rect 675477 759928 676292 759930
rect 675477 759872 675482 759928
rect 675538 759872 676292 759928
rect 675477 759870 676292 759872
rect 675477 759867 675543 759870
rect 32397 759658 32463 759661
rect 41822 759658 41828 759660
rect 32397 759656 41828 759658
rect 32397 759600 32402 759656
rect 32458 759600 41828 759656
rect 32397 759598 41828 759600
rect 32397 759595 32463 759598
rect 41822 759596 41828 759598
rect 41892 759596 41898 759660
rect 675477 759522 675543 759525
rect 675477 759520 676292 759522
rect 675477 759464 675482 759520
rect 675538 759464 676292 759520
rect 675477 759462 676292 759464
rect 675477 759459 675543 759462
rect 675477 759114 675543 759117
rect 675477 759112 676292 759114
rect 675477 759056 675482 759112
rect 675538 759056 676292 759112
rect 675477 759054 676292 759056
rect 675477 759051 675543 759054
rect 675477 758706 675543 758709
rect 675477 758704 676292 758706
rect 675477 758648 675482 758704
rect 675538 758648 676292 758704
rect 675477 758646 676292 758648
rect 675477 758643 675543 758646
rect 40401 758298 40467 758301
rect 42425 758298 42491 758301
rect 40401 758296 42491 758298
rect 40401 758240 40406 758296
rect 40462 758240 42430 758296
rect 42486 758240 42491 758296
rect 40401 758238 42491 758240
rect 40401 758235 40467 758238
rect 42425 758235 42491 758238
rect 675477 758298 675543 758301
rect 675477 758296 676292 758298
rect 675477 758240 675482 758296
rect 675538 758240 676292 758296
rect 675477 758238 676292 758240
rect 675477 758235 675543 758238
rect 675293 757890 675359 757893
rect 675293 757888 676292 757890
rect 675293 757832 675298 757888
rect 675354 757832 676292 757888
rect 675293 757830 676292 757832
rect 675293 757827 675359 757830
rect 39297 757754 39363 757757
rect 41638 757754 41644 757756
rect 39297 757752 41644 757754
rect 39297 757696 39302 757752
rect 39358 757696 41644 757752
rect 39297 757694 41644 757696
rect 39297 757691 39363 757694
rect 41638 757692 41644 757694
rect 41708 757692 41714 757756
rect 675477 757482 675543 757485
rect 675477 757480 676292 757482
rect 675477 757424 675482 757480
rect 675538 757424 676292 757480
rect 675477 757422 676292 757424
rect 675477 757419 675543 757422
rect 41413 757346 41479 757349
rect 41413 757344 41522 757346
rect 41413 757288 41418 757344
rect 41474 757288 41522 757344
rect 41413 757283 41522 757288
rect 41462 756666 41522 757283
rect 676949 757074 677015 757077
rect 676949 757072 677028 757074
rect 676949 757016 676954 757072
rect 677010 757016 677028 757072
rect 676949 757014 677028 757016
rect 676949 757011 677015 757014
rect 41781 756666 41847 756669
rect 41462 756664 41847 756666
rect 41462 756608 41786 756664
rect 41842 756608 41847 756664
rect 41462 756606 41847 756608
rect 41781 756603 41847 756606
rect 680997 756666 681063 756669
rect 680997 756664 681076 756666
rect 680997 756608 681002 756664
rect 681058 756608 681076 756664
rect 680997 756606 681076 756608
rect 680997 756603 681063 756606
rect 679617 756258 679683 756261
rect 679604 756256 679683 756258
rect 679604 756200 679622 756256
rect 679678 756200 679683 756256
rect 679604 756198 679683 756200
rect 679617 756195 679683 756198
rect 675845 755850 675911 755853
rect 675845 755848 676292 755850
rect 675845 755792 675850 755848
rect 675906 755792 676292 755848
rect 675845 755790 676292 755792
rect 675845 755787 675911 755790
rect 682377 755442 682443 755445
rect 682364 755440 682443 755442
rect 682364 755384 682382 755440
rect 682438 755384 682443 755440
rect 682364 755382 682443 755384
rect 682377 755379 682443 755382
rect 675477 755034 675543 755037
rect 675477 755032 676292 755034
rect 675477 754976 675482 755032
rect 675538 754976 676292 755032
rect 675477 754974 676292 754976
rect 675477 754971 675543 754974
rect 675477 754626 675543 754629
rect 675477 754624 676292 754626
rect 675477 754568 675482 754624
rect 675538 754568 676292 754624
rect 675477 754566 676292 754568
rect 675477 754563 675543 754566
rect 62113 754354 62179 754357
rect 62113 754352 64492 754354
rect 62113 754296 62118 754352
rect 62174 754296 64492 754352
rect 62113 754294 64492 754296
rect 62113 754291 62179 754294
rect 684033 754218 684099 754221
rect 684020 754216 684099 754218
rect 684020 754160 684038 754216
rect 684094 754160 684099 754216
rect 684020 754158 684099 754160
rect 684033 754155 684099 754158
rect 42057 754082 42123 754085
rect 43437 754082 43503 754085
rect 42057 754080 43503 754082
rect 42057 754024 42062 754080
rect 42118 754024 43442 754080
rect 43498 754024 43503 754080
rect 42057 754022 43503 754024
rect 42057 754019 42123 754022
rect 43437 754019 43503 754022
rect 675886 753748 675892 753812
rect 675956 753810 675962 753812
rect 675956 753750 676292 753810
rect 675956 753748 675962 753750
rect 675477 753402 675543 753405
rect 675477 753400 676292 753402
rect 675477 753344 675482 753400
rect 675538 753344 676292 753400
rect 675477 753342 676292 753344
rect 675477 753339 675543 753342
rect 42057 752994 42123 752997
rect 43805 752994 43871 752997
rect 42057 752992 43871 752994
rect 42057 752936 42062 752992
rect 42118 752936 43810 752992
rect 43866 752936 43871 752992
rect 42057 752934 43871 752936
rect 42057 752931 42123 752934
rect 43805 752931 43871 752934
rect 675477 752994 675543 752997
rect 675477 752992 676292 752994
rect 675477 752936 675482 752992
rect 675538 752936 676292 752992
rect 675477 752934 676292 752936
rect 675477 752931 675543 752934
rect 683389 752586 683455 752589
rect 683389 752584 683468 752586
rect 683389 752528 683394 752584
rect 683450 752528 683468 752584
rect 683389 752526 683468 752528
rect 683389 752523 683455 752526
rect 672993 752314 673059 752317
rect 675845 752314 675911 752317
rect 672993 752312 675911 752314
rect 672993 752256 672998 752312
rect 673054 752256 675850 752312
rect 675906 752256 675911 752312
rect 672993 752254 675911 752256
rect 672993 752251 673059 752254
rect 675845 752251 675911 752254
rect 683205 752178 683271 752181
rect 683205 752176 683284 752178
rect 683205 752120 683210 752176
rect 683266 752120 683284 752176
rect 683205 752118 683284 752120
rect 683205 752115 683271 752118
rect 675477 751770 675543 751773
rect 675477 751768 676292 751770
rect 675477 751712 675482 751768
rect 675538 751712 676292 751768
rect 675477 751710 676292 751712
rect 675477 751707 675543 751710
rect 42241 751636 42307 751637
rect 42190 751572 42196 751636
rect 42260 751634 42307 751636
rect 42260 751632 42352 751634
rect 42302 751576 42352 751632
rect 42260 751574 42352 751576
rect 42260 751572 42307 751574
rect 42241 751571 42307 751572
rect 675477 751362 675543 751365
rect 675477 751360 676292 751362
rect 675477 751304 675482 751360
rect 675538 751304 676292 751360
rect 675477 751302 676292 751304
rect 675477 751299 675543 751302
rect 40902 751028 40908 751092
rect 40972 751090 40978 751092
rect 41781 751090 41847 751093
rect 40972 751088 41847 751090
rect 40972 751032 41786 751088
rect 41842 751032 41847 751088
rect 40972 751030 41847 751032
rect 40972 751028 40978 751030
rect 41781 751027 41847 751030
rect 674925 751090 674991 751093
rect 676070 751090 676076 751092
rect 674925 751088 676076 751090
rect 674925 751032 674930 751088
rect 674986 751032 676076 751088
rect 674925 751030 676076 751032
rect 674925 751027 674991 751030
rect 676070 751028 676076 751030
rect 676140 751028 676146 751092
rect 683070 750753 683130 750924
rect 683070 750748 683179 750753
rect 683070 750692 683118 750748
rect 683174 750692 683179 750748
rect 683070 750687 683179 750692
rect 42190 750484 42196 750548
rect 42260 750546 42266 750548
rect 42609 750546 42675 750549
rect 42260 750544 42675 750546
rect 42260 750488 42614 750544
rect 42670 750488 42675 750544
rect 683070 750516 683130 750687
rect 42260 750486 42675 750488
rect 42260 750484 42266 750486
rect 42609 750483 42675 750486
rect 40718 750348 40724 750412
rect 40788 750410 40794 750412
rect 41781 750410 41847 750413
rect 40788 750408 41847 750410
rect 40788 750352 41786 750408
rect 41842 750352 41847 750408
rect 40788 750350 41847 750352
rect 40788 750348 40794 750350
rect 41781 750347 41847 750350
rect 652017 750138 652083 750141
rect 650164 750136 652083 750138
rect 650164 750080 652022 750136
rect 652078 750080 652083 750136
rect 650164 750078 652083 750080
rect 652017 750075 652083 750078
rect 675477 750138 675543 750141
rect 675477 750136 676292 750138
rect 675477 750080 675482 750136
rect 675538 750080 676292 750136
rect 675477 750078 676292 750080
rect 675477 750075 675543 750078
rect 40534 749396 40540 749460
rect 40604 749458 40610 749460
rect 42425 749458 42491 749461
rect 40604 749456 42491 749458
rect 40604 749400 42430 749456
rect 42486 749400 42491 749456
rect 40604 749398 42491 749400
rect 40604 749396 40610 749398
rect 42425 749395 42491 749398
rect 41822 745588 41828 745652
rect 41892 745650 41898 745652
rect 42241 745650 42307 745653
rect 41892 745648 42307 745650
rect 41892 745592 42246 745648
rect 42302 745592 42307 745648
rect 41892 745590 42307 745592
rect 41892 745588 41898 745590
rect 42241 745587 42307 745590
rect 41638 745044 41644 745108
rect 41708 745106 41714 745108
rect 42425 745106 42491 745109
rect 41708 745104 42491 745106
rect 41708 745048 42430 745104
rect 42486 745048 42491 745104
rect 41708 745046 42491 745048
rect 41708 745044 41714 745046
rect 42425 745043 42491 745046
rect 41454 743684 41460 743748
rect 41524 743746 41530 743748
rect 41781 743746 41847 743749
rect 41524 743744 41847 743746
rect 41524 743688 41786 743744
rect 41842 743688 41847 743744
rect 41524 743686 41847 743688
rect 41524 743684 41530 743686
rect 41781 743683 41847 743686
rect 675569 743068 675635 743069
rect 675518 743066 675524 743068
rect 675478 743006 675524 743066
rect 675588 743064 675635 743068
rect 675630 743008 675635 743064
rect 675518 743004 675524 743006
rect 675588 743004 675635 743008
rect 675569 743003 675635 743004
rect 62113 741298 62179 741301
rect 62113 741296 64492 741298
rect 62113 741240 62118 741296
rect 62174 741240 64492 741296
rect 62113 741238 64492 741240
rect 62113 741235 62179 741238
rect 674414 738652 674420 738716
rect 674484 738714 674490 738716
rect 675385 738714 675451 738717
rect 674484 738712 675451 738714
rect 674484 738656 675390 738712
rect 675446 738656 675451 738712
rect 674484 738654 675451 738656
rect 674484 738652 674490 738654
rect 675385 738651 675451 738654
rect 674598 738108 674604 738172
rect 674668 738170 674674 738172
rect 675109 738170 675175 738173
rect 674668 738168 675175 738170
rect 674668 738112 675114 738168
rect 675170 738112 675175 738168
rect 674668 738110 675175 738112
rect 674668 738108 674674 738110
rect 675109 738107 675175 738110
rect 651649 736810 651715 736813
rect 650164 736808 651715 736810
rect 650164 736752 651654 736808
rect 651710 736752 651715 736808
rect 650164 736750 651715 736752
rect 651649 736747 651715 736750
rect 669589 735178 669655 735181
rect 675334 735178 675340 735180
rect 669589 735176 675340 735178
rect 669589 735120 669594 735176
rect 669650 735120 675340 735176
rect 669589 735118 675340 735120
rect 669589 735115 669655 735118
rect 675334 735116 675340 735118
rect 675404 735116 675410 735180
rect 673453 734906 673519 734909
rect 675477 734906 675543 734909
rect 673453 734904 675543 734906
rect 673453 734848 673458 734904
rect 673514 734848 675482 734904
rect 675538 734848 675543 734904
rect 673453 734846 675543 734848
rect 673453 734843 673519 734846
rect 675477 734843 675543 734846
rect 670417 734498 670483 734501
rect 675477 734498 675543 734501
rect 670417 734496 675543 734498
rect 670417 734440 670422 734496
rect 670478 734440 675482 734496
rect 675538 734440 675543 734496
rect 670417 734438 675543 734440
rect 670417 734435 670483 734438
rect 675477 734435 675543 734438
rect 671245 734226 671311 734229
rect 675477 734226 675543 734229
rect 671245 734224 675543 734226
rect 671245 734168 671250 734224
rect 671306 734168 675482 734224
rect 675538 734168 675543 734224
rect 671245 734166 675543 734168
rect 671245 734163 671311 734166
rect 675477 734163 675543 734166
rect 675293 733682 675359 733685
rect 676806 733682 676812 733684
rect 675293 733680 676812 733682
rect 675293 733624 675298 733680
rect 675354 733624 676812 733680
rect 675293 733622 676812 733624
rect 675293 733619 675359 733622
rect 676806 733620 676812 733622
rect 676876 733620 676882 733684
rect 673821 732730 673887 732733
rect 675385 732730 675451 732733
rect 673821 732728 675451 732730
rect 673821 732672 673826 732728
rect 673882 732672 675390 732728
rect 675446 732672 675451 732728
rect 673821 732670 675451 732672
rect 673821 732667 673887 732670
rect 675385 732667 675451 732670
rect 47761 731370 47827 731373
rect 41492 731368 47827 731370
rect 41492 731312 47766 731368
rect 47822 731312 47827 731368
rect 41492 731310 47827 731312
rect 47761 731307 47827 731310
rect 42425 730962 42491 730965
rect 41492 730960 42491 730962
rect 41492 730904 42430 730960
rect 42486 730904 42491 730960
rect 41492 730902 42491 730904
rect 42425 730899 42491 730902
rect 41137 730554 41203 730557
rect 41124 730552 41203 730554
rect 41124 730496 41142 730552
rect 41198 730496 41203 730552
rect 41124 730494 41203 730496
rect 41137 730491 41203 730494
rect 43069 730146 43135 730149
rect 41492 730144 43135 730146
rect 41492 730088 43074 730144
rect 43130 730088 43135 730144
rect 41492 730086 43135 730088
rect 43069 730083 43135 730086
rect 672809 730146 672875 730149
rect 675385 730146 675451 730149
rect 672809 730144 675451 730146
rect 672809 730088 672814 730144
rect 672870 730088 675390 730144
rect 675446 730088 675451 730144
rect 672809 730086 675451 730088
rect 672809 730083 672875 730086
rect 675385 730083 675451 730086
rect 45001 729738 45067 729741
rect 41492 729736 45067 729738
rect 41492 729680 45006 729736
rect 45062 729680 45067 729736
rect 41492 729678 45067 729680
rect 45001 729675 45067 729678
rect 42885 729330 42951 729333
rect 41492 729328 42951 729330
rect 41492 729272 42890 729328
rect 42946 729272 42951 729328
rect 41492 729270 42951 729272
rect 42885 729267 42951 729270
rect 45185 728922 45251 728925
rect 41492 728920 45251 728922
rect 41492 728864 45190 728920
rect 45246 728864 45251 728920
rect 41492 728862 45251 728864
rect 45185 728859 45251 728862
rect 668577 728786 668643 728789
rect 675385 728786 675451 728789
rect 668577 728784 675451 728786
rect 668577 728728 668582 728784
rect 668638 728728 675390 728784
rect 675446 728728 675451 728784
rect 668577 728726 675451 728728
rect 668577 728723 668643 728726
rect 675385 728723 675451 728726
rect 40861 728684 40927 728687
rect 40861 728682 40970 728684
rect 40861 728626 40866 728682
rect 40922 728626 40970 728682
rect 40861 728621 40970 728626
rect 40910 728484 40970 728621
rect 62113 728242 62179 728245
rect 62113 728240 64492 728242
rect 62113 728184 62118 728240
rect 62174 728184 64492 728240
rect 62113 728182 64492 728184
rect 62113 728179 62179 728182
rect 43069 728106 43135 728109
rect 41492 728104 43135 728106
rect 41492 728048 43074 728104
rect 43130 728048 43135 728104
rect 41492 728046 43135 728048
rect 43069 728043 43135 728046
rect 674557 728106 674623 728109
rect 676029 728106 676095 728109
rect 674557 728104 676095 728106
rect 674557 728048 674562 728104
rect 674618 728048 676034 728104
rect 676090 728048 676095 728104
rect 674557 728046 676095 728048
rect 674557 728043 674623 728046
rect 676029 728043 676095 728046
rect 41278 727463 41338 727668
rect 41045 727460 41111 727463
rect 41045 727458 41154 727460
rect 41045 727402 41050 727458
rect 41106 727402 41154 727458
rect 41045 727397 41154 727402
rect 41278 727458 41387 727463
rect 41278 727402 41326 727458
rect 41382 727402 41387 727458
rect 41278 727400 41387 727402
rect 41321 727397 41387 727400
rect 41094 727260 41154 727397
rect 41137 726882 41203 726885
rect 41124 726880 41203 726882
rect 41124 726824 41142 726880
rect 41198 726824 41203 726880
rect 41124 726822 41203 726824
rect 41137 726819 41203 726822
rect 41278 726239 41338 726444
rect 40953 726236 41019 726239
rect 40910 726234 41019 726236
rect 40910 726178 40958 726234
rect 41014 726178 41019 726234
rect 40910 726173 41019 726178
rect 41278 726234 41387 726239
rect 41278 726178 41326 726234
rect 41382 726178 41387 726234
rect 41278 726176 41387 726178
rect 41321 726173 41387 726176
rect 40910 726036 40970 726173
rect 673637 725930 673703 725933
rect 674598 725930 674604 725932
rect 673637 725928 674604 725930
rect 673637 725872 673642 725928
rect 673698 725872 674604 725928
rect 673637 725870 674604 725872
rect 673637 725867 673703 725870
rect 674598 725868 674604 725870
rect 674668 725868 674674 725932
rect 41781 725796 41847 725797
rect 41781 725794 41828 725796
rect 41736 725792 41828 725794
rect 41736 725736 41786 725792
rect 41736 725734 41828 725736
rect 41781 725732 41828 725734
rect 41892 725732 41898 725796
rect 41781 725731 41847 725732
rect 41321 725658 41387 725661
rect 41308 725656 41387 725658
rect 41308 725600 41326 725656
rect 41382 725600 41387 725656
rect 41308 725598 41387 725600
rect 41321 725595 41387 725598
rect 37917 725250 37983 725253
rect 37917 725248 37996 725250
rect 37917 725192 37922 725248
rect 37978 725192 37996 725248
rect 37917 725190 37996 725192
rect 37917 725187 37983 725190
rect 35157 724842 35223 724845
rect 35157 724840 35236 724842
rect 35157 724784 35162 724840
rect 35218 724784 35236 724840
rect 35157 724782 35236 724784
rect 35157 724779 35223 724782
rect 33041 724434 33107 724437
rect 33028 724432 33107 724434
rect 33028 724376 33046 724432
rect 33102 724376 33107 724432
rect 33028 724374 33107 724376
rect 33041 724371 33107 724374
rect 33734 723791 33794 723996
rect 33734 723786 33843 723791
rect 33734 723730 33782 723786
rect 33838 723730 33843 723786
rect 33734 723728 33843 723730
rect 33777 723725 33843 723728
rect 43253 723618 43319 723621
rect 41492 723616 43319 723618
rect 41492 723560 43258 723616
rect 43314 723560 43319 723616
rect 41492 723558 43319 723560
rect 43253 723555 43319 723558
rect 651649 723482 651715 723485
rect 650164 723480 651715 723482
rect 650164 723424 651654 723480
rect 651710 723424 651715 723480
rect 650164 723422 651715 723424
rect 651649 723419 651715 723422
rect 40677 723210 40743 723213
rect 674281 723210 674347 723213
rect 675845 723210 675911 723213
rect 40677 723208 40756 723210
rect 40677 723152 40682 723208
rect 40738 723152 40756 723208
rect 40677 723150 40756 723152
rect 674281 723208 675911 723210
rect 674281 723152 674286 723208
rect 674342 723152 675850 723208
rect 675906 723152 675911 723208
rect 674281 723150 675911 723152
rect 40677 723147 40743 723150
rect 674281 723147 674347 723150
rect 675845 723147 675911 723150
rect 44357 722802 44423 722805
rect 41492 722800 44423 722802
rect 41492 722744 44362 722800
rect 44418 722744 44423 722800
rect 41492 722742 44423 722744
rect 44357 722739 44423 722742
rect 41781 722394 41847 722397
rect 41492 722392 41847 722394
rect 41492 722336 41786 722392
rect 41842 722336 41847 722392
rect 41492 722334 41847 722336
rect 41781 722331 41847 722334
rect 40726 721772 40786 721956
rect 40718 721708 40724 721772
rect 40788 721708 40794 721772
rect 40902 721708 40908 721772
rect 40972 721708 40978 721772
rect 41137 721770 41203 721773
rect 41638 721770 41644 721772
rect 41137 721768 41644 721770
rect 41137 721712 41142 721768
rect 41198 721712 41644 721768
rect 41137 721710 41644 721712
rect 40910 721548 40970 721708
rect 41137 721707 41203 721710
rect 41638 721708 41644 721710
rect 41708 721708 41714 721772
rect 675201 721578 675267 721581
rect 676070 721578 676076 721580
rect 675201 721576 676076 721578
rect 675201 721520 675206 721576
rect 675262 721520 676076 721576
rect 675201 721518 676076 721520
rect 675201 721515 675267 721518
rect 676070 721516 676076 721518
rect 676140 721516 676146 721580
rect 46381 721170 46447 721173
rect 41492 721168 46447 721170
rect 41492 721112 46386 721168
rect 46442 721112 46447 721168
rect 41492 721110 46447 721112
rect 46381 721107 46447 721110
rect 31710 720357 31770 720732
rect 31710 720352 31819 720357
rect 31710 720324 31758 720352
rect 31740 720296 31758 720324
rect 31814 720296 31819 720352
rect 31740 720294 31819 720296
rect 31753 720291 31819 720294
rect 43437 719946 43503 719949
rect 41492 719944 43503 719946
rect 41492 719888 43442 719944
rect 43498 719888 43503 719944
rect 41492 719886 43503 719888
rect 43437 719883 43503 719886
rect 40534 718524 40540 718588
rect 40604 718586 40610 718588
rect 41781 718586 41847 718589
rect 40604 718584 41847 718586
rect 40604 718528 41786 718584
rect 41842 718528 41847 718584
rect 40604 718526 41847 718528
rect 40604 718524 40610 718526
rect 41781 718523 41847 718526
rect 33041 716818 33107 716821
rect 41822 716818 41828 716820
rect 33041 716816 41828 716818
rect 33041 716760 33046 716816
rect 33102 716760 41828 716816
rect 33041 716758 41828 716760
rect 33041 716755 33107 716758
rect 41822 716756 41828 716758
rect 41892 716756 41898 716820
rect 675477 716546 675543 716549
rect 675477 716544 676292 716546
rect 675477 716488 675482 716544
rect 675538 716488 676292 716544
rect 675477 716486 676292 716488
rect 675477 716483 675543 716486
rect 675293 716138 675359 716141
rect 675293 716136 676292 716138
rect 675293 716080 675298 716136
rect 675354 716080 676292 716136
rect 675293 716078 676292 716080
rect 675293 716075 675359 716078
rect 675477 715730 675543 715733
rect 675477 715728 676292 715730
rect 675477 715672 675482 715728
rect 675538 715672 676292 715728
rect 675477 715670 676292 715672
rect 675477 715667 675543 715670
rect 62113 715322 62179 715325
rect 674833 715322 674899 715325
rect 62113 715320 64492 715322
rect 62113 715264 62118 715320
rect 62174 715264 64492 715320
rect 62113 715262 64492 715264
rect 674833 715320 676292 715322
rect 674833 715264 674838 715320
rect 674894 715264 676292 715320
rect 674833 715262 676292 715264
rect 62113 715259 62179 715262
rect 674833 715259 674899 715262
rect 39205 715186 39271 715189
rect 42333 715186 42399 715189
rect 39205 715184 42399 715186
rect 39205 715128 39210 715184
rect 39266 715128 42338 715184
rect 42394 715128 42399 715184
rect 39205 715126 42399 715128
rect 39205 715123 39271 715126
rect 42333 715123 42399 715126
rect 42517 715186 42583 715189
rect 42517 715184 42626 715186
rect 42517 715128 42522 715184
rect 42578 715128 42626 715184
rect 42517 715123 42626 715128
rect 42566 714780 42626 715123
rect 675477 714914 675543 714917
rect 675477 714912 676292 714914
rect 675477 714856 675482 714912
rect 675538 714856 676292 714912
rect 675477 714854 676292 714856
rect 675477 714851 675543 714854
rect 42558 714716 42564 714780
rect 42628 714716 42634 714780
rect 41321 714506 41387 714509
rect 42517 714506 42583 714509
rect 41321 714504 42583 714506
rect 41321 714448 41326 714504
rect 41382 714448 42522 714504
rect 42578 714448 42583 714504
rect 41321 714446 42583 714448
rect 41321 714443 41387 714446
rect 42517 714443 42583 714446
rect 675477 714506 675543 714509
rect 675477 714504 676292 714506
rect 675477 714448 675482 714504
rect 675538 714448 676292 714504
rect 675477 714446 676292 714448
rect 675477 714443 675543 714446
rect 40033 714234 40099 714237
rect 40350 714234 40356 714236
rect 40033 714232 40356 714234
rect 40033 714176 40038 714232
rect 40094 714176 40356 714232
rect 40033 714174 40356 714176
rect 40033 714171 40099 714174
rect 40350 714172 40356 714174
rect 40420 714172 40426 714236
rect 41505 714234 41571 714237
rect 42374 714234 42380 714236
rect 41505 714232 42380 714234
rect 41505 714176 41510 714232
rect 41566 714176 42380 714232
rect 41505 714174 42380 714176
rect 41505 714171 41571 714174
rect 42374 714172 42380 714174
rect 42444 714172 42450 714236
rect 675477 714098 675543 714101
rect 675477 714096 676292 714098
rect 675477 714040 675482 714096
rect 675538 714040 676292 714096
rect 675477 714038 676292 714040
rect 675477 714035 675543 714038
rect 41781 713962 41847 713965
rect 42006 713962 42012 713964
rect 41781 713960 42012 713962
rect 41781 713904 41786 713960
rect 41842 713904 42012 713960
rect 41781 713902 42012 713904
rect 41781 713899 41847 713902
rect 42006 713900 42012 713902
rect 42076 713900 42082 713964
rect 675477 713690 675543 713693
rect 675477 713688 676292 713690
rect 675477 713632 675482 713688
rect 675538 713632 676292 713688
rect 675477 713630 676292 713632
rect 675477 713627 675543 713630
rect 677685 713492 677751 713493
rect 677685 713488 677732 713492
rect 677796 713490 677802 713492
rect 677685 713432 677690 713488
rect 677685 713428 677732 713432
rect 677796 713430 677842 713490
rect 677796 713428 677802 713430
rect 677685 713427 677751 713428
rect 675477 713282 675543 713285
rect 675477 713280 676292 713282
rect 675477 713224 675482 713280
rect 675538 713224 676292 713280
rect 675477 713222 676292 713224
rect 675477 713219 675543 713222
rect 675477 712874 675543 712877
rect 675477 712872 676292 712874
rect 675477 712816 675482 712872
rect 675538 712816 676292 712872
rect 675477 712814 676292 712816
rect 675477 712811 675543 712814
rect 675477 712466 675543 712469
rect 675477 712464 676292 712466
rect 675477 712408 675482 712464
rect 675538 712408 676292 712464
rect 675477 712406 676292 712408
rect 675477 712403 675543 712406
rect 40350 712132 40356 712196
rect 40420 712194 40426 712196
rect 41781 712194 41847 712197
rect 40420 712192 41847 712194
rect 40420 712136 41786 712192
rect 41842 712136 41847 712192
rect 40420 712134 41847 712136
rect 40420 712132 40426 712134
rect 41781 712131 41847 712134
rect 675477 712058 675543 712061
rect 675477 712056 676292 712058
rect 675477 712000 675482 712056
rect 675538 712000 676292 712056
rect 675477 711998 676292 712000
rect 675477 711995 675543 711998
rect 42149 711650 42215 711653
rect 42558 711650 42564 711652
rect 42149 711648 42564 711650
rect 42149 711592 42154 711648
rect 42210 711592 42564 711648
rect 42149 711590 42564 711592
rect 42149 711587 42215 711590
rect 42558 711588 42564 711590
rect 42628 711588 42634 711652
rect 676029 711650 676095 711653
rect 676029 711648 676292 711650
rect 676029 711592 676034 711648
rect 676090 711592 676292 711648
rect 676029 711590 676292 711592
rect 676029 711587 676095 711590
rect 675477 711242 675543 711245
rect 675477 711240 676292 711242
rect 675477 711184 675482 711240
rect 675538 711184 676292 711240
rect 675477 711182 676292 711184
rect 675477 711179 675543 711182
rect 683113 710834 683179 710837
rect 683100 710832 683179 710834
rect 683100 710776 683118 710832
rect 683174 710776 683179 710832
rect 683100 710774 683179 710776
rect 683113 710771 683179 710774
rect 669405 710698 669471 710701
rect 675845 710698 675911 710701
rect 669405 710696 675911 710698
rect 669405 710640 669410 710696
rect 669466 710640 675850 710696
rect 675906 710640 675911 710696
rect 669405 710638 675911 710640
rect 669405 710635 669471 710638
rect 675845 710635 675911 710638
rect 42006 710364 42012 710428
rect 42076 710426 42082 710428
rect 42241 710426 42307 710429
rect 42076 710424 42307 710426
rect 42076 710368 42246 710424
rect 42302 710368 42307 710424
rect 42076 710366 42307 710368
rect 42076 710364 42082 710366
rect 42241 710363 42307 710366
rect 675477 710426 675543 710429
rect 675477 710424 676292 710426
rect 675477 710368 675482 710424
rect 675538 710368 676292 710424
rect 675477 710366 676292 710368
rect 675477 710363 675543 710366
rect 651649 710290 651715 710293
rect 650164 710288 651715 710290
rect 650164 710232 651654 710288
rect 651710 710232 651715 710288
rect 650164 710230 651715 710232
rect 651649 710227 651715 710230
rect 675293 710018 675359 710021
rect 675293 710016 676292 710018
rect 675293 709960 675298 710016
rect 675354 709960 676292 710016
rect 675293 709958 676292 709960
rect 675293 709955 675359 709958
rect 675477 709610 675543 709613
rect 675477 709608 676292 709610
rect 675477 709552 675482 709608
rect 675538 709552 676292 709608
rect 675477 709550 676292 709552
rect 675477 709547 675543 709550
rect 40718 709412 40724 709476
rect 40788 709474 40794 709476
rect 40788 709414 42258 709474
rect 40788 709412 40794 709414
rect 42198 709205 42258 709414
rect 42198 709200 42307 709205
rect 42198 709144 42246 709200
rect 42302 709144 42307 709200
rect 42198 709142 42307 709144
rect 42241 709139 42307 709142
rect 674230 709140 674236 709204
rect 674300 709202 674306 709204
rect 674300 709142 676292 709202
rect 674300 709140 674306 709142
rect 675477 708794 675543 708797
rect 675477 708792 676292 708794
rect 675477 708736 675482 708792
rect 675538 708736 676292 708792
rect 675477 708734 676292 708736
rect 675477 708731 675543 708734
rect 40902 708460 40908 708524
rect 40972 708522 40978 708524
rect 41781 708522 41847 708525
rect 40972 708520 41847 708522
rect 40972 708464 41786 708520
rect 41842 708464 41847 708520
rect 40972 708462 41847 708464
rect 40972 708460 40978 708462
rect 41781 708459 41847 708462
rect 675477 708386 675543 708389
rect 675477 708384 676292 708386
rect 675477 708328 675482 708384
rect 675538 708328 676292 708384
rect 675477 708326 676292 708328
rect 675477 708323 675543 708326
rect 683481 707978 683547 707981
rect 683468 707976 683547 707978
rect 683468 707920 683486 707976
rect 683542 707920 683547 707976
rect 683468 707918 683547 707920
rect 683481 707915 683547 707918
rect 42057 707842 42123 707845
rect 44357 707842 44423 707845
rect 42057 707840 44423 707842
rect 42057 707784 42062 707840
rect 42118 707784 44362 707840
rect 44418 707784 44423 707840
rect 42057 707782 44423 707784
rect 42057 707779 42123 707782
rect 44357 707779 44423 707782
rect 675477 707570 675543 707573
rect 675477 707568 676292 707570
rect 675477 707512 675482 707568
rect 675538 707512 676292 707568
rect 675477 707510 676292 707512
rect 675477 707507 675543 707510
rect 40534 707236 40540 707300
rect 40604 707298 40610 707300
rect 42425 707298 42491 707301
rect 40604 707296 42491 707298
rect 40604 707240 42430 707296
rect 42486 707240 42491 707296
rect 40604 707238 42491 707240
rect 40604 707236 40610 707238
rect 42425 707235 42491 707238
rect 674465 707162 674531 707165
rect 674465 707160 676292 707162
rect 674465 707104 674470 707160
rect 674526 707104 676292 707160
rect 674465 707102 676292 707104
rect 674465 707099 674531 707102
rect 683297 706754 683363 706757
rect 683284 706752 683363 706754
rect 683284 706696 683302 706752
rect 683358 706696 683363 706752
rect 683284 706694 683363 706696
rect 683297 706691 683363 706694
rect 42057 706618 42123 706621
rect 42374 706618 42380 706620
rect 42057 706616 42380 706618
rect 42057 706560 42062 706616
rect 42118 706560 42380 706616
rect 42057 706558 42380 706560
rect 42057 706555 42123 706558
rect 42374 706556 42380 706558
rect 42444 706556 42450 706620
rect 675477 706346 675543 706349
rect 675477 706344 676292 706346
rect 675477 706288 675482 706344
rect 675538 706288 676292 706344
rect 675477 706286 676292 706288
rect 675477 706283 675543 706286
rect 677182 705530 677242 705908
rect 683113 705530 683179 705533
rect 677182 705528 683179 705530
rect 677182 705500 683118 705528
rect 677212 705472 683118 705500
rect 683174 705472 683179 705528
rect 677212 705470 683179 705472
rect 683113 705467 683179 705470
rect 675477 705122 675543 705125
rect 675477 705120 676292 705122
rect 675477 705064 675482 705120
rect 675538 705064 676292 705120
rect 675477 705062 676292 705064
rect 675477 705059 675543 705062
rect 41454 702476 41460 702540
rect 41524 702538 41530 702540
rect 42609 702538 42675 702541
rect 41524 702536 42675 702538
rect 41524 702480 42614 702536
rect 42670 702480 42675 702536
rect 41524 702478 42675 702480
rect 41524 702476 41530 702478
rect 42609 702475 42675 702478
rect 62113 702266 62179 702269
rect 62113 702264 64492 702266
rect 62113 702208 62118 702264
rect 62174 702208 64492 702264
rect 62113 702206 64492 702208
rect 62113 702203 62179 702206
rect 41638 701388 41644 701452
rect 41708 701450 41714 701452
rect 42425 701450 42491 701453
rect 41708 701448 42491 701450
rect 41708 701392 42430 701448
rect 42486 701392 42491 701448
rect 41708 701390 42491 701392
rect 41708 701388 41714 701390
rect 42425 701387 42491 701390
rect 41822 701116 41828 701180
rect 41892 701178 41898 701180
rect 42241 701178 42307 701181
rect 41892 701176 42307 701178
rect 41892 701120 42246 701176
rect 42302 701120 42307 701176
rect 41892 701118 42307 701120
rect 41892 701116 41898 701118
rect 42241 701115 42307 701118
rect 651649 696962 651715 696965
rect 650164 696960 651715 696962
rect 650164 696904 651654 696960
rect 651710 696904 651715 696960
rect 650164 696902 651715 696904
rect 651649 696899 651715 696902
rect 675385 696828 675451 696829
rect 675334 696826 675340 696828
rect 675294 696766 675340 696826
rect 675404 696824 675451 696828
rect 675446 696768 675451 696824
rect 675334 696764 675340 696766
rect 675404 696764 675451 696768
rect 675385 696763 675451 696764
rect 674046 694588 674052 694652
rect 674116 694650 674122 694652
rect 675109 694650 675175 694653
rect 674116 694648 675175 694650
rect 674116 694592 675114 694648
rect 675170 694592 675175 694648
rect 674116 694590 675175 694592
rect 674116 694588 674122 694590
rect 675109 694587 675175 694590
rect 674925 694106 674991 694109
rect 676990 694106 676996 694108
rect 674925 694104 676996 694106
rect 674925 694048 674930 694104
rect 674986 694048 676996 694104
rect 674925 694046 676996 694048
rect 674925 694043 674991 694046
rect 676990 694044 676996 694046
rect 677060 694044 677066 694108
rect 674598 692956 674604 693020
rect 674668 693018 674674 693020
rect 675109 693018 675175 693021
rect 674668 693016 675175 693018
rect 674668 692960 675114 693016
rect 675170 692960 675175 693016
rect 674668 692958 675175 692960
rect 674668 692956 674674 692958
rect 675109 692955 675175 692958
rect 62113 689210 62179 689213
rect 62113 689208 64492 689210
rect 62113 689152 62118 689208
rect 62174 689152 64492 689208
rect 62113 689150 64492 689152
rect 62113 689147 62179 689150
rect 668761 688666 668827 688669
rect 675109 688666 675175 688669
rect 668761 688664 675175 688666
rect 668761 688608 668766 688664
rect 668822 688608 675114 688664
rect 675170 688608 675175 688664
rect 668761 688606 675175 688608
rect 668761 688603 668827 688606
rect 675109 688603 675175 688606
rect 40953 688394 41019 688397
rect 40910 688392 41019 688394
rect 40910 688336 40958 688392
rect 41014 688336 41019 688392
rect 40910 688331 41019 688336
rect 40910 688092 40970 688331
rect 43437 687714 43503 687717
rect 41492 687712 43503 687714
rect 41492 687656 43442 687712
rect 43498 687656 43503 687712
rect 41492 687654 43503 687656
rect 43437 687651 43503 687654
rect 42517 687306 42583 687309
rect 41492 687304 42583 687306
rect 41492 687248 42522 687304
rect 42578 687248 42583 687304
rect 41492 687246 42583 687248
rect 42517 687243 42583 687246
rect 41137 686898 41203 686901
rect 41124 686896 41203 686898
rect 41124 686840 41142 686896
rect 41198 686840 41203 686896
rect 41124 686838 41203 686840
rect 41137 686835 41203 686838
rect 44265 686490 44331 686493
rect 41492 686488 44331 686490
rect 41492 686432 44270 686488
rect 44326 686432 44331 686488
rect 41492 686430 44331 686432
rect 44265 686427 44331 686430
rect 41278 685915 41338 686052
rect 40861 685912 40927 685915
rect 40861 685910 40970 685912
rect 40861 685854 40866 685910
rect 40922 685854 40970 685910
rect 40861 685849 40970 685854
rect 41278 685910 41387 685915
rect 41278 685854 41326 685910
rect 41382 685854 41387 685910
rect 675334 685890 675340 685948
rect 41278 685852 41387 685854
rect 41321 685849 41387 685852
rect 675296 685884 675340 685890
rect 675404 685884 675410 685948
rect 40910 685644 40970 685849
rect 675296 685830 675402 685884
rect 675296 685677 675356 685830
rect 675293 685672 675359 685677
rect 675293 685616 675298 685672
rect 675354 685616 675359 685672
rect 675293 685611 675359 685616
rect 41137 685266 41203 685269
rect 41124 685264 41203 685266
rect 41124 685208 41142 685264
rect 41198 685208 41203 685264
rect 41124 685206 41203 685208
rect 41137 685203 41203 685206
rect 669037 685130 669103 685133
rect 675477 685130 675543 685133
rect 669037 685128 675543 685130
rect 669037 685072 669042 685128
rect 669098 685072 675482 685128
rect 675538 685072 675543 685128
rect 669037 685070 675543 685072
rect 669037 685067 669103 685070
rect 675477 685067 675543 685070
rect 41492 684798 41844 684858
rect 40769 684688 40835 684691
rect 40726 684686 40835 684688
rect 40726 684630 40774 684686
rect 40830 684630 40835 684686
rect 40726 684625 40835 684630
rect 40726 684420 40786 684625
rect 41784 684586 41844 684798
rect 43069 684586 43135 684589
rect 41784 684584 43135 684586
rect 41784 684528 43074 684584
rect 43130 684528 43135 684584
rect 41784 684526 43135 684528
rect 43069 684523 43135 684526
rect 674833 684314 674899 684317
rect 675477 684314 675543 684317
rect 674833 684312 675543 684314
rect 674833 684256 674838 684312
rect 674894 684256 675482 684312
rect 675538 684256 675543 684312
rect 674833 684254 675543 684256
rect 674833 684251 674899 684254
rect 675477 684251 675543 684254
rect 41137 684042 41203 684045
rect 41124 684040 41203 684042
rect 41124 683984 41142 684040
rect 41198 683984 41203 684040
rect 41124 683982 41203 683984
rect 41137 683979 41203 683982
rect 40953 683634 41019 683637
rect 651649 683634 651715 683637
rect 40940 683632 41019 683634
rect 40940 683576 40958 683632
rect 41014 683576 41019 683632
rect 40940 683574 41019 683576
rect 650164 683632 651715 683634
rect 650164 683576 651654 683632
rect 651710 683576 651715 683632
rect 650164 683574 651715 683576
rect 40953 683571 41019 683574
rect 651649 683571 651715 683574
rect 41321 683226 41387 683229
rect 41308 683224 41387 683226
rect 41308 683168 41326 683224
rect 41382 683168 41387 683224
rect 41308 683166 41387 683168
rect 41321 683163 41387 683166
rect 673637 683090 673703 683093
rect 675845 683090 675911 683093
rect 673637 683088 675911 683090
rect 673637 683032 673642 683088
rect 673698 683032 675850 683088
rect 675906 683032 675911 683088
rect 673637 683030 675911 683032
rect 673637 683027 673703 683030
rect 675845 683027 675911 683030
rect 41321 682818 41387 682821
rect 41308 682816 41387 682818
rect 41308 682760 41326 682816
rect 41382 682760 41387 682816
rect 41308 682758 41387 682760
rect 41321 682755 41387 682758
rect 673453 682818 673519 682821
rect 676029 682818 676095 682821
rect 673453 682816 676095 682818
rect 673453 682760 673458 682816
rect 673514 682760 676034 682816
rect 676090 682760 676095 682816
rect 673453 682758 676095 682760
rect 673453 682755 673519 682758
rect 676029 682755 676095 682758
rect 34421 682410 34487 682413
rect 41781 682412 41847 682413
rect 34421 682408 34500 682410
rect 34421 682352 34426 682408
rect 34482 682352 34500 682408
rect 34421 682350 34500 682352
rect 41781 682408 41828 682412
rect 41892 682410 41898 682412
rect 41781 682352 41786 682408
rect 34421 682347 34487 682350
rect 41781 682348 41828 682352
rect 41892 682350 41938 682410
rect 41892 682348 41898 682350
rect 41781 682347 41847 682348
rect 40677 682002 40743 682005
rect 40677 682000 40756 682002
rect 40677 681944 40682 682000
rect 40738 681944 40756 682000
rect 40677 681942 40756 681944
rect 40677 681939 40743 681942
rect 676070 681804 676076 681868
rect 676140 681866 676146 681868
rect 680997 681866 681063 681869
rect 676140 681864 681063 681866
rect 676140 681808 681002 681864
rect 681058 681808 681063 681864
rect 676140 681806 681063 681808
rect 676140 681804 676146 681806
rect 680997 681803 681063 681806
rect 36537 681594 36603 681597
rect 36524 681592 36603 681594
rect 36524 681536 36542 681592
rect 36598 681536 36603 681592
rect 36524 681534 36603 681536
rect 36537 681531 36603 681534
rect 32397 681186 32463 681189
rect 32397 681184 32476 681186
rect 32397 681128 32402 681184
rect 32458 681128 32476 681184
rect 32397 681126 32476 681128
rect 32397 681123 32463 681126
rect 31017 680778 31083 680781
rect 31004 680776 31083 680778
rect 31004 680720 31022 680776
rect 31078 680720 31083 680776
rect 31004 680718 31083 680720
rect 31017 680715 31083 680718
rect 43253 680642 43319 680645
rect 41784 680640 43319 680642
rect 41784 680608 43258 680640
rect 41462 680584 43258 680608
rect 43314 680584 43319 680640
rect 41462 680582 43319 680584
rect 41462 680548 41844 680582
rect 43253 680579 43319 680582
rect 41462 680340 41522 680548
rect 41781 680372 41847 680373
rect 41781 680368 41828 680372
rect 41892 680370 41898 680372
rect 41781 680312 41786 680368
rect 41781 680308 41828 680312
rect 41892 680310 41938 680370
rect 41892 680308 41898 680310
rect 41781 680307 41847 680308
rect 44633 679962 44699 679965
rect 41492 679960 44699 679962
rect 41492 679904 44638 679960
rect 44694 679904 44699 679960
rect 41492 679902 44699 679904
rect 44633 679899 44699 679902
rect 45185 679554 45251 679557
rect 41492 679552 45251 679554
rect 41492 679496 45190 679552
rect 45246 679496 45251 679552
rect 41492 679494 45251 679496
rect 45185 679491 45251 679494
rect 40542 678992 40602 679116
rect 40534 678928 40540 678992
rect 40604 678928 40610 678992
rect 40718 678928 40724 678992
rect 40788 678928 40794 678992
rect 40726 678708 40786 678928
rect 43437 678330 43503 678333
rect 41492 678328 43503 678330
rect 41492 678272 43442 678328
rect 43498 678272 43503 678328
rect 41492 678270 43503 678272
rect 43437 678267 43503 678270
rect 45001 677922 45067 677925
rect 41492 677920 45067 677922
rect 41492 677864 45006 677920
rect 45062 677864 45067 677920
rect 41492 677862 45067 677864
rect 45001 677859 45067 677862
rect 41094 677109 41154 677484
rect 41094 677104 41203 677109
rect 41094 677076 41142 677104
rect 41124 677048 41142 677076
rect 41198 677048 41203 677104
rect 41124 677046 41203 677048
rect 41137 677043 41203 677046
rect 42057 676698 42123 676701
rect 41492 676696 42123 676698
rect 41492 676640 42062 676696
rect 42118 676640 42123 676696
rect 41492 676638 42123 676640
rect 42057 676635 42123 676638
rect 62113 676154 62179 676157
rect 62113 676152 64492 676154
rect 62113 676096 62118 676152
rect 62174 676096 64492 676152
rect 62113 676094 64492 676096
rect 62113 676091 62179 676094
rect 40677 675610 40743 675613
rect 42057 675610 42123 675613
rect 40677 675608 42123 675610
rect 40677 675552 40682 675608
rect 40738 675552 42062 675608
rect 42118 675552 42123 675608
rect 40677 675550 42123 675552
rect 40677 675547 40743 675550
rect 42057 675547 42123 675550
rect 674414 674052 674420 674116
rect 674484 674114 674490 674116
rect 684033 674114 684099 674117
rect 674484 674112 684099 674114
rect 674484 674056 684038 674112
rect 684094 674056 684099 674112
rect 674484 674054 684099 674056
rect 674484 674052 674490 674054
rect 684033 674051 684099 674054
rect 32397 672754 32463 672757
rect 41822 672754 41828 672756
rect 32397 672752 41828 672754
rect 32397 672696 32402 672752
rect 32458 672696 41828 672752
rect 32397 672694 41828 672696
rect 32397 672691 32463 672694
rect 41822 672692 41828 672694
rect 41892 672692 41898 672756
rect 41137 672482 41203 672485
rect 42333 672482 42399 672485
rect 41137 672480 42399 672482
rect 41137 672424 41142 672480
rect 41198 672424 42338 672480
rect 42394 672424 42399 672480
rect 41137 672422 42399 672424
rect 41137 672419 41203 672422
rect 42333 672419 42399 672422
rect 675477 671394 675543 671397
rect 675477 671392 676292 671394
rect 675477 671336 675482 671392
rect 675538 671336 676292 671392
rect 675477 671334 676292 671336
rect 675477 671331 675543 671334
rect 40401 671258 40467 671261
rect 41086 671258 41092 671260
rect 40401 671256 41092 671258
rect 40401 671200 40406 671256
rect 40462 671200 41092 671256
rect 40401 671198 41092 671200
rect 40401 671195 40467 671198
rect 41086 671196 41092 671198
rect 41156 671196 41162 671260
rect 39757 670986 39823 670989
rect 40902 670986 40908 670988
rect 39757 670984 40908 670986
rect 39757 670928 39762 670984
rect 39818 670928 40908 670984
rect 39757 670926 40908 670928
rect 39757 670923 39823 670926
rect 40902 670924 40908 670926
rect 40972 670924 40978 670988
rect 675477 670986 675543 670989
rect 675477 670984 676292 670986
rect 675477 670928 675482 670984
rect 675538 670928 676292 670984
rect 675477 670926 676292 670928
rect 675477 670923 675543 670926
rect 675477 670578 675543 670581
rect 675477 670576 676292 670578
rect 675477 670520 675482 670576
rect 675538 670520 676292 670576
rect 675477 670518 676292 670520
rect 675477 670515 675543 670518
rect 651649 670442 651715 670445
rect 650164 670440 651715 670442
rect 650164 670384 651654 670440
rect 651710 670384 651715 670440
rect 650164 670382 651715 670384
rect 651649 670379 651715 670382
rect 675477 670170 675543 670173
rect 675477 670168 676292 670170
rect 675477 670112 675482 670168
rect 675538 670112 676292 670168
rect 675477 670110 676292 670112
rect 675477 670107 675543 670110
rect 674833 669762 674899 669765
rect 674833 669760 676292 669762
rect 674833 669704 674838 669760
rect 674894 669704 676292 669760
rect 674833 669702 676292 669704
rect 674833 669699 674899 669702
rect 675477 669354 675543 669357
rect 675477 669352 676292 669354
rect 675477 669296 675482 669352
rect 675538 669296 676292 669352
rect 675477 669294 676292 669296
rect 675477 669291 675543 669294
rect 674005 668946 674071 668949
rect 674005 668944 676292 668946
rect 674005 668888 674010 668944
rect 674066 668888 676292 668944
rect 674005 668886 676292 668888
rect 674005 668883 674071 668886
rect 675477 668538 675543 668541
rect 675477 668536 676292 668538
rect 675477 668480 675482 668536
rect 675538 668480 676292 668536
rect 675477 668478 676292 668480
rect 675477 668475 675543 668478
rect 671846 668070 676292 668130
rect 40902 667932 40908 667996
rect 40972 667994 40978 667996
rect 42609 667994 42675 667997
rect 40972 667992 42675 667994
rect 40972 667936 42614 667992
rect 42670 667936 42675 667992
rect 40972 667934 42675 667936
rect 40972 667932 40978 667934
rect 42609 667931 42675 667934
rect 671846 667861 671906 668070
rect 671797 667856 671906 667861
rect 671797 667800 671802 667856
rect 671858 667800 671906 667856
rect 671797 667798 671906 667800
rect 671797 667795 671863 667798
rect 42149 667722 42215 667725
rect 43621 667722 43687 667725
rect 42149 667720 43687 667722
rect 42149 667664 42154 667720
rect 42210 667664 43626 667720
rect 43682 667664 43687 667720
rect 42149 667662 43687 667664
rect 42149 667659 42215 667662
rect 43621 667659 43687 667662
rect 675477 667722 675543 667725
rect 675477 667720 676292 667722
rect 675477 667664 675482 667720
rect 675538 667664 676292 667720
rect 675477 667662 676292 667664
rect 675477 667659 675543 667662
rect 41086 667388 41092 667452
rect 41156 667450 41162 667452
rect 42425 667450 42491 667453
rect 41156 667448 42491 667450
rect 41156 667392 42430 667448
rect 42486 667392 42491 667448
rect 41156 667390 42491 667392
rect 41156 667388 41162 667390
rect 42425 667387 42491 667390
rect 675477 667314 675543 667317
rect 675477 667312 676292 667314
rect 675477 667256 675482 667312
rect 675538 667256 676292 667312
rect 675477 667254 676292 667256
rect 675477 667251 675543 667254
rect 680997 667042 681063 667045
rect 680997 667040 681106 667042
rect 680997 666984 681002 667040
rect 681058 666984 681106 667040
rect 680997 666979 681106 666984
rect 681046 666876 681106 666979
rect 676990 666572 676996 666636
rect 677060 666572 677066 666636
rect 40718 666436 40724 666500
rect 40788 666498 40794 666500
rect 42006 666498 42012 666500
rect 40788 666438 42012 666498
rect 40788 666436 40794 666438
rect 42006 666436 42012 666438
rect 42076 666436 42082 666500
rect 676998 666468 677058 666572
rect 42149 666362 42215 666365
rect 44633 666362 44699 666365
rect 42149 666360 44699 666362
rect 42149 666304 42154 666360
rect 42210 666304 44638 666360
rect 44694 666304 44699 666360
rect 42149 666302 44699 666304
rect 42149 666299 42215 666302
rect 44633 666299 44699 666302
rect 675477 666090 675543 666093
rect 675477 666088 676292 666090
rect 675477 666032 675482 666088
rect 675538 666032 676292 666088
rect 675477 666030 676292 666032
rect 675477 666027 675543 666030
rect 675477 665682 675543 665685
rect 675477 665680 676292 665682
rect 675477 665624 675482 665680
rect 675538 665624 676292 665680
rect 675477 665622 676292 665624
rect 675477 665619 675543 665622
rect 676806 665348 676812 665412
rect 676876 665348 676882 665412
rect 676814 665244 676874 665348
rect 675661 664866 675727 664869
rect 675661 664864 676292 664866
rect 675661 664808 675666 664864
rect 675722 664808 676292 664864
rect 675661 664806 676292 664808
rect 675661 664803 675727 664806
rect 675477 664458 675543 664461
rect 675477 664456 676292 664458
rect 675477 664400 675482 664456
rect 675538 664400 676292 664456
rect 675477 664398 676292 664400
rect 675477 664395 675543 664398
rect 41965 664052 42031 664053
rect 41965 664048 42012 664052
rect 42076 664050 42082 664052
rect 674833 664050 674899 664053
rect 41965 663992 41970 664048
rect 41965 663988 42012 663992
rect 42076 663990 42122 664050
rect 674833 664048 676292 664050
rect 674833 663992 674838 664048
rect 674894 663992 676292 664048
rect 674833 663990 676292 663992
rect 42076 663988 42082 663990
rect 41965 663987 42031 663988
rect 674833 663987 674899 663990
rect 684033 663778 684099 663781
rect 683990 663776 684099 663778
rect 683990 663720 684038 663776
rect 684094 663720 684099 663776
rect 683990 663715 684099 663720
rect 683990 663612 684050 663715
rect 672901 663506 672967 663509
rect 675845 663506 675911 663509
rect 672901 663504 675911 663506
rect 672901 663448 672906 663504
rect 672962 663448 675850 663504
rect 675906 663448 675911 663504
rect 672901 663446 675911 663448
rect 672901 663443 672967 663446
rect 675845 663443 675911 663446
rect 675477 663234 675543 663237
rect 675477 663232 676292 663234
rect 675477 663176 675482 663232
rect 675538 663176 676292 663232
rect 675477 663174 676292 663176
rect 675477 663171 675543 663174
rect 62113 663098 62179 663101
rect 62113 663096 64492 663098
rect 62113 663040 62118 663096
rect 62174 663040 64492 663096
rect 62113 663038 64492 663040
rect 62113 663035 62179 663038
rect 42057 662826 42123 662829
rect 41370 662824 42123 662826
rect 41370 662768 42062 662824
rect 42118 662768 42123 662824
rect 41370 662766 42123 662768
rect 40534 662628 40540 662692
rect 40604 662690 40610 662692
rect 41370 662690 41430 662766
rect 42057 662763 42123 662766
rect 675477 662826 675543 662829
rect 675477 662824 676292 662826
rect 675477 662768 675482 662824
rect 675538 662768 676292 662824
rect 675477 662766 676292 662768
rect 675477 662763 675543 662766
rect 40604 662630 41430 662690
rect 40604 662628 40610 662630
rect 683205 662554 683271 662557
rect 683205 662552 683314 662554
rect 683205 662496 683210 662552
rect 683266 662496 683314 662552
rect 683205 662491 683314 662496
rect 683254 662388 683314 662491
rect 683389 662146 683455 662149
rect 683389 662144 683498 662146
rect 683389 662088 683394 662144
rect 683450 662088 683498 662144
rect 683389 662083 683498 662088
rect 683438 661980 683498 662083
rect 675477 661602 675543 661605
rect 675477 661600 676292 661602
rect 675477 661544 675482 661600
rect 675538 661544 676292 661600
rect 675477 661542 676292 661544
rect 675477 661539 675543 661542
rect 675477 661194 675543 661197
rect 675477 661192 676292 661194
rect 675477 661136 675482 661192
rect 675538 661136 676292 661192
rect 675477 661134 676292 661136
rect 675477 661131 675543 661134
rect 683070 660109 683130 660756
rect 683070 660104 683179 660109
rect 683070 660048 683118 660104
rect 683174 660048 683179 660104
rect 683070 660046 683179 660048
rect 683113 660043 683179 660046
rect 675477 659970 675543 659973
rect 675477 659968 676292 659970
rect 675477 659912 675482 659968
rect 675538 659912 676292 659968
rect 675477 659910 676292 659912
rect 675477 659907 675543 659910
rect 41454 659636 41460 659700
rect 41524 659698 41530 659700
rect 42701 659698 42767 659701
rect 41524 659696 42767 659698
rect 41524 659640 42706 659696
rect 42762 659640 42767 659696
rect 41524 659638 42767 659640
rect 41524 659636 41530 659638
rect 42701 659635 42767 659638
rect 41638 658548 41644 658612
rect 41708 658610 41714 658612
rect 42425 658610 42491 658613
rect 41708 658608 42491 658610
rect 41708 658552 42430 658608
rect 42486 658552 42491 658608
rect 41708 658550 42491 658552
rect 41708 658548 41714 658550
rect 42425 658547 42491 658550
rect 41822 658276 41828 658340
rect 41892 658338 41898 658340
rect 42149 658338 42215 658341
rect 41892 658336 42215 658338
rect 41892 658280 42154 658336
rect 42210 658280 42215 658336
rect 41892 658278 42215 658280
rect 41892 658276 41898 658278
rect 42149 658275 42215 658278
rect 651649 657114 651715 657117
rect 650164 657112 651715 657114
rect 650164 657056 651654 657112
rect 651710 657056 651715 657112
rect 650164 657054 651715 657056
rect 651649 657051 651715 657054
rect 675569 652900 675635 652901
rect 675518 652898 675524 652900
rect 675478 652838 675524 652898
rect 675588 652896 675635 652900
rect 675630 652840 675635 652896
rect 675518 652836 675524 652838
rect 675588 652836 675635 652840
rect 675569 652835 675635 652836
rect 675201 650180 675267 650181
rect 675150 650178 675156 650180
rect 675110 650118 675156 650178
rect 675220 650176 675267 650180
rect 675262 650120 675267 650176
rect 675150 650116 675156 650118
rect 675220 650116 675267 650120
rect 675201 650115 675267 650116
rect 62113 650042 62179 650045
rect 62113 650040 64492 650042
rect 62113 649984 62118 650040
rect 62174 649984 64492 650040
rect 62113 649982 64492 649984
rect 62113 649979 62179 649982
rect 674230 648892 674236 648956
rect 674300 648954 674306 648956
rect 675385 648954 675451 648957
rect 674300 648952 675451 648954
rect 674300 648896 675390 648952
rect 675446 648896 675451 648952
rect 674300 648894 675451 648896
rect 674300 648892 674306 648894
rect 675385 648891 675451 648894
rect 675150 647940 675156 648004
rect 675220 648002 675226 648004
rect 675385 648002 675451 648005
rect 675220 648000 675451 648002
rect 675220 647944 675390 648000
rect 675446 647944 675451 648000
rect 675220 647942 675451 647944
rect 675220 647940 675226 647942
rect 675385 647939 675451 647942
rect 670785 647458 670851 647461
rect 675661 647458 675727 647461
rect 670785 647456 675727 647458
rect 670785 647400 670790 647456
rect 670846 647400 675666 647456
rect 675722 647400 675727 647456
rect 670785 647398 675727 647400
rect 670785 647395 670851 647398
rect 675661 647395 675727 647398
rect 38837 646098 38903 646101
rect 47761 646098 47827 646101
rect 38837 646096 47827 646098
rect 38837 646040 38842 646096
rect 38898 646040 47766 646096
rect 47822 646040 47827 646096
rect 38837 646038 47827 646040
rect 38837 646035 38903 646038
rect 47761 646035 47827 646038
rect 41229 645690 41295 645693
rect 43805 645690 43871 645693
rect 41229 645688 43871 645690
rect 41229 645632 41234 645688
rect 41290 645632 43810 645688
rect 43866 645632 43871 645688
rect 41229 645630 43871 645632
rect 41229 645627 41295 645630
rect 43805 645627 43871 645630
rect 35574 644741 35634 644912
rect 35525 644736 35634 644741
rect 35801 644738 35867 644741
rect 35525 644680 35530 644736
rect 35586 644680 35634 644736
rect 35525 644678 35634 644680
rect 35758 644736 35867 644738
rect 35758 644680 35806 644736
rect 35862 644680 35867 644736
rect 35525 644675 35591 644678
rect 35758 644675 35867 644680
rect 39665 644738 39731 644741
rect 44449 644738 44515 644741
rect 39665 644736 44515 644738
rect 39665 644680 39670 644736
rect 39726 644680 44454 644736
rect 44510 644680 44515 644736
rect 39665 644678 44515 644680
rect 39665 644675 39731 644678
rect 44449 644675 44515 644678
rect 674005 644738 674071 644741
rect 675385 644738 675451 644741
rect 674005 644736 675451 644738
rect 674005 644680 674010 644736
rect 674066 644680 675390 644736
rect 675446 644680 675451 644736
rect 674005 644678 675451 644680
rect 674005 644675 674071 644678
rect 675385 644675 675451 644678
rect 35758 644504 35818 644675
rect 673729 644330 673795 644333
rect 675385 644330 675451 644333
rect 673729 644328 675451 644330
rect 673729 644272 673734 644328
rect 673790 644272 675390 644328
rect 675446 644272 675451 644328
rect 673729 644270 675451 644272
rect 673729 644267 673795 644270
rect 675385 644267 675451 644270
rect 35390 643925 35450 644096
rect 35341 643920 35450 643925
rect 674925 643924 674991 643925
rect 674925 643922 674972 643924
rect 35341 643864 35346 643920
rect 35402 643864 35450 643920
rect 35341 643862 35450 643864
rect 674880 643920 674972 643922
rect 674880 643864 674930 643920
rect 674880 643862 674972 643864
rect 35341 643859 35407 643862
rect 674925 643860 674972 643862
rect 675036 643860 675042 643924
rect 674925 643859 674991 643860
rect 651649 643786 651715 643789
rect 650164 643784 651715 643786
rect 650164 643728 651654 643784
rect 651710 643728 651715 643784
rect 650164 643726 651715 643728
rect 651649 643723 651715 643726
rect 35574 643517 35634 643688
rect 35525 643512 35634 643517
rect 35801 643514 35867 643517
rect 35525 643456 35530 643512
rect 35586 643456 35634 643512
rect 35525 643454 35634 643456
rect 35758 643512 35867 643514
rect 35758 643456 35806 643512
rect 35862 643456 35867 643512
rect 35525 643451 35591 643454
rect 35758 643451 35867 643456
rect 673913 643514 673979 643517
rect 675385 643514 675451 643517
rect 673913 643512 675451 643514
rect 673913 643456 673918 643512
rect 673974 643456 675390 643512
rect 675446 643456 675451 643512
rect 673913 643454 675451 643456
rect 673913 643451 673979 643454
rect 675385 643451 675451 643454
rect 35758 643280 35818 643451
rect 35390 642701 35450 642872
rect 35390 642696 35499 642701
rect 35390 642640 35438 642696
rect 35494 642640 35499 642696
rect 35390 642638 35499 642640
rect 35433 642635 35499 642638
rect 35574 642293 35634 642464
rect 35574 642288 35683 642293
rect 35574 642232 35622 642288
rect 35678 642232 35683 642288
rect 35574 642230 35683 642232
rect 35617 642227 35683 642230
rect 39021 642290 39087 642293
rect 43069 642290 43135 642293
rect 39021 642288 43135 642290
rect 39021 642232 39026 642288
rect 39082 642232 43074 642288
rect 43130 642232 43135 642288
rect 39021 642230 43135 642232
rect 39021 642227 39087 642230
rect 43069 642227 43135 642230
rect 669589 642154 669655 642157
rect 675385 642154 675451 642157
rect 669589 642152 675451 642154
rect 669589 642096 669594 642152
rect 669650 642096 675390 642152
rect 675446 642096 675451 642152
rect 669589 642094 675451 642096
rect 669589 642091 669655 642094
rect 675385 642091 675451 642094
rect 35758 641885 35818 642056
rect 35758 641880 35867 641885
rect 35758 641824 35806 641880
rect 35862 641824 35867 641880
rect 35758 641822 35867 641824
rect 35801 641819 35867 641822
rect 35390 641477 35450 641648
rect 35341 641472 35450 641477
rect 35341 641416 35346 641472
rect 35402 641416 35450 641472
rect 35341 641414 35450 641416
rect 39757 641474 39823 641477
rect 44265 641474 44331 641477
rect 39757 641472 44331 641474
rect 39757 641416 39762 641472
rect 39818 641416 44270 641472
rect 44326 641416 44331 641472
rect 39757 641414 44331 641416
rect 35341 641411 35407 641414
rect 39757 641411 39823 641414
rect 44265 641411 44331 641414
rect 35574 641069 35634 641240
rect 35525 641064 35634 641069
rect 35801 641066 35867 641069
rect 35525 641008 35530 641064
rect 35586 641008 35634 641064
rect 35525 641006 35634 641008
rect 35758 641064 35867 641066
rect 35758 641008 35806 641064
rect 35862 641008 35867 641064
rect 35525 641003 35591 641006
rect 35758 641003 35867 641008
rect 40309 641066 40375 641069
rect 44633 641066 44699 641069
rect 40309 641064 44699 641066
rect 40309 641008 40314 641064
rect 40370 641008 44638 641064
rect 44694 641008 44699 641064
rect 40309 641006 44699 641008
rect 40309 641003 40375 641006
rect 44633 641003 44699 641006
rect 35758 640832 35818 641003
rect 41454 640596 41460 640660
rect 41524 640596 41530 640660
rect 41462 640424 41522 640596
rect 675661 640386 675727 640389
rect 675661 640384 675770 640386
rect 675661 640328 675666 640384
rect 675722 640328 675770 640384
rect 675661 640323 675770 640328
rect 39849 640250 39915 640253
rect 42885 640250 42951 640253
rect 39849 640248 42951 640250
rect 39849 640192 39854 640248
rect 39910 640192 42890 640248
rect 42946 640192 42951 640248
rect 39849 640190 42951 640192
rect 675710 640250 675770 640323
rect 676806 640250 676812 640252
rect 675710 640190 676812 640250
rect 39849 640187 39915 640190
rect 42885 640187 42951 640190
rect 676806 640188 676812 640190
rect 676876 640188 676882 640252
rect 34470 639845 34530 640016
rect 34421 639840 34530 639845
rect 34421 639784 34426 639840
rect 34482 639784 34530 639840
rect 34421 639782 34530 639784
rect 34421 639779 34487 639782
rect 35574 639437 35634 639608
rect 35525 639432 35634 639437
rect 35801 639434 35867 639437
rect 35525 639376 35530 639432
rect 35586 639376 35634 639432
rect 35525 639374 35634 639376
rect 35758 639432 35867 639434
rect 35758 639376 35806 639432
rect 35862 639376 35867 639432
rect 35525 639371 35591 639374
rect 35758 639371 35867 639376
rect 35758 639200 35818 639371
rect 33734 638621 33794 638792
rect 33734 638616 33843 638621
rect 33734 638560 33782 638616
rect 33838 638560 33843 638616
rect 33734 638558 33843 638560
rect 33777 638555 33843 638558
rect 32446 638213 32506 638384
rect 32397 638208 32506 638213
rect 32397 638152 32402 638208
rect 32458 638152 32506 638208
rect 32397 638150 32506 638152
rect 32397 638147 32463 638150
rect 674966 638148 674972 638212
rect 675036 638210 675042 638212
rect 675477 638210 675543 638213
rect 675036 638208 675543 638210
rect 675036 638152 675482 638208
rect 675538 638152 675543 638208
rect 675036 638150 675543 638152
rect 675036 638148 675042 638150
rect 675477 638147 675543 638150
rect 35758 637805 35818 637976
rect 675293 637938 675359 637941
rect 675845 637938 675911 637941
rect 675293 637936 675911 637938
rect 675293 637880 675298 637936
rect 675354 637880 675850 637936
rect 675906 637880 675911 637936
rect 675293 637878 675911 637880
rect 675293 637875 675359 637878
rect 675845 637875 675911 637878
rect 35525 637802 35591 637805
rect 35525 637800 35634 637802
rect 35525 637744 35530 637800
rect 35586 637744 35634 637800
rect 35525 637739 35634 637744
rect 35758 637800 35867 637805
rect 35758 637744 35806 637800
rect 35862 637744 35867 637800
rect 35758 637742 35867 637744
rect 35801 637739 35867 637742
rect 41505 637802 41571 637805
rect 44449 637802 44515 637805
rect 41505 637800 44515 637802
rect 41505 637744 41510 637800
rect 41566 637744 44454 637800
rect 44510 637744 44515 637800
rect 41505 637742 44515 637744
rect 41505 637739 41571 637742
rect 44449 637739 44515 637742
rect 35574 637568 35634 637739
rect 675201 637666 675267 637669
rect 675518 637666 675524 637668
rect 675201 637664 675524 637666
rect 675201 637608 675206 637664
rect 675262 637608 675524 637664
rect 675201 637606 675524 637608
rect 675201 637603 675267 637606
rect 675518 637604 675524 637606
rect 675588 637604 675594 637668
rect 40033 637394 40099 637397
rect 41638 637394 41644 637396
rect 40033 637392 41644 637394
rect 40033 637336 40038 637392
rect 40094 637336 41644 637392
rect 40033 637334 41644 637336
rect 40033 637331 40099 637334
rect 41638 637332 41644 637334
rect 41708 637332 41714 637396
rect 40542 636988 40602 637160
rect 62113 637122 62179 637125
rect 62113 637120 64492 637122
rect 62113 637064 62118 637120
rect 62174 637064 64492 637120
rect 62113 637062 64492 637064
rect 62113 637059 62179 637062
rect 40534 636924 40540 636988
rect 40604 636924 40610 636988
rect 674046 636788 674052 636852
rect 674116 636850 674122 636852
rect 683389 636850 683455 636853
rect 674116 636848 683455 636850
rect 674116 636792 683394 636848
rect 683450 636792 683455 636848
rect 674116 636790 683455 636792
rect 674116 636788 674122 636790
rect 683389 636787 683455 636790
rect 35758 636581 35818 636752
rect 35758 636576 35867 636581
rect 35758 636520 35806 636576
rect 35862 636520 35867 636576
rect 35758 636518 35867 636520
rect 35801 636515 35867 636518
rect 675477 636578 675543 636581
rect 683205 636578 683271 636581
rect 675477 636576 683271 636578
rect 675477 636520 675482 636576
rect 675538 636520 683210 636576
rect 683266 636520 683271 636576
rect 675477 636518 683271 636520
rect 675477 636515 675543 636518
rect 683205 636515 683271 636518
rect 40910 636172 40970 636344
rect 40902 636108 40908 636172
rect 40972 636108 40978 636172
rect 41321 636170 41387 636173
rect 43989 636170 44055 636173
rect 41321 636168 44055 636170
rect 41321 636112 41326 636168
rect 41382 636112 43994 636168
rect 44050 636112 44055 636168
rect 41321 636110 44055 636112
rect 41321 636107 41387 636110
rect 43989 636107 44055 636110
rect 40726 635764 40786 635936
rect 40718 635700 40724 635764
rect 40788 635700 40794 635764
rect 35574 635357 35634 635528
rect 35574 635352 35683 635357
rect 35574 635296 35622 635352
rect 35678 635296 35683 635352
rect 35574 635294 35683 635296
rect 35617 635291 35683 635294
rect 40217 635354 40283 635357
rect 41822 635354 41828 635356
rect 40217 635352 41828 635354
rect 40217 635296 40222 635352
rect 40278 635296 41828 635352
rect 40217 635294 41828 635296
rect 40217 635291 40283 635294
rect 41822 635292 41828 635294
rect 41892 635292 41898 635356
rect 35758 634949 35818 635120
rect 35758 634944 35867 634949
rect 35758 634888 35806 634944
rect 35862 634888 35867 634944
rect 35758 634886 35867 634888
rect 35801 634883 35867 634886
rect 39757 634946 39823 634949
rect 43805 634946 43871 634949
rect 39757 634944 43871 634946
rect 39757 634888 39762 634944
rect 39818 634888 43810 634944
rect 43866 634888 43871 634944
rect 39757 634886 43871 634888
rect 39757 634883 39823 634886
rect 43805 634883 43871 634886
rect 35574 634541 35634 634712
rect 35574 634536 35683 634541
rect 35574 634480 35622 634536
rect 35678 634480 35683 634536
rect 35574 634478 35683 634480
rect 35617 634475 35683 634478
rect 41462 633858 41522 634304
rect 42333 633858 42399 633861
rect 41462 633856 42399 633858
rect 41462 633800 42338 633856
rect 42394 633800 42399 633856
rect 41462 633798 42399 633800
rect 42333 633795 42399 633798
rect 35801 633722 35867 633725
rect 35758 633720 35867 633722
rect 35758 633664 35806 633720
rect 35862 633664 35867 633720
rect 35758 633659 35867 633664
rect 35758 633488 35818 633659
rect 39297 631410 39363 631413
rect 45185 631410 45251 631413
rect 675201 631412 675267 631413
rect 675150 631410 675156 631412
rect 39297 631408 45251 631410
rect 39297 631352 39302 631408
rect 39358 631352 45190 631408
rect 45246 631352 45251 631408
rect 39297 631350 45251 631352
rect 675110 631350 675156 631410
rect 675220 631408 675267 631412
rect 675262 631352 675267 631408
rect 39297 631347 39363 631350
rect 45185 631347 45251 631350
rect 675150 631348 675156 631350
rect 675220 631348 675267 631352
rect 675201 631347 675267 631348
rect 675385 631410 675451 631413
rect 676070 631410 676076 631412
rect 675385 631408 676076 631410
rect 675385 631352 675390 631408
rect 675446 631352 676076 631408
rect 675385 631350 676076 631352
rect 675385 631347 675451 631350
rect 676070 631348 676076 631350
rect 676140 631348 676146 631412
rect 652017 630594 652083 630597
rect 650164 630592 652083 630594
rect 650164 630536 652022 630592
rect 652078 630536 652083 630592
rect 650164 630534 652083 630536
rect 652017 630531 652083 630534
rect 42190 626724 42196 626788
rect 42260 626786 42266 626788
rect 42701 626786 42767 626789
rect 42260 626784 42767 626786
rect 42260 626728 42706 626784
rect 42762 626728 42767 626784
rect 42260 626726 42767 626728
rect 42260 626724 42266 626726
rect 42701 626723 42767 626726
rect 675293 626378 675359 626381
rect 675293 626376 676292 626378
rect 675293 626320 675298 626376
rect 675354 626320 676292 626376
rect 675293 626318 676292 626320
rect 675293 626315 675359 626318
rect 675109 625970 675175 625973
rect 675109 625968 676292 625970
rect 675109 625912 675114 625968
rect 675170 625912 676292 625968
rect 675109 625910 676292 625912
rect 675109 625907 675175 625910
rect 675477 625562 675543 625565
rect 675477 625560 676292 625562
rect 675477 625504 675482 625560
rect 675538 625504 676292 625560
rect 675477 625502 676292 625504
rect 675477 625499 675543 625502
rect 40902 625228 40908 625292
rect 40972 625290 40978 625292
rect 42006 625290 42012 625292
rect 40972 625230 42012 625290
rect 40972 625228 40978 625230
rect 42006 625228 42012 625230
rect 42076 625228 42082 625292
rect 675293 625154 675359 625157
rect 675293 625152 676292 625154
rect 675293 625096 675298 625152
rect 675354 625096 676292 625152
rect 675293 625094 676292 625096
rect 675293 625091 675359 625094
rect 675109 624746 675175 624749
rect 675109 624744 676292 624746
rect 675109 624688 675114 624744
rect 675170 624688 676292 624744
rect 675109 624686 676292 624688
rect 675109 624683 675175 624686
rect 675477 624338 675543 624341
rect 675477 624336 676292 624338
rect 675477 624280 675482 624336
rect 675538 624280 676292 624336
rect 675477 624278 676292 624280
rect 675477 624275 675543 624278
rect 62113 624066 62179 624069
rect 62113 624064 64492 624066
rect 62113 624008 62118 624064
rect 62174 624008 64492 624064
rect 62113 624006 64492 624008
rect 62113 624003 62179 624006
rect 675477 623930 675543 623933
rect 675477 623928 676292 623930
rect 675477 623872 675482 623928
rect 675538 623872 676292 623928
rect 675477 623870 676292 623872
rect 675477 623867 675543 623870
rect 674598 623596 674604 623660
rect 674668 623658 674674 623660
rect 675293 623658 675359 623661
rect 674668 623656 675359 623658
rect 674668 623600 675298 623656
rect 675354 623600 675359 623656
rect 674668 623598 675359 623600
rect 674668 623596 674674 623598
rect 675293 623595 675359 623598
rect 676397 623658 676463 623661
rect 683389 623658 683455 623661
rect 676397 623656 683455 623658
rect 676397 623600 676402 623656
rect 676458 623600 683394 623656
rect 683450 623600 683455 623656
rect 676397 623598 683455 623600
rect 676397 623595 676463 623598
rect 683389 623595 683455 623598
rect 675477 623522 675543 623525
rect 675477 623520 676292 623522
rect 675477 623464 675482 623520
rect 675538 623464 676292 623520
rect 675477 623462 676292 623464
rect 675477 623459 675543 623462
rect 42149 623386 42215 623389
rect 43989 623386 44055 623389
rect 42149 623384 44055 623386
rect 42149 623328 42154 623384
rect 42210 623328 43994 623384
rect 44050 623328 44055 623384
rect 42149 623326 44055 623328
rect 42149 623323 42215 623326
rect 43989 623323 44055 623326
rect 675293 623114 675359 623117
rect 675293 623112 676292 623114
rect 675293 623056 675298 623112
rect 675354 623056 676292 623112
rect 675293 623054 676292 623056
rect 675293 623051 675359 623054
rect 675477 622706 675543 622709
rect 675477 622704 676292 622706
rect 675477 622648 675482 622704
rect 675538 622648 676292 622704
rect 675477 622646 676292 622648
rect 675477 622643 675543 622646
rect 675293 622298 675359 622301
rect 675293 622296 676292 622298
rect 675293 622240 675298 622296
rect 675354 622240 676292 622296
rect 675293 622238 676292 622240
rect 675293 622235 675359 622238
rect 679617 622026 679683 622029
rect 679574 622024 679683 622026
rect 679574 621968 679622 622024
rect 679678 621968 679683 622024
rect 679574 621963 679683 621968
rect 679574 621860 679634 621963
rect 682377 621618 682443 621621
rect 682334 621616 682443 621618
rect 682334 621560 682382 621616
rect 682438 621560 682443 621616
rect 682334 621555 682443 621560
rect 41965 621484 42031 621485
rect 41965 621480 42012 621484
rect 42076 621482 42082 621484
rect 41965 621424 41970 621480
rect 41965 621420 42012 621424
rect 42076 621422 42122 621482
rect 682334 621452 682394 621555
rect 42076 621420 42082 621422
rect 41965 621419 42031 621420
rect 675477 621074 675543 621077
rect 675477 621072 676292 621074
rect 675477 621016 675482 621072
rect 675538 621016 676292 621072
rect 675477 621014 676292 621016
rect 675477 621011 675543 621014
rect 683205 620802 683271 620805
rect 683205 620800 683314 620802
rect 683205 620744 683210 620800
rect 683266 620744 683314 620800
rect 683205 620739 683314 620744
rect 683254 620636 683314 620739
rect 41965 620258 42031 620261
rect 42190 620258 42196 620260
rect 41965 620256 42196 620258
rect 41965 620200 41970 620256
rect 42026 620200 42196 620256
rect 41965 620198 42196 620200
rect 41965 620195 42031 620198
rect 42190 620196 42196 620198
rect 42260 620196 42266 620260
rect 675477 620258 675543 620261
rect 675477 620256 676292 620258
rect 675477 620200 675482 620256
rect 675538 620200 676292 620256
rect 675477 620198 676292 620200
rect 675477 620195 675543 620198
rect 40718 619788 40724 619852
rect 40788 619850 40794 619852
rect 42241 619850 42307 619853
rect 40788 619848 42307 619850
rect 40788 619792 42246 619848
rect 42302 619792 42307 619848
rect 40788 619790 42307 619792
rect 40788 619788 40794 619790
rect 42241 619787 42307 619790
rect 675293 619850 675359 619853
rect 675293 619848 676292 619850
rect 675293 619792 675298 619848
rect 675354 619792 676292 619848
rect 675293 619790 676292 619792
rect 675293 619787 675359 619790
rect 675477 619442 675543 619445
rect 675477 619440 676292 619442
rect 675477 619384 675482 619440
rect 675538 619384 676292 619440
rect 675477 619382 676292 619384
rect 675477 619379 675543 619382
rect 683573 619170 683639 619173
rect 683573 619168 683682 619170
rect 683573 619112 683578 619168
rect 683634 619112 683682 619168
rect 683573 619107 683682 619112
rect 40534 618972 40540 619036
rect 40604 619034 40610 619036
rect 42425 619034 42491 619037
rect 40604 619032 42491 619034
rect 40604 618976 42430 619032
rect 42486 618976 42491 619032
rect 683622 619004 683682 619107
rect 40604 618974 42491 618976
rect 40604 618972 40610 618974
rect 42425 618971 42491 618974
rect 41822 618700 41828 618764
rect 41892 618762 41898 618764
rect 42701 618762 42767 618765
rect 41892 618760 42767 618762
rect 41892 618704 42706 618760
rect 42762 618704 42767 618760
rect 41892 618702 42767 618704
rect 41892 618700 41898 618702
rect 42701 618699 42767 618702
rect 674465 618626 674531 618629
rect 674465 618624 676292 618626
rect 674465 618568 674470 618624
rect 674526 618568 676292 618624
rect 674465 618566 676292 618568
rect 674465 618563 674531 618566
rect 675477 618218 675543 618221
rect 675477 618216 676292 618218
rect 675477 618160 675482 618216
rect 675538 618160 676292 618216
rect 675477 618158 676292 618160
rect 675477 618155 675543 618158
rect 674281 617810 674347 617813
rect 674281 617808 676292 617810
rect 674281 617752 674286 617808
rect 674342 617752 676292 617808
rect 674281 617750 676292 617752
rect 674281 617747 674347 617750
rect 683389 617538 683455 617541
rect 683389 617536 683498 617538
rect 683389 617480 683394 617536
rect 683450 617480 683498 617536
rect 683389 617475 683498 617480
rect 683438 617372 683498 617475
rect 651649 617266 651715 617269
rect 650164 617264 651715 617266
rect 650164 617208 651654 617264
rect 651710 617208 651715 617264
rect 650164 617206 651715 617208
rect 651649 617203 651715 617206
rect 669037 617266 669103 617269
rect 675845 617266 675911 617269
rect 669037 617264 675911 617266
rect 669037 617208 669042 617264
rect 669098 617208 675850 617264
rect 675906 617208 675911 617264
rect 669037 617206 675911 617208
rect 669037 617203 669103 617206
rect 675845 617203 675911 617206
rect 674649 616994 674715 616997
rect 674649 616992 676292 616994
rect 674649 616936 674654 616992
rect 674710 616936 676292 616992
rect 674649 616934 676292 616936
rect 674649 616931 674715 616934
rect 671470 616796 671476 616860
rect 671540 616858 671546 616860
rect 671889 616858 671955 616861
rect 671540 616856 671955 616858
rect 671540 616800 671894 616856
rect 671950 616800 671955 616856
rect 671540 616798 671955 616800
rect 671540 616796 671546 616798
rect 671889 616795 671955 616798
rect 675477 616586 675543 616589
rect 675477 616584 676292 616586
rect 675477 616528 675482 616584
rect 675538 616528 676292 616584
rect 675477 616526 676292 616528
rect 675477 616523 675543 616526
rect 675293 616178 675359 616181
rect 675293 616176 676292 616178
rect 675293 616120 675298 616176
rect 675354 616120 676292 616176
rect 675293 616118 676292 616120
rect 675293 616115 675359 616118
rect 41454 615980 41460 616044
rect 41524 616042 41530 616044
rect 42241 616042 42307 616045
rect 41524 616040 42307 616042
rect 41524 615984 42246 616040
rect 42302 615984 42307 616040
rect 41524 615982 42307 615984
rect 41524 615980 41530 615982
rect 42241 615979 42307 615982
rect 683070 615501 683130 615740
rect 683070 615498 683179 615501
rect 683070 615496 683260 615498
rect 683070 615440 683118 615496
rect 683174 615440 683260 615496
rect 683070 615438 683260 615440
rect 683070 615435 683179 615438
rect 683070 615332 683130 615435
rect 675477 614954 675543 614957
rect 675477 614952 676292 614954
rect 675477 614896 675482 614952
rect 675538 614896 676292 614952
rect 675477 614894 676292 614896
rect 675477 614891 675543 614894
rect 41781 612780 41847 612781
rect 41781 612776 41828 612780
rect 41892 612778 41898 612780
rect 41781 612720 41786 612776
rect 41781 612716 41828 612720
rect 41892 612718 41938 612778
rect 41892 612716 41898 612718
rect 41781 612715 41847 612716
rect 62113 611010 62179 611013
rect 62113 611008 64492 611010
rect 62113 610952 62118 611008
rect 62174 610952 64492 611008
rect 62113 610950 64492 610952
rect 62113 610947 62179 610950
rect 671521 608700 671587 608701
rect 671470 608636 671476 608700
rect 671540 608698 671587 608700
rect 671540 608696 671632 608698
rect 671582 608640 671632 608696
rect 671540 608638 671632 608640
rect 671540 608636 671587 608638
rect 671521 608635 671587 608636
rect 674414 604420 674420 604484
rect 674484 604482 674490 604484
rect 675109 604482 675175 604485
rect 674484 604480 675175 604482
rect 674484 604424 675114 604480
rect 675170 604424 675175 604480
rect 674484 604422 675175 604424
rect 674484 604420 674490 604422
rect 675109 604419 675175 604422
rect 652017 603938 652083 603941
rect 650164 603936 652083 603938
rect 650164 603880 652022 603936
rect 652078 603880 652083 603936
rect 650164 603878 652083 603880
rect 652017 603875 652083 603878
rect 674598 602924 674604 602988
rect 674668 602986 674674 602988
rect 675109 602986 675175 602989
rect 674668 602984 675175 602986
rect 674668 602928 675114 602984
rect 675170 602928 675175 602984
rect 674668 602926 675175 602928
rect 674668 602924 674674 602926
rect 675109 602923 675175 602926
rect 35801 601762 35867 601765
rect 35788 601760 35867 601762
rect 35788 601704 35806 601760
rect 35862 601704 35867 601760
rect 35788 601702 35867 601704
rect 35801 601699 35867 601702
rect 47761 601354 47827 601357
rect 41492 601352 47827 601354
rect 41492 601296 47766 601352
rect 47822 601296 47827 601352
rect 41492 601294 47827 601296
rect 47761 601291 47827 601294
rect 42609 600946 42675 600949
rect 41492 600944 42675 600946
rect 41492 600888 42614 600944
rect 42670 600888 42675 600944
rect 41492 600886 42675 600888
rect 42609 600883 42675 600886
rect 44633 600538 44699 600541
rect 41492 600536 44699 600538
rect 41492 600480 44638 600536
rect 44694 600480 44699 600536
rect 41492 600478 44699 600480
rect 44633 600475 44699 600478
rect 44081 600130 44147 600133
rect 41492 600128 44147 600130
rect 41492 600072 44086 600128
rect 44142 600072 44147 600128
rect 41492 600070 44147 600072
rect 44081 600067 44147 600070
rect 673545 599858 673611 599861
rect 675477 599858 675543 599861
rect 673545 599856 675543 599858
rect 673545 599800 673550 599856
rect 673606 599800 675482 599856
rect 675538 599800 675543 599856
rect 673545 599798 675543 599800
rect 673545 599795 673611 599798
rect 675477 599795 675543 599798
rect 44265 599722 44331 599725
rect 41492 599720 44331 599722
rect 41492 599664 44270 599720
rect 44326 599664 44331 599720
rect 41492 599662 44331 599664
rect 44265 599659 44331 599662
rect 41321 599314 41387 599317
rect 41308 599312 41387 599314
rect 41308 599256 41326 599312
rect 41382 599256 41387 599312
rect 41308 599254 41387 599256
rect 41321 599251 41387 599254
rect 43161 598906 43227 598909
rect 41492 598904 43227 598906
rect 41492 598848 43166 598904
rect 43222 598848 43227 598904
rect 41492 598846 43227 598848
rect 43161 598843 43227 598846
rect 40861 598498 40927 598501
rect 40861 598496 40940 598498
rect 40861 598440 40866 598496
rect 40922 598440 40940 598496
rect 40861 598438 40940 598440
rect 40861 598435 40927 598438
rect 41094 597855 41154 598060
rect 62113 597954 62179 597957
rect 62113 597952 64492 597954
rect 62113 597896 62118 597952
rect 62174 597896 64492 597952
rect 62113 597894 64492 597896
rect 62113 597891 62179 597894
rect 41045 597850 41154 597855
rect 41321 597852 41387 597855
rect 41045 597794 41050 597850
rect 41106 597794 41154 597850
rect 41045 597792 41154 597794
rect 41278 597850 41387 597852
rect 41278 597794 41326 597850
rect 41382 597794 41387 597850
rect 41045 597789 41111 597792
rect 41278 597789 41387 597794
rect 41278 597652 41338 597789
rect 41137 597274 41203 597277
rect 41124 597272 41203 597274
rect 41124 597216 41142 597272
rect 41198 597216 41203 597272
rect 41124 597214 41203 597216
rect 41137 597211 41203 597214
rect 41321 596866 41387 596869
rect 41308 596864 41387 596866
rect 41308 596808 41326 596864
rect 41382 596808 41387 596864
rect 41308 596806 41387 596808
rect 41321 596803 41387 596806
rect 42006 596458 42012 596460
rect 41492 596398 42012 596458
rect 42006 596396 42012 596398
rect 42076 596396 42082 596460
rect 41321 596050 41387 596053
rect 41308 596048 41387 596050
rect 41308 595992 41326 596048
rect 41382 595992 41387 596048
rect 41308 595990 41387 595992
rect 41321 595987 41387 595990
rect 41781 596052 41847 596053
rect 41781 596048 41828 596052
rect 41892 596050 41898 596052
rect 41781 595992 41786 596048
rect 41781 595988 41828 595992
rect 41892 595990 41938 596050
rect 41892 595988 41898 595990
rect 41781 595987 41847 595988
rect 33041 595642 33107 595645
rect 33028 595640 33107 595642
rect 33028 595584 33046 595640
rect 33102 595584 33107 595640
rect 33028 595582 33107 595584
rect 33041 595579 33107 595582
rect 35157 595234 35223 595237
rect 35157 595232 35236 595234
rect 35157 595176 35162 595232
rect 35218 595176 35236 595232
rect 35157 595174 35236 595176
rect 35157 595171 35223 595174
rect 34421 594826 34487 594829
rect 34421 594824 34500 594826
rect 34421 594768 34426 594824
rect 34482 594768 34500 594824
rect 34421 594766 34500 594768
rect 34421 594763 34487 594766
rect 31017 594418 31083 594421
rect 31004 594416 31083 594418
rect 31004 594360 31022 594416
rect 31078 594360 31083 594416
rect 31004 594358 31083 594360
rect 31017 594355 31083 594358
rect 41781 594010 41847 594013
rect 41492 594008 41847 594010
rect 41492 593952 41786 594008
rect 41842 593952 41847 594008
rect 41492 593950 41847 593952
rect 41781 593947 41847 593950
rect 36537 593602 36603 593605
rect 36524 593600 36603 593602
rect 36524 593544 36542 593600
rect 36598 593544 36603 593600
rect 36524 593542 36603 593544
rect 36537 593539 36603 593542
rect 669037 593602 669103 593605
rect 675385 593602 675451 593605
rect 669037 593600 675451 593602
rect 669037 593544 669042 593600
rect 669098 593544 675390 593600
rect 675446 593544 675451 593600
rect 669037 593542 675451 593544
rect 669037 593539 669103 593542
rect 675385 593539 675451 593542
rect 43253 593194 43319 593197
rect 41492 593192 43319 593194
rect 41492 593136 43258 593192
rect 43314 593136 43319 593192
rect 41492 593134 43319 593136
rect 43253 593131 43319 593134
rect 41781 592920 41847 592925
rect 41781 592864 41786 592920
rect 41842 592864 41847 592920
rect 41781 592859 41847 592864
rect 674097 592922 674163 592925
rect 675845 592922 675911 592925
rect 674097 592920 675911 592922
rect 674097 592864 674102 592920
rect 674158 592864 675850 592920
rect 675906 592864 675911 592920
rect 674097 592862 675911 592864
rect 674097 592859 674163 592862
rect 675845 592859 675911 592862
rect 676070 592860 676076 592924
rect 676140 592922 676146 592924
rect 678237 592922 678303 592925
rect 676140 592920 678303 592922
rect 676140 592864 678242 592920
rect 678298 592864 678303 592920
rect 676140 592862 678303 592864
rect 676140 592860 676146 592862
rect 678237 592859 678303 592862
rect 41462 592752 41522 592756
rect 41784 592752 41844 592859
rect 41462 592692 41844 592752
rect 675150 592588 675156 592652
rect 675220 592650 675226 592652
rect 676029 592650 676095 592653
rect 675220 592648 676095 592650
rect 675220 592592 676034 592648
rect 676090 592592 676095 592648
rect 675220 592590 676095 592592
rect 675220 592588 675226 592590
rect 676029 592587 676095 592590
rect 41781 592378 41847 592381
rect 41492 592376 41847 592378
rect 41492 592320 41786 592376
rect 41842 592320 41847 592376
rect 41492 592318 41847 592320
rect 41781 592315 41847 592318
rect 44633 591970 44699 591973
rect 41492 591968 44699 591970
rect 41492 591912 44638 591968
rect 44694 591912 44699 591968
rect 41492 591910 44699 591912
rect 44633 591907 44699 591910
rect 43805 591562 43871 591565
rect 41492 591560 43871 591562
rect 41492 591504 43810 591560
rect 43866 591504 43871 591560
rect 41492 591502 43871 591504
rect 43805 591499 43871 591502
rect 39990 590749 40050 591124
rect 39941 590744 40050 590749
rect 651649 590746 651715 590749
rect 39941 590688 39946 590744
rect 40002 590716 40050 590744
rect 650164 590744 651715 590746
rect 40002 590688 40020 590716
rect 39941 590686 40020 590688
rect 650164 590688 651654 590744
rect 651710 590688 651715 590744
rect 650164 590686 651715 590688
rect 39941 590683 40007 590686
rect 651649 590683 651715 590686
rect 47761 590338 47827 590341
rect 41492 590336 47827 590338
rect 41492 590280 47766 590336
rect 47822 590280 47827 590336
rect 41492 590278 47827 590280
rect 47761 590275 47827 590278
rect 40769 589660 40835 589661
rect 40718 589658 40724 589660
rect 40678 589598 40724 589658
rect 40788 589656 40835 589660
rect 40830 589600 40835 589656
rect 40718 589596 40724 589598
rect 40788 589596 40835 589600
rect 40769 589595 40835 589596
rect 40902 589460 40908 589524
rect 40972 589522 40978 589524
rect 41781 589522 41847 589525
rect 40972 589520 41847 589522
rect 40972 589464 41786 589520
rect 41842 589464 41847 589520
rect 40972 589462 41847 589464
rect 40972 589460 40978 589462
rect 41781 589459 41847 589462
rect 40585 589388 40651 589389
rect 40534 589386 40540 589388
rect 40494 589326 40540 589386
rect 40604 589384 40651 589388
rect 40646 589328 40651 589384
rect 40534 589324 40540 589326
rect 40604 589324 40651 589328
rect 40585 589323 40651 589324
rect 34421 587210 34487 587213
rect 41822 587210 41828 587212
rect 34421 587208 41828 587210
rect 34421 587152 34426 587208
rect 34482 587152 41828 587208
rect 34421 587150 41828 587152
rect 34421 587147 34487 587150
rect 41822 587148 41828 587150
rect 41892 587148 41898 587212
rect 674833 586258 674899 586261
rect 676070 586258 676076 586260
rect 674833 586256 676076 586258
rect 674833 586200 674838 586256
rect 674894 586200 676076 586256
rect 674833 586198 676076 586200
rect 674833 586195 674899 586198
rect 676070 586196 676076 586198
rect 676140 586196 676146 586260
rect 40125 584898 40191 584901
rect 41086 584898 41092 584900
rect 40125 584896 41092 584898
rect 40125 584840 40130 584896
rect 40186 584840 41092 584896
rect 40125 584838 41092 584840
rect 40125 584835 40191 584838
rect 41086 584836 41092 584838
rect 41156 584836 41162 584900
rect 41413 584898 41479 584901
rect 42006 584898 42012 584900
rect 41413 584896 42012 584898
rect 41413 584840 41418 584896
rect 41474 584840 42012 584896
rect 41413 584838 42012 584840
rect 41413 584835 41479 584838
rect 42006 584836 42012 584838
rect 42076 584836 42082 584900
rect 62113 584898 62179 584901
rect 62113 584896 64492 584898
rect 62113 584840 62118 584896
rect 62174 584840 64492 584896
rect 62113 584838 64492 584840
rect 62113 584835 62179 584838
rect 39389 584626 39455 584629
rect 40350 584626 40356 584628
rect 39389 584624 40356 584626
rect 39389 584568 39394 584624
rect 39450 584568 40356 584624
rect 39389 584566 40356 584568
rect 39389 584563 39455 584566
rect 40350 584564 40356 584566
rect 40420 584564 40426 584628
rect 41597 584626 41663 584629
rect 42558 584626 42564 584628
rect 41597 584624 42564 584626
rect 41597 584568 41602 584624
rect 41658 584568 42564 584624
rect 41597 584566 42564 584568
rect 41597 584563 41663 584566
rect 42558 584564 42564 584566
rect 42628 584564 42634 584628
rect 41781 584354 41847 584357
rect 41781 584352 41890 584354
rect 41781 584296 41786 584352
rect 41842 584296 41890 584352
rect 41781 584291 41890 584296
rect 41830 583949 41890 584291
rect 41781 583944 41890 583949
rect 41781 583888 41786 583944
rect 41842 583888 41890 583944
rect 41781 583886 41890 583888
rect 41781 583883 41847 583886
rect 41965 582588 42031 582589
rect 41965 582584 42012 582588
rect 42076 582586 42082 582588
rect 41965 582528 41970 582584
rect 41965 582524 42012 582528
rect 42076 582526 42122 582586
rect 42076 582524 42082 582526
rect 41965 582523 42031 582524
rect 42149 581226 42215 581229
rect 43437 581226 43503 581229
rect 42149 581224 43503 581226
rect 42149 581168 42154 581224
rect 42210 581168 43442 581224
rect 43498 581168 43503 581224
rect 42149 581166 43503 581168
rect 42149 581163 42215 581166
rect 43437 581163 43503 581166
rect 675477 581090 675543 581093
rect 675477 581088 676292 581090
rect 675477 581032 675482 581088
rect 675538 581032 676292 581088
rect 675477 581030 676292 581032
rect 675477 581027 675543 581030
rect 675293 580682 675359 580685
rect 675293 580680 676292 580682
rect 675293 580624 675298 580680
rect 675354 580624 676292 580680
rect 675293 580622 676292 580624
rect 675293 580619 675359 580622
rect 41086 580484 41092 580548
rect 41156 580546 41162 580548
rect 42609 580546 42675 580549
rect 41156 580544 42675 580546
rect 41156 580488 42614 580544
rect 42670 580488 42675 580544
rect 41156 580486 42675 580488
rect 41156 580484 41162 580486
rect 42609 580483 42675 580486
rect 40350 580212 40356 580276
rect 40420 580274 40426 580276
rect 41781 580274 41847 580277
rect 40420 580272 41847 580274
rect 40420 580216 41786 580272
rect 41842 580216 41847 580272
rect 40420 580214 41847 580216
rect 40420 580212 40426 580214
rect 41781 580211 41847 580214
rect 675477 580274 675543 580277
rect 675477 580272 676292 580274
rect 675477 580216 675482 580272
rect 675538 580216 676292 580272
rect 675477 580214 676292 580216
rect 675477 580211 675543 580214
rect 40902 579940 40908 580004
rect 40972 580002 40978 580004
rect 42241 580002 42307 580005
rect 40972 580000 42307 580002
rect 40972 579944 42246 580000
rect 42302 579944 42307 580000
rect 40972 579942 42307 579944
rect 40972 579940 40978 579942
rect 42241 579939 42307 579942
rect 674741 579866 674807 579869
rect 674741 579864 676292 579866
rect 674741 579808 674746 579864
rect 674802 579808 676292 579864
rect 674741 579806 676292 579808
rect 674741 579803 674807 579806
rect 675477 579458 675543 579461
rect 675477 579456 676292 579458
rect 675477 579400 675482 579456
rect 675538 579400 676292 579456
rect 675477 579398 676292 579400
rect 675477 579395 675543 579398
rect 675477 579050 675543 579053
rect 675477 579048 676292 579050
rect 675477 578992 675482 579048
rect 675538 578992 676292 579048
rect 675477 578990 676292 578992
rect 675477 578987 675543 578990
rect 675477 578642 675543 578645
rect 675477 578640 676292 578642
rect 675477 578584 675482 578640
rect 675538 578584 676292 578640
rect 675477 578582 676292 578584
rect 675477 578579 675543 578582
rect 42057 578234 42123 578237
rect 43253 578234 43319 578237
rect 42057 578232 43319 578234
rect 42057 578176 42062 578232
rect 42118 578176 43258 578232
rect 43314 578176 43319 578232
rect 42057 578174 43319 578176
rect 42057 578171 42123 578174
rect 43253 578171 43319 578174
rect 675293 578234 675359 578237
rect 675293 578232 676292 578234
rect 675293 578176 675298 578232
rect 675354 578176 676292 578232
rect 675293 578174 676292 578176
rect 675293 578171 675359 578174
rect 675293 577826 675359 577829
rect 675293 577824 676292 577826
rect 675293 577768 675298 577824
rect 675354 577768 676292 577824
rect 675293 577766 676292 577768
rect 675293 577763 675359 577766
rect 651649 577418 651715 577421
rect 650164 577416 651715 577418
rect 650164 577360 651654 577416
rect 651710 577360 651715 577416
rect 650164 577358 651715 577360
rect 651649 577355 651715 577358
rect 675293 577418 675359 577421
rect 675293 577416 676292 577418
rect 675293 577360 675298 577416
rect 675354 577360 676292 577416
rect 675293 577358 676292 577360
rect 675293 577355 675359 577358
rect 675293 577010 675359 577013
rect 675293 577008 676292 577010
rect 675293 576952 675298 577008
rect 675354 576952 676292 577008
rect 675293 576950 676292 576952
rect 675293 576947 675359 576950
rect 42333 576602 42399 576605
rect 42558 576602 42564 576604
rect 42333 576600 42564 576602
rect 42333 576544 42338 576600
rect 42394 576544 42564 576600
rect 42333 576542 42564 576544
rect 42333 576539 42399 576542
rect 42558 576540 42564 576542
rect 42628 576540 42634 576604
rect 675477 576602 675543 576605
rect 675477 576600 676292 576602
rect 675477 576544 675482 576600
rect 675538 576544 676292 576600
rect 675477 576542 676292 576544
rect 675477 576539 675543 576542
rect 676806 576404 676812 576468
rect 676876 576404 676882 576468
rect 676814 576164 676874 576404
rect 676029 575786 676095 575789
rect 676029 575784 676292 575786
rect 676029 575728 676034 575784
rect 676090 575728 676292 575784
rect 676029 575726 676292 575728
rect 676029 575723 676095 575726
rect 42057 575650 42123 575653
rect 41370 575648 42123 575650
rect 41370 575592 42062 575648
rect 42118 575592 42123 575648
rect 41370 575590 42123 575592
rect 40534 575452 40540 575516
rect 40604 575514 40610 575516
rect 41370 575514 41430 575590
rect 42057 575587 42123 575590
rect 678237 575650 678303 575653
rect 678237 575648 678346 575650
rect 678237 575592 678242 575648
rect 678298 575592 678346 575648
rect 678237 575587 678346 575592
rect 40604 575454 41430 575514
rect 40604 575452 40610 575454
rect 678286 575348 678346 575587
rect 675293 574970 675359 574973
rect 675293 574968 676292 574970
rect 675293 574912 675298 574968
rect 675354 574912 676292 574968
rect 675293 574910 676292 574912
rect 675293 574907 675359 574910
rect 40718 574636 40724 574700
rect 40788 574698 40794 574700
rect 41781 574698 41847 574701
rect 40788 574696 41847 574698
rect 40788 574640 41786 574696
rect 41842 574640 41847 574696
rect 40788 574638 41847 574640
rect 40788 574636 40794 574638
rect 41781 574635 41847 574638
rect 673637 574562 673703 574565
rect 673637 574560 676292 574562
rect 673637 574504 673642 574560
rect 673698 574504 676292 574560
rect 673637 574502 676292 574504
rect 673637 574499 673703 574502
rect 675477 574154 675543 574157
rect 675477 574152 676292 574154
rect 675477 574096 675482 574152
rect 675538 574096 676292 574152
rect 675477 574094 676292 574096
rect 675477 574091 675543 574094
rect 41454 573956 41460 574020
rect 41524 574018 41530 574020
rect 42701 574018 42767 574021
rect 41524 574016 42767 574018
rect 41524 573960 42706 574016
rect 42762 573960 42767 574016
rect 41524 573958 42767 573960
rect 41524 573956 41530 573958
rect 42701 573955 42767 573958
rect 675477 573746 675543 573749
rect 675477 573744 676292 573746
rect 675477 573688 675482 573744
rect 675538 573688 676292 573744
rect 675477 573686 676292 573688
rect 675477 573683 675543 573686
rect 674230 573276 674236 573340
rect 674300 573338 674306 573340
rect 674300 573278 676292 573338
rect 674300 573276 674306 573278
rect 675477 572930 675543 572933
rect 675477 572928 676292 572930
rect 675477 572872 675482 572928
rect 675538 572872 676292 572928
rect 675477 572870 676292 572872
rect 675477 572867 675543 572870
rect 675477 572522 675543 572525
rect 675477 572520 676292 572522
rect 675477 572464 675482 572520
rect 675538 572464 676292 572520
rect 675477 572462 676292 572464
rect 675477 572459 675543 572462
rect 41822 572188 41828 572252
rect 41892 572250 41898 572252
rect 42241 572250 42307 572253
rect 41892 572248 42307 572250
rect 41892 572192 42246 572248
rect 42302 572192 42307 572248
rect 41892 572190 42307 572192
rect 41892 572188 41898 572190
rect 42241 572187 42307 572190
rect 675477 572114 675543 572117
rect 675477 572112 676292 572114
rect 675477 572056 675482 572112
rect 675538 572056 676292 572112
rect 675477 572054 676292 572056
rect 675477 572051 675543 572054
rect 41638 571916 41644 571980
rect 41708 571978 41714 571980
rect 42425 571978 42491 571981
rect 41708 571976 42491 571978
rect 41708 571920 42430 571976
rect 42486 571920 42491 571976
rect 41708 571918 42491 571920
rect 41708 571916 41714 571918
rect 42425 571915 42491 571918
rect 683205 571978 683271 571981
rect 683205 571976 683314 571978
rect 683205 571920 683210 571976
rect 683266 571920 683314 571976
rect 683205 571915 683314 571920
rect 62113 571842 62179 571845
rect 62113 571840 64492 571842
rect 62113 571784 62118 571840
rect 62174 571784 64492 571840
rect 62113 571782 64492 571784
rect 62113 571779 62179 571782
rect 683254 571676 683314 571915
rect 674925 571570 674991 571573
rect 676990 571570 676996 571572
rect 674925 571568 676996 571570
rect 674925 571512 674930 571568
rect 674986 571512 676996 571568
rect 674925 571510 676996 571512
rect 674925 571507 674991 571510
rect 676990 571508 676996 571510
rect 677060 571508 677066 571572
rect 683438 571165 683498 571268
rect 683389 571160 683498 571165
rect 683389 571104 683394 571160
rect 683450 571104 683498 571160
rect 683389 571102 683498 571104
rect 683389 571099 683455 571102
rect 675477 570890 675543 570893
rect 675477 570888 676292 570890
rect 675477 570832 675482 570888
rect 675538 570832 676292 570888
rect 675477 570830 676292 570832
rect 675477 570827 675543 570830
rect 682886 570346 682946 570452
rect 683113 570346 683179 570349
rect 682886 570344 683179 570346
rect 682886 570288 683118 570344
rect 683174 570288 683179 570344
rect 682886 570286 683179 570288
rect 682886 570044 682946 570286
rect 683113 570283 683179 570286
rect 675477 569666 675543 569669
rect 675477 569664 676292 569666
rect 675477 569608 675482 569664
rect 675538 569608 676292 569664
rect 675477 569606 676292 569608
rect 675477 569603 675543 569606
rect 651649 564090 651715 564093
rect 650164 564088 651715 564090
rect 650164 564032 651654 564088
rect 651710 564032 651715 564088
rect 650164 564030 651715 564032
rect 651649 564027 651715 564030
rect 675385 561916 675451 561917
rect 675334 561914 675340 561916
rect 675294 561854 675340 561914
rect 675404 561912 675451 561916
rect 675446 561856 675451 561912
rect 675334 561852 675340 561854
rect 675404 561852 675451 561856
rect 675385 561851 675451 561852
rect 675477 559468 675543 559469
rect 675477 559464 675524 559468
rect 675588 559466 675594 559468
rect 675477 559408 675482 559464
rect 675477 559404 675524 559408
rect 675588 559406 675634 559466
rect 675588 559404 675594 559406
rect 675477 559403 675543 559404
rect 675753 559058 675819 559061
rect 676806 559058 676812 559060
rect 675753 559056 676812 559058
rect 675753 559000 675758 559056
rect 675814 559000 676812 559056
rect 675753 558998 676812 559000
rect 675753 558995 675819 558998
rect 676806 558996 676812 558998
rect 676876 558996 676882 559060
rect 62113 558786 62179 558789
rect 62113 558784 64492 558786
rect 62113 558728 62118 558784
rect 62174 558728 64492 558784
rect 62113 558726 64492 558728
rect 62113 558723 62179 558726
rect 43805 558514 43871 558517
rect 41492 558512 43871 558514
rect 41492 558456 43810 558512
rect 43866 558456 43871 558512
rect 41492 558454 43871 558456
rect 43805 558451 43871 558454
rect 43437 558106 43503 558109
rect 41492 558104 43503 558106
rect 41492 558048 43442 558104
rect 43498 558048 43503 558104
rect 41492 558046 43503 558048
rect 43437 558043 43503 558046
rect 41321 557698 41387 557701
rect 41308 557696 41387 557698
rect 41308 557640 41326 557696
rect 41382 557640 41387 557696
rect 41308 557638 41387 557640
rect 41321 557635 41387 557638
rect 44173 557290 44239 557293
rect 41492 557288 44239 557290
rect 41492 557232 44178 557288
rect 44234 557232 44239 557288
rect 41492 557230 44239 557232
rect 44173 557227 44239 557230
rect 44633 556882 44699 556885
rect 41492 556880 44699 556882
rect 41492 556824 44638 556880
rect 44694 556824 44699 556880
rect 41492 556822 44699 556824
rect 44633 556819 44699 556822
rect 44449 556474 44515 556477
rect 41492 556472 44515 556474
rect 41492 556416 44454 556472
rect 44510 556416 44515 556472
rect 41492 556414 44515 556416
rect 44449 556411 44515 556414
rect 40585 556066 40651 556069
rect 40572 556064 40651 556066
rect 40572 556008 40590 556064
rect 40646 556008 40651 556064
rect 40572 556006 40651 556008
rect 40585 556003 40651 556006
rect 41137 555658 41203 555661
rect 41124 555656 41203 555658
rect 41124 555600 41142 555656
rect 41198 555600 41203 555656
rect 41124 555598 41203 555600
rect 41137 555595 41203 555598
rect 42793 555250 42859 555253
rect 41492 555248 42859 555250
rect 41492 555192 42798 555248
rect 42854 555192 42859 555248
rect 41492 555190 42859 555192
rect 42793 555187 42859 555190
rect 41045 555080 41111 555083
rect 41045 555078 41154 555080
rect 41045 555022 41050 555078
rect 41106 555022 41154 555078
rect 41045 555017 41154 555022
rect 41094 554812 41154 555017
rect 43161 554434 43227 554437
rect 41492 554432 43227 554434
rect 41492 554376 43166 554432
rect 43222 554376 43227 554432
rect 41492 554374 43227 554376
rect 43161 554371 43227 554374
rect 42374 554026 42380 554028
rect 41492 553966 42380 554026
rect 42374 553964 42380 553966
rect 42444 553964 42450 554028
rect 672809 554026 672875 554029
rect 675477 554026 675543 554029
rect 672809 554024 675543 554026
rect 672809 553968 672814 554024
rect 672870 553968 675482 554024
rect 675538 553968 675543 554024
rect 672809 553966 675543 553968
rect 672809 553963 672875 553966
rect 675477 553963 675543 553966
rect 39990 553413 40050 553588
rect 39990 553408 40099 553413
rect 40953 553410 41019 553413
rect 39990 553352 40038 553408
rect 40094 553352 40099 553408
rect 39990 553350 40099 553352
rect 40033 553347 40099 553350
rect 40910 553408 41019 553410
rect 40910 553352 40958 553408
rect 41014 553352 41019 553408
rect 40910 553347 41019 553352
rect 40910 553180 40970 553347
rect 42190 552802 42196 552804
rect 41492 552742 42196 552802
rect 42190 552740 42196 552742
rect 42260 552740 42266 552804
rect 45553 552394 45619 552397
rect 41492 552392 45619 552394
rect 41492 552336 45558 552392
rect 45614 552336 45619 552392
rect 41492 552334 45619 552336
rect 45553 552331 45619 552334
rect 29637 551986 29703 551989
rect 29637 551984 29716 551986
rect 29637 551928 29642 551984
rect 29698 551928 29716 551984
rect 29637 551926 29716 551928
rect 29637 551923 29703 551926
rect 43805 551578 43871 551581
rect 41492 551576 43871 551578
rect 41492 551520 43810 551576
rect 43866 551520 43871 551576
rect 41492 551518 43871 551520
rect 43805 551515 43871 551518
rect 45185 551170 45251 551173
rect 41492 551168 45251 551170
rect 41492 551112 45190 551168
rect 45246 551112 45251 551168
rect 41492 551110 45251 551112
rect 45185 551107 45251 551110
rect 651649 550898 651715 550901
rect 650164 550896 651715 550898
rect 650164 550840 651654 550896
rect 651710 550840 651715 550896
rect 650164 550838 651715 550840
rect 651649 550835 651715 550838
rect 43989 550762 44055 550765
rect 41492 550760 44055 550762
rect 41492 550704 43994 550760
rect 44050 550704 44055 550760
rect 41492 550702 44055 550704
rect 43989 550699 44055 550702
rect 41822 550456 41828 550492
rect 41278 550428 41828 550456
rect 41892 550428 41898 550492
rect 41278 550396 41890 550428
rect 41278 550324 41338 550396
rect 675150 550292 675156 550356
rect 675220 550354 675226 550356
rect 675385 550354 675451 550357
rect 675220 550352 675451 550354
rect 675220 550296 675390 550352
rect 675446 550296 675451 550352
rect 675220 550294 675451 550296
rect 675220 550292 675226 550294
rect 675385 550291 675451 550294
rect 41873 549946 41939 549949
rect 41492 549944 41939 549946
rect 41492 549888 41878 549944
rect 41934 549888 41939 549944
rect 41492 549886 41939 549888
rect 41873 549883 41939 549886
rect 675017 549810 675083 549813
rect 675017 549808 675540 549810
rect 675017 549752 675022 549808
rect 675078 549752 675540 549808
rect 675017 549750 675540 549752
rect 675017 549747 675083 549750
rect 42057 549538 42123 549541
rect 41492 549536 42123 549538
rect 41492 549480 42062 549536
rect 42118 549480 42123 549536
rect 41492 549478 42123 549480
rect 42057 549475 42123 549478
rect 675480 549269 675540 549750
rect 675477 549264 675543 549269
rect 675477 549208 675482 549264
rect 675538 549208 675543 549264
rect 675477 549203 675543 549208
rect 42701 549130 42767 549133
rect 41492 549128 42767 549130
rect 41492 549072 42706 549128
rect 42762 549072 42767 549128
rect 41492 549070 42767 549072
rect 42701 549067 42767 549070
rect 45369 548722 45435 548725
rect 41492 548720 45435 548722
rect 41492 548664 45374 548720
rect 45430 548664 45435 548720
rect 41492 548662 45435 548664
rect 45369 548659 45435 548662
rect 42333 548314 42399 548317
rect 41492 548312 42399 548314
rect 41492 548256 42338 548312
rect 42394 548256 42399 548312
rect 41492 548254 42399 548256
rect 42333 548251 42399 548254
rect 675477 547908 675543 547909
rect 675477 547906 675524 547908
rect 675432 547904 675524 547906
rect 28766 547498 28826 547890
rect 675432 547848 675482 547904
rect 675432 547846 675524 547848
rect 675477 547844 675524 547846
rect 675588 547844 675594 547908
rect 675477 547843 675543 547844
rect 675334 547572 675340 547636
rect 675404 547634 675410 547636
rect 675753 547634 675819 547637
rect 675404 547632 675819 547634
rect 675404 547576 675758 547632
rect 675814 547576 675819 547632
rect 675404 547574 675819 547576
rect 675404 547572 675410 547574
rect 675753 547571 675819 547574
rect 31753 547498 31819 547501
rect 28766 547496 31819 547498
rect 28766 547468 31758 547496
rect 28796 547440 31758 547468
rect 31814 547440 31819 547496
rect 28796 547438 31819 547440
rect 31753 547435 31819 547438
rect 674741 547362 674807 547365
rect 675937 547362 676003 547365
rect 674741 547360 676003 547362
rect 674741 547304 674746 547360
rect 674802 547304 675942 547360
rect 675998 547304 676003 547360
rect 674741 547302 676003 547304
rect 674741 547299 674807 547302
rect 675937 547299 676003 547302
rect 43437 547090 43503 547093
rect 41492 547088 43503 547090
rect 41492 547032 43442 547088
rect 43498 547032 43503 547088
rect 41492 547030 43503 547032
rect 43437 547027 43503 547030
rect 673545 547090 673611 547093
rect 675937 547090 676003 547093
rect 673545 547088 676003 547090
rect 673545 547032 673550 547088
rect 673606 547032 675942 547088
rect 675998 547032 676003 547088
rect 673545 547030 676003 547032
rect 673545 547027 673611 547030
rect 675937 547027 676003 547030
rect 674557 546818 674623 546821
rect 676121 546818 676187 546821
rect 674557 546816 676187 546818
rect 674557 546760 674562 546816
rect 674618 546760 676126 546816
rect 676182 546760 676187 546816
rect 674557 546758 676187 546760
rect 674557 546755 674623 546758
rect 676121 546755 676187 546758
rect 41321 546410 41387 546413
rect 41638 546410 41644 546412
rect 41321 546408 41644 546410
rect 41321 546352 41326 546408
rect 41382 546352 41644 546408
rect 41321 546350 41644 546352
rect 41321 546347 41387 546350
rect 41638 546348 41644 546350
rect 41708 546348 41714 546412
rect 41454 546076 41460 546140
rect 41524 546138 41530 546140
rect 42374 546138 42380 546140
rect 41524 546078 42380 546138
rect 41524 546076 41530 546078
rect 42374 546076 42380 546078
rect 42444 546076 42450 546140
rect 40902 545804 40908 545868
rect 40972 545866 40978 545868
rect 41822 545866 41828 545868
rect 40972 545806 41828 545866
rect 40972 545804 40978 545806
rect 41822 545804 41828 545806
rect 41892 545804 41898 545868
rect 62113 545866 62179 545869
rect 675201 545868 675267 545869
rect 62113 545864 64492 545866
rect 62113 545808 62118 545864
rect 62174 545808 64492 545864
rect 62113 545806 64492 545808
rect 62113 545803 62179 545806
rect 675150 545804 675156 545868
rect 675220 545866 675267 545868
rect 675220 545864 675312 545866
rect 675262 545808 675312 545864
rect 675220 545806 675312 545808
rect 675220 545804 675267 545806
rect 675201 545803 675267 545804
rect 40718 545532 40724 545596
rect 40788 545594 40794 545596
rect 41873 545594 41939 545597
rect 40788 545592 41939 545594
rect 40788 545536 41878 545592
rect 41934 545536 41939 545592
rect 40788 545534 41939 545536
rect 40788 545532 40794 545534
rect 41873 545531 41939 545534
rect 40534 545260 40540 545324
rect 40604 545322 40610 545324
rect 42057 545322 42123 545325
rect 40604 545320 42123 545322
rect 40604 545264 42062 545320
rect 42118 545264 42123 545320
rect 40604 545262 42123 545264
rect 40604 545260 40610 545262
rect 42057 545259 42123 545262
rect 676070 545124 676076 545188
rect 676140 545186 676146 545188
rect 682377 545186 682443 545189
rect 676140 545184 682443 545186
rect 676140 545128 682382 545184
rect 682438 545128 682443 545184
rect 676140 545126 682443 545128
rect 676140 545124 676146 545126
rect 682377 545123 682443 545126
rect 40902 538188 40908 538252
rect 40972 538250 40978 538252
rect 42241 538250 42307 538253
rect 40972 538248 42307 538250
rect 40972 538192 42246 538248
rect 42302 538192 42307 538248
rect 40972 538190 42307 538192
rect 40972 538188 40978 538190
rect 42241 538187 42307 538190
rect 42057 537978 42123 537981
rect 43621 537978 43687 537981
rect 42057 537976 43687 537978
rect 42057 537920 42062 537976
rect 42118 537920 43626 537976
rect 43682 537920 43687 537976
rect 42057 537918 43687 537920
rect 42057 537915 42123 537918
rect 43621 537915 43687 537918
rect 652017 537570 652083 537573
rect 650164 537568 652083 537570
rect 650164 537512 652022 537568
rect 652078 537512 652083 537568
rect 650164 537510 652083 537512
rect 652017 537507 652083 537510
rect 42425 537026 42491 537029
rect 41370 537024 42491 537026
rect 41370 536968 42430 537024
rect 42486 536968 42491 537024
rect 41370 536966 42491 536968
rect 40718 536828 40724 536892
rect 40788 536890 40794 536892
rect 41370 536890 41430 536966
rect 42425 536963 42491 536966
rect 40788 536830 41430 536890
rect 40788 536828 40794 536830
rect 675477 536074 675543 536077
rect 676262 536074 676322 536112
rect 675477 536072 676322 536074
rect 675477 536016 675482 536072
rect 675538 536016 676322 536072
rect 675477 536014 676322 536016
rect 675477 536011 675543 536014
rect 675477 535530 675543 535533
rect 676262 535530 676322 535704
rect 675477 535528 676322 535530
rect 675477 535472 675482 535528
rect 675538 535472 676322 535528
rect 675477 535470 676322 535472
rect 675477 535467 675543 535470
rect 674557 535122 674623 535125
rect 676262 535122 676322 535296
rect 674557 535120 676322 535122
rect 674557 535064 674562 535120
rect 674618 535064 676322 535120
rect 674557 535062 676322 535064
rect 674557 535059 674623 535062
rect 675477 534850 675543 534853
rect 676262 534850 676322 534888
rect 675477 534848 676322 534850
rect 675477 534792 675482 534848
rect 675538 534792 676322 534848
rect 675477 534790 676322 534792
rect 675477 534787 675543 534790
rect 675477 534442 675543 534445
rect 676262 534442 676322 534480
rect 675477 534440 676322 534442
rect 675477 534384 675482 534440
rect 675538 534384 676322 534440
rect 675477 534382 676322 534384
rect 675477 534379 675543 534382
rect 674741 534170 674807 534173
rect 674741 534168 676322 534170
rect 674741 534112 674746 534168
rect 674802 534112 676322 534168
rect 674741 534110 676322 534112
rect 674741 534107 674807 534110
rect 676262 534072 676322 534110
rect 674557 533626 674623 533629
rect 676262 533626 676322 533664
rect 674557 533624 676322 533626
rect 674557 533568 674562 533624
rect 674618 533568 676322 533624
rect 674557 533566 676322 533568
rect 674557 533563 674623 533566
rect 40534 533292 40540 533356
rect 40604 533354 40610 533356
rect 42241 533354 42307 533357
rect 40604 533352 42307 533354
rect 40604 533296 42246 533352
rect 42302 533296 42307 533352
rect 40604 533294 42307 533296
rect 40604 533292 40610 533294
rect 42241 533291 42307 533294
rect 675477 533218 675543 533221
rect 676262 533218 676322 533256
rect 675477 533216 676322 533218
rect 675477 533160 675482 533216
rect 675538 533160 676322 533216
rect 675477 533158 676322 533160
rect 675477 533155 675543 533158
rect 675937 532878 676003 532881
rect 675937 532876 676292 532878
rect 675937 532820 675942 532876
rect 675998 532820 676292 532876
rect 675937 532818 676292 532820
rect 675937 532815 676003 532818
rect 62757 532810 62823 532813
rect 62757 532808 64492 532810
rect 62757 532752 62762 532808
rect 62818 532752 64492 532808
rect 62757 532750 64492 532752
rect 62757 532747 62823 532750
rect 41822 532612 41828 532676
rect 41892 532674 41898 532676
rect 42425 532674 42491 532677
rect 41892 532672 42491 532674
rect 41892 532616 42430 532672
rect 42486 532616 42491 532672
rect 41892 532614 42491 532616
rect 41892 532612 41898 532614
rect 42425 532611 42491 532614
rect 675477 532402 675543 532405
rect 676262 532402 676322 532440
rect 675477 532400 676322 532402
rect 675477 532344 675482 532400
rect 675538 532344 676322 532400
rect 675477 532342 676322 532344
rect 675477 532339 675543 532342
rect 674741 531994 674807 531997
rect 676262 531994 676322 532032
rect 674741 531992 676322 531994
rect 674741 531936 674746 531992
rect 674802 531936 676322 531992
rect 674741 531934 676322 531936
rect 674741 531931 674807 531934
rect 675477 531586 675543 531589
rect 676262 531586 676322 531624
rect 675477 531584 676322 531586
rect 675477 531528 675482 531584
rect 675538 531528 676322 531584
rect 675477 531526 676322 531528
rect 675477 531523 675543 531526
rect 676990 531388 676996 531452
rect 677060 531388 677066 531452
rect 676998 531216 677058 531388
rect 675477 530770 675543 530773
rect 676262 530770 676322 530808
rect 675477 530768 676322 530770
rect 675477 530712 675482 530768
rect 675538 530712 676322 530768
rect 675477 530710 676322 530712
rect 675477 530707 675543 530710
rect 682377 530634 682443 530637
rect 682334 530632 682443 530634
rect 682334 530576 682382 530632
rect 682438 530576 682443 530632
rect 682334 530571 682443 530576
rect 682334 530400 682394 530571
rect 675477 529954 675543 529957
rect 676262 529954 676322 529992
rect 675477 529952 676322 529954
rect 675477 529896 675482 529952
rect 675538 529896 676322 529952
rect 675477 529894 676322 529896
rect 675477 529891 675543 529894
rect 41638 529756 41644 529820
rect 41708 529818 41714 529820
rect 42609 529818 42675 529821
rect 41708 529816 42675 529818
rect 41708 529760 42614 529816
rect 42670 529760 42675 529816
rect 41708 529758 42675 529760
rect 41708 529756 41714 529758
rect 42609 529755 42675 529758
rect 675477 529410 675543 529413
rect 676262 529410 676322 529584
rect 675477 529408 676322 529410
rect 675477 529352 675482 529408
rect 675538 529352 676322 529408
rect 675477 529350 676322 529352
rect 675477 529347 675543 529350
rect 675477 529138 675543 529141
rect 676262 529138 676322 529176
rect 675477 529136 676322 529138
rect 675477 529080 675482 529136
rect 675538 529080 676322 529136
rect 675477 529078 676322 529080
rect 675477 529075 675543 529078
rect 674414 528804 674420 528868
rect 674484 528866 674490 528868
rect 674484 528806 676322 528866
rect 674484 528804 674490 528806
rect 676262 528768 676322 528806
rect 675477 528322 675543 528325
rect 676262 528322 676322 528360
rect 675477 528320 676322 528322
rect 675477 528264 675482 528320
rect 675538 528264 676322 528320
rect 675477 528262 676322 528264
rect 675477 528259 675543 528262
rect 683389 528186 683455 528189
rect 683389 528184 683498 528186
rect 683389 528128 683394 528184
rect 683450 528128 683498 528184
rect 683389 528123 683498 528128
rect 683438 527952 683498 528123
rect 41454 527580 41460 527644
rect 41524 527642 41530 527644
rect 41781 527642 41847 527645
rect 41524 527640 41847 527642
rect 41524 527584 41786 527640
rect 41842 527584 41847 527640
rect 41524 527582 41847 527584
rect 41524 527580 41530 527582
rect 41781 527579 41847 527582
rect 675477 527642 675543 527645
rect 675477 527640 676322 527642
rect 675477 527584 675482 527640
rect 675538 527584 676322 527640
rect 675477 527582 676322 527584
rect 675477 527579 675543 527582
rect 676262 527544 676322 527582
rect 674598 527036 674604 527100
rect 674668 527098 674674 527100
rect 676262 527098 676322 527136
rect 674668 527038 676322 527098
rect 674668 527036 674674 527038
rect 683205 526962 683271 526965
rect 683205 526960 683314 526962
rect 683205 526904 683210 526960
rect 683266 526904 683314 526960
rect 683205 526899 683314 526904
rect 683254 526728 683314 526899
rect 675477 526146 675543 526149
rect 676262 526146 676322 526320
rect 675477 526144 676322 526146
rect 675477 526088 675482 526144
rect 675538 526088 676322 526144
rect 675477 526086 676322 526088
rect 675477 526083 675543 526086
rect 673862 525812 673868 525876
rect 673932 525874 673938 525876
rect 676262 525874 676322 525912
rect 673932 525814 676322 525874
rect 673932 525812 673938 525814
rect 683113 525738 683179 525741
rect 683070 525736 683179 525738
rect 683070 525680 683118 525736
rect 683174 525680 683179 525736
rect 683070 525675 683179 525680
rect 683070 525096 683130 525675
rect 675477 524650 675543 524653
rect 676262 524650 676322 524688
rect 675477 524648 676322 524650
rect 675477 524592 675482 524648
rect 675538 524592 676322 524648
rect 675477 524590 676322 524592
rect 675477 524587 675543 524590
rect 651649 524242 651715 524245
rect 650164 524240 651715 524242
rect 650164 524184 651654 524240
rect 651710 524184 651715 524240
rect 650164 524182 651715 524184
rect 651649 524179 651715 524182
rect 40677 522746 40743 522749
rect 42517 522746 42583 522749
rect 40677 522744 42583 522746
rect 40677 522688 40682 522744
rect 40738 522688 42522 522744
rect 42578 522688 42583 522744
rect 40677 522686 42583 522688
rect 40677 522683 40743 522686
rect 42517 522683 42583 522686
rect 62113 519754 62179 519757
rect 62113 519752 64492 519754
rect 62113 519696 62118 519752
rect 62174 519696 64492 519752
rect 62113 519694 64492 519696
rect 62113 519691 62179 519694
rect 651649 511050 651715 511053
rect 650164 511048 651715 511050
rect 650164 510992 651654 511048
rect 651710 510992 651715 511048
rect 650164 510990 651715 510992
rect 651649 510987 651715 510990
rect 675109 508874 675175 508877
rect 676121 508874 676187 508877
rect 675109 508872 676187 508874
rect 675109 508816 675114 508872
rect 675170 508816 676126 508872
rect 676182 508816 676187 508872
rect 675109 508814 676187 508816
rect 675109 508811 675175 508814
rect 676121 508811 676187 508814
rect 62113 506698 62179 506701
rect 62113 506696 64492 506698
rect 62113 506640 62118 506696
rect 62174 506640 64492 506696
rect 62113 506638 64492 506640
rect 62113 506635 62179 506638
rect 676806 500924 676812 500988
rect 676876 500986 676882 500988
rect 683297 500986 683363 500989
rect 676876 500984 683363 500986
rect 676876 500928 683302 500984
rect 683358 500928 683363 500984
rect 676876 500926 683363 500928
rect 676876 500924 676882 500926
rect 683297 500923 683363 500926
rect 651649 497722 651715 497725
rect 650164 497720 651715 497722
rect 650164 497664 651654 497720
rect 651710 497664 651715 497720
rect 650164 497662 651715 497664
rect 651649 497659 651715 497662
rect 62113 493642 62179 493645
rect 62113 493640 64492 493642
rect 62113 493584 62118 493640
rect 62174 493584 64492 493640
rect 62113 493582 64492 493584
rect 62113 493579 62179 493582
rect 674741 492146 674807 492149
rect 674741 492144 676292 492146
rect 674741 492088 674746 492144
rect 674802 492088 676292 492144
rect 674741 492086 676292 492088
rect 674741 492083 674807 492086
rect 675109 491738 675175 491741
rect 675109 491736 676292 491738
rect 675109 491680 675114 491736
rect 675170 491680 676292 491736
rect 675109 491678 676292 491680
rect 675109 491675 675175 491678
rect 675477 491330 675543 491333
rect 675477 491328 676292 491330
rect 675477 491272 675482 491328
rect 675538 491272 676292 491328
rect 675477 491270 676292 491272
rect 675477 491267 675543 491270
rect 675477 490922 675543 490925
rect 675477 490920 676292 490922
rect 675477 490864 675482 490920
rect 675538 490864 676292 490920
rect 675477 490862 676292 490864
rect 675477 490859 675543 490862
rect 677409 490514 677475 490517
rect 677396 490512 677475 490514
rect 677396 490456 677414 490512
rect 677470 490456 677475 490512
rect 677396 490454 677475 490456
rect 677409 490451 677475 490454
rect 674557 490106 674623 490109
rect 674557 490104 676292 490106
rect 674557 490048 674562 490104
rect 674618 490048 676292 490104
rect 674557 490046 676292 490048
rect 674557 490043 674623 490046
rect 677225 489698 677291 489701
rect 677212 489696 677291 489698
rect 677212 489640 677230 489696
rect 677286 489640 677291 489696
rect 677212 489638 677291 489640
rect 677225 489635 677291 489638
rect 675937 489290 676003 489293
rect 675937 489288 676292 489290
rect 675937 489232 675942 489288
rect 675998 489232 676292 489288
rect 675937 489230 676292 489232
rect 675937 489227 676003 489230
rect 676029 488882 676095 488885
rect 676029 488880 676292 488882
rect 676029 488824 676034 488880
rect 676090 488824 676292 488880
rect 676029 488822 676292 488824
rect 676029 488819 676095 488822
rect 675477 488474 675543 488477
rect 675477 488472 676292 488474
rect 675477 488416 675482 488472
rect 675538 488416 676292 488472
rect 675477 488414 676292 488416
rect 675477 488411 675543 488414
rect 675937 488066 676003 488069
rect 675937 488064 676292 488066
rect 675937 488008 675942 488064
rect 675998 488008 676292 488064
rect 675937 488006 676292 488008
rect 675937 488003 676003 488006
rect 675753 487658 675819 487661
rect 675753 487656 676292 487658
rect 675753 487600 675758 487656
rect 675814 487600 676292 487656
rect 675753 487598 676292 487600
rect 675753 487595 675819 487598
rect 679617 487250 679683 487253
rect 679604 487248 679683 487250
rect 679604 487192 679622 487248
rect 679678 487192 679683 487248
rect 679604 487190 679683 487192
rect 679617 487187 679683 487190
rect 675293 486842 675359 486845
rect 675293 486840 676292 486842
rect 675293 486784 675298 486840
rect 675354 486784 676292 486840
rect 675293 486782 676292 486784
rect 675293 486779 675359 486782
rect 675477 486434 675543 486437
rect 675477 486432 676292 486434
rect 675477 486376 675482 486432
rect 675538 486376 676292 486432
rect 675477 486374 676292 486376
rect 675477 486371 675543 486374
rect 675477 486026 675543 486029
rect 675477 486024 676292 486026
rect 675477 485968 675482 486024
rect 675538 485968 676292 486024
rect 675477 485966 676292 485968
rect 675477 485963 675543 485966
rect 675477 485618 675543 485621
rect 675477 485616 676292 485618
rect 675477 485560 675482 485616
rect 675538 485560 676292 485616
rect 675477 485558 676292 485560
rect 675477 485555 675543 485558
rect 674741 485210 674807 485213
rect 674741 485208 676292 485210
rect 674741 485152 674746 485208
rect 674802 485152 676292 485208
rect 674741 485150 676292 485152
rect 674741 485147 674807 485150
rect 683297 484802 683363 484805
rect 683284 484800 683363 484802
rect 683284 484744 683302 484800
rect 683358 484744 683363 484800
rect 683284 484742 683363 484744
rect 683297 484739 683363 484742
rect 651649 484530 651715 484533
rect 650164 484528 651715 484530
rect 650164 484472 651654 484528
rect 651710 484472 651715 484528
rect 650164 484470 651715 484472
rect 651649 484467 651715 484470
rect 675477 484394 675543 484397
rect 675477 484392 676292 484394
rect 675477 484336 675482 484392
rect 675538 484336 676292 484392
rect 675477 484334 676292 484336
rect 675477 484331 675543 484334
rect 675293 483986 675359 483989
rect 675293 483984 676292 483986
rect 675293 483928 675298 483984
rect 675354 483928 676292 483984
rect 675293 483926 676292 483928
rect 675293 483923 675359 483926
rect 675293 483578 675359 483581
rect 675293 483576 676292 483578
rect 675293 483520 675298 483576
rect 675354 483520 676292 483576
rect 675293 483518 676292 483520
rect 675293 483515 675359 483518
rect 674097 483170 674163 483173
rect 674097 483168 676292 483170
rect 674097 483112 674102 483168
rect 674158 483112 676292 483168
rect 674097 483110 676292 483112
rect 674097 483107 674163 483110
rect 674373 482762 674439 482765
rect 674373 482760 676292 482762
rect 674373 482704 674378 482760
rect 674434 482704 676292 482760
rect 674373 482702 676292 482704
rect 674373 482699 674439 482702
rect 675477 482354 675543 482357
rect 675477 482352 676292 482354
rect 675477 482296 675482 482352
rect 675538 482296 676292 482352
rect 675477 482294 676292 482296
rect 675477 482291 675543 482294
rect 675477 481946 675543 481949
rect 675477 481944 676292 481946
rect 675477 481888 675482 481944
rect 675538 481888 676292 481944
rect 675477 481886 676292 481888
rect 675477 481883 675543 481886
rect 674925 481538 674991 481541
rect 674925 481536 676292 481538
rect 674925 481480 674930 481536
rect 674986 481508 676292 481536
rect 674986 481480 676322 481508
rect 674925 481478 676322 481480
rect 674925 481475 674991 481478
rect 676262 481100 676322 481478
rect 675477 480722 675543 480725
rect 675477 480720 676292 480722
rect 675477 480664 675482 480720
rect 675538 480664 676292 480720
rect 675477 480662 676292 480664
rect 675477 480659 675543 480662
rect 62113 480586 62179 480589
rect 62113 480584 64492 480586
rect 62113 480528 62118 480584
rect 62174 480528 64492 480584
rect 62113 480526 64492 480528
rect 62113 480523 62179 480526
rect 651649 471202 651715 471205
rect 650164 471200 651715 471202
rect 650164 471144 651654 471200
rect 651710 471144 651715 471200
rect 650164 471142 651715 471144
rect 651649 471139 651715 471142
rect 62113 467530 62179 467533
rect 62113 467528 64492 467530
rect 62113 467472 62118 467528
rect 62174 467472 64492 467528
rect 62113 467470 64492 467472
rect 62113 467467 62179 467470
rect 651649 457874 651715 457877
rect 650164 457872 651715 457874
rect 650164 457816 651654 457872
rect 651710 457816 651715 457872
rect 650164 457814 651715 457816
rect 651649 457811 651715 457814
rect 62757 454610 62823 454613
rect 62757 454608 64492 454610
rect 62757 454552 62762 454608
rect 62818 454552 64492 454608
rect 62757 454550 64492 454552
rect 62757 454547 62823 454550
rect 651649 444546 651715 444549
rect 650164 444544 651715 444546
rect 650164 444488 651654 444544
rect 651710 444488 651715 444544
rect 650164 444486 651715 444488
rect 651649 444483 651715 444486
rect 62113 441554 62179 441557
rect 62113 441552 64492 441554
rect 62113 441496 62118 441552
rect 62174 441496 64492 441552
rect 62113 441494 64492 441496
rect 62113 441491 62179 441494
rect 652017 431354 652083 431357
rect 650164 431352 652083 431354
rect 650164 431296 652022 431352
rect 652078 431296 652083 431352
rect 650164 431294 652083 431296
rect 652017 431291 652083 431294
rect 40677 431218 40743 431221
rect 40677 431216 40786 431218
rect 40677 431160 40682 431216
rect 40738 431160 40786 431216
rect 40677 431155 40786 431160
rect 41454 431156 41460 431220
rect 41524 431218 41530 431220
rect 42885 431218 42951 431221
rect 41524 431216 42951 431218
rect 41524 431160 42890 431216
rect 42946 431160 42951 431216
rect 41524 431158 42951 431160
rect 41524 431156 41530 431158
rect 42885 431155 42951 431158
rect 40726 430916 40786 431155
rect 41321 430538 41387 430541
rect 41308 430536 41387 430538
rect 41308 430480 41326 430536
rect 41382 430480 41387 430536
rect 41308 430478 41387 430480
rect 41321 430475 41387 430478
rect 41137 430130 41203 430133
rect 41124 430128 41203 430130
rect 41124 430072 41142 430128
rect 41198 430072 41203 430128
rect 41124 430070 41203 430072
rect 41137 430067 41203 430070
rect 40910 429487 40970 429692
rect 40910 429482 41019 429487
rect 41321 429484 41387 429487
rect 40910 429426 40958 429482
rect 41014 429426 41019 429482
rect 40910 429424 41019 429426
rect 40953 429421 41019 429424
rect 41278 429482 41387 429484
rect 41278 429426 41326 429482
rect 41382 429426 41387 429482
rect 41278 429421 41387 429426
rect 41278 429284 41338 429421
rect 44265 428906 44331 428909
rect 41492 428904 44331 428906
rect 41492 428848 44270 428904
rect 44326 428848 44331 428904
rect 41492 428846 44331 428848
rect 44265 428843 44331 428846
rect 62113 428498 62179 428501
rect 41492 428438 41890 428498
rect 41454 428198 41460 428262
rect 41524 428198 41530 428262
rect 41830 428226 41890 428438
rect 62113 428496 64492 428498
rect 62113 428440 62118 428496
rect 62174 428440 64492 428496
rect 62113 428438 64492 428440
rect 62113 428435 62179 428438
rect 42977 428226 43043 428229
rect 41830 428224 43043 428226
rect 41462 428060 41522 428198
rect 41830 428168 42982 428224
rect 43038 428168 43043 428224
rect 41830 428166 43043 428168
rect 42977 428163 43043 428166
rect 41137 427682 41203 427685
rect 41124 427680 41203 427682
rect 41124 427624 41142 427680
rect 41198 427624 41203 427680
rect 41124 427622 41203 427624
rect 41137 427619 41203 427622
rect 43161 427274 43227 427277
rect 41492 427272 43227 427274
rect 41492 427216 43166 427272
rect 43222 427216 43227 427272
rect 41492 427214 43227 427216
rect 43161 427211 43227 427214
rect 44173 426866 44239 426869
rect 41492 426864 44239 426866
rect 41492 426808 44178 426864
rect 44234 426808 44239 426864
rect 41492 426806 44239 426808
rect 44173 426803 44239 426806
rect 41822 426458 41828 426460
rect 41492 426398 41828 426458
rect 41822 426396 41828 426398
rect 41892 426396 41898 426460
rect 41137 426050 41203 426053
rect 41124 426048 41203 426050
rect 41124 425992 41142 426048
rect 41198 425992 41203 426048
rect 41124 425990 41203 425992
rect 41137 425987 41203 425990
rect 41822 425642 41828 425644
rect 41492 425582 41828 425642
rect 41822 425580 41828 425582
rect 41892 425580 41898 425644
rect 40769 425234 40835 425237
rect 40756 425232 40835 425234
rect 40756 425176 40774 425232
rect 40830 425176 40835 425232
rect 40756 425174 40835 425176
rect 40769 425171 40835 425174
rect 45553 424826 45619 424829
rect 41492 424824 45619 424826
rect 41492 424768 45558 424824
rect 45614 424768 45619 424824
rect 41492 424766 45619 424768
rect 45553 424763 45619 424766
rect 41965 424418 42031 424421
rect 41492 424416 42031 424418
rect 41492 424360 41970 424416
rect 42026 424360 42031 424416
rect 41492 424358 42031 424360
rect 41965 424355 42031 424358
rect 46933 424010 46999 424013
rect 41492 424008 46999 424010
rect 41492 423952 46938 424008
rect 46994 423952 46999 424008
rect 41492 423950 46999 423952
rect 46933 423947 46999 423950
rect 43345 423602 43411 423605
rect 41492 423600 43411 423602
rect 41492 423544 43350 423600
rect 43406 423544 43411 423600
rect 41492 423542 43411 423544
rect 43345 423539 43411 423542
rect 42793 423194 42859 423197
rect 41492 423192 42859 423194
rect 41492 423136 42798 423192
rect 42854 423136 42859 423192
rect 41492 423134 42859 423136
rect 42793 423131 42859 423134
rect 43161 422786 43227 422789
rect 41492 422784 43227 422786
rect 41492 422728 43166 422784
rect 43222 422728 43227 422784
rect 41492 422726 43227 422728
rect 43161 422723 43227 422726
rect 40726 422312 40786 422348
rect 40718 422248 40724 422312
rect 40788 422248 40794 422312
rect 42006 421970 42012 421972
rect 41492 421910 42012 421970
rect 42006 421908 42012 421910
rect 42076 421908 42082 421972
rect 45369 421562 45435 421565
rect 41492 421560 45435 421562
rect 41492 421504 45374 421560
rect 45430 421504 45435 421560
rect 41492 421502 45435 421504
rect 45369 421499 45435 421502
rect 44357 421290 44423 421293
rect 41784 421288 44423 421290
rect 41784 421232 44362 421288
rect 44418 421232 44423 421288
rect 41784 421230 44423 421232
rect 41784 421154 41844 421230
rect 44357 421227 44423 421230
rect 41492 421094 41844 421154
rect 45185 420746 45251 420749
rect 41492 420744 45251 420746
rect 41492 420688 45190 420744
rect 45246 420688 45251 420744
rect 41492 420686 45251 420688
rect 45185 420683 45251 420686
rect 41462 419930 41522 420308
rect 42241 419930 42307 419933
rect 41462 419928 42307 419930
rect 41462 419900 42246 419928
rect 41492 419872 42246 419900
rect 42302 419872 42307 419928
rect 41492 419870 42307 419872
rect 42241 419867 42307 419870
rect 42609 419522 42675 419525
rect 41492 419520 42675 419522
rect 41492 419464 42614 419520
rect 42670 419464 42675 419520
rect 41492 419462 42675 419464
rect 42609 419459 42675 419462
rect 40534 418644 40540 418708
rect 40604 418706 40610 418708
rect 42006 418706 42012 418708
rect 40604 418646 42012 418706
rect 40604 418644 40610 418646
rect 42006 418644 42012 418646
rect 42076 418644 42082 418708
rect 40769 418434 40835 418437
rect 41822 418434 41828 418436
rect 40769 418432 41828 418434
rect 40769 418376 40774 418432
rect 40830 418376 41828 418432
rect 40769 418374 41828 418376
rect 40769 418371 40835 418374
rect 41822 418372 41828 418374
rect 41892 418372 41898 418436
rect 41137 418026 41203 418029
rect 42425 418026 42491 418029
rect 651649 418026 651715 418029
rect 41137 418024 42491 418026
rect 41137 417968 41142 418024
rect 41198 417968 42430 418024
rect 42486 417968 42491 418024
rect 41137 417966 42491 417968
rect 650164 418024 651715 418026
rect 650164 417968 651654 418024
rect 651710 417968 651715 418024
rect 650164 417966 651715 417968
rect 41137 417963 41203 417966
rect 42425 417963 42491 417966
rect 651649 417963 651715 417966
rect 62113 415442 62179 415445
rect 62113 415440 64492 415442
rect 62113 415384 62118 415440
rect 62174 415384 64492 415440
rect 62113 415382 64492 415384
rect 62113 415379 62179 415382
rect 40718 407492 40724 407556
rect 40788 407554 40794 407556
rect 41781 407554 41847 407557
rect 40788 407552 41847 407554
rect 40788 407496 41786 407552
rect 41842 407496 41847 407552
rect 40788 407494 41847 407496
rect 40788 407492 40794 407494
rect 41781 407491 41847 407494
rect 651649 404698 651715 404701
rect 650164 404696 651715 404698
rect 650164 404640 651654 404696
rect 651710 404640 651715 404696
rect 650164 404638 651715 404640
rect 651649 404635 651715 404638
rect 40534 403820 40540 403884
rect 40604 403882 40610 403884
rect 41781 403882 41847 403885
rect 40604 403880 41847 403882
rect 40604 403824 41786 403880
rect 41842 403824 41847 403880
rect 40604 403822 41847 403824
rect 40604 403820 40610 403822
rect 41781 403819 41847 403822
rect 675293 403882 675359 403885
rect 675293 403880 676292 403882
rect 675293 403824 675298 403880
rect 675354 403824 676292 403880
rect 675293 403822 676292 403824
rect 675293 403819 675359 403822
rect 675477 403474 675543 403477
rect 675477 403472 676292 403474
rect 675477 403416 675482 403472
rect 675538 403416 676292 403472
rect 675477 403414 676292 403416
rect 675477 403411 675543 403414
rect 675477 403066 675543 403069
rect 675477 403064 676292 403066
rect 675477 403008 675482 403064
rect 675538 403008 676292 403064
rect 675477 403006 676292 403008
rect 675477 403003 675543 403006
rect 677409 402930 677475 402933
rect 677366 402928 677475 402930
rect 677366 402872 677414 402928
rect 677470 402872 677475 402928
rect 677366 402867 677475 402872
rect 677366 402628 677426 402867
rect 62113 402386 62179 402389
rect 62113 402384 64492 402386
rect 62113 402328 62118 402384
rect 62174 402328 64492 402384
rect 62113 402326 64492 402328
rect 62113 402323 62179 402326
rect 674649 402250 674715 402253
rect 674649 402248 676292 402250
rect 674649 402192 674654 402248
rect 674710 402192 676292 402248
rect 674649 402190 676292 402192
rect 674649 402187 674715 402190
rect 677225 402114 677291 402117
rect 677182 402112 677291 402114
rect 677182 402056 677230 402112
rect 677286 402056 677291 402112
rect 677182 402051 677291 402056
rect 41781 401980 41847 401981
rect 41781 401976 41828 401980
rect 41892 401978 41898 401980
rect 41781 401920 41786 401976
rect 41781 401916 41828 401920
rect 41892 401918 41938 401978
rect 41892 401916 41898 401918
rect 41781 401915 41847 401916
rect 677182 401812 677242 402051
rect 675477 401434 675543 401437
rect 675477 401432 676292 401434
rect 675477 401376 675482 401432
rect 675538 401376 676292 401432
rect 675477 401374 676292 401376
rect 675477 401371 675543 401374
rect 676029 401026 676095 401029
rect 676029 401024 676292 401026
rect 676029 400968 676034 401024
rect 676090 400968 676292 401024
rect 676029 400966 676292 400968
rect 676029 400963 676095 400966
rect 675477 400618 675543 400621
rect 675477 400616 676292 400618
rect 675477 400560 675482 400616
rect 675538 400560 676292 400616
rect 675477 400558 676292 400560
rect 675477 400555 675543 400558
rect 675845 400210 675911 400213
rect 675845 400208 676292 400210
rect 675845 400152 675850 400208
rect 675906 400152 676292 400208
rect 675845 400150 676292 400152
rect 675845 400147 675911 400150
rect 41454 400012 41460 400076
rect 41524 400074 41530 400076
rect 41781 400074 41847 400077
rect 41524 400072 41847 400074
rect 41524 400016 41786 400072
rect 41842 400016 41847 400072
rect 41524 400014 41847 400016
rect 41524 400012 41530 400014
rect 41781 400011 41847 400014
rect 675477 399802 675543 399805
rect 675477 399800 676292 399802
rect 675477 399744 675482 399800
rect 675538 399744 676292 399800
rect 675477 399742 676292 399744
rect 675477 399739 675543 399742
rect 675661 399394 675727 399397
rect 675661 399392 676292 399394
rect 675661 399336 675666 399392
rect 675722 399336 676292 399392
rect 675661 399334 676292 399336
rect 675661 399331 675727 399334
rect 41781 398852 41847 398853
rect 41781 398848 41828 398852
rect 41892 398850 41898 398852
rect 41781 398792 41786 398848
rect 41781 398788 41828 398792
rect 41892 398790 41938 398850
rect 41892 398788 41898 398790
rect 676070 398788 676076 398852
rect 676140 398850 676146 398852
rect 676262 398850 676322 398956
rect 676140 398790 676322 398850
rect 676140 398788 676146 398790
rect 41781 398787 41847 398788
rect 676262 398445 676322 398548
rect 676213 398440 676322 398445
rect 676213 398384 676218 398440
rect 676274 398384 676322 398440
rect 676213 398382 676322 398384
rect 676213 398379 676279 398382
rect 675109 398170 675175 398173
rect 675109 398168 676292 398170
rect 675109 398112 675114 398168
rect 675170 398112 676292 398168
rect 675109 398110 676292 398112
rect 675109 398107 675175 398110
rect 681046 397629 681106 397732
rect 680997 397624 681106 397629
rect 680997 397568 681002 397624
rect 681058 397568 681106 397624
rect 680997 397566 681106 397568
rect 680997 397563 681063 397566
rect 675293 397354 675359 397357
rect 675293 397352 676292 397354
rect 675293 397296 675298 397352
rect 675354 397296 676292 397352
rect 675293 397294 676292 397296
rect 675293 397291 675359 397294
rect 676262 396812 676322 396916
rect 676254 396748 676260 396812
rect 676324 396748 676330 396812
rect 675477 396538 675543 396541
rect 675477 396536 676292 396538
rect 675477 396480 675482 396536
rect 675538 396480 676292 396536
rect 675477 396478 676292 396480
rect 675477 396475 675543 396478
rect 674281 396130 674347 396133
rect 674281 396128 676292 396130
rect 674281 396072 674286 396128
rect 674342 396072 676292 396128
rect 674281 396070 676292 396072
rect 674281 396067 674347 396070
rect 674465 395722 674531 395725
rect 674465 395720 676292 395722
rect 674465 395664 674470 395720
rect 674526 395664 676292 395720
rect 674465 395662 676292 395664
rect 674465 395659 674531 395662
rect 676630 395180 676690 395284
rect 676622 395116 676628 395180
rect 676692 395116 676698 395180
rect 676446 394772 676506 394876
rect 676438 394708 676444 394772
rect 676508 394708 676514 394772
rect 672942 394572 672948 394636
rect 673012 394634 673018 394636
rect 673269 394634 673335 394637
rect 673012 394632 673335 394634
rect 673012 394576 673274 394632
rect 673330 394576 673335 394632
rect 673012 394574 673335 394576
rect 673012 394572 673018 394574
rect 673269 394571 673335 394574
rect 675477 394498 675543 394501
rect 675477 394496 676292 394498
rect 675477 394440 675482 394496
rect 675538 394440 676292 394496
rect 675477 394438 676292 394440
rect 675477 394435 675543 394438
rect 675477 394090 675543 394093
rect 675477 394088 676292 394090
rect 675477 394032 675482 394088
rect 675538 394032 676292 394088
rect 675477 394030 676292 394032
rect 675477 394027 675543 394030
rect 674097 393682 674163 393685
rect 674097 393680 676292 393682
rect 674097 393624 674102 393680
rect 674158 393624 676292 393680
rect 674097 393622 676292 393624
rect 674097 393619 674163 393622
rect 683070 392733 683130 393244
rect 683021 392728 683130 392733
rect 683021 392672 683026 392728
rect 683082 392672 683130 392728
rect 683021 392670 683130 392672
rect 683021 392667 683087 392670
rect 675477 392458 675543 392461
rect 675477 392456 676292 392458
rect 675477 392400 675482 392456
rect 675538 392400 676292 392456
rect 675477 392398 676292 392400
rect 675477 392395 675543 392398
rect 651649 391506 651715 391509
rect 650164 391504 651715 391506
rect 650164 391448 651654 391504
rect 651710 391448 651715 391504
rect 650164 391446 651715 391448
rect 651649 391443 651715 391446
rect 675886 389812 675892 389876
rect 675956 389874 675962 389876
rect 683021 389874 683087 389877
rect 675956 389872 683087 389874
rect 675956 389816 683026 389872
rect 683082 389816 683087 389872
rect 675956 389814 683087 389816
rect 675956 389812 675962 389814
rect 683021 389811 683087 389814
rect 62113 389330 62179 389333
rect 62113 389328 64492 389330
rect 62113 389272 62118 389328
rect 62174 389272 64492 389328
rect 62113 389270 64492 389272
rect 62113 389267 62179 389270
rect 675702 388452 675708 388516
rect 675772 388514 675778 388516
rect 680997 388514 681063 388517
rect 675772 388512 681063 388514
rect 675772 388456 681002 388512
rect 681058 388456 681063 388512
rect 675772 388454 681063 388456
rect 675772 388452 675778 388454
rect 680997 388451 681063 388454
rect 35390 387565 35450 387668
rect 35341 387560 35450 387565
rect 35341 387504 35346 387560
rect 35402 387504 35450 387560
rect 35341 387502 35450 387504
rect 39941 387562 40007 387565
rect 43621 387562 43687 387565
rect 39941 387560 43687 387562
rect 39941 387504 39946 387560
rect 40002 387504 43626 387560
rect 43682 387504 43687 387560
rect 39941 387502 43687 387504
rect 35341 387499 35407 387502
rect 39941 387499 40007 387502
rect 43621 387499 43687 387502
rect 35574 387157 35634 387260
rect 35525 387152 35634 387157
rect 35801 387154 35867 387157
rect 35525 387096 35530 387152
rect 35586 387096 35634 387152
rect 35525 387094 35634 387096
rect 35758 387152 35867 387154
rect 35758 387096 35806 387152
rect 35862 387096 35867 387152
rect 35525 387091 35591 387094
rect 35758 387091 35867 387096
rect 40125 387154 40191 387157
rect 43989 387154 44055 387157
rect 40125 387152 44055 387154
rect 40125 387096 40130 387152
rect 40186 387096 43994 387152
rect 44050 387096 44055 387152
rect 40125 387094 44055 387096
rect 40125 387091 40191 387094
rect 43989 387091 44055 387094
rect 35758 386852 35818 387091
rect 40309 386746 40375 386749
rect 47945 386746 48011 386749
rect 40309 386744 48011 386746
rect 40309 386688 40314 386744
rect 40370 386688 47950 386744
rect 48006 386688 48011 386744
rect 40309 386686 48011 386688
rect 40309 386683 40375 386686
rect 47945 386683 48011 386686
rect 35758 386341 35818 386444
rect 35758 386336 35867 386341
rect 35758 386280 35806 386336
rect 35862 386280 35867 386336
rect 35758 386278 35867 386280
rect 35801 386275 35867 386278
rect 35390 385933 35450 386036
rect 35341 385928 35450 385933
rect 35341 385872 35346 385928
rect 35402 385872 35450 385928
rect 35341 385870 35450 385872
rect 35341 385867 35407 385870
rect 35574 385525 35634 385628
rect 35525 385520 35634 385525
rect 35801 385522 35867 385525
rect 35525 385464 35530 385520
rect 35586 385464 35634 385520
rect 35525 385462 35634 385464
rect 35758 385520 35867 385522
rect 35758 385464 35806 385520
rect 35862 385464 35867 385520
rect 35525 385459 35591 385462
rect 35758 385459 35867 385464
rect 35758 385220 35818 385459
rect 39573 385114 39639 385117
rect 43069 385114 43135 385117
rect 39573 385112 43135 385114
rect 39573 385056 39578 385112
rect 39634 385056 43074 385112
rect 43130 385056 43135 385112
rect 39573 385054 43135 385056
rect 39573 385051 39639 385054
rect 43069 385051 43135 385054
rect 675753 384978 675819 384981
rect 676254 384978 676260 384980
rect 675753 384976 676260 384978
rect 675753 384920 675758 384976
rect 675814 384920 676260 384976
rect 675753 384918 676260 384920
rect 675753 384915 675819 384918
rect 676254 384916 676260 384918
rect 676324 384916 676330 384980
rect 35574 384709 35634 384812
rect 35574 384704 35683 384709
rect 35574 384648 35622 384704
rect 35678 384648 35683 384704
rect 35574 384646 35683 384648
rect 35617 384643 35683 384646
rect 35758 384301 35818 384404
rect 35758 384296 35867 384301
rect 35758 384240 35806 384296
rect 35862 384240 35867 384296
rect 35758 384238 35867 384240
rect 35801 384235 35867 384238
rect 35758 383893 35818 383996
rect 35758 383888 35867 383893
rect 35758 383832 35806 383888
rect 35862 383832 35867 383888
rect 35758 383830 35867 383832
rect 35801 383827 35867 383830
rect 39665 383890 39731 383893
rect 43989 383890 44055 383893
rect 39665 383888 44055 383890
rect 39665 383832 39670 383888
rect 39726 383832 43994 383888
rect 44050 383832 44055 383888
rect 39665 383830 44055 383832
rect 39665 383827 39731 383830
rect 43989 383827 44055 383830
rect 35390 383485 35450 383588
rect 35341 383480 35450 383485
rect 35341 383424 35346 383480
rect 35402 383424 35450 383480
rect 35341 383422 35450 383424
rect 35341 383419 35407 383422
rect 35574 383077 35634 383180
rect 35525 383072 35634 383077
rect 35801 383074 35867 383077
rect 35525 383016 35530 383072
rect 35586 383016 35634 383072
rect 35525 383014 35634 383016
rect 35758 383072 35867 383074
rect 35758 383016 35806 383072
rect 35862 383016 35867 383072
rect 35525 383011 35591 383014
rect 35758 383011 35867 383016
rect 35758 382772 35818 383011
rect 35758 382261 35818 382364
rect 35758 382256 35867 382261
rect 35758 382200 35806 382256
rect 35862 382200 35867 382256
rect 35758 382198 35867 382200
rect 35801 382195 35867 382198
rect 40033 382258 40099 382261
rect 41454 382258 41460 382260
rect 40033 382256 41460 382258
rect 40033 382200 40038 382256
rect 40094 382200 41460 382256
rect 40033 382198 41460 382200
rect 40033 382195 40099 382198
rect 41454 382196 41460 382198
rect 41524 382196 41530 382260
rect 35574 381853 35634 381956
rect 35574 381848 35683 381853
rect 35574 381792 35622 381848
rect 35678 381792 35683 381848
rect 35574 381790 35683 381792
rect 35617 381787 35683 381790
rect 41413 381850 41479 381853
rect 44173 381850 44239 381853
rect 41413 381848 44239 381850
rect 41413 381792 41418 381848
rect 41474 381792 44178 381848
rect 44234 381792 44239 381848
rect 41413 381790 44239 381792
rect 41413 381787 41479 381790
rect 44173 381787 44239 381790
rect 32446 381445 32506 381548
rect 32397 381440 32506 381445
rect 35801 381442 35867 381445
rect 32397 381384 32402 381440
rect 32458 381384 32506 381440
rect 32397 381382 32506 381384
rect 35758 381440 35867 381442
rect 35758 381384 35806 381440
rect 35862 381384 35867 381440
rect 32397 381379 32463 381382
rect 35758 381379 35867 381384
rect 35758 381140 35818 381379
rect 35574 380629 35634 380732
rect 35574 380624 35683 380629
rect 35574 380568 35622 380624
rect 35678 380568 35683 380624
rect 35574 380566 35683 380568
rect 35617 380563 35683 380566
rect 39849 380626 39915 380629
rect 42793 380626 42859 380629
rect 39849 380624 42859 380626
rect 39849 380568 39854 380624
rect 39910 380568 42798 380624
rect 42854 380568 42859 380624
rect 39849 380566 42859 380568
rect 39849 380563 39915 380566
rect 42793 380563 42859 380566
rect 675753 380626 675819 380629
rect 676438 380626 676444 380628
rect 675753 380624 676444 380626
rect 675753 380568 675758 380624
rect 675814 380568 676444 380624
rect 675753 380566 676444 380568
rect 675753 380563 675819 380566
rect 676438 380564 676444 380566
rect 676508 380564 676514 380628
rect 35390 380221 35450 380324
rect 35390 380216 35499 380221
rect 35801 380218 35867 380221
rect 35390 380160 35438 380216
rect 35494 380160 35499 380216
rect 35390 380158 35499 380160
rect 35433 380155 35499 380158
rect 35758 380216 35867 380218
rect 35758 380160 35806 380216
rect 35862 380160 35867 380216
rect 35758 380155 35867 380160
rect 40033 380218 40099 380221
rect 41638 380218 41644 380220
rect 40033 380216 41644 380218
rect 40033 380160 40038 380216
rect 40094 380160 41644 380216
rect 40033 380158 41644 380160
rect 40033 380155 40099 380158
rect 41638 380156 41644 380158
rect 41708 380156 41714 380220
rect 35758 379916 35818 380155
rect 41045 379810 41111 379813
rect 45369 379810 45435 379813
rect 41045 379808 45435 379810
rect 41045 379752 41050 379808
rect 41106 379752 45374 379808
rect 45430 379752 45435 379808
rect 41045 379750 45435 379752
rect 41045 379747 41111 379750
rect 45369 379747 45435 379750
rect 40910 379404 40970 379508
rect 40902 379340 40908 379404
rect 40972 379340 40978 379404
rect 35758 378997 35818 379100
rect 35758 378992 35867 378997
rect 35758 378936 35806 378992
rect 35862 378936 35867 378992
rect 35758 378934 35867 378936
rect 35801 378931 35867 378934
rect 40217 378994 40283 378997
rect 41822 378994 41828 378996
rect 40217 378992 41828 378994
rect 40217 378936 40222 378992
rect 40278 378936 41828 378992
rect 40217 378934 41828 378936
rect 40217 378931 40283 378934
rect 41822 378932 41828 378934
rect 41892 378932 41898 378996
rect 675753 378724 675819 378725
rect 675702 378722 675708 378724
rect 40542 378588 40602 378692
rect 675662 378662 675708 378722
rect 675772 378720 675819 378724
rect 675814 378664 675819 378720
rect 675702 378660 675708 378662
rect 675772 378660 675819 378664
rect 675753 378659 675819 378660
rect 40534 378524 40540 378588
rect 40604 378524 40610 378588
rect 40726 378180 40786 378284
rect 40718 378116 40724 378180
rect 40788 378116 40794 378180
rect 41505 378178 41571 378181
rect 44541 378178 44607 378181
rect 651649 378178 651715 378181
rect 41505 378176 44607 378178
rect 41505 378120 41510 378176
rect 41566 378120 44546 378176
rect 44602 378120 44607 378176
rect 41505 378118 44607 378120
rect 650164 378176 651715 378178
rect 650164 378120 651654 378176
rect 651710 378120 651715 378176
rect 650164 378118 651715 378120
rect 41505 378115 41571 378118
rect 44541 378115 44607 378118
rect 651649 378115 651715 378118
rect 672533 378042 672599 378045
rect 674782 378042 674788 378044
rect 672533 378040 674788 378042
rect 672533 377984 672538 378040
rect 672594 377984 674788 378040
rect 672533 377982 674788 377984
rect 672533 377979 672599 377982
rect 674782 377980 674788 377982
rect 674852 377980 674858 378044
rect 35574 377773 35634 377876
rect 35574 377768 35683 377773
rect 35574 377712 35622 377768
rect 35678 377712 35683 377768
rect 35574 377710 35683 377712
rect 35617 377707 35683 377710
rect 39757 377770 39823 377773
rect 43437 377770 43503 377773
rect 39757 377768 43503 377770
rect 39757 377712 39762 377768
rect 39818 377712 43442 377768
rect 43498 377712 43503 377768
rect 39757 377710 43503 377712
rect 39757 377707 39823 377710
rect 43437 377707 43503 377710
rect 35758 377365 35818 377468
rect 35758 377360 35867 377365
rect 35758 377304 35806 377360
rect 35862 377304 35867 377360
rect 35758 377302 35867 377304
rect 35801 377299 35867 377302
rect 39573 377362 39639 377365
rect 43621 377362 43687 377365
rect 39573 377360 43687 377362
rect 39573 377304 39578 377360
rect 39634 377304 43626 377360
rect 43682 377304 43687 377360
rect 39573 377302 43687 377304
rect 39573 377299 39639 377302
rect 43621 377299 43687 377302
rect 675753 377362 675819 377365
rect 676622 377362 676628 377364
rect 675753 377360 676628 377362
rect 675753 377304 675758 377360
rect 675814 377304 676628 377360
rect 675753 377302 676628 377304
rect 675753 377299 675819 377302
rect 676622 377300 676628 377302
rect 676692 377300 676698 377364
rect 28766 376549 28826 377060
rect 41505 376954 41571 376957
rect 44357 376954 44423 376957
rect 41505 376952 44423 376954
rect 41505 376896 41510 376952
rect 41566 376896 44362 376952
rect 44418 376896 44423 376952
rect 41505 376894 44423 376896
rect 41505 376891 41571 376894
rect 44357 376891 44423 376894
rect 28766 376544 28875 376549
rect 28766 376488 28814 376544
rect 28870 376488 28875 376544
rect 28766 376486 28875 376488
rect 28809 376483 28875 376486
rect 62113 376274 62179 376277
rect 62113 376272 64492 376274
rect 35758 376141 35818 376244
rect 62113 376216 62118 376272
rect 62174 376216 64492 376272
rect 62113 376214 64492 376216
rect 62113 376211 62179 376214
rect 35758 376136 35867 376141
rect 35758 376080 35806 376136
rect 35862 376080 35867 376136
rect 35758 376078 35867 376080
rect 35801 376075 35867 376078
rect 675293 375050 675359 375053
rect 676070 375050 676076 375052
rect 675293 375048 676076 375050
rect 675293 374992 675298 375048
rect 675354 374992 676076 375048
rect 675293 374990 676076 374992
rect 675293 374987 675359 374990
rect 676070 374988 676076 374990
rect 676140 374988 676146 375052
rect 675661 373010 675727 373013
rect 675886 373010 675892 373012
rect 675661 373008 675892 373010
rect 675661 372952 675666 373008
rect 675722 372952 675892 373008
rect 675661 372950 675892 372952
rect 675661 372947 675727 372950
rect 675886 372948 675892 372950
rect 675956 372948 675962 373012
rect 674782 372540 674788 372604
rect 674852 372602 674858 372604
rect 675109 372602 675175 372605
rect 674852 372600 675175 372602
rect 674852 372544 675114 372600
rect 675170 372544 675175 372600
rect 674852 372542 675175 372544
rect 674852 372540 674858 372542
rect 675109 372539 675175 372542
rect 42057 369746 42123 369749
rect 42793 369746 42859 369749
rect 42057 369744 42859 369746
rect 42057 369688 42062 369744
rect 42118 369688 42798 369744
rect 42854 369688 42859 369744
rect 42057 369686 42859 369688
rect 42057 369683 42123 369686
rect 42793 369683 42859 369686
rect 40902 365604 40908 365668
rect 40972 365666 40978 365668
rect 41781 365666 41847 365669
rect 40972 365664 41847 365666
rect 40972 365608 41786 365664
rect 41842 365608 41847 365664
rect 40972 365606 41847 365608
rect 40972 365604 40978 365606
rect 41781 365603 41847 365606
rect 42057 364986 42123 364989
rect 44357 364986 44423 364989
rect 42057 364984 44423 364986
rect 42057 364928 42062 364984
rect 42118 364928 44362 364984
rect 44418 364928 44423 364984
rect 42057 364926 44423 364928
rect 42057 364923 42123 364926
rect 44357 364923 44423 364926
rect 651649 364850 651715 364853
rect 650164 364848 651715 364850
rect 650164 364792 651654 364848
rect 651710 364792 651715 364848
rect 650164 364790 651715 364792
rect 651649 364787 651715 364790
rect 40718 363700 40724 363764
rect 40788 363762 40794 363764
rect 41781 363762 41847 363765
rect 40788 363760 41847 363762
rect 40788 363704 41786 363760
rect 41842 363704 41847 363760
rect 40788 363702 41847 363704
rect 40788 363700 40794 363702
rect 41781 363699 41847 363702
rect 62941 363354 63007 363357
rect 62941 363352 64492 363354
rect 62941 363296 62946 363352
rect 63002 363296 64492 363352
rect 62941 363294 64492 363296
rect 62941 363291 63007 363294
rect 40534 360572 40540 360636
rect 40604 360634 40610 360636
rect 41781 360634 41847 360637
rect 40604 360632 41847 360634
rect 40604 360576 41786 360632
rect 41842 360576 41847 360632
rect 40604 360574 41847 360576
rect 40604 360572 40610 360574
rect 41781 360571 41847 360574
rect 41873 358732 41939 358733
rect 41822 358730 41828 358732
rect 41782 358670 41828 358730
rect 41892 358728 41939 358732
rect 41934 358672 41939 358728
rect 41822 358668 41828 358670
rect 41892 358668 41939 358672
rect 41873 358667 41939 358668
rect 675293 358730 675359 358733
rect 675293 358728 676292 358730
rect 675293 358672 675298 358728
rect 675354 358672 676292 358728
rect 675293 358670 676292 358672
rect 675293 358667 675359 358670
rect 675109 358322 675175 358325
rect 675109 358320 676292 358322
rect 675109 358264 675114 358320
rect 675170 358264 676292 358320
rect 675109 358262 676292 358264
rect 675109 358259 675175 358262
rect 675477 357914 675543 357917
rect 675477 357912 676292 357914
rect 675477 357856 675482 357912
rect 675538 357856 676292 357912
rect 675477 357854 676292 357856
rect 675477 357851 675543 357854
rect 674649 357506 674715 357509
rect 674649 357504 676292 357506
rect 674649 357448 674654 357504
rect 674710 357448 676292 357504
rect 674649 357446 676292 357448
rect 674649 357443 674715 357446
rect 675477 357098 675543 357101
rect 675477 357096 676292 357098
rect 675477 357040 675482 357096
rect 675538 357040 676292 357096
rect 675477 357038 676292 357040
rect 675477 357035 675543 357038
rect 41454 356900 41460 356964
rect 41524 356962 41530 356964
rect 41781 356962 41847 356965
rect 41524 356960 41847 356962
rect 41524 356904 41786 356960
rect 41842 356904 41847 356960
rect 41524 356902 41847 356904
rect 41524 356900 41530 356902
rect 41781 356899 41847 356902
rect 674741 356690 674807 356693
rect 674741 356688 676292 356690
rect 674741 356632 674746 356688
rect 674802 356632 676292 356688
rect 674741 356630 676292 356632
rect 674741 356627 674807 356630
rect 674649 356282 674715 356285
rect 674649 356280 676292 356282
rect 674649 356224 674654 356280
rect 674710 356224 676292 356280
rect 674649 356222 676292 356224
rect 674649 356219 674715 356222
rect 675477 355874 675543 355877
rect 675477 355872 676292 355874
rect 675477 355816 675482 355872
rect 675538 355816 676292 355872
rect 675477 355814 676292 355816
rect 675477 355811 675543 355814
rect 41965 355740 42031 355741
rect 41965 355736 42012 355740
rect 42076 355738 42082 355740
rect 41965 355680 41970 355736
rect 41965 355676 42012 355680
rect 42076 355678 42122 355738
rect 42076 355676 42082 355678
rect 41965 355675 42031 355676
rect 675293 355466 675359 355469
rect 675293 355464 676292 355466
rect 675293 355408 675298 355464
rect 675354 355408 676292 355464
rect 675293 355406 676292 355408
rect 675293 355403 675359 355406
rect 675477 355058 675543 355061
rect 675477 355056 676292 355058
rect 675477 355000 675482 355056
rect 675538 355000 676292 355056
rect 675477 354998 676292 355000
rect 675477 354995 675543 354998
rect 675109 354650 675175 354653
rect 675109 354648 676292 354650
rect 675109 354592 675114 354648
rect 675170 354592 676292 354648
rect 675109 354590 676292 354592
rect 675109 354587 675175 354590
rect 675334 354180 675340 354244
rect 675404 354242 675410 354244
rect 675404 354182 676292 354242
rect 675404 354180 675410 354182
rect 675293 353834 675359 353837
rect 675293 353832 676292 353834
rect 675293 353776 675298 353832
rect 675354 353776 676292 353832
rect 675293 353774 676292 353776
rect 675293 353771 675359 353774
rect 675477 353426 675543 353429
rect 675477 353424 676292 353426
rect 675477 353368 675482 353424
rect 675538 353368 676292 353424
rect 675477 353366 676292 353368
rect 675477 353363 675543 353366
rect 675518 352956 675524 353020
rect 675588 353018 675594 353020
rect 675588 352958 676292 353018
rect 675588 352956 675594 352958
rect 675477 352610 675543 352613
rect 675477 352608 676292 352610
rect 675477 352552 675482 352608
rect 675538 352552 676292 352608
rect 675477 352550 676292 352552
rect 675477 352547 675543 352550
rect 675702 352140 675708 352204
rect 675772 352202 675778 352204
rect 675772 352142 676292 352202
rect 675772 352140 675778 352142
rect 675886 351732 675892 351796
rect 675956 351794 675962 351796
rect 675956 351734 676292 351794
rect 675956 351732 675962 351734
rect 651649 351658 651715 351661
rect 650164 351656 651715 351658
rect 650164 351600 651654 351656
rect 651710 351600 651715 351656
rect 650164 351598 651715 351600
rect 651649 351595 651715 351598
rect 675293 351386 675359 351389
rect 675293 351384 676292 351386
rect 675293 351328 675298 351384
rect 675354 351328 676292 351384
rect 675293 351326 676292 351328
rect 675293 351323 675359 351326
rect 675886 350916 675892 350980
rect 675956 350978 675962 350980
rect 675956 350918 676292 350978
rect 675956 350916 675962 350918
rect 675477 350570 675543 350573
rect 675477 350568 676292 350570
rect 675477 350512 675482 350568
rect 675538 350512 676292 350568
rect 675477 350510 676292 350512
rect 675477 350507 675543 350510
rect 62757 350298 62823 350301
rect 62757 350296 64492 350298
rect 62757 350240 62762 350296
rect 62818 350240 64492 350296
rect 62757 350238 64492 350240
rect 62757 350235 62823 350238
rect 675886 350100 675892 350164
rect 675956 350162 675962 350164
rect 675956 350102 676292 350162
rect 675956 350100 675962 350102
rect 674465 349754 674531 349757
rect 674465 349752 676292 349754
rect 674465 349696 674470 349752
rect 674526 349696 676292 349752
rect 674465 349694 676292 349696
rect 674465 349691 674531 349694
rect 675477 349346 675543 349349
rect 675477 349344 676292 349346
rect 675477 349288 675482 349344
rect 675538 349288 676292 349344
rect 675477 349286 676292 349288
rect 675477 349283 675543 349286
rect 675477 348938 675543 348941
rect 675477 348936 676292 348938
rect 675477 348880 675482 348936
rect 675538 348880 676292 348936
rect 675477 348878 676292 348880
rect 675477 348875 675543 348878
rect 674281 348530 674347 348533
rect 674281 348528 676292 348530
rect 674281 348472 674286 348528
rect 674342 348472 676292 348528
rect 674281 348470 676292 348472
rect 674281 348467 674347 348470
rect 683070 347717 683130 348092
rect 683070 347712 683179 347717
rect 683070 347684 683118 347712
rect 683100 347656 683118 347684
rect 683174 347656 683179 347712
rect 683100 347654 683179 347656
rect 683113 347651 683179 347654
rect 675477 347306 675543 347309
rect 675477 347304 676292 347306
rect 675477 347248 675482 347304
rect 675538 347248 676292 347304
rect 675477 347246 676292 347248
rect 675477 347243 675543 347246
rect 40401 345810 40467 345813
rect 45185 345810 45251 345813
rect 40401 345808 45251 345810
rect 40401 345752 40406 345808
rect 40462 345752 45190 345808
rect 45246 345752 45251 345808
rect 40401 345750 45251 345752
rect 40401 345747 40467 345750
rect 45185 345747 45251 345750
rect 675334 345476 675340 345540
rect 675404 345538 675410 345540
rect 675886 345538 675892 345540
rect 675404 345478 675892 345538
rect 675404 345476 675410 345478
rect 675886 345476 675892 345478
rect 675956 345476 675962 345540
rect 671797 345268 671863 345269
rect 671797 345266 671844 345268
rect 671752 345264 671844 345266
rect 671752 345208 671802 345264
rect 671752 345206 671844 345208
rect 671797 345204 671844 345206
rect 671908 345204 671914 345268
rect 671797 345203 671863 345204
rect 39757 344994 39823 344997
rect 43989 344994 44055 344997
rect 39757 344992 44055 344994
rect 39757 344936 39762 344992
rect 39818 344936 43994 344992
rect 44050 344936 44055 344992
rect 39757 344934 44055 344936
rect 39757 344931 39823 344934
rect 43989 344931 44055 344934
rect 670969 344994 671035 344997
rect 671286 344994 671292 344996
rect 670969 344992 671292 344994
rect 670969 344936 670974 344992
rect 671030 344936 671292 344992
rect 670969 344934 671292 344936
rect 670969 344931 671035 344934
rect 671286 344932 671292 344934
rect 671356 344932 671362 344996
rect 39573 344722 39639 344725
rect 43805 344722 43871 344725
rect 39573 344720 43871 344722
rect 39573 344664 39578 344720
rect 39634 344664 43810 344720
rect 43866 344664 43871 344720
rect 39573 344662 43871 344664
rect 39573 344659 39639 344662
rect 43805 344659 43871 344662
rect 35390 344317 35450 344556
rect 35341 344312 35450 344317
rect 35617 344314 35683 344317
rect 35341 344256 35346 344312
rect 35402 344256 35450 344312
rect 35341 344254 35450 344256
rect 35574 344312 35683 344314
rect 35574 344256 35622 344312
rect 35678 344256 35683 344312
rect 35341 344251 35407 344254
rect 35574 344251 35683 344256
rect 35574 344148 35634 344251
rect 35801 343906 35867 343909
rect 35758 343904 35867 343906
rect 35758 343848 35806 343904
rect 35862 343848 35867 343904
rect 35758 343843 35867 343848
rect 35758 343740 35818 343843
rect 39573 343498 39639 343501
rect 43253 343498 43319 343501
rect 39573 343496 43319 343498
rect 39573 343440 39578 343496
rect 39634 343440 43258 343496
rect 43314 343440 43319 343496
rect 39573 343438 43319 343440
rect 39573 343435 39639 343438
rect 43253 343435 43319 343438
rect 35390 343093 35450 343332
rect 35341 343088 35450 343093
rect 35341 343032 35346 343088
rect 35402 343032 35450 343088
rect 35341 343030 35450 343032
rect 39941 343090 40007 343093
rect 42977 343090 43043 343093
rect 39941 343088 43043 343090
rect 39941 343032 39946 343088
rect 40002 343032 42982 343088
rect 43038 343032 43043 343088
rect 39941 343030 43043 343032
rect 35341 343027 35407 343030
rect 39941 343027 40007 343030
rect 42977 343027 43043 343030
rect 35574 342685 35634 342924
rect 35525 342680 35634 342685
rect 35801 342682 35867 342685
rect 35525 342624 35530 342680
rect 35586 342624 35634 342680
rect 35525 342622 35634 342624
rect 35758 342680 35867 342682
rect 35758 342624 35806 342680
rect 35862 342624 35867 342680
rect 35525 342619 35591 342622
rect 35758 342619 35867 342624
rect 35758 342516 35818 342619
rect 40309 342274 40375 342277
rect 43253 342274 43319 342277
rect 40309 342272 43319 342274
rect 40309 342216 40314 342272
rect 40370 342216 43258 342272
rect 43314 342216 43319 342272
rect 40309 342214 43319 342216
rect 40309 342211 40375 342214
rect 43253 342211 43319 342214
rect 669221 342138 669287 342141
rect 675845 342138 675911 342141
rect 669221 342136 675911 342138
rect 35574 341869 35634 342108
rect 669221 342080 669226 342136
rect 669282 342080 675850 342136
rect 675906 342080 675911 342136
rect 669221 342078 675911 342080
rect 669221 342075 669287 342078
rect 675845 342075 675911 342078
rect 35574 341864 35683 341869
rect 35574 341808 35622 341864
rect 35678 341808 35683 341864
rect 35574 341806 35683 341808
rect 35617 341803 35683 341806
rect 35758 341461 35818 341700
rect 35758 341456 35867 341461
rect 35758 341400 35806 341456
rect 35862 341400 35867 341456
rect 35758 341398 35867 341400
rect 35801 341395 35867 341398
rect 35574 341053 35634 341292
rect 35574 341048 35683 341053
rect 35574 340992 35622 341048
rect 35678 340992 35683 341048
rect 35574 340990 35683 340992
rect 35617 340987 35683 340990
rect 40309 341050 40375 341053
rect 42885 341050 42951 341053
rect 40309 341048 42951 341050
rect 40309 340992 40314 341048
rect 40370 340992 42890 341048
rect 42946 340992 42951 341048
rect 40309 340990 42951 340992
rect 40309 340987 40375 340990
rect 42885 340987 42951 340990
rect 35758 340645 35818 340884
rect 35758 340640 35867 340645
rect 35758 340584 35806 340640
rect 35862 340584 35867 340640
rect 35758 340582 35867 340584
rect 35801 340579 35867 340582
rect 35574 340237 35634 340476
rect 671838 340444 671844 340508
rect 671908 340506 671914 340508
rect 673269 340506 673335 340509
rect 671908 340504 673335 340506
rect 671908 340448 673274 340504
rect 673330 340448 673335 340504
rect 671908 340446 673335 340448
rect 671908 340444 671914 340446
rect 673269 340443 673335 340446
rect 675753 340370 675819 340373
rect 676622 340370 676628 340372
rect 675753 340368 676628 340370
rect 675753 340312 675758 340368
rect 675814 340312 676628 340368
rect 675753 340310 676628 340312
rect 675753 340307 675819 340310
rect 676622 340308 676628 340310
rect 676692 340308 676698 340372
rect 35574 340232 35683 340237
rect 35574 340176 35622 340232
rect 35678 340176 35683 340232
rect 35574 340174 35683 340176
rect 35617 340171 35683 340174
rect 41462 339828 41522 340068
rect 41454 339764 41460 339828
rect 41524 339764 41530 339828
rect 41278 339554 41338 339660
rect 41822 339554 41828 339556
rect 41278 339494 41828 339554
rect 41822 339492 41828 339494
rect 41892 339492 41898 339556
rect 675661 339418 675727 339421
rect 675886 339418 675892 339420
rect 675661 339416 675892 339418
rect 675661 339360 675666 339416
rect 675722 339360 675892 339416
rect 675661 339358 675892 339360
rect 675661 339355 675727 339358
rect 675886 339356 675892 339358
rect 675956 339356 675962 339420
rect 35574 339013 35634 339252
rect 35574 339008 35683 339013
rect 35574 338952 35622 339008
rect 35678 338952 35683 339008
rect 35574 338950 35683 338952
rect 35617 338947 35683 338950
rect 39573 339010 39639 339013
rect 44173 339010 44239 339013
rect 39573 339008 44239 339010
rect 39573 338952 39578 339008
rect 39634 338952 44178 339008
rect 44234 338952 44239 339008
rect 39573 338950 44239 338952
rect 39573 338947 39639 338950
rect 44173 338947 44239 338950
rect 35801 338602 35867 338605
rect 35758 338600 35867 338602
rect 35758 338544 35806 338600
rect 35862 338544 35867 338600
rect 35758 338539 35867 338544
rect 41462 338602 41522 338844
rect 41638 338602 41644 338604
rect 41462 338542 41644 338602
rect 41638 338540 41644 338542
rect 41708 338540 41714 338604
rect 35758 338436 35818 338539
rect 651649 338330 651715 338333
rect 650164 338328 651715 338330
rect 650164 338272 651654 338328
rect 651710 338272 651715 338328
rect 650164 338270 651715 338272
rect 651649 338267 651715 338270
rect 41505 338194 41571 338197
rect 47025 338194 47091 338197
rect 41505 338192 47091 338194
rect 41505 338136 41510 338192
rect 41566 338136 47030 338192
rect 47086 338136 47091 338192
rect 41505 338134 47091 338136
rect 41505 338131 41571 338134
rect 47025 338131 47091 338134
rect 35758 337789 35818 338028
rect 35758 337784 35867 337789
rect 675569 337788 675635 337789
rect 675518 337786 675524 337788
rect 35758 337728 35806 337784
rect 35862 337728 35867 337784
rect 35758 337726 35867 337728
rect 675478 337726 675524 337786
rect 675588 337784 675635 337788
rect 675630 337728 675635 337784
rect 35801 337723 35867 337726
rect 675518 337724 675524 337726
rect 675588 337724 675635 337728
rect 675569 337723 675635 337724
rect 40542 337380 40602 337620
rect 40534 337316 40540 337380
rect 40604 337316 40610 337380
rect 62113 337242 62179 337245
rect 62113 337240 64492 337242
rect 35574 336973 35634 337212
rect 62113 337184 62118 337240
rect 62174 337184 64492 337240
rect 62113 337182 64492 337184
rect 62113 337179 62179 337182
rect 35525 336968 35634 336973
rect 35801 336970 35867 336973
rect 35525 336912 35530 336968
rect 35586 336912 35634 336968
rect 35525 336910 35634 336912
rect 35758 336968 35867 336970
rect 35758 336912 35806 336968
rect 35862 336912 35867 336968
rect 35525 336907 35591 336910
rect 35758 336907 35867 336912
rect 40033 336970 40099 336973
rect 43437 336970 43503 336973
rect 40033 336968 43503 336970
rect 40033 336912 40038 336968
rect 40094 336912 43442 336968
rect 43498 336912 43503 336968
rect 40033 336910 43503 336912
rect 40033 336907 40099 336910
rect 43437 336907 43503 336910
rect 35758 336804 35818 336907
rect 675753 336698 675819 336701
rect 676438 336698 676444 336700
rect 675753 336696 676444 336698
rect 675753 336640 675758 336696
rect 675814 336640 676444 336696
rect 675753 336638 676444 336640
rect 675753 336635 675819 336638
rect 676438 336636 676444 336638
rect 676508 336636 676514 336700
rect 35617 336154 35683 336157
rect 40726 336156 40786 336396
rect 35574 336152 35683 336154
rect 35574 336096 35622 336152
rect 35678 336096 35683 336152
rect 35574 336091 35683 336096
rect 40718 336092 40724 336156
rect 40788 336092 40794 336156
rect 35574 335988 35634 336091
rect 35801 335746 35867 335749
rect 35758 335744 35867 335746
rect 35758 335688 35806 335744
rect 35862 335688 35867 335744
rect 35758 335683 35867 335688
rect 35758 335580 35818 335683
rect 39665 335338 39731 335341
rect 43989 335338 44055 335341
rect 39665 335336 44055 335338
rect 39665 335280 39670 335336
rect 39726 335280 43994 335336
rect 44050 335280 44055 335336
rect 39665 335278 44055 335280
rect 39665 335275 39731 335278
rect 43989 335275 44055 335278
rect 35390 334933 35450 335172
rect 35390 334928 35499 334933
rect 35801 334930 35867 334933
rect 35390 334872 35438 334928
rect 35494 334872 35499 334928
rect 35390 334870 35499 334872
rect 35433 334867 35499 334870
rect 35758 334928 35867 334930
rect 35758 334872 35806 334928
rect 35862 334872 35867 334928
rect 35758 334867 35867 334872
rect 40309 334930 40375 334933
rect 43621 334930 43687 334933
rect 40309 334928 43687 334930
rect 40309 334872 40314 334928
rect 40370 334872 43626 334928
rect 43682 334872 43687 334928
rect 40309 334870 43687 334872
rect 40309 334867 40375 334870
rect 43621 334867 43687 334870
rect 35758 334764 35818 334867
rect 35617 334522 35683 334525
rect 35574 334520 35683 334522
rect 35574 334464 35622 334520
rect 35678 334464 35683 334520
rect 35574 334459 35683 334464
rect 35574 334356 35634 334459
rect 39573 334114 39639 334117
rect 44633 334114 44699 334117
rect 39573 334112 44699 334114
rect 39573 334056 39578 334112
rect 39634 334056 44638 334112
rect 44694 334056 44699 334112
rect 39573 334054 44699 334056
rect 39573 334051 39639 334054
rect 44633 334051 44699 334054
rect 35574 333301 35634 333948
rect 40309 333706 40375 333709
rect 44449 333706 44515 333709
rect 40309 333704 44515 333706
rect 40309 333648 40314 333704
rect 40370 333648 44454 333704
rect 44510 333648 44515 333704
rect 40309 333646 44515 333648
rect 40309 333643 40375 333646
rect 44449 333643 44515 333646
rect 35574 333296 35683 333301
rect 35574 333240 35622 333296
rect 35678 333240 35683 333296
rect 35574 333238 35683 333240
rect 35617 333235 35683 333238
rect 35758 332893 35818 333132
rect 35758 332888 35867 332893
rect 35758 332832 35806 332888
rect 35862 332832 35867 332888
rect 35758 332830 35867 332832
rect 35801 332827 35867 332830
rect 675753 332346 675819 332349
rect 676254 332346 676260 332348
rect 675753 332344 676260 332346
rect 675753 332288 675758 332344
rect 675814 332288 676260 332344
rect 675753 332286 676260 332288
rect 675753 332283 675819 332286
rect 676254 332284 676260 332286
rect 676324 332284 676330 332348
rect 39573 330578 39639 330581
rect 45553 330578 45619 330581
rect 39573 330576 45619 330578
rect 39573 330520 39578 330576
rect 39634 330520 45558 330576
rect 45614 330520 45619 330576
rect 39573 330518 45619 330520
rect 39573 330515 39639 330518
rect 45553 330515 45619 330518
rect 675753 326906 675819 326909
rect 676070 326906 676076 326908
rect 675753 326904 676076 326906
rect 675753 326848 675758 326904
rect 675814 326848 676076 326904
rect 675753 326846 676076 326848
rect 675753 326843 675819 326846
rect 676070 326844 676076 326846
rect 676140 326844 676146 326908
rect 651649 325002 651715 325005
rect 650164 325000 651715 325002
rect 650164 324944 651654 325000
rect 651710 324944 651715 325000
rect 650164 324942 651715 324944
rect 651649 324939 651715 324942
rect 41781 324868 41847 324869
rect 41781 324864 41828 324868
rect 41892 324866 41898 324868
rect 41781 324808 41786 324864
rect 41781 324804 41828 324808
rect 41892 324806 41938 324866
rect 41892 324804 41898 324806
rect 41781 324803 41847 324804
rect 62113 324186 62179 324189
rect 62113 324184 64492 324186
rect 62113 324128 62118 324184
rect 62174 324128 64492 324184
rect 62113 324126 64492 324128
rect 62113 324123 62179 324126
rect 40718 322764 40724 322828
rect 40788 322826 40794 322828
rect 41781 322826 41847 322829
rect 40788 322824 41847 322826
rect 40788 322768 41786 322824
rect 41842 322768 41847 322824
rect 40788 322766 41847 322768
rect 40788 322764 40794 322766
rect 41781 322763 41847 322766
rect 41781 315620 41847 315621
rect 41781 315616 41828 315620
rect 41892 315618 41898 315620
rect 41781 315560 41786 315616
rect 41781 315556 41828 315560
rect 41892 315558 41938 315618
rect 41892 315556 41898 315558
rect 41781 315555 41847 315556
rect 41454 313652 41460 313716
rect 41524 313714 41530 313716
rect 41781 313714 41847 313717
rect 41524 313712 41847 313714
rect 41524 313656 41786 313712
rect 41842 313656 41847 313712
rect 41524 313654 41847 313656
rect 41524 313652 41530 313654
rect 41781 313651 41847 313654
rect 675477 313714 675543 313717
rect 675477 313712 676292 313714
rect 675477 313656 675482 313712
rect 675538 313656 676292 313712
rect 675477 313654 676292 313656
rect 675477 313651 675543 313654
rect 675477 313306 675543 313309
rect 675477 313304 676292 313306
rect 675477 313248 675482 313304
rect 675538 313248 676292 313304
rect 675477 313246 676292 313248
rect 675477 313243 675543 313246
rect 40534 312972 40540 313036
rect 40604 313034 40610 313036
rect 41781 313034 41847 313037
rect 40604 313032 41847 313034
rect 40604 312976 41786 313032
rect 41842 312976 41847 313032
rect 40604 312974 41847 312976
rect 40604 312972 40610 312974
rect 41781 312971 41847 312974
rect 675293 312898 675359 312901
rect 675293 312896 676292 312898
rect 675293 312840 675298 312896
rect 675354 312840 676292 312896
rect 675293 312838 676292 312840
rect 675293 312835 675359 312838
rect 675477 312490 675543 312493
rect 675477 312488 676292 312490
rect 675477 312432 675482 312488
rect 675538 312432 676292 312488
rect 675477 312430 676292 312432
rect 675477 312427 675543 312430
rect 675477 312082 675543 312085
rect 675477 312080 676292 312082
rect 675477 312024 675482 312080
rect 675538 312024 676292 312080
rect 675477 312022 676292 312024
rect 675477 312019 675543 312022
rect 652017 311810 652083 311813
rect 650164 311808 652083 311810
rect 650164 311752 652022 311808
rect 652078 311752 652083 311808
rect 650164 311750 652083 311752
rect 652017 311747 652083 311750
rect 674649 311674 674715 311677
rect 674649 311672 676292 311674
rect 674649 311616 674654 311672
rect 674710 311616 676292 311672
rect 674649 311614 676292 311616
rect 674649 311611 674715 311614
rect 675477 311266 675543 311269
rect 675477 311264 676292 311266
rect 675477 311208 675482 311264
rect 675538 311208 676292 311264
rect 675477 311206 676292 311208
rect 675477 311203 675543 311206
rect 62113 311130 62179 311133
rect 62113 311128 64492 311130
rect 62113 311072 62118 311128
rect 62174 311072 64492 311128
rect 62113 311070 64492 311072
rect 62113 311067 62179 311070
rect 675293 310858 675359 310861
rect 675293 310856 676292 310858
rect 675293 310800 675298 310856
rect 675354 310800 676292 310856
rect 675293 310798 676292 310800
rect 675293 310795 675359 310798
rect 675293 310450 675359 310453
rect 675293 310448 676292 310450
rect 675293 310392 675298 310448
rect 675354 310392 676292 310448
rect 675293 310390 676292 310392
rect 675293 310387 675359 310390
rect 675477 310042 675543 310045
rect 675477 310040 676292 310042
rect 675477 309984 675482 310040
rect 675538 309984 676292 310040
rect 675477 309982 676292 309984
rect 675477 309979 675543 309982
rect 675477 309634 675543 309637
rect 675477 309632 676292 309634
rect 675477 309576 675482 309632
rect 675538 309576 676292 309632
rect 675477 309574 676292 309576
rect 675477 309571 675543 309574
rect 675477 309226 675543 309229
rect 675477 309224 676292 309226
rect 675477 309168 675482 309224
rect 675538 309168 676292 309224
rect 675477 309166 676292 309168
rect 675477 309163 675543 309166
rect 675886 308756 675892 308820
rect 675956 308818 675962 308820
rect 675956 308758 676292 308818
rect 675956 308756 675962 308758
rect 676029 308410 676095 308413
rect 676029 308408 676292 308410
rect 676029 308352 676034 308408
rect 676090 308352 676292 308408
rect 676029 308350 676292 308352
rect 676029 308347 676095 308350
rect 675017 308002 675083 308005
rect 675017 308000 676292 308002
rect 675017 307944 675022 308000
rect 675078 307944 676292 308000
rect 675017 307942 676292 307944
rect 675017 307939 675083 307942
rect 675017 307594 675083 307597
rect 675017 307592 676292 307594
rect 675017 307536 675022 307592
rect 675078 307536 676292 307592
rect 675017 307534 676292 307536
rect 675017 307531 675083 307534
rect 678237 307186 678303 307189
rect 678237 307184 678316 307186
rect 678237 307128 678242 307184
rect 678298 307128 678316 307184
rect 678237 307126 678316 307128
rect 678237 307123 678303 307126
rect 680997 306778 681063 306781
rect 680997 306776 681076 306778
rect 680997 306720 681002 306776
rect 681058 306720 681076 306776
rect 680997 306718 681076 306720
rect 680997 306715 681063 306718
rect 674465 306370 674531 306373
rect 674465 306368 676292 306370
rect 674465 306312 674470 306368
rect 674526 306312 676292 306368
rect 674465 306310 676292 306312
rect 674465 306307 674531 306310
rect 676397 305962 676463 305965
rect 676397 305960 676476 305962
rect 676397 305904 676402 305960
rect 676458 305904 676476 305960
rect 676397 305902 676476 305904
rect 676397 305899 676463 305902
rect 675477 305554 675543 305557
rect 675477 305552 676292 305554
rect 675477 305496 675482 305552
rect 675538 305496 676292 305552
rect 675477 305494 676292 305496
rect 675477 305491 675543 305494
rect 676032 305086 676292 305146
rect 676032 304978 676092 305086
rect 676032 304916 676076 304978
rect 676070 304914 676076 304916
rect 676140 304914 676146 304978
rect 676029 304738 676095 304741
rect 676029 304736 676292 304738
rect 676029 304680 676034 304736
rect 676090 304680 676292 304736
rect 676029 304678 676292 304680
rect 676029 304675 676095 304678
rect 674649 304330 674715 304333
rect 674649 304328 676292 304330
rect 674649 304272 674654 304328
rect 674710 304272 676292 304328
rect 674649 304270 676292 304272
rect 674649 304267 674715 304270
rect 675477 303922 675543 303925
rect 675477 303920 676292 303922
rect 675477 303864 675482 303920
rect 675538 303864 676292 303920
rect 675477 303862 676292 303864
rect 675477 303859 675543 303862
rect 675477 303514 675543 303517
rect 675477 303512 676292 303514
rect 675477 303456 675482 303512
rect 675538 303456 676292 303512
rect 675477 303454 676292 303456
rect 675477 303451 675543 303454
rect 676029 302972 676095 302973
rect 676029 302970 676076 302972
rect 675984 302968 676076 302970
rect 675984 302912 676034 302968
rect 675984 302910 676076 302912
rect 676029 302908 676076 302910
rect 676140 302908 676146 302972
rect 676029 302907 676095 302908
rect 677182 302698 677242 303076
rect 683113 302698 683179 302701
rect 677182 302696 683179 302698
rect 677182 302668 683118 302696
rect 677212 302640 683118 302668
rect 683174 302640 683179 302696
rect 677212 302638 683179 302640
rect 683113 302635 683179 302638
rect 675477 302290 675543 302293
rect 675477 302288 676292 302290
rect 675477 302232 675482 302288
rect 675538 302232 676292 302288
rect 675477 302230 676292 302232
rect 675477 302227 675543 302230
rect 43805 301610 43871 301613
rect 41094 301608 43871 301610
rect 41094 301552 43810 301608
rect 43866 301552 43871 301608
rect 41094 301550 43871 301552
rect 41094 301308 41154 301550
rect 43805 301547 43871 301550
rect 676397 301612 676463 301613
rect 676397 301608 676444 301612
rect 676508 301610 676514 301612
rect 676397 301552 676402 301608
rect 676397 301548 676444 301552
rect 676508 301550 676554 301610
rect 676508 301548 676514 301550
rect 676397 301547 676463 301548
rect 45369 300930 45435 300933
rect 41492 300928 45435 300930
rect 41492 300872 45374 300928
rect 45430 300872 45435 300928
rect 41492 300870 45435 300872
rect 45369 300867 45435 300870
rect 675477 300658 675543 300661
rect 676213 300658 676279 300661
rect 675477 300656 676279 300658
rect 675477 300600 675482 300656
rect 675538 300600 676218 300656
rect 676274 300600 676279 300656
rect 675477 300598 676279 300600
rect 675477 300595 675543 300598
rect 676213 300595 676279 300598
rect 48129 300522 48195 300525
rect 41492 300520 48195 300522
rect 41492 300464 48134 300520
rect 48190 300464 48195 300520
rect 41492 300462 48195 300464
rect 48129 300459 48195 300462
rect 43253 300114 43319 300117
rect 41492 300112 43319 300114
rect 41492 300056 43258 300112
rect 43314 300056 43319 300112
rect 41492 300054 43319 300056
rect 43253 300051 43319 300054
rect 44541 299706 44607 299709
rect 41492 299704 44607 299706
rect 41492 299648 44546 299704
rect 44602 299648 44607 299704
rect 41492 299646 44607 299648
rect 44541 299643 44607 299646
rect 675886 299372 675892 299436
rect 675956 299434 675962 299436
rect 680353 299434 680419 299437
rect 675956 299432 680419 299434
rect 675956 299376 680358 299432
rect 680414 299376 680419 299432
rect 675956 299374 680419 299376
rect 675956 299372 675962 299374
rect 680353 299371 680419 299374
rect 41137 299298 41203 299301
rect 41124 299296 41203 299298
rect 41124 299240 41142 299296
rect 41198 299240 41203 299296
rect 41124 299238 41203 299240
rect 41137 299235 41203 299238
rect 42701 298890 42767 298893
rect 41492 298888 42767 298890
rect 41492 298832 42706 298888
rect 42762 298832 42767 298888
rect 41492 298830 42767 298832
rect 42701 298827 42767 298830
rect 40953 298482 41019 298485
rect 652201 298482 652267 298485
rect 40940 298480 41019 298482
rect 40940 298424 40958 298480
rect 41014 298424 41019 298480
rect 40940 298422 41019 298424
rect 650164 298480 652267 298482
rect 650164 298424 652206 298480
rect 652262 298424 652267 298480
rect 650164 298422 652267 298424
rect 40953 298419 41019 298422
rect 652201 298419 652267 298422
rect 62113 298210 62179 298213
rect 62113 298208 64492 298210
rect 62113 298152 62118 298208
rect 62174 298152 64492 298208
rect 62113 298150 64492 298152
rect 62113 298147 62179 298150
rect 40953 298074 41019 298077
rect 40940 298072 41019 298074
rect 40940 298016 40958 298072
rect 41014 298016 41019 298072
rect 40940 298014 41019 298016
rect 40953 298011 41019 298014
rect 44173 297666 44239 297669
rect 41492 297664 44239 297666
rect 41492 297608 44178 297664
rect 44234 297608 44239 297664
rect 41492 297606 44239 297608
rect 44173 297603 44239 297606
rect 675702 297332 675708 297396
rect 675772 297394 675778 297396
rect 678237 297394 678303 297397
rect 675772 297392 678303 297394
rect 675772 297336 678242 297392
rect 678298 297336 678303 297392
rect 675772 297334 678303 297336
rect 675772 297332 675778 297334
rect 678237 297331 678303 297334
rect 43253 297258 43319 297261
rect 41492 297256 43319 297258
rect 41492 297200 43258 297256
rect 43314 297200 43319 297256
rect 41492 297198 43319 297200
rect 43253 297195 43319 297198
rect 41822 296850 41828 296852
rect 41492 296790 41828 296850
rect 41822 296788 41828 296790
rect 41892 296788 41898 296852
rect 675518 296516 675524 296580
rect 675588 296578 675594 296580
rect 675845 296578 675911 296581
rect 675588 296576 675911 296578
rect 675588 296520 675850 296576
rect 675906 296520 675911 296576
rect 675588 296518 675911 296520
rect 675588 296516 675594 296518
rect 675845 296515 675911 296518
rect 42006 296442 42012 296444
rect 41492 296382 42012 296442
rect 42006 296380 42012 296382
rect 42076 296380 42082 296444
rect 45553 296034 45619 296037
rect 41492 296032 45619 296034
rect 41492 295976 45558 296032
rect 45614 295976 45619 296032
rect 41492 295974 45619 295976
rect 45553 295971 45619 295974
rect 42057 295626 42123 295629
rect 41492 295624 42123 295626
rect 41492 295568 42062 295624
rect 42118 295568 42123 295624
rect 41492 295566 42123 295568
rect 42057 295563 42123 295566
rect 675569 295356 675635 295357
rect 675518 295292 675524 295356
rect 675588 295354 675635 295356
rect 675588 295352 675680 295354
rect 675630 295296 675680 295352
rect 675588 295294 675680 295296
rect 675588 295292 675635 295294
rect 675569 295291 675635 295292
rect 41781 295218 41847 295221
rect 41492 295216 41847 295218
rect 41492 295160 41786 295216
rect 41842 295160 41847 295216
rect 41492 295158 41847 295160
rect 41781 295155 41847 295158
rect 41781 294946 41847 294949
rect 45737 294946 45803 294949
rect 41781 294944 45803 294946
rect 41781 294888 41786 294944
rect 41842 294888 45742 294944
rect 45798 294888 45803 294944
rect 41781 294886 45803 294888
rect 41781 294883 41847 294886
rect 45737 294883 45803 294886
rect 35157 294810 35223 294813
rect 35157 294808 35236 294810
rect 35157 294752 35162 294808
rect 35218 294752 35236 294808
rect 35157 294750 35236 294752
rect 35157 294747 35223 294750
rect 45921 294402 45987 294405
rect 41492 294400 45987 294402
rect 41492 294344 45926 294400
rect 45982 294344 45987 294400
rect 41492 294342 45987 294344
rect 45921 294339 45987 294342
rect 43069 293994 43135 293997
rect 41492 293992 43135 293994
rect 41492 293936 43074 293992
rect 43130 293936 43135 293992
rect 41492 293934 43135 293936
rect 43069 293931 43135 293934
rect 41781 293586 41847 293589
rect 41492 293584 41847 293586
rect 41492 293528 41786 293584
rect 41842 293528 41847 293584
rect 41492 293526 41847 293528
rect 41781 293523 41847 293526
rect 43989 293178 44055 293181
rect 41492 293176 44055 293178
rect 41492 293120 43994 293176
rect 44050 293120 44055 293176
rect 41492 293118 44055 293120
rect 43989 293115 44055 293118
rect 40493 292592 40559 292593
rect 40726 292592 40786 292740
rect 40493 292590 40540 292592
rect 40448 292588 40540 292590
rect 40448 292532 40498 292588
rect 40448 292530 40540 292532
rect 40493 292528 40540 292530
rect 40604 292528 40610 292592
rect 40718 292528 40724 292592
rect 40788 292528 40794 292592
rect 40902 292528 40908 292592
rect 40972 292528 40978 292592
rect 40493 292527 40559 292528
rect 40910 292332 40970 292528
rect 41822 292300 41828 292364
rect 41892 292362 41898 292364
rect 42057 292362 42123 292365
rect 41892 292360 42123 292362
rect 41892 292304 42062 292360
rect 42118 292304 42123 292360
rect 41892 292302 42123 292304
rect 41892 292300 41898 292302
rect 42057 292299 42123 292302
rect 41492 291894 41844 291954
rect 41784 291818 41844 291894
rect 44173 291818 44239 291821
rect 41784 291816 44239 291818
rect 41784 291760 44178 291816
rect 44234 291760 44239 291816
rect 41784 291758 44239 291760
rect 44173 291755 44239 291758
rect 44357 291546 44423 291549
rect 41492 291544 44423 291546
rect 41492 291488 44362 291544
rect 44418 291488 44423 291544
rect 41492 291486 44423 291488
rect 44357 291483 44423 291486
rect 675753 291546 675819 291549
rect 676438 291546 676444 291548
rect 675753 291544 676444 291546
rect 675753 291488 675758 291544
rect 675814 291488 676444 291544
rect 675753 291486 676444 291488
rect 675753 291483 675819 291486
rect 676438 291484 676444 291486
rect 676508 291484 676514 291548
rect 42885 291138 42951 291141
rect 41492 291136 42951 291138
rect 41492 291080 42890 291136
rect 42946 291080 42951 291136
rect 41492 291078 42951 291080
rect 42885 291075 42951 291078
rect 675753 291002 675819 291005
rect 676254 291002 676260 291004
rect 675753 291000 676260 291002
rect 675753 290944 675758 291000
rect 675814 290944 676260 291000
rect 675753 290942 676260 290944
rect 675753 290939 675819 290942
rect 676254 290940 676260 290942
rect 676324 290940 676330 291004
rect 41137 290730 41203 290733
rect 41124 290728 41203 290730
rect 41124 290672 41142 290728
rect 41198 290672 41203 290728
rect 41124 290670 41203 290672
rect 41137 290667 41203 290670
rect 40953 290322 41019 290325
rect 40940 290320 41019 290322
rect 40940 290264 40958 290320
rect 41014 290264 41019 290320
rect 40940 290262 41019 290264
rect 40953 290259 41019 290262
rect 41781 290050 41847 290053
rect 43805 290050 43871 290053
rect 41781 290048 43871 290050
rect 41781 289992 41786 290048
rect 41842 289992 43810 290048
rect 43866 289992 43871 290048
rect 41781 289990 43871 289992
rect 41781 289987 41847 289990
rect 43805 289987 43871 289990
rect 41278 289833 41338 289884
rect 41278 289828 41387 289833
rect 41278 289772 41326 289828
rect 41382 289772 41387 289828
rect 41278 289770 41387 289772
rect 41321 289767 41387 289770
rect 675753 287058 675819 287061
rect 676622 287058 676628 287060
rect 675753 287056 676628 287058
rect 675753 287000 675758 287056
rect 675814 287000 676628 287056
rect 675753 286998 676628 287000
rect 675753 286995 675819 286998
rect 676622 286996 676628 286998
rect 676692 286996 676698 287060
rect 673361 286514 673427 286517
rect 675385 286514 675451 286517
rect 673361 286512 675451 286514
rect 673361 286456 673366 286512
rect 673422 286456 675390 286512
rect 675446 286456 675451 286512
rect 673361 286454 675451 286456
rect 673361 286451 673427 286454
rect 675385 286451 675451 286454
rect 673085 285562 673151 285565
rect 675109 285562 675175 285565
rect 673085 285560 675175 285562
rect 673085 285504 673090 285560
rect 673146 285504 675114 285560
rect 675170 285504 675175 285560
rect 673085 285502 675175 285504
rect 673085 285499 673151 285502
rect 675109 285499 675175 285502
rect 651649 285290 651715 285293
rect 650164 285288 651715 285290
rect 650164 285232 651654 285288
rect 651710 285232 651715 285288
rect 650164 285230 651715 285232
rect 651649 285227 651715 285230
rect 62757 285154 62823 285157
rect 62757 285152 64492 285154
rect 62757 285096 62762 285152
rect 62818 285096 64492 285152
rect 62757 285094 64492 285096
rect 62757 285091 62823 285094
rect 675753 283658 675819 283661
rect 676070 283658 676076 283660
rect 675753 283656 676076 283658
rect 675753 283600 675758 283656
rect 675814 283600 676076 283656
rect 675753 283598 676076 283600
rect 675753 283595 675819 283598
rect 676070 283596 676076 283598
rect 676140 283596 676146 283660
rect 675661 282842 675727 282845
rect 675886 282842 675892 282844
rect 675661 282840 675892 282842
rect 675661 282784 675666 282840
rect 675722 282784 675892 282840
rect 675661 282782 675892 282784
rect 675661 282779 675727 282782
rect 675886 282780 675892 282782
rect 675956 282780 675962 282844
rect 675661 281620 675727 281621
rect 675661 281616 675708 281620
rect 675772 281618 675778 281620
rect 675661 281560 675666 281616
rect 675661 281556 675708 281560
rect 675772 281558 675818 281618
rect 675772 281556 675778 281558
rect 675661 281555 675727 281556
rect 41965 281484 42031 281485
rect 41965 281480 42012 281484
rect 42076 281482 42082 281484
rect 41965 281424 41970 281480
rect 41965 281420 42012 281424
rect 42076 281422 42122 281482
rect 42076 281420 42082 281422
rect 41965 281419 42031 281420
rect 670969 278762 671035 278765
rect 671286 278762 671292 278764
rect 670969 278760 671292 278762
rect 670969 278704 670974 278760
rect 671030 278704 671292 278760
rect 670969 278702 671292 278704
rect 670969 278699 671035 278702
rect 671286 278700 671292 278702
rect 671356 278700 671362 278764
rect 672533 278762 672599 278765
rect 672942 278762 672948 278764
rect 672533 278760 672948 278762
rect 672533 278704 672538 278760
rect 672594 278704 672948 278760
rect 672533 278702 672948 278704
rect 672533 278699 672599 278702
rect 672942 278700 672948 278702
rect 673012 278700 673018 278764
rect 673862 278564 673868 278628
rect 673932 278564 673938 278628
rect 48957 278082 49023 278085
rect 644657 278082 644723 278085
rect 48957 278080 644723 278082
rect 48957 278024 48962 278080
rect 49018 278024 644662 278080
rect 644718 278024 644723 278080
rect 48957 278022 644723 278024
rect 48957 278019 49023 278022
rect 644657 278019 644723 278022
rect 40902 277884 40908 277948
rect 40972 277946 40978 277948
rect 42241 277946 42307 277949
rect 40972 277944 42307 277946
rect 40972 277888 42246 277944
rect 42302 277888 42307 277944
rect 40972 277886 42307 277888
rect 40972 277884 40978 277886
rect 42241 277883 42307 277886
rect 673870 277676 673930 278564
rect 673862 277612 673868 277676
rect 673932 277612 673938 277676
rect 475745 277538 475811 277541
rect 476665 277538 476731 277541
rect 475745 277536 476731 277538
rect 475745 277480 475750 277536
rect 475806 277480 476670 277536
rect 476726 277480 476731 277536
rect 475745 277478 476731 277480
rect 475745 277475 475811 277478
rect 476665 277475 476731 277478
rect 40718 277340 40724 277404
rect 40788 277402 40794 277404
rect 41781 277402 41847 277405
rect 40788 277400 41847 277402
rect 40788 277344 41786 277400
rect 41842 277344 41847 277400
rect 40788 277342 41847 277344
rect 40788 277340 40794 277342
rect 41781 277339 41847 277342
rect 475561 277266 475627 277269
rect 476389 277266 476455 277269
rect 475561 277264 476455 277266
rect 475561 277208 475566 277264
rect 475622 277208 476394 277264
rect 476450 277208 476455 277264
rect 475561 277206 476455 277208
rect 475561 277203 475627 277206
rect 476389 277203 476455 277206
rect 499389 277266 499455 277269
rect 502517 277266 502583 277269
rect 499389 277264 502583 277266
rect 499389 277208 499394 277264
rect 499450 277208 502522 277264
rect 502578 277208 502583 277264
rect 499389 277206 502583 277208
rect 499389 277203 499455 277206
rect 502517 277203 502583 277206
rect 509417 277266 509483 277269
rect 512177 277266 512243 277269
rect 509417 277264 512243 277266
rect 509417 277208 509422 277264
rect 509478 277208 512182 277264
rect 512238 277208 512243 277264
rect 509417 277206 512243 277208
rect 509417 277203 509483 277206
rect 512177 277203 512243 277206
rect 42057 277130 42123 277133
rect 44173 277130 44239 277133
rect 42057 277128 44239 277130
rect 42057 277072 42062 277128
rect 42118 277072 44178 277128
rect 44234 277072 44239 277128
rect 42057 277070 44239 277072
rect 42057 277067 42123 277070
rect 44173 277067 44239 277070
rect 56041 276994 56107 276997
rect 653029 276994 653095 276997
rect 56041 276992 653095 276994
rect 56041 276936 56046 276992
rect 56102 276936 653034 276992
rect 653090 276936 653095 276992
rect 56041 276934 653095 276936
rect 56041 276931 56107 276934
rect 653029 276931 653095 276934
rect 53465 276722 53531 276725
rect 656893 276722 656959 276725
rect 53465 276720 656959 276722
rect 53465 276664 53470 276720
rect 53526 276664 656898 276720
rect 656954 276664 656959 276720
rect 53465 276662 656959 276664
rect 53465 276659 53531 276662
rect 656893 276659 656959 276662
rect 42057 276586 42123 276589
rect 45737 276586 45803 276589
rect 42057 276584 45803 276586
rect 42057 276528 42062 276584
rect 42118 276528 45742 276584
rect 45798 276528 45803 276584
rect 42057 276526 45803 276528
rect 42057 276523 42123 276526
rect 45737 276523 45803 276526
rect 475745 276450 475811 276453
rect 485865 276450 485931 276453
rect 475745 276448 485931 276450
rect 475745 276392 475750 276448
rect 475806 276392 485870 276448
rect 485926 276392 485931 276448
rect 475745 276390 485931 276392
rect 475745 276387 475811 276390
rect 485865 276387 485931 276390
rect 493133 276450 493199 276453
rect 508865 276450 508931 276453
rect 493133 276448 508931 276450
rect 493133 276392 493138 276448
rect 493194 276392 508870 276448
rect 508926 276392 508931 276448
rect 493133 276390 508931 276392
rect 493133 276387 493199 276390
rect 508865 276387 508931 276390
rect 509049 276450 509115 276453
rect 509233 276450 509299 276453
rect 509049 276448 509299 276450
rect 509049 276392 509054 276448
rect 509110 276392 509238 276448
rect 509294 276392 509299 276448
rect 509049 276390 509299 276392
rect 509049 276387 509115 276390
rect 509233 276387 509299 276390
rect 469949 276042 470015 276045
rect 473905 276042 473971 276045
rect 469949 276040 473971 276042
rect 469949 275984 469954 276040
rect 470010 275984 473910 276040
rect 473966 275984 473971 276040
rect 469949 275982 473971 275984
rect 469949 275979 470015 275982
rect 473905 275979 473971 275982
rect 486049 276042 486115 276045
rect 492213 276042 492279 276045
rect 486049 276040 492279 276042
rect 486049 275984 486054 276040
rect 486110 275984 492218 276040
rect 492274 275984 492279 276040
rect 486049 275982 492279 275984
rect 486049 275979 486115 275982
rect 492213 275979 492279 275982
rect 480989 275906 481055 275909
rect 480210 275904 481055 275906
rect 480210 275848 480994 275904
rect 481050 275848 481055 275904
rect 480210 275846 481055 275848
rect 470501 275770 470567 275773
rect 471421 275770 471487 275773
rect 470501 275768 471487 275770
rect 470501 275712 470506 275768
rect 470562 275712 471426 275768
rect 471482 275712 471487 275768
rect 470501 275710 471487 275712
rect 470501 275707 470567 275710
rect 471421 275707 471487 275710
rect 473905 275770 473971 275773
rect 480210 275770 480270 275846
rect 480989 275843 481055 275846
rect 484117 275906 484183 275909
rect 485865 275906 485931 275909
rect 484117 275904 485931 275906
rect 484117 275848 484122 275904
rect 484178 275848 485870 275904
rect 485926 275848 485931 275904
rect 484117 275846 485931 275848
rect 484117 275843 484183 275846
rect 485865 275843 485931 275846
rect 492581 275906 492647 275909
rect 499389 275906 499455 275909
rect 492581 275904 499455 275906
rect 492581 275848 492586 275904
rect 492642 275848 499394 275904
rect 499450 275848 499455 275904
rect 492581 275846 499455 275848
rect 492581 275843 492647 275846
rect 499389 275843 499455 275846
rect 473905 275768 480270 275770
rect 473905 275712 473910 275768
rect 473966 275712 480270 275768
rect 473905 275710 480270 275712
rect 487337 275770 487403 275773
rect 490741 275770 490807 275773
rect 487337 275768 490807 275770
rect 487337 275712 487342 275768
rect 487398 275712 490746 275768
rect 490802 275712 490807 275768
rect 487337 275710 490807 275712
rect 473905 275707 473971 275710
rect 487337 275707 487403 275710
rect 490741 275707 490807 275710
rect 445477 275498 445543 275501
rect 541065 275498 541131 275501
rect 445477 275496 541131 275498
rect 445477 275440 445482 275496
rect 445538 275440 541070 275496
rect 541126 275440 541131 275496
rect 445477 275438 541131 275440
rect 445477 275435 445543 275438
rect 541065 275435 541131 275438
rect 461577 275226 461643 275229
rect 466545 275226 466611 275229
rect 461577 275224 466611 275226
rect 461577 275168 461582 275224
rect 461638 275168 466550 275224
rect 466606 275168 466611 275224
rect 461577 275166 466611 275168
rect 461577 275163 461643 275166
rect 466545 275163 466611 275166
rect 481265 275226 481331 275229
rect 619081 275226 619147 275229
rect 481265 275224 619147 275226
rect 481265 275168 481270 275224
rect 481326 275168 619086 275224
rect 619142 275168 619147 275224
rect 481265 275166 619147 275168
rect 481265 275163 481331 275166
rect 619081 275163 619147 275166
rect 466453 274954 466519 274957
rect 469765 274954 469831 274957
rect 466453 274952 469831 274954
rect 466453 274896 466458 274952
rect 466514 274896 469770 274952
rect 469826 274896 469831 274952
rect 466453 274894 469831 274896
rect 466453 274891 466519 274894
rect 469765 274891 469831 274894
rect 484301 274954 484367 274957
rect 486693 274954 486759 274957
rect 484301 274952 486759 274954
rect 484301 274896 484306 274952
rect 484362 274896 486698 274952
rect 486754 274896 486759 274952
rect 484301 274894 486759 274896
rect 484301 274891 484367 274894
rect 486693 274891 486759 274894
rect 494145 274954 494211 274957
rect 498929 274954 498995 274957
rect 494145 274952 498995 274954
rect 494145 274896 494150 274952
rect 494206 274896 498934 274952
rect 498990 274896 498995 274952
rect 494145 274894 498995 274896
rect 494145 274891 494211 274894
rect 498929 274891 498995 274894
rect 499389 274954 499455 274957
rect 499665 274954 499731 274957
rect 499389 274952 499731 274954
rect 499389 274896 499394 274952
rect 499450 274896 499670 274952
rect 499726 274896 499731 274952
rect 499389 274894 499731 274896
rect 499389 274891 499455 274894
rect 499665 274891 499731 274894
rect 486693 274682 486759 274685
rect 494973 274682 495039 274685
rect 486693 274680 495039 274682
rect 486693 274624 486698 274680
rect 486754 274624 494978 274680
rect 495034 274624 495039 274680
rect 486693 274622 495039 274624
rect 486693 274619 486759 274622
rect 494973 274619 495039 274622
rect 495249 274682 495315 274685
rect 497181 274682 497247 274685
rect 495249 274680 497247 274682
rect 495249 274624 495254 274680
rect 495310 274624 497186 274680
rect 497242 274624 497247 274680
rect 495249 274622 497247 274624
rect 495249 274619 495315 274622
rect 497181 274619 497247 274622
rect 466407 274546 466473 274549
rect 472157 274546 472223 274549
rect 466407 274544 472223 274546
rect 466407 274488 466412 274544
rect 466468 274488 472162 274544
rect 472218 274488 472223 274544
rect 466407 274486 472223 274488
rect 466407 274483 466473 274486
rect 472157 274483 472223 274486
rect 475377 274546 475443 274549
rect 480345 274546 480411 274549
rect 475377 274544 480411 274546
rect 475377 274488 475382 274544
rect 475438 274488 480350 274544
rect 480406 274488 480411 274544
rect 475377 274486 480411 274488
rect 475377 274483 475443 274486
rect 480345 274483 480411 274486
rect 481449 274410 481515 274413
rect 486417 274410 486483 274413
rect 481449 274408 486483 274410
rect 481449 274352 481454 274408
rect 481510 274352 486422 274408
rect 486478 274352 486483 274408
rect 481449 274350 486483 274352
rect 481449 274347 481515 274350
rect 486417 274347 486483 274350
rect 486877 274410 486943 274413
rect 495249 274410 495315 274413
rect 486877 274408 495315 274410
rect 486877 274352 486882 274408
rect 486938 274352 495254 274408
rect 495310 274352 495315 274408
rect 486877 274350 495315 274352
rect 486877 274347 486943 274350
rect 495249 274347 495315 274350
rect 454585 274138 454651 274141
rect 569493 274138 569559 274141
rect 454585 274136 569559 274138
rect 454585 274080 454590 274136
rect 454646 274080 569498 274136
rect 569554 274080 569559 274136
rect 454585 274078 569559 274080
rect 454585 274075 454651 274078
rect 569493 274075 569559 274078
rect 434437 274002 434503 274005
rect 435357 274002 435423 274005
rect 434437 274000 435423 274002
rect 434437 273944 434442 274000
rect 434498 273944 435362 274000
rect 435418 273944 435423 274000
rect 434437 273942 435423 273944
rect 434437 273939 434503 273942
rect 435357 273939 435423 273942
rect 448145 274002 448211 274005
rect 451365 274002 451431 274005
rect 448145 274000 451431 274002
rect 448145 273944 448150 274000
rect 448206 273944 451370 274000
rect 451426 273944 451431 274000
rect 448145 273942 451431 273944
rect 448145 273939 448211 273942
rect 451365 273939 451431 273942
rect 487061 273866 487127 273869
rect 488717 273866 488783 273869
rect 487061 273864 488783 273866
rect 487061 273808 487066 273864
rect 487122 273808 488722 273864
rect 488778 273808 488783 273864
rect 487061 273806 488783 273808
rect 487061 273803 487127 273806
rect 488717 273803 488783 273806
rect 489361 273866 489427 273869
rect 632145 273866 632211 273869
rect 489361 273864 632211 273866
rect 489361 273808 489366 273864
rect 489422 273808 632150 273864
rect 632206 273808 632211 273864
rect 489361 273806 632211 273808
rect 489361 273803 489427 273806
rect 632145 273803 632211 273806
rect 460749 273730 460815 273733
rect 466545 273730 466611 273733
rect 460749 273728 466611 273730
rect 460749 273672 460754 273728
rect 460810 273672 466550 273728
rect 466606 273672 466611 273728
rect 460749 273670 466611 273672
rect 460749 273667 460815 273670
rect 466545 273667 466611 273670
rect 497457 273594 497523 273597
rect 505277 273594 505343 273597
rect 497457 273592 505343 273594
rect 497457 273536 497462 273592
rect 497518 273536 505282 273592
rect 505338 273536 505343 273592
rect 497457 273534 505343 273536
rect 497457 273531 497523 273534
rect 505277 273531 505343 273534
rect 40534 273396 40540 273460
rect 40604 273458 40610 273460
rect 41781 273458 41847 273461
rect 40604 273456 41847 273458
rect 40604 273400 41786 273456
rect 41842 273400 41847 273456
rect 40604 273398 41847 273400
rect 40604 273396 40610 273398
rect 41781 273395 41847 273398
rect 494881 273322 494947 273325
rect 500861 273322 500927 273325
rect 494881 273320 500927 273322
rect 494881 273264 494886 273320
rect 494942 273264 500866 273320
rect 500922 273264 500927 273320
rect 494881 273262 500927 273264
rect 494881 273259 494947 273262
rect 500861 273259 500927 273262
rect 449709 273186 449775 273189
rect 460933 273186 460999 273189
rect 449709 273184 460999 273186
rect 449709 273128 449714 273184
rect 449770 273128 460938 273184
rect 460994 273128 460999 273184
rect 449709 273126 460999 273128
rect 449709 273123 449775 273126
rect 460933 273123 460999 273126
rect 436921 273050 436987 273053
rect 438209 273050 438275 273053
rect 436921 273048 438275 273050
rect 436921 272992 436926 273048
rect 436982 272992 438214 273048
rect 438270 272992 438275 273048
rect 436921 272990 438275 272992
rect 436921 272987 436987 272990
rect 438209 272987 438275 272990
rect 445385 273050 445451 273053
rect 447225 273050 447291 273053
rect 445385 273048 447291 273050
rect 445385 272992 445390 273048
rect 445446 272992 447230 273048
rect 447286 272992 447291 273048
rect 445385 272990 447291 272992
rect 445385 272987 445451 272990
rect 447225 272987 447291 272990
rect 495893 273050 495959 273053
rect 507853 273050 507919 273053
rect 495893 273048 507919 273050
rect 495893 272992 495898 273048
rect 495954 272992 507858 273048
rect 507914 272992 507919 273048
rect 495893 272990 507919 272992
rect 495893 272987 495959 272990
rect 507853 272987 507919 272990
rect 433149 272778 433215 272781
rect 437289 272778 437355 272781
rect 433149 272776 437355 272778
rect 433149 272720 433154 272776
rect 433210 272720 437294 272776
rect 437350 272720 437355 272776
rect 433149 272718 437355 272720
rect 433149 272715 433215 272718
rect 437289 272715 437355 272718
rect 456609 272778 456675 272781
rect 457437 272778 457503 272781
rect 476757 272778 476823 272781
rect 456609 272776 457503 272778
rect 456609 272720 456614 272776
rect 456670 272720 457442 272776
rect 457498 272720 457503 272776
rect 456609 272718 457503 272720
rect 456609 272715 456675 272718
rect 457437 272715 457503 272718
rect 466686 272776 476823 272778
rect 466686 272720 476762 272776
rect 476818 272720 476823 272776
rect 466686 272718 476823 272720
rect 466269 272506 466335 272509
rect 466686 272506 466746 272718
rect 476757 272715 476823 272718
rect 491017 272778 491083 272781
rect 511349 272778 511415 272781
rect 491017 272776 511415 272778
rect 491017 272720 491022 272776
rect 491078 272720 511354 272776
rect 511410 272720 511415 272776
rect 491017 272718 511415 272720
rect 491017 272715 491083 272718
rect 511349 272715 511415 272718
rect 593137 272506 593203 272509
rect 466269 272504 466746 272506
rect 466269 272448 466274 272504
rect 466330 272448 466746 272504
rect 466269 272446 466746 272448
rect 476070 272504 593203 272506
rect 476070 272448 593142 272504
rect 593198 272448 593203 272504
rect 476070 272446 593203 272448
rect 466269 272443 466335 272446
rect 41781 272372 41847 272373
rect 41781 272368 41828 272372
rect 41892 272370 41898 272372
rect 427813 272370 427879 272373
rect 430941 272370 431007 272373
rect 41781 272312 41786 272368
rect 41781 272308 41828 272312
rect 41892 272310 41938 272370
rect 427813 272368 431007 272370
rect 427813 272312 427818 272368
rect 427874 272312 430946 272368
rect 431002 272312 431007 272368
rect 427813 272310 431007 272312
rect 41892 272308 41898 272310
rect 41781 272307 41847 272308
rect 427813 272307 427879 272310
rect 430941 272307 431007 272310
rect 446765 272370 446831 272373
rect 447409 272370 447475 272373
rect 446765 272368 447475 272370
rect 446765 272312 446770 272368
rect 446826 272312 447414 272368
rect 447470 272312 447475 272368
rect 446765 272310 447475 272312
rect 446765 272307 446831 272310
rect 447409 272307 447475 272310
rect 447593 272370 447659 272373
rect 454401 272370 454467 272373
rect 447593 272368 454467 272370
rect 447593 272312 447598 272368
rect 447654 272312 454406 272368
rect 454462 272312 454467 272368
rect 447593 272310 454467 272312
rect 447593 272307 447659 272310
rect 454401 272307 454467 272310
rect 464889 272234 464955 272237
rect 476070 272234 476130 272446
rect 593137 272443 593203 272446
rect 464889 272232 476130 272234
rect 464889 272176 464894 272232
rect 464950 272176 476130 272232
rect 464889 272174 476130 272176
rect 476757 272234 476823 272237
rect 485865 272234 485931 272237
rect 476757 272232 485931 272234
rect 476757 272176 476762 272232
rect 476818 272176 485870 272232
rect 485926 272176 485931 272232
rect 476757 272174 485931 272176
rect 464889 272171 464955 272174
rect 476757 272171 476823 272174
rect 485865 272171 485931 272174
rect 486049 272234 486115 272237
rect 495893 272234 495959 272237
rect 486049 272232 495959 272234
rect 486049 272176 486054 272232
rect 486110 272176 495898 272232
rect 495954 272176 495959 272232
rect 486049 272174 495959 272176
rect 486049 272171 486115 272174
rect 495893 272171 495959 272174
rect 441521 272098 441587 272101
rect 443361 272098 443427 272101
rect 441521 272096 443427 272098
rect 441521 272040 441526 272096
rect 441582 272040 443366 272096
rect 443422 272040 443427 272096
rect 441521 272038 443427 272040
rect 441521 272035 441587 272038
rect 443361 272035 443427 272038
rect 427077 271962 427143 271965
rect 427905 271962 427971 271965
rect 427077 271960 427971 271962
rect 427077 271904 427082 271960
rect 427138 271904 427910 271960
rect 427966 271904 427971 271960
rect 427077 271902 427971 271904
rect 427077 271899 427143 271902
rect 427905 271899 427971 271902
rect 458633 271962 458699 271965
rect 466269 271962 466335 271965
rect 458633 271960 466335 271962
rect 458633 271904 458638 271960
rect 458694 271904 466274 271960
rect 466330 271904 466335 271960
rect 458633 271902 466335 271904
rect 458633 271899 458699 271902
rect 466269 271899 466335 271902
rect 485773 271962 485839 271965
rect 492949 271962 493015 271965
rect 485773 271960 493015 271962
rect 485773 271904 485778 271960
rect 485834 271904 492954 271960
rect 493010 271904 493015 271960
rect 485773 271902 493015 271904
rect 485773 271899 485839 271902
rect 492949 271899 493015 271902
rect 428181 271690 428247 271693
rect 429377 271690 429443 271693
rect 428181 271688 429443 271690
rect 428181 271632 428186 271688
rect 428242 271632 429382 271688
rect 429438 271632 429443 271688
rect 428181 271630 429443 271632
rect 428181 271627 428247 271630
rect 429377 271627 429443 271630
rect 431769 271690 431835 271693
rect 539869 271690 539935 271693
rect 431769 271688 539935 271690
rect 431769 271632 431774 271688
rect 431830 271632 539874 271688
rect 539930 271632 539935 271688
rect 431769 271630 539935 271632
rect 431769 271627 431835 271630
rect 539869 271627 539935 271630
rect 429101 271418 429167 271421
rect 433517 271418 433583 271421
rect 429101 271416 433583 271418
rect 429101 271360 429106 271416
rect 429162 271360 433522 271416
rect 433578 271360 433583 271416
rect 429101 271358 433583 271360
rect 429101 271355 429167 271358
rect 433517 271355 433583 271358
rect 441153 271418 441219 271421
rect 442717 271418 442783 271421
rect 441153 271416 442783 271418
rect 441153 271360 441158 271416
rect 441214 271360 442722 271416
rect 442778 271360 442783 271416
rect 441153 271358 442783 271360
rect 441153 271355 441219 271358
rect 442717 271355 442783 271358
rect 462773 271418 462839 271421
rect 466545 271418 466611 271421
rect 462773 271416 466611 271418
rect 462773 271360 462778 271416
rect 462834 271360 466550 271416
rect 466606 271360 466611 271416
rect 462773 271358 466611 271360
rect 462773 271355 462839 271358
rect 466545 271355 466611 271358
rect 466729 271418 466795 271421
rect 485865 271418 485931 271421
rect 626165 271418 626231 271421
rect 466729 271416 485931 271418
rect 466729 271360 466734 271416
rect 466790 271360 485870 271416
rect 485926 271360 485931 271416
rect 466729 271358 485931 271360
rect 466729 271355 466795 271358
rect 485865 271355 485931 271358
rect 495390 271416 626231 271418
rect 495390 271360 626170 271416
rect 626226 271360 626231 271416
rect 495390 271358 626231 271360
rect 456609 271282 456675 271285
rect 461853 271282 461919 271285
rect 456609 271280 461919 271282
rect 456609 271224 456614 271280
rect 456670 271224 461858 271280
rect 461914 271224 461919 271280
rect 456609 271222 461919 271224
rect 456609 271219 456675 271222
rect 461853 271219 461919 271222
rect 412633 271146 412699 271149
rect 418981 271146 419047 271149
rect 412633 271144 419047 271146
rect 412633 271088 412638 271144
rect 412694 271088 418986 271144
rect 419042 271088 419047 271144
rect 412633 271086 419047 271088
rect 412633 271083 412699 271086
rect 418981 271083 419047 271086
rect 439497 271146 439563 271149
rect 444741 271146 444807 271149
rect 439497 271144 444807 271146
rect 439497 271088 439502 271144
rect 439558 271088 444746 271144
rect 444802 271088 444807 271144
rect 439497 271086 444807 271088
rect 439497 271083 439563 271086
rect 444741 271083 444807 271086
rect 446121 271146 446187 271149
rect 495390 271146 495450 271358
rect 626165 271355 626231 271358
rect 446121 271144 447150 271146
rect 446121 271088 446126 271144
rect 446182 271088 447150 271144
rect 446121 271086 447150 271088
rect 446121 271083 446187 271086
rect 431401 271010 431467 271013
rect 432965 271010 433031 271013
rect 431401 271008 433031 271010
rect 431401 270952 431406 271008
rect 431462 270952 432970 271008
rect 433026 270952 433031 271008
rect 431401 270950 433031 270952
rect 447090 271010 447150 271086
rect 485730 271086 495450 271146
rect 495801 271146 495867 271149
rect 496353 271146 496419 271149
rect 495801 271144 496419 271146
rect 495801 271088 495806 271144
rect 495862 271088 496358 271144
rect 496414 271088 496419 271144
rect 495801 271086 496419 271088
rect 457437 271010 457503 271013
rect 447090 271008 457503 271010
rect 447090 270952 457442 271008
rect 457498 270952 457503 271008
rect 447090 270950 457503 270952
rect 431401 270947 431467 270950
rect 432965 270947 433031 270950
rect 457437 270947 457503 270950
rect 485497 271010 485563 271013
rect 485730 271010 485790 271086
rect 495801 271083 495867 271086
rect 496353 271083 496419 271086
rect 496721 271146 496787 271149
rect 642725 271146 642791 271149
rect 496721 271144 642791 271146
rect 496721 271088 496726 271144
rect 496782 271088 642730 271144
rect 642786 271088 642791 271144
rect 496721 271086 642791 271088
rect 496721 271083 496787 271086
rect 642725 271083 642791 271086
rect 485497 271008 485790 271010
rect 485497 270952 485502 271008
rect 485558 270952 485790 271008
rect 485497 270950 485790 270952
rect 485497 270947 485563 270950
rect 493961 270874 494027 270877
rect 496537 270874 496603 270877
rect 493961 270872 496603 270874
rect 493961 270816 493966 270872
rect 494022 270816 496542 270872
rect 496598 270816 496603 270872
rect 493961 270814 496603 270816
rect 493961 270811 494027 270814
rect 496537 270811 496603 270814
rect 412081 270738 412147 270741
rect 412725 270738 412791 270741
rect 412081 270736 412791 270738
rect 412081 270680 412086 270736
rect 412142 270680 412730 270736
rect 412786 270680 412791 270736
rect 412081 270678 412791 270680
rect 412081 270675 412147 270678
rect 412725 270675 412791 270678
rect 418889 270738 418955 270741
rect 423305 270738 423371 270741
rect 418889 270736 423371 270738
rect 418889 270680 418894 270736
rect 418950 270680 423310 270736
rect 423366 270680 423371 270736
rect 418889 270678 423371 270680
rect 418889 270675 418955 270678
rect 423305 270675 423371 270678
rect 472249 270738 472315 270741
rect 486877 270738 486943 270741
rect 472249 270736 486943 270738
rect 472249 270680 472254 270736
rect 472310 270680 486882 270736
rect 486938 270680 486943 270736
rect 472249 270678 486943 270680
rect 472249 270675 472315 270678
rect 486877 270675 486943 270678
rect 403985 270602 404051 270605
rect 408493 270602 408559 270605
rect 403985 270600 408559 270602
rect 403985 270544 403990 270600
rect 404046 270544 408498 270600
rect 408554 270544 408559 270600
rect 403985 270542 408559 270544
rect 403985 270539 404051 270542
rect 408493 270539 408559 270542
rect 417233 270602 417299 270605
rect 418245 270602 418311 270605
rect 417233 270600 418311 270602
rect 417233 270544 417238 270600
rect 417294 270544 418250 270600
rect 418306 270544 418311 270600
rect 417233 270542 418311 270544
rect 417233 270539 417299 270542
rect 418245 270539 418311 270542
rect 456609 270602 456675 270605
rect 459921 270602 459987 270605
rect 456609 270600 459987 270602
rect 456609 270544 456614 270600
rect 456670 270544 459926 270600
rect 459982 270544 459987 270600
rect 456609 270542 459987 270544
rect 456609 270539 456675 270542
rect 459921 270539 459987 270542
rect 495433 270602 495499 270605
rect 504173 270602 504239 270605
rect 495433 270600 504239 270602
rect 495433 270544 495438 270600
rect 495494 270544 504178 270600
rect 504234 270544 504239 270600
rect 495433 270542 504239 270544
rect 495433 270539 495499 270542
rect 504173 270539 504239 270542
rect 41454 270404 41460 270468
rect 41524 270466 41530 270468
rect 41781 270466 41847 270469
rect 41524 270464 41847 270466
rect 41524 270408 41786 270464
rect 41842 270408 41847 270464
rect 41524 270406 41847 270408
rect 41524 270404 41530 270406
rect 41781 270403 41847 270406
rect 409505 270466 409571 270469
rect 412449 270466 412515 270469
rect 409505 270464 412515 270466
rect 409505 270408 409510 270464
rect 409566 270408 412454 270464
rect 412510 270408 412515 270464
rect 409505 270406 412515 270408
rect 409505 270403 409571 270406
rect 412449 270403 412515 270406
rect 384941 270330 385007 270333
rect 386597 270330 386663 270333
rect 384941 270328 386663 270330
rect 384941 270272 384946 270328
rect 385002 270272 386602 270328
rect 386658 270272 386663 270328
rect 384941 270270 386663 270272
rect 384941 270267 385007 270270
rect 386597 270267 386663 270270
rect 459001 270330 459067 270333
rect 582741 270330 582807 270333
rect 459001 270328 582807 270330
rect 459001 270272 459006 270328
rect 459062 270272 582746 270328
rect 582802 270272 582807 270328
rect 459001 270270 582807 270272
rect 459001 270267 459067 270270
rect 582741 270267 582807 270270
rect 448697 270194 448763 270197
rect 456609 270194 456675 270197
rect 448697 270192 456675 270194
rect 448697 270136 448702 270192
rect 448758 270136 456614 270192
rect 456670 270136 456675 270192
rect 448697 270134 456675 270136
rect 448697 270131 448763 270134
rect 456609 270131 456675 270134
rect 412449 270058 412515 270061
rect 412725 270058 412791 270061
rect 412449 270056 412791 270058
rect 412449 270000 412454 270056
rect 412510 270000 412730 270056
rect 412786 270000 412791 270056
rect 412449 269998 412791 270000
rect 412449 269995 412515 269998
rect 412725 269995 412791 269998
rect 427813 270058 427879 270061
rect 434805 270058 434871 270061
rect 427813 270056 434871 270058
rect 427813 270000 427818 270056
rect 427874 270000 434810 270056
rect 434866 270000 434871 270056
rect 427813 269998 434871 270000
rect 427813 269995 427879 269998
rect 434805 269995 434871 269998
rect 475745 270058 475811 270061
rect 477861 270058 477927 270061
rect 475745 270056 477927 270058
rect 475745 270000 475750 270056
rect 475806 270000 477866 270056
rect 477922 270000 477927 270056
rect 475745 269998 477927 270000
rect 475745 269995 475811 269998
rect 477861 269995 477927 269998
rect 479977 270058 480043 270061
rect 484853 270058 484919 270061
rect 479977 270056 484919 270058
rect 479977 270000 479982 270056
rect 480038 270000 484858 270056
rect 484914 270000 484919 270056
rect 479977 269998 484919 270000
rect 479977 269995 480043 269998
rect 484853 269995 484919 269998
rect 488349 270058 488415 270061
rect 630673 270058 630739 270061
rect 488349 270056 630739 270058
rect 488349 270000 488354 270056
rect 488410 270000 630678 270056
rect 630734 270000 630739 270056
rect 488349 269998 630739 270000
rect 488349 269995 488415 269998
rect 630673 269995 630739 269998
rect 400121 269786 400187 269789
rect 488533 269786 488599 269789
rect 400121 269784 488599 269786
rect 400121 269728 400126 269784
rect 400182 269728 488538 269784
rect 488594 269728 488599 269784
rect 400121 269726 488599 269728
rect 400121 269723 400187 269726
rect 488533 269723 488599 269726
rect 494697 269786 494763 269789
rect 640609 269786 640675 269789
rect 494697 269784 640675 269786
rect 494697 269728 494702 269784
rect 494758 269728 640614 269784
rect 640670 269728 640675 269784
rect 494697 269726 640675 269728
rect 494697 269723 494763 269726
rect 640609 269723 640675 269726
rect 382181 269650 382247 269653
rect 384481 269650 384547 269653
rect 382181 269648 384547 269650
rect 382181 269592 382186 269648
rect 382242 269592 384486 269648
rect 384542 269592 384547 269648
rect 382181 269590 384547 269592
rect 382181 269587 382247 269590
rect 384481 269587 384547 269590
rect 420729 269514 420795 269517
rect 427445 269514 427511 269517
rect 420729 269512 427511 269514
rect 420729 269456 420734 269512
rect 420790 269456 427450 269512
rect 427506 269456 427511 269512
rect 420729 269454 427511 269456
rect 420729 269451 420795 269454
rect 427445 269451 427511 269454
rect 429561 269514 429627 269517
rect 535453 269514 535519 269517
rect 429561 269512 535519 269514
rect 429561 269456 429566 269512
rect 429622 269456 535458 269512
rect 535514 269456 535519 269512
rect 429561 269454 535519 269456
rect 429561 269451 429627 269454
rect 535453 269451 535519 269454
rect 393405 269242 393471 269245
rect 402421 269242 402487 269245
rect 393405 269240 402487 269242
rect 393405 269184 393410 269240
rect 393466 269184 402426 269240
rect 402482 269184 402487 269240
rect 393405 269182 402487 269184
rect 393405 269179 393471 269182
rect 402421 269179 402487 269182
rect 427629 269242 427695 269245
rect 427997 269242 428063 269245
rect 427629 269240 428063 269242
rect 427629 269184 427634 269240
rect 427690 269184 428002 269240
rect 428058 269184 428063 269240
rect 427629 269182 428063 269184
rect 427629 269179 427695 269182
rect 427997 269179 428063 269182
rect 466269 269242 466335 269245
rect 466453 269242 466519 269245
rect 466269 269240 466519 269242
rect 466269 269184 466274 269240
rect 466330 269184 466458 269240
rect 466514 269184 466519 269240
rect 466269 269182 466519 269184
rect 466269 269179 466335 269182
rect 466453 269179 466519 269182
rect 469673 269242 469739 269245
rect 476481 269242 476547 269245
rect 469673 269240 476547 269242
rect 469673 269184 469678 269240
rect 469734 269184 476486 269240
rect 476542 269184 476547 269240
rect 469673 269182 476547 269184
rect 469673 269179 469739 269182
rect 476481 269179 476547 269182
rect 476665 269242 476731 269245
rect 484117 269242 484183 269245
rect 476665 269240 484183 269242
rect 476665 269184 476670 269240
rect 476726 269184 484122 269240
rect 484178 269184 484183 269240
rect 476665 269182 484183 269184
rect 476665 269179 476731 269182
rect 484117 269179 484183 269182
rect 486601 269242 486667 269245
rect 491569 269242 491635 269245
rect 486601 269240 491635 269242
rect 486601 269184 486606 269240
rect 486662 269184 491574 269240
rect 491630 269184 491635 269240
rect 486601 269182 491635 269184
rect 486601 269179 486667 269182
rect 491569 269179 491635 269182
rect 493225 269242 493291 269245
rect 495525 269242 495591 269245
rect 493225 269240 495591 269242
rect 493225 269184 493230 269240
rect 493286 269184 495530 269240
rect 495586 269184 495591 269240
rect 493225 269182 495591 269184
rect 493225 269179 493291 269182
rect 495525 269179 495591 269182
rect 456425 268970 456491 268973
rect 462313 268970 462379 268973
rect 456425 268968 462379 268970
rect 456425 268912 456430 268968
rect 456486 268912 462318 268968
rect 462374 268912 462379 268968
rect 456425 268910 462379 268912
rect 456425 268907 456491 268910
rect 462313 268907 462379 268910
rect 484669 268970 484735 268973
rect 486417 268970 486483 268973
rect 484669 268968 486483 268970
rect 484669 268912 484674 268968
rect 484730 268912 486422 268968
rect 486478 268912 486483 268968
rect 484669 268910 486483 268912
rect 484669 268907 484735 268910
rect 486417 268907 486483 268910
rect 437289 268698 437355 268701
rect 438853 268698 438919 268701
rect 437289 268696 438919 268698
rect 437289 268640 437294 268696
rect 437350 268640 438858 268696
rect 438914 268640 438919 268696
rect 437289 268638 438919 268640
rect 437289 268635 437355 268638
rect 438853 268635 438919 268638
rect 446765 268698 446831 268701
rect 448513 268698 448579 268701
rect 446765 268696 448579 268698
rect 446765 268640 446770 268696
rect 446826 268640 448518 268696
rect 448574 268640 448579 268696
rect 446765 268638 448579 268640
rect 446765 268635 446831 268638
rect 448513 268635 448579 268638
rect 461025 268698 461091 268701
rect 462497 268698 462563 268701
rect 461025 268696 462563 268698
rect 461025 268640 461030 268696
rect 461086 268640 462502 268696
rect 462558 268640 462563 268696
rect 461025 268638 462563 268640
rect 461025 268635 461091 268638
rect 462497 268635 462563 268638
rect 466729 268698 466795 268701
rect 471421 268698 471487 268701
rect 466729 268696 471487 268698
rect 466729 268640 466734 268696
rect 466790 268640 471426 268696
rect 471482 268640 471487 268696
rect 466729 268638 471487 268640
rect 466729 268635 466795 268638
rect 471421 268635 471487 268638
rect 484853 268698 484919 268701
rect 486233 268698 486299 268701
rect 484853 268696 486299 268698
rect 484853 268640 484858 268696
rect 484914 268640 486238 268696
rect 486294 268640 486299 268696
rect 484853 268638 486299 268640
rect 484853 268635 484919 268638
rect 486233 268635 486299 268638
rect 490189 268698 490255 268701
rect 493041 268698 493107 268701
rect 490189 268696 493107 268698
rect 490189 268640 490194 268696
rect 490250 268640 493046 268696
rect 493102 268640 493107 268696
rect 490189 268638 493107 268640
rect 490189 268635 490255 268638
rect 493041 268635 493107 268638
rect 495065 268698 495131 268701
rect 495525 268698 495591 268701
rect 495065 268696 495591 268698
rect 495065 268640 495070 268696
rect 495126 268640 495530 268696
rect 495586 268640 495591 268696
rect 495065 268638 495591 268640
rect 495065 268635 495131 268638
rect 495525 268635 495591 268638
rect 504909 268698 504975 268701
rect 506473 268698 506539 268701
rect 504909 268696 506539 268698
rect 504909 268640 504914 268696
rect 504970 268640 506478 268696
rect 506534 268640 506539 268696
rect 504909 268638 506539 268640
rect 504909 268635 504975 268638
rect 506473 268635 506539 268638
rect 675477 268698 675543 268701
rect 675477 268696 676292 268698
rect 675477 268640 675482 268696
rect 675538 268640 676292 268696
rect 675477 268638 676292 268640
rect 675477 268635 675543 268638
rect 436921 268426 436987 268429
rect 547873 268426 547939 268429
rect 436921 268424 547939 268426
rect 436921 268368 436926 268424
rect 436982 268368 547878 268424
rect 547934 268368 547939 268424
rect 436921 268366 547939 268368
rect 436921 268363 436987 268366
rect 547873 268363 547939 268366
rect 675477 268290 675543 268293
rect 675477 268288 676292 268290
rect 675477 268232 675482 268288
rect 675538 268232 676292 268288
rect 675477 268230 676292 268232
rect 675477 268227 675543 268230
rect 417049 268154 417115 268157
rect 418061 268154 418127 268157
rect 417049 268152 418127 268154
rect 417049 268096 417054 268152
rect 417110 268096 418066 268152
rect 418122 268096 418127 268152
rect 417049 268094 418127 268096
rect 417049 268091 417115 268094
rect 418061 268091 418127 268094
rect 427629 268154 427695 268157
rect 427813 268154 427879 268157
rect 427629 268152 427879 268154
rect 427629 268096 427634 268152
rect 427690 268096 427818 268152
rect 427874 268096 427879 268152
rect 427629 268094 427879 268096
rect 427629 268091 427695 268094
rect 427813 268091 427879 268094
rect 474089 268154 474155 268157
rect 476205 268154 476271 268157
rect 474089 268152 476271 268154
rect 474089 268096 474094 268152
rect 474150 268096 476210 268152
rect 476266 268096 476271 268152
rect 474089 268094 476271 268096
rect 474089 268091 474155 268094
rect 476205 268091 476271 268094
rect 485037 268154 485103 268157
rect 494513 268154 494579 268157
rect 504909 268154 504975 268157
rect 485037 268152 486066 268154
rect 485037 268096 485042 268152
rect 485098 268096 486066 268152
rect 485037 268094 486066 268096
rect 485037 268091 485103 268094
rect 486006 268021 486066 268094
rect 494513 268152 504975 268154
rect 494513 268096 494518 268152
rect 494574 268096 504914 268152
rect 504970 268096 504975 268152
rect 494513 268094 504975 268096
rect 494513 268091 494579 268094
rect 504909 268091 504975 268094
rect 436553 268018 436619 268021
rect 442993 268018 443059 268021
rect 436553 268016 443059 268018
rect 436553 267960 436558 268016
rect 436614 267960 442998 268016
rect 443054 267960 443059 268016
rect 436553 267958 443059 267960
rect 436553 267955 436619 267958
rect 442993 267955 443059 267958
rect 456609 268018 456675 268021
rect 461577 268018 461643 268021
rect 456609 268016 461643 268018
rect 456609 267960 456614 268016
rect 456670 267960 461582 268016
rect 461638 267960 461643 268016
rect 456609 267958 461643 267960
rect 486006 268016 486115 268021
rect 486006 267960 486054 268016
rect 486110 267960 486115 268016
rect 486006 267958 486115 267960
rect 456609 267955 456675 267958
rect 461577 267955 461643 267958
rect 486049 267955 486115 267958
rect 491569 268018 491635 268021
rect 491569 268016 493058 268018
rect 491569 267960 491574 268016
rect 491630 267960 493058 268016
rect 491569 267958 493058 267960
rect 491569 267955 491635 267958
rect 415485 267882 415551 267885
rect 417785 267882 417851 267885
rect 415485 267880 417851 267882
rect 415485 267824 415490 267880
rect 415546 267824 417790 267880
rect 417846 267824 417851 267880
rect 415485 267822 417851 267824
rect 415485 267819 415551 267822
rect 417785 267819 417851 267822
rect 475745 267882 475811 267885
rect 485681 267882 485747 267885
rect 475745 267880 485747 267882
rect 475745 267824 475750 267880
rect 475806 267824 485686 267880
rect 485742 267824 485747 267880
rect 475745 267822 485747 267824
rect 492998 267882 493058 267958
rect 502149 267882 502215 267885
rect 492998 267880 502215 267882
rect 492998 267824 502154 267880
rect 502210 267824 502215 267880
rect 492998 267822 502215 267824
rect 475745 267819 475811 267822
rect 485681 267819 485747 267822
rect 502149 267819 502215 267822
rect 675477 267882 675543 267885
rect 675477 267880 676292 267882
rect 675477 267824 675482 267880
rect 675538 267824 676292 267880
rect 675477 267822 676292 267824
rect 675477 267819 675543 267822
rect 364149 267746 364215 267749
rect 366357 267746 366423 267749
rect 418337 267746 418403 267749
rect 364149 267744 366423 267746
rect 364149 267688 364154 267744
rect 364210 267688 366362 267744
rect 366418 267688 366423 267744
rect 364149 267686 366423 267688
rect 364149 267683 364215 267686
rect 366357 267683 366423 267686
rect 417926 267744 418403 267746
rect 417926 267688 418342 267744
rect 418398 267688 418403 267744
rect 417926 267686 418403 267688
rect 411989 267610 412055 267613
rect 412725 267610 412791 267613
rect 411989 267608 412791 267610
rect 411989 267552 411994 267608
rect 412050 267552 412730 267608
rect 412786 267552 412791 267608
rect 411989 267550 412791 267552
rect 411989 267547 412055 267550
rect 412725 267547 412791 267550
rect 415117 267610 415183 267613
rect 417926 267610 417986 267686
rect 418337 267683 418403 267686
rect 433241 267746 433307 267749
rect 437289 267746 437355 267749
rect 433241 267744 437355 267746
rect 433241 267688 433246 267744
rect 433302 267688 437294 267744
rect 437350 267688 437355 267744
rect 433241 267686 437355 267688
rect 433241 267683 433307 267686
rect 437289 267683 437355 267686
rect 485865 267746 485931 267749
rect 492765 267746 492831 267749
rect 485865 267744 492831 267746
rect 485865 267688 485870 267744
rect 485926 267688 492770 267744
rect 492826 267688 492831 267744
rect 485865 267686 492831 267688
rect 485865 267683 485931 267686
rect 492765 267683 492831 267686
rect 415117 267608 417986 267610
rect 415117 267552 415122 267608
rect 415178 267552 417986 267608
rect 415117 267550 417986 267552
rect 421097 267610 421163 267613
rect 424225 267610 424291 267613
rect 421097 267608 424291 267610
rect 421097 267552 421102 267608
rect 421158 267552 424230 267608
rect 424286 267552 424291 267608
rect 421097 267550 424291 267552
rect 415117 267547 415183 267550
rect 421097 267547 421163 267550
rect 424225 267547 424291 267550
rect 424961 267610 425027 267613
rect 427905 267610 427971 267613
rect 424961 267608 427971 267610
rect 424961 267552 424966 267608
rect 425022 267552 427910 267608
rect 427966 267552 427971 267608
rect 424961 267550 427971 267552
rect 424961 267547 425027 267550
rect 427905 267547 427971 267550
rect 446765 267610 446831 267613
rect 447409 267610 447475 267613
rect 446765 267608 447475 267610
rect 446765 267552 446770 267608
rect 446826 267552 447414 267608
rect 447470 267552 447475 267608
rect 446765 267550 447475 267552
rect 446765 267547 446831 267550
rect 447409 267547 447475 267550
rect 475745 267610 475811 267613
rect 476113 267610 476179 267613
rect 475745 267608 476179 267610
rect 475745 267552 475750 267608
rect 475806 267552 476118 267608
rect 476174 267552 476179 267608
rect 475745 267550 476179 267552
rect 475745 267547 475811 267550
rect 476113 267547 476179 267550
rect 476297 267610 476363 267613
rect 482277 267610 482343 267613
rect 476297 267608 482343 267610
rect 476297 267552 476302 267608
rect 476358 267552 482282 267608
rect 482338 267552 482343 267608
rect 476297 267550 482343 267552
rect 476297 267547 476363 267550
rect 482277 267547 482343 267550
rect 499941 267610 500007 267613
rect 578877 267610 578943 267613
rect 499941 267608 578943 267610
rect 499941 267552 499946 267608
rect 500002 267552 578882 267608
rect 578938 267552 578943 267608
rect 499941 267550 578943 267552
rect 499941 267547 500007 267550
rect 578877 267547 578943 267550
rect 377673 267474 377739 267477
rect 379513 267474 379579 267477
rect 377673 267472 379579 267474
rect 377673 267416 377678 267472
rect 377734 267416 379518 267472
rect 379574 267416 379579 267472
rect 377673 267414 379579 267416
rect 377673 267411 377739 267414
rect 379513 267411 379579 267414
rect 675477 267474 675543 267477
rect 675477 267472 676292 267474
rect 675477 267416 675482 267472
rect 675538 267416 676292 267472
rect 675477 267414 676292 267416
rect 675477 267411 675543 267414
rect 412633 267338 412699 267341
rect 416313 267338 416379 267341
rect 412633 267336 416379 267338
rect 412633 267280 412638 267336
rect 412694 267280 416318 267336
rect 416374 267280 416379 267336
rect 412633 267278 416379 267280
rect 412633 267275 412699 267278
rect 416313 267275 416379 267278
rect 419257 267338 419323 267341
rect 518893 267338 518959 267341
rect 419257 267336 518959 267338
rect 419257 267280 419262 267336
rect 419318 267280 518898 267336
rect 518954 267280 518959 267336
rect 419257 267278 518959 267280
rect 419257 267275 419323 267278
rect 518893 267275 518959 267278
rect 401133 267202 401199 267205
rect 402605 267202 402671 267205
rect 401133 267200 402671 267202
rect 401133 267144 401138 267200
rect 401194 267144 402610 267200
rect 402666 267144 402671 267200
rect 401133 267142 402671 267144
rect 401133 267139 401199 267142
rect 402605 267139 402671 267142
rect 383653 267066 383719 267069
rect 384665 267066 384731 267069
rect 383653 267064 384731 267066
rect 383653 267008 383658 267064
rect 383714 267008 384670 267064
rect 384726 267008 384731 267064
rect 383653 267006 384731 267008
rect 383653 267003 383719 267006
rect 384665 267003 384731 267006
rect 388989 267066 389055 267069
rect 393313 267066 393379 267069
rect 388989 267064 393379 267066
rect 388989 267008 388994 267064
rect 389050 267008 393318 267064
rect 393374 267008 393379 267064
rect 388989 267006 393379 267008
rect 388989 267003 389055 267006
rect 393313 267003 393379 267006
rect 446765 267066 446831 267069
rect 447225 267066 447291 267069
rect 446765 267064 447291 267066
rect 446765 267008 446770 267064
rect 446826 267008 447230 267064
rect 447286 267008 447291 267064
rect 446765 267006 447291 267008
rect 446765 267003 446831 267006
rect 447225 267003 447291 267006
rect 450905 267066 450971 267069
rect 457253 267066 457319 267069
rect 450905 267064 457319 267066
rect 450905 267008 450910 267064
rect 450966 267008 457258 267064
rect 457314 267008 457319 267064
rect 450905 267006 457319 267008
rect 450905 267003 450971 267006
rect 457253 267003 457319 267006
rect 466269 267066 466335 267069
rect 466729 267066 466795 267069
rect 466269 267064 466795 267066
rect 466269 267008 466274 267064
rect 466330 267008 466734 267064
rect 466790 267008 466795 267064
rect 466269 267006 466795 267008
rect 466269 267003 466335 267006
rect 466729 267003 466795 267006
rect 474641 267066 474707 267069
rect 476205 267066 476271 267069
rect 474641 267064 476271 267066
rect 474641 267008 474646 267064
rect 474702 267008 476210 267064
rect 476266 267008 476271 267064
rect 474641 267006 476271 267008
rect 474641 267003 474707 267006
rect 476205 267003 476271 267006
rect 485589 267066 485655 267069
rect 490005 267066 490071 267069
rect 485589 267064 490071 267066
rect 485589 267008 485594 267064
rect 485650 267008 490010 267064
rect 490066 267008 490071 267064
rect 485589 267006 490071 267008
rect 485589 267003 485655 267006
rect 490005 267003 490071 267006
rect 498009 267066 498075 267069
rect 504817 267066 504883 267069
rect 585777 267066 585843 267069
rect 498009 267064 504883 267066
rect 498009 267008 498014 267064
rect 498070 267008 504822 267064
rect 504878 267008 504883 267064
rect 498009 267006 504883 267008
rect 498009 267003 498075 267006
rect 504817 267003 504883 267006
rect 505050 267064 585843 267066
rect 505050 267008 585782 267064
rect 585838 267008 585843 267064
rect 505050 267006 585843 267008
rect 428549 266930 428615 266933
rect 437289 266930 437355 266933
rect 428549 266928 437355 266930
rect 428549 266872 428554 266928
rect 428610 266872 437294 266928
rect 437350 266872 437355 266928
rect 428549 266870 437355 266872
rect 428549 266867 428615 266870
rect 437289 266867 437355 266870
rect 490189 266930 490255 266933
rect 491201 266930 491267 266933
rect 490189 266928 491267 266930
rect 490189 266872 490194 266928
rect 490250 266872 491206 266928
rect 491262 266872 491267 266928
rect 490189 266870 491267 266872
rect 490189 266867 490255 266870
rect 491201 266867 491267 266870
rect 446581 266794 446647 266797
rect 454769 266794 454835 266797
rect 446581 266792 454835 266794
rect 446581 266736 446586 266792
rect 446642 266736 454774 266792
rect 454830 266736 454835 266792
rect 446581 266734 454835 266736
rect 446581 266731 446647 266734
rect 454769 266731 454835 266734
rect 457161 266794 457227 266797
rect 462773 266794 462839 266797
rect 457161 266792 462839 266794
rect 457161 266736 457166 266792
rect 457222 266736 462778 266792
rect 462834 266736 462839 266792
rect 457161 266734 462839 266736
rect 457161 266731 457227 266734
rect 462773 266731 462839 266734
rect 463601 266794 463667 266797
rect 466545 266794 466611 266797
rect 463601 266792 466611 266794
rect 463601 266736 463606 266792
rect 463662 266736 466550 266792
rect 466606 266736 466611 266792
rect 463601 266734 466611 266736
rect 463601 266731 463667 266734
rect 466545 266731 466611 266734
rect 492121 266794 492187 266797
rect 499941 266794 500007 266797
rect 505050 266794 505110 267006
rect 585777 267003 585843 267006
rect 675293 267066 675359 267069
rect 675293 267064 676292 267066
rect 675293 267008 675298 267064
rect 675354 267008 676292 267064
rect 675293 267006 676292 267008
rect 675293 267003 675359 267006
rect 492121 266792 500007 266794
rect 492121 266736 492126 266792
rect 492182 266736 499946 266792
rect 500002 266736 500007 266792
rect 492121 266734 500007 266736
rect 492121 266731 492187 266734
rect 499941 266731 500007 266734
rect 500174 266734 505110 266794
rect 436737 266522 436803 266525
rect 437933 266522 437999 266525
rect 436737 266520 437999 266522
rect 436737 266464 436742 266520
rect 436798 266464 437938 266520
rect 437994 266464 437999 266520
rect 436737 266462 437999 266464
rect 436737 266459 436803 266462
rect 437933 266459 437999 266462
rect 483289 266522 483355 266525
rect 500174 266522 500234 266734
rect 675477 266658 675543 266661
rect 675477 266656 676292 266658
rect 675477 266600 675482 266656
rect 675538 266600 676292 266656
rect 675477 266598 676292 266600
rect 675477 266595 675543 266598
rect 483289 266520 500234 266522
rect 483289 266464 483294 266520
rect 483350 266464 500234 266520
rect 483289 266462 500234 266464
rect 504725 266522 504791 266525
rect 507117 266522 507183 266525
rect 504725 266520 507183 266522
rect 504725 266464 504730 266520
rect 504786 266464 507122 266520
rect 507178 266464 507183 266520
rect 504725 266462 507183 266464
rect 483289 266459 483355 266462
rect 504725 266459 504791 266462
rect 507117 266459 507183 266462
rect 441705 266386 441771 266389
rect 442901 266386 442967 266389
rect 441705 266384 442967 266386
rect 441705 266328 441710 266384
rect 441766 266328 442906 266384
rect 442962 266328 442967 266384
rect 441705 266326 442967 266328
rect 441705 266323 441771 266326
rect 442901 266323 442967 266326
rect 466545 266386 466611 266389
rect 473905 266386 473971 266389
rect 466545 266384 473971 266386
rect 466545 266328 466550 266384
rect 466606 266328 473910 266384
rect 473966 266328 473971 266384
rect 466545 266326 473971 266328
rect 466545 266323 466611 266326
rect 473905 266323 473971 266326
rect 435081 266250 435147 266253
rect 437749 266250 437815 266253
rect 435081 266248 437815 266250
rect 435081 266192 435086 266248
rect 435142 266192 437754 266248
rect 437810 266192 437815 266248
rect 435081 266190 437815 266192
rect 435081 266187 435147 266190
rect 437749 266187 437815 266190
rect 675477 266250 675543 266253
rect 675477 266248 676292 266250
rect 675477 266192 675482 266248
rect 675538 266192 676292 266248
rect 675477 266190 676292 266192
rect 675477 266187 675543 266190
rect 462681 266114 462747 266117
rect 589273 266114 589339 266117
rect 462681 266112 589339 266114
rect 462681 266056 462686 266112
rect 462742 266056 589278 266112
rect 589334 266056 589339 266112
rect 462681 266054 589339 266056
rect 462681 266051 462747 266054
rect 589273 266051 589339 266054
rect 461393 265842 461459 265845
rect 462129 265842 462195 265845
rect 461393 265840 462195 265842
rect 461393 265784 461398 265840
rect 461454 265784 462134 265840
rect 462190 265784 462195 265840
rect 461393 265782 462195 265784
rect 461393 265779 461459 265782
rect 462129 265779 462195 265782
rect 481817 265842 481883 265845
rect 619633 265842 619699 265845
rect 481817 265840 619699 265842
rect 481817 265784 481822 265840
rect 481878 265784 619638 265840
rect 619694 265784 619699 265840
rect 481817 265782 619699 265784
rect 481817 265779 481883 265782
rect 619633 265779 619699 265782
rect 675293 265842 675359 265845
rect 675293 265840 676292 265842
rect 675293 265784 675298 265840
rect 675354 265784 676292 265840
rect 675293 265782 676292 265784
rect 675293 265779 675359 265782
rect 54845 265570 54911 265573
rect 658457 265570 658523 265573
rect 54845 265568 658523 265570
rect 54845 265512 54850 265568
rect 54906 265512 658462 265568
rect 658518 265512 658523 265568
rect 54845 265510 658523 265512
rect 54845 265507 54911 265510
rect 658457 265507 658523 265510
rect 675477 265434 675543 265437
rect 675477 265432 676292 265434
rect 675477 265376 675482 265432
rect 675538 265376 676292 265432
rect 675477 265374 676292 265376
rect 675477 265371 675543 265374
rect 479241 265298 479307 265301
rect 485589 265298 485655 265301
rect 479241 265296 485655 265298
rect 479241 265240 479246 265296
rect 479302 265240 485594 265296
rect 485650 265240 485655 265296
rect 479241 265238 485655 265240
rect 479241 265235 479307 265238
rect 485589 265235 485655 265238
rect 675477 265026 675543 265029
rect 675477 265024 676292 265026
rect 675477 264968 675482 265024
rect 675538 264968 676292 265024
rect 675477 264966 676292 264968
rect 675477 264963 675543 264966
rect 675477 264618 675543 264621
rect 675477 264616 676292 264618
rect 675477 264560 675482 264616
rect 675538 264560 676292 264616
rect 675477 264558 676292 264560
rect 675477 264555 675543 264558
rect 674782 264148 674788 264212
rect 674852 264210 674858 264212
rect 674852 264150 676292 264210
rect 674852 264148 674858 264150
rect 676070 263604 676076 263668
rect 676140 263666 676146 263668
rect 676262 263666 676322 263772
rect 676140 263606 676322 263666
rect 676140 263604 676146 263606
rect 676262 263261 676322 263364
rect 676213 263256 676322 263261
rect 676213 263200 676218 263256
rect 676274 263200 676322 263256
rect 676213 263198 676322 263200
rect 676213 263195 676279 263198
rect 676446 262853 676506 262956
rect 676397 262848 676506 262853
rect 676397 262792 676402 262848
rect 676458 262792 676506 262848
rect 676397 262790 676506 262792
rect 676397 262787 676463 262790
rect 511533 262714 511599 262717
rect 508484 262712 511599 262714
rect 508484 262656 511538 262712
rect 511594 262656 511599 262712
rect 508484 262654 511599 262656
rect 511533 262651 511599 262654
rect 675477 262578 675543 262581
rect 675477 262576 676292 262578
rect 675477 262520 675482 262576
rect 675538 262520 676292 262576
rect 675477 262518 676292 262520
rect 675477 262515 675543 262518
rect 675477 262170 675543 262173
rect 675477 262168 676292 262170
rect 675477 262112 675482 262168
rect 675538 262112 676292 262168
rect 675477 262110 676292 262112
rect 675477 262107 675543 262110
rect 676998 261628 677058 261732
rect 676990 261564 676996 261628
rect 677060 261564 677066 261628
rect 674465 261354 674531 261357
rect 674465 261352 676292 261354
rect 674465 261296 674470 261352
rect 674526 261296 676292 261352
rect 674465 261294 676292 261296
rect 674465 261291 674531 261294
rect 674833 261082 674899 261085
rect 675845 261082 675911 261085
rect 674833 261080 675911 261082
rect 674833 261024 674838 261080
rect 674894 261024 675850 261080
rect 675906 261024 675911 261080
rect 674833 261022 675911 261024
rect 674833 261019 674899 261022
rect 675845 261019 675911 261022
rect 676814 260812 676874 260916
rect 676806 260748 676812 260812
rect 676876 260748 676882 260812
rect 675477 260538 675543 260541
rect 675477 260536 676292 260538
rect 675477 260480 675482 260536
rect 675538 260480 676292 260536
rect 675477 260478 676292 260480
rect 675477 260475 675543 260478
rect 510981 260266 511047 260269
rect 508484 260264 511047 260266
rect 508484 260208 510986 260264
rect 511042 260208 511047 260264
rect 508484 260206 511047 260208
rect 510981 260203 511047 260206
rect 675477 260130 675543 260133
rect 675477 260128 676292 260130
rect 675477 260072 675482 260128
rect 675538 260072 676292 260128
rect 675477 260070 676292 260072
rect 675477 260067 675543 260070
rect 675477 259722 675543 259725
rect 675477 259720 676292 259722
rect 675477 259664 675482 259720
rect 675538 259664 676292 259720
rect 675477 259662 676292 259664
rect 675477 259659 675543 259662
rect 40033 259450 40099 259453
rect 46749 259450 46815 259453
rect 40033 259448 46815 259450
rect 40033 259392 40038 259448
rect 40094 259392 46754 259448
rect 46810 259392 46815 259448
rect 40033 259390 46815 259392
rect 40033 259387 40099 259390
rect 46749 259387 46815 259390
rect 674649 259314 674715 259317
rect 674649 259312 676292 259314
rect 674649 259256 674654 259312
rect 674710 259256 676292 259312
rect 674649 259254 676292 259256
rect 674649 259251 674715 259254
rect 40401 258906 40467 258909
rect 44541 258906 44607 258909
rect 40401 258904 44607 258906
rect 40401 258848 40406 258904
rect 40462 258848 44546 258904
rect 44602 258848 44607 258904
rect 40401 258846 44607 258848
rect 40401 258843 40467 258846
rect 44541 258843 44607 258846
rect 675477 258906 675543 258909
rect 675477 258904 676292 258906
rect 675477 258848 675482 258904
rect 675538 258848 676292 258904
rect 675477 258846 676292 258848
rect 675477 258843 675543 258846
rect 675477 258498 675543 258501
rect 675477 258496 676292 258498
rect 675477 258440 675482 258496
rect 675538 258440 676292 258496
rect 675477 258438 676292 258440
rect 675477 258435 675543 258438
rect 35801 258090 35867 258093
rect 35788 258088 35867 258090
rect 35788 258032 35806 258088
rect 35862 258032 35867 258088
rect 35788 258030 35867 258032
rect 35801 258027 35867 258030
rect 39573 257954 39639 257957
rect 43621 257954 43687 257957
rect 39573 257952 43687 257954
rect 39573 257896 39578 257952
rect 39634 257896 43626 257952
rect 43682 257896 43687 257952
rect 39573 257894 43687 257896
rect 39573 257891 39639 257894
rect 43621 257891 43687 257894
rect 510797 257818 510863 257821
rect 508484 257816 510863 257818
rect 508484 257760 510802 257816
rect 510858 257760 510863 257816
rect 508484 257758 510863 257760
rect 510797 257755 510863 257758
rect 35574 257549 35634 257652
rect 683070 257549 683130 258060
rect 35574 257544 35683 257549
rect 35574 257488 35622 257544
rect 35678 257488 35683 257544
rect 35574 257486 35683 257488
rect 35617 257483 35683 257486
rect 39941 257546 40007 257549
rect 43253 257546 43319 257549
rect 39941 257544 43319 257546
rect 39941 257488 39946 257544
rect 40002 257488 43258 257544
rect 43314 257488 43319 257544
rect 39941 257486 43319 257488
rect 683070 257544 683179 257549
rect 683070 257488 683118 257544
rect 683174 257488 683179 257544
rect 683070 257486 683179 257488
rect 39941 257483 40007 257486
rect 43253 257483 43319 257486
rect 683113 257483 683179 257486
rect 675477 257274 675543 257277
rect 675477 257272 676292 257274
rect 35758 257141 35818 257244
rect 675477 257216 675482 257272
rect 675538 257216 676292 257272
rect 675477 257214 676292 257216
rect 675477 257211 675543 257214
rect 35758 257136 35867 257141
rect 35758 257080 35806 257136
rect 35862 257080 35867 257136
rect 35758 257078 35867 257080
rect 35801 257075 35867 257078
rect 35758 256733 35818 256836
rect 35758 256728 35867 256733
rect 35758 256672 35806 256728
rect 35862 256672 35867 256728
rect 35758 256670 35867 256672
rect 35801 256667 35867 256670
rect 40309 256730 40375 256733
rect 45185 256730 45251 256733
rect 40309 256728 45251 256730
rect 40309 256672 40314 256728
rect 40370 256672 45190 256728
rect 45246 256672 45251 256728
rect 40309 256670 45251 256672
rect 40309 256667 40375 256670
rect 45185 256667 45251 256670
rect 35758 256325 35818 256428
rect 35758 256320 35867 256325
rect 35758 256264 35806 256320
rect 35862 256264 35867 256320
rect 35758 256262 35867 256264
rect 35801 256259 35867 256262
rect 35574 255917 35634 256020
rect 35574 255912 35683 255917
rect 35574 255856 35622 255912
rect 35678 255856 35683 255912
rect 35574 255854 35683 255856
rect 35617 255851 35683 255854
rect 35758 255509 35818 255612
rect 35758 255504 35867 255509
rect 35758 255448 35806 255504
rect 35862 255448 35867 255504
rect 35758 255446 35867 255448
rect 35801 255443 35867 255446
rect 511533 255370 511599 255373
rect 508484 255368 511599 255370
rect 508484 255312 511538 255368
rect 511594 255312 511599 255368
rect 508484 255310 511599 255312
rect 511533 255307 511599 255310
rect 35390 255101 35450 255204
rect 35341 255096 35450 255101
rect 35341 255040 35346 255096
rect 35402 255040 35450 255096
rect 35341 255038 35450 255040
rect 41413 255098 41479 255101
rect 44173 255098 44239 255101
rect 41413 255096 44239 255098
rect 41413 255040 41418 255096
rect 41474 255040 44178 255096
rect 44234 255040 44239 255096
rect 41413 255038 44239 255040
rect 35341 255035 35407 255038
rect 41413 255035 41479 255038
rect 44173 255035 44239 255038
rect 35206 254693 35266 254796
rect 35157 254688 35266 254693
rect 35157 254632 35162 254688
rect 35218 254632 35266 254688
rect 35157 254630 35266 254632
rect 35157 254627 35223 254630
rect 35758 254285 35818 254388
rect 35525 254282 35591 254285
rect 35525 254280 35634 254282
rect 35525 254224 35530 254280
rect 35586 254224 35634 254280
rect 35525 254219 35634 254224
rect 35758 254280 35867 254285
rect 35758 254224 35806 254280
rect 35862 254224 35867 254280
rect 35758 254222 35867 254224
rect 35801 254219 35867 254222
rect 35574 253980 35634 254219
rect 675017 254010 675083 254013
rect 675845 254010 675911 254013
rect 675017 254008 675911 254010
rect 675017 253952 675022 254008
rect 675078 253952 675850 254008
rect 675906 253952 675911 254008
rect 675017 253950 675911 253952
rect 675017 253947 675083 253950
rect 675845 253947 675911 253950
rect 35758 253469 35818 253572
rect 35758 253464 35867 253469
rect 35758 253408 35806 253464
rect 35862 253408 35867 253464
rect 35758 253406 35867 253408
rect 35801 253403 35867 253406
rect 35574 253061 35634 253164
rect 35574 253056 35683 253061
rect 35574 253000 35622 253056
rect 35678 253000 35683 253056
rect 35574 252998 35683 253000
rect 35617 252995 35683 252998
rect 39297 253058 39363 253061
rect 42885 253058 42951 253061
rect 39297 253056 42951 253058
rect 39297 253000 39302 253056
rect 39358 253000 42890 253056
rect 42946 253000 42951 253056
rect 39297 252998 42951 253000
rect 39297 252995 39363 252998
rect 42885 252995 42951 252998
rect 511901 252922 511967 252925
rect 508484 252920 511967 252922
rect 508484 252864 511906 252920
rect 511962 252864 511967 252920
rect 508484 252862 511967 252864
rect 511901 252859 511967 252862
rect 35758 252653 35818 252756
rect 35758 252648 35867 252653
rect 35758 252592 35806 252648
rect 35862 252592 35867 252648
rect 35758 252590 35867 252592
rect 35801 252587 35867 252590
rect 41505 252650 41571 252653
rect 46933 252650 46999 252653
rect 41505 252648 46999 252650
rect 41505 252592 41510 252648
rect 41566 252592 46938 252648
rect 46994 252592 46999 252648
rect 41505 252590 46999 252592
rect 41505 252587 41571 252590
rect 46933 252587 46999 252590
rect 35758 252245 35818 252348
rect 35758 252240 35867 252245
rect 35758 252184 35806 252240
rect 35862 252184 35867 252240
rect 35758 252182 35867 252184
rect 35801 252179 35867 252182
rect 40585 252242 40651 252245
rect 42517 252242 42583 252245
rect 40585 252240 42583 252242
rect 40585 252184 40590 252240
rect 40646 252184 42522 252240
rect 42578 252184 42583 252240
rect 40585 252182 42583 252184
rect 40585 252179 40651 252182
rect 42517 252179 42583 252182
rect 35574 251837 35634 251940
rect 35574 251832 35683 251837
rect 35574 251776 35622 251832
rect 35678 251776 35683 251832
rect 35574 251774 35683 251776
rect 35617 251771 35683 251774
rect 41321 251834 41387 251837
rect 45185 251834 45251 251837
rect 41321 251832 45251 251834
rect 41321 251776 41326 251832
rect 41382 251776 45190 251832
rect 45246 251776 45251 251832
rect 41321 251774 45251 251776
rect 41321 251771 41387 251774
rect 45185 251771 45251 251774
rect 35758 251429 35818 251532
rect 35758 251424 35867 251429
rect 35758 251368 35806 251424
rect 35862 251368 35867 251424
rect 35758 251366 35867 251368
rect 35801 251363 35867 251366
rect 41505 251426 41571 251429
rect 45829 251426 45895 251429
rect 41505 251424 45895 251426
rect 41505 251368 41510 251424
rect 41566 251368 45834 251424
rect 45890 251368 45895 251424
rect 41505 251366 45895 251368
rect 41505 251363 41571 251366
rect 45829 251363 45895 251366
rect 35390 251021 35450 251124
rect 35390 251016 35499 251021
rect 35390 250960 35438 251016
rect 35494 250960 35499 251016
rect 35390 250958 35499 250960
rect 35433 250955 35499 250958
rect 35574 250613 35634 250716
rect 35574 250608 35683 250613
rect 35574 250552 35622 250608
rect 35678 250552 35683 250608
rect 35574 250550 35683 250552
rect 35617 250547 35683 250550
rect 510797 250474 510863 250477
rect 508484 250472 510863 250474
rect 508484 250416 510802 250472
rect 510858 250416 510863 250472
rect 508484 250414 510863 250416
rect 510797 250411 510863 250414
rect 35758 250205 35818 250308
rect 35758 250200 35867 250205
rect 35758 250144 35806 250200
rect 35862 250144 35867 250200
rect 35758 250142 35867 250144
rect 35801 250139 35867 250142
rect 39389 250202 39455 250205
rect 43069 250202 43135 250205
rect 39389 250200 43135 250202
rect 39389 250144 39394 250200
rect 39450 250144 43074 250200
rect 43130 250144 43135 250200
rect 39389 250142 43135 250144
rect 39389 250139 39455 250142
rect 43069 250139 43135 250142
rect 40726 249796 40786 249900
rect 673913 249796 673979 249797
rect 40718 249732 40724 249796
rect 40788 249732 40794 249796
rect 673862 249794 673868 249796
rect 673822 249734 673868 249794
rect 673932 249792 673979 249796
rect 673974 249736 673979 249792
rect 673862 249732 673868 249734
rect 673932 249732 673979 249736
rect 674782 249732 674788 249796
rect 674852 249732 674858 249796
rect 675201 249794 675267 249797
rect 676070 249794 676076 249796
rect 675201 249792 676076 249794
rect 675201 249736 675206 249792
rect 675262 249736 676076 249792
rect 675201 249734 676076 249736
rect 673913 249731 673979 249732
rect 674790 249522 674850 249732
rect 675201 249731 675267 249734
rect 676070 249732 676076 249734
rect 676140 249732 676146 249796
rect 675569 249522 675635 249525
rect 674790 249520 675635 249522
rect 40542 249388 40602 249492
rect 674790 249464 675574 249520
rect 675630 249464 675635 249520
rect 674790 249462 675635 249464
rect 675569 249459 675635 249462
rect 40534 249324 40540 249388
rect 40604 249324 40610 249388
rect 35574 248981 35634 249084
rect 35525 248976 35634 248981
rect 35801 248978 35867 248981
rect 35525 248920 35530 248976
rect 35586 248920 35634 248976
rect 35525 248918 35634 248920
rect 35758 248976 35867 248978
rect 35758 248920 35806 248976
rect 35862 248920 35867 248976
rect 35525 248915 35591 248918
rect 35758 248915 35867 248920
rect 40125 248978 40191 248981
rect 43253 248978 43319 248981
rect 40125 248976 43319 248978
rect 40125 248920 40130 248976
rect 40186 248920 43258 248976
rect 43314 248920 43319 248976
rect 40125 248918 43319 248920
rect 40125 248915 40191 248918
rect 43253 248915 43319 248918
rect 35758 248676 35818 248915
rect 39941 248570 40007 248573
rect 43621 248570 43687 248573
rect 39941 248568 43687 248570
rect 39941 248512 39946 248568
rect 40002 248512 43626 248568
rect 43682 248512 43687 248568
rect 39941 248510 43687 248512
rect 39941 248507 40007 248510
rect 43621 248507 43687 248510
rect 675385 248298 675451 248301
rect 676990 248298 676996 248300
rect 675385 248296 676996 248298
rect 35574 248165 35634 248268
rect 675385 248240 675390 248296
rect 675446 248240 676996 248296
rect 675385 248238 676996 248240
rect 675385 248235 675451 248238
rect 676990 248236 676996 248238
rect 677060 248236 677066 248300
rect 35574 248160 35683 248165
rect 35574 248104 35622 248160
rect 35678 248104 35683 248160
rect 35574 248102 35683 248104
rect 35617 248099 35683 248102
rect 40125 248162 40191 248165
rect 44541 248162 44607 248165
rect 40125 248160 44607 248162
rect 40125 248104 40130 248160
rect 40186 248104 44546 248160
rect 44602 248104 44607 248160
rect 40125 248102 44607 248104
rect 40125 248099 40191 248102
rect 44541 248099 44607 248102
rect 510981 248026 511047 248029
rect 508484 248024 511047 248026
rect 508484 247968 510986 248024
rect 511042 247968 511047 248024
rect 508484 247966 511047 247968
rect 510981 247963 511047 247966
rect 35390 247757 35450 247860
rect 35390 247752 35499 247757
rect 35390 247696 35438 247752
rect 35494 247696 35499 247752
rect 35390 247694 35499 247696
rect 35433 247691 35499 247694
rect 41505 247754 41571 247757
rect 42149 247754 42215 247757
rect 41505 247752 42215 247754
rect 41505 247696 41510 247752
rect 41566 247696 42154 247752
rect 42210 247696 42215 247752
rect 41505 247694 42215 247696
rect 41505 247691 41571 247694
rect 42149 247691 42215 247694
rect 35758 247349 35818 247452
rect 35758 247344 35867 247349
rect 35758 247288 35806 247344
rect 35862 247288 35867 247344
rect 35758 247286 35867 247288
rect 35801 247283 35867 247286
rect 40125 247346 40191 247349
rect 44357 247346 44423 247349
rect 40125 247344 44423 247346
rect 40125 247288 40130 247344
rect 40186 247288 44362 247344
rect 44418 247288 44423 247344
rect 40125 247286 44423 247288
rect 40125 247283 40191 247286
rect 44357 247283 44423 247286
rect 35574 246941 35634 247044
rect 35574 246936 35683 246941
rect 35574 246880 35622 246936
rect 35678 246880 35683 246936
rect 35574 246878 35683 246880
rect 35617 246875 35683 246878
rect 41505 246938 41571 246941
rect 42057 246938 42123 246941
rect 41505 246936 42123 246938
rect 41505 246880 41510 246936
rect 41566 246880 42062 246936
rect 42118 246880 42123 246936
rect 41505 246878 42123 246880
rect 41505 246875 41571 246878
rect 42057 246875 42123 246878
rect 675753 246666 675819 246669
rect 676806 246666 676812 246668
rect 675753 246664 676812 246666
rect 41462 246530 41522 246636
rect 675753 246608 675758 246664
rect 675814 246608 676812 246664
rect 675753 246606 676812 246608
rect 675753 246603 675819 246606
rect 676806 246604 676812 246606
rect 676876 246604 676882 246668
rect 41462 246470 51090 246530
rect 41045 246122 41111 246125
rect 46013 246122 46079 246125
rect 41045 246120 46079 246122
rect 41045 246064 41050 246120
rect 41106 246064 46018 246120
rect 46074 246064 46079 246120
rect 41045 246062 46079 246064
rect 41045 246059 41111 246062
rect 46013 246059 46079 246062
rect 51030 245714 51090 246470
rect 666870 246060 666876 246124
rect 666940 246122 666946 246124
rect 667381 246122 667447 246125
rect 666940 246120 667447 246122
rect 666940 246064 667386 246120
rect 667442 246064 667447 246120
rect 666940 246062 667447 246064
rect 666940 246060 666946 246062
rect 667381 246059 667447 246062
rect 666502 245924 666508 245988
rect 666572 245986 666578 245988
rect 666737 245986 666803 245989
rect 668117 245988 668183 245989
rect 668117 245986 668164 245988
rect 666572 245984 666803 245986
rect 666572 245928 666742 245984
rect 666798 245928 666803 245984
rect 666572 245926 666803 245928
rect 668072 245984 668164 245986
rect 668072 245928 668122 245984
rect 668072 245926 668164 245928
rect 666572 245924 666578 245926
rect 666737 245923 666803 245926
rect 668117 245924 668164 245926
rect 668228 245924 668234 245988
rect 668117 245923 668183 245924
rect 131757 245714 131823 245717
rect 51030 245712 131823 245714
rect 51030 245656 131762 245712
rect 131818 245656 131823 245712
rect 51030 245654 131823 245656
rect 131757 245651 131823 245654
rect 666686 245652 666692 245716
rect 666756 245714 666762 245716
rect 666921 245714 666987 245717
rect 668301 245716 668367 245717
rect 668301 245714 668348 245716
rect 666756 245712 666987 245714
rect 666756 245656 666926 245712
rect 666982 245656 666987 245712
rect 666756 245654 666987 245656
rect 668256 245712 668348 245714
rect 668256 245656 668306 245712
rect 668256 245654 668348 245656
rect 666756 245652 666762 245654
rect 666921 245651 666987 245654
rect 668301 245652 668348 245654
rect 668412 245652 668418 245716
rect 671889 245714 671955 245717
rect 675385 245714 675451 245717
rect 671889 245712 675451 245714
rect 671889 245656 671894 245712
rect 671950 245656 675390 245712
rect 675446 245656 675451 245712
rect 671889 245654 675451 245656
rect 668301 245651 668367 245652
rect 671889 245651 671955 245654
rect 675385 245651 675451 245654
rect 39573 245578 39639 245581
rect 47117 245578 47183 245581
rect 511257 245578 511323 245581
rect 39573 245576 47183 245578
rect 39573 245520 39578 245576
rect 39634 245520 47122 245576
rect 47178 245520 47183 245576
rect 39573 245518 47183 245520
rect 508484 245576 511323 245578
rect 508484 245520 511262 245576
rect 511318 245520 511323 245576
rect 508484 245518 511323 245520
rect 39573 245515 39639 245518
rect 47117 245515 47183 245518
rect 511257 245515 511323 245518
rect 675293 243268 675359 243269
rect 675293 243266 675340 243268
rect 675248 243264 675340 243266
rect 675248 243208 675298 243264
rect 675248 243206 675340 243208
rect 675293 243204 675340 243206
rect 675404 243204 675410 243268
rect 675293 243203 675359 243204
rect 511901 243130 511967 243133
rect 508484 243128 511967 243130
rect 508484 243072 511906 243128
rect 511962 243072 511967 243128
rect 508484 243070 511967 243072
rect 511901 243067 511967 243070
rect 674557 242722 674623 242725
rect 675477 242722 675543 242725
rect 674557 242720 675543 242722
rect 674557 242664 674562 242720
rect 674618 242664 675482 242720
rect 675538 242664 675543 242720
rect 674557 242662 675543 242664
rect 674557 242659 674623 242662
rect 675477 242659 675543 242662
rect 669129 242042 669195 242045
rect 675477 242042 675543 242045
rect 669129 242040 675543 242042
rect 669129 241984 669134 242040
rect 669190 241984 675482 242040
rect 675538 241984 675543 242040
rect 669129 241982 675543 241984
rect 669129 241979 669195 241982
rect 675477 241979 675543 241982
rect 672901 241770 672967 241773
rect 675109 241770 675175 241773
rect 672901 241768 675175 241770
rect 672901 241712 672906 241768
rect 672962 241712 675114 241768
rect 675170 241712 675175 241768
rect 672901 241710 675175 241712
rect 672901 241707 672967 241710
rect 675109 241707 675175 241710
rect 511073 240682 511139 240685
rect 508484 240680 511139 240682
rect 508484 240624 511078 240680
rect 511134 240624 511139 240680
rect 508484 240622 511139 240624
rect 511073 240619 511139 240622
rect 675385 238644 675451 238645
rect 675334 238642 675340 238644
rect 675294 238582 675340 238642
rect 675404 238640 675451 238644
rect 675446 238584 675451 238640
rect 675334 238580 675340 238582
rect 675404 238580 675451 238584
rect 675385 238579 675451 238580
rect 42241 238506 42307 238509
rect 46013 238506 46079 238509
rect 42241 238504 46079 238506
rect 42241 238448 42246 238504
rect 42302 238448 46018 238504
rect 46074 238448 46079 238504
rect 42241 238446 46079 238448
rect 42241 238443 42307 238446
rect 46013 238443 46079 238446
rect 511257 238234 511323 238237
rect 508484 238232 511323 238234
rect 508484 238176 511262 238232
rect 511318 238176 511323 238232
rect 508484 238174 511323 238176
rect 511257 238171 511323 238174
rect 42374 237356 42380 237420
rect 42444 237418 42450 237420
rect 42701 237418 42767 237421
rect 42444 237416 42767 237418
rect 42444 237360 42706 237416
rect 42762 237360 42767 237416
rect 42444 237358 42767 237360
rect 42444 237356 42450 237358
rect 42701 237355 42767 237358
rect 40718 236540 40724 236604
rect 40788 236602 40794 236604
rect 41781 236602 41847 236605
rect 40788 236600 41847 236602
rect 40788 236544 41786 236600
rect 41842 236544 41847 236600
rect 40788 236542 41847 236544
rect 40788 236540 40794 236542
rect 41781 236539 41847 236542
rect 510889 235786 510955 235789
rect 508484 235784 510955 235786
rect 508484 235728 510894 235784
rect 510950 235728 510955 235784
rect 508484 235726 510955 235728
rect 510889 235723 510955 235726
rect 40534 234500 40540 234564
rect 40604 234562 40610 234564
rect 41781 234562 41847 234565
rect 40604 234560 41847 234562
rect 40604 234504 41786 234560
rect 41842 234504 41847 234560
rect 40604 234502 41847 234504
rect 40604 234500 40610 234502
rect 41781 234499 41847 234502
rect 507534 233069 507594 233308
rect 507485 233064 507594 233069
rect 507485 233008 507490 233064
rect 507546 233008 507594 233064
rect 507485 233006 507594 233008
rect 507485 233003 507551 233006
rect 147121 231298 147187 231301
rect 148685 231298 148751 231301
rect 147121 231296 148751 231298
rect 147121 231240 147126 231296
rect 147182 231240 148690 231296
rect 148746 231240 148751 231296
rect 147121 231238 148751 231240
rect 147121 231235 147187 231238
rect 148685 231235 148751 231238
rect 148869 231298 148935 231301
rect 153009 231298 153075 231301
rect 148869 231296 153075 231298
rect 148869 231240 148874 231296
rect 148930 231240 153014 231296
rect 153070 231240 153075 231296
rect 148869 231238 153075 231240
rect 148869 231235 148935 231238
rect 153009 231235 153075 231238
rect 157609 231162 157675 231165
rect 169293 231162 169359 231165
rect 157609 231160 169359 231162
rect 157609 231104 157614 231160
rect 157670 231104 169298 231160
rect 169354 231104 169359 231160
rect 157609 231102 169359 231104
rect 157609 231099 157675 231102
rect 169293 231099 169359 231102
rect 147806 230964 147812 231028
rect 147876 231026 147882 231028
rect 149421 231026 149487 231029
rect 147876 231024 149487 231026
rect 147876 230968 149426 231024
rect 149482 230968 149487 231024
rect 147876 230966 149487 230968
rect 147876 230964 147882 230966
rect 149421 230963 149487 230966
rect 176837 231026 176903 231029
rect 178309 231026 178375 231029
rect 176837 231024 178375 231026
rect 176837 230968 176842 231024
rect 176898 230968 178314 231024
rect 178370 230968 178375 231024
rect 176837 230966 178375 230968
rect 176837 230963 176903 230966
rect 178309 230963 178375 230966
rect 144269 230890 144335 230893
rect 147305 230890 147371 230893
rect 144269 230888 147371 230890
rect 144269 230832 144274 230888
rect 144330 230832 147310 230888
rect 147366 230832 147371 230888
rect 144269 230830 147371 230832
rect 144269 230827 144335 230830
rect 147305 230827 147371 230830
rect 159817 230754 159883 230757
rect 167821 230754 167887 230757
rect 159817 230752 167887 230754
rect 159817 230696 159822 230752
rect 159878 230696 167826 230752
rect 167882 230696 167887 230752
rect 159817 230694 167887 230696
rect 159817 230691 159883 230694
rect 167821 230691 167887 230694
rect 176009 230754 176075 230757
rect 177573 230754 177639 230757
rect 176009 230752 177639 230754
rect 176009 230696 176014 230752
rect 176070 230696 177578 230752
rect 177634 230696 177639 230752
rect 176009 230694 177639 230696
rect 176009 230691 176075 230694
rect 177573 230691 177639 230694
rect 132861 230618 132927 230621
rect 147305 230618 147371 230621
rect 132861 230616 147371 230618
rect 132861 230560 132866 230616
rect 132922 230560 147310 230616
rect 147366 230560 147371 230616
rect 132861 230558 147371 230560
rect 132861 230555 132927 230558
rect 147305 230555 147371 230558
rect 148685 230618 148751 230621
rect 159541 230618 159607 230621
rect 148685 230616 159607 230618
rect 148685 230560 148690 230616
rect 148746 230560 159546 230616
rect 159602 230560 159607 230616
rect 148685 230558 159607 230560
rect 148685 230555 148751 230558
rect 159541 230555 159607 230558
rect 147806 230482 147812 230484
rect 147630 230422 147812 230482
rect 79317 230346 79383 230349
rect 140773 230346 140839 230349
rect 79317 230344 140839 230346
rect 79317 230288 79322 230344
rect 79378 230288 140778 230344
rect 140834 230288 140839 230344
rect 79317 230286 140839 230288
rect 79317 230283 79383 230286
rect 140773 230283 140839 230286
rect 147029 230346 147095 230349
rect 147630 230346 147690 230422
rect 147806 230420 147812 230422
rect 147876 230420 147882 230484
rect 147029 230344 147690 230346
rect 147029 230288 147034 230344
rect 147090 230288 147690 230344
rect 147029 230286 147690 230288
rect 151721 230346 151787 230349
rect 153285 230346 153351 230349
rect 151721 230344 153351 230346
rect 151721 230288 151726 230344
rect 151782 230288 153290 230344
rect 153346 230288 153351 230344
rect 151721 230286 153351 230288
rect 147029 230283 147095 230286
rect 151721 230283 151787 230286
rect 153285 230283 153351 230286
rect 167177 230346 167243 230349
rect 176377 230346 176443 230349
rect 167177 230344 176443 230346
rect 167177 230288 167182 230344
rect 167238 230288 176382 230344
rect 176438 230288 176443 230344
rect 167177 230286 176443 230288
rect 167177 230283 167243 230286
rect 176377 230283 176443 230286
rect 186129 230346 186195 230349
rect 189165 230346 189231 230349
rect 186129 230344 189231 230346
rect 186129 230288 186134 230344
rect 186190 230288 189170 230344
rect 189226 230288 189231 230344
rect 186129 230286 189231 230288
rect 186129 230283 186195 230286
rect 189165 230283 189231 230286
rect 193029 230346 193095 230349
rect 194593 230346 194659 230349
rect 193029 230344 194659 230346
rect 193029 230288 193034 230344
rect 193090 230288 194598 230344
rect 194654 230288 194659 230344
rect 193029 230286 194659 230288
rect 193029 230283 193095 230286
rect 194593 230283 194659 230286
rect 495433 230346 495499 230349
rect 499849 230346 499915 230349
rect 495433 230344 499915 230346
rect 495433 230288 495438 230344
rect 495494 230288 499854 230344
rect 499910 230288 499915 230344
rect 495433 230286 499915 230288
rect 495433 230283 495499 230286
rect 499849 230283 499915 230286
rect 54661 230074 54727 230077
rect 654317 230074 654383 230077
rect 54661 230072 654383 230074
rect 54661 230016 54666 230072
rect 54722 230016 654322 230072
rect 654378 230016 654383 230072
rect 54661 230014 654383 230016
rect 54661 230011 54727 230014
rect 654317 230011 654383 230014
rect 45001 229802 45067 229805
rect 648613 229802 648679 229805
rect 45001 229800 648679 229802
rect 45001 229744 45006 229800
rect 45062 229744 648618 229800
rect 648674 229744 648679 229800
rect 45001 229742 648679 229744
rect 45001 229739 45067 229742
rect 648613 229739 648679 229742
rect 140773 229530 140839 229533
rect 151905 229530 151971 229533
rect 140773 229528 151971 229530
rect 140773 229472 140778 229528
rect 140834 229472 151910 229528
rect 151966 229472 151971 229528
rect 140773 229470 151971 229472
rect 140773 229467 140839 229470
rect 151905 229467 151971 229470
rect 154113 229530 154179 229533
rect 157609 229530 157675 229533
rect 154113 229528 157675 229530
rect 154113 229472 154118 229528
rect 154174 229472 157614 229528
rect 157670 229472 157675 229528
rect 154113 229470 157675 229472
rect 154113 229467 154179 229470
rect 157609 229467 157675 229470
rect 169201 229530 169267 229533
rect 176561 229530 176627 229533
rect 169201 229528 176627 229530
rect 169201 229472 169206 229528
rect 169262 229472 176566 229528
rect 176622 229472 176627 229528
rect 169201 229470 176627 229472
rect 169201 229467 169267 229470
rect 176561 229467 176627 229470
rect 184841 229530 184907 229533
rect 186129 229530 186195 229533
rect 184841 229528 186195 229530
rect 184841 229472 184846 229528
rect 184902 229472 186134 229528
rect 186190 229472 186195 229528
rect 184841 229470 186195 229472
rect 184841 229467 184907 229470
rect 186129 229467 186195 229470
rect 490189 229530 490255 229533
rect 495617 229530 495683 229533
rect 499665 229530 499731 229533
rect 490189 229528 495450 229530
rect 490189 229472 490194 229528
rect 490250 229472 495450 229528
rect 490189 229470 495450 229472
rect 490189 229467 490255 229470
rect 200113 229394 200179 229397
rect 201401 229394 201467 229397
rect 200113 229392 201467 229394
rect 200113 229336 200118 229392
rect 200174 229336 201406 229392
rect 201462 229336 201467 229392
rect 200113 229334 201467 229336
rect 200113 229331 200179 229334
rect 201401 229331 201467 229334
rect 455873 229394 455939 229397
rect 458817 229394 458883 229397
rect 455873 229392 458883 229394
rect 455873 229336 455878 229392
rect 455934 229336 458822 229392
rect 458878 229336 458883 229392
rect 455873 229334 458883 229336
rect 455873 229331 455939 229334
rect 458817 229331 458883 229334
rect 480161 229394 480227 229397
rect 480529 229394 480595 229397
rect 480161 229392 480595 229394
rect 480161 229336 480166 229392
rect 480222 229336 480534 229392
rect 480590 229336 480595 229392
rect 480161 229334 480595 229336
rect 480161 229331 480227 229334
rect 480529 229331 480595 229334
rect 487337 229394 487403 229397
rect 487337 229392 489930 229394
rect 487337 229336 487342 229392
rect 487398 229336 489930 229392
rect 487337 229334 489930 229336
rect 487337 229331 487403 229334
rect 166349 229258 166415 229261
rect 172329 229258 172395 229261
rect 166349 229256 172395 229258
rect 166349 229200 166354 229256
rect 166410 229200 172334 229256
rect 172390 229200 172395 229256
rect 166349 229198 172395 229200
rect 166349 229195 166415 229198
rect 172329 229195 172395 229198
rect 147489 229122 147555 229125
rect 149973 229122 150039 229125
rect 147489 229120 150039 229122
rect 147489 229064 147494 229120
rect 147550 229064 149978 229120
rect 150034 229064 150039 229120
rect 147489 229062 150039 229064
rect 147489 229059 147555 229062
rect 149973 229059 150039 229062
rect 156321 229122 156387 229125
rect 158161 229122 158227 229125
rect 156321 229120 158227 229122
rect 156321 229064 156326 229120
rect 156382 229064 158166 229120
rect 158222 229064 158227 229120
rect 156321 229062 158227 229064
rect 489870 229122 489930 229334
rect 495390 229258 495450 229470
rect 495617 229528 499731 229530
rect 495617 229472 495622 229528
rect 495678 229472 499670 229528
rect 499726 229472 499731 229528
rect 495617 229470 499731 229472
rect 495617 229467 495683 229470
rect 499665 229467 499731 229470
rect 495893 229258 495959 229261
rect 495390 229256 495959 229258
rect 495390 229200 495898 229256
rect 495954 229200 495959 229256
rect 495390 229198 495959 229200
rect 495893 229195 495959 229198
rect 490189 229122 490255 229125
rect 489870 229120 490255 229122
rect 489870 229064 490194 229120
rect 490250 229064 490255 229120
rect 489870 229062 490255 229064
rect 156321 229059 156387 229062
rect 158161 229059 158227 229062
rect 490189 229059 490255 229062
rect 164785 228986 164851 228989
rect 166993 228986 167059 228989
rect 164785 228984 167059 228986
rect 164785 228928 164790 228984
rect 164846 228928 166998 228984
rect 167054 228928 167059 228984
rect 164785 228926 167059 228928
rect 164785 228923 164851 228926
rect 166993 228923 167059 228926
rect 147305 228850 147371 228853
rect 150985 228850 151051 228853
rect 147305 228848 151051 228850
rect 147305 228792 147310 228848
rect 147366 228792 150990 228848
rect 151046 228792 151051 228848
rect 147305 228790 151051 228792
rect 147305 228787 147371 228790
rect 150985 228787 151051 228790
rect 151353 228850 151419 228853
rect 152917 228850 152983 228853
rect 151353 228848 152983 228850
rect 151353 228792 151358 228848
rect 151414 228792 152922 228848
rect 152978 228792 152983 228848
rect 151353 228790 152983 228792
rect 151353 228787 151419 228790
rect 152917 228787 152983 228790
rect 167177 228850 167243 228853
rect 174905 228850 174971 228853
rect 167177 228848 174971 228850
rect 167177 228792 167182 228848
rect 167238 228792 174910 228848
rect 174966 228792 174971 228848
rect 167177 228790 174971 228792
rect 167177 228787 167243 228790
rect 174905 228787 174971 228790
rect 179045 228850 179111 228853
rect 183277 228850 183343 228853
rect 179045 228848 183343 228850
rect 179045 228792 179050 228848
rect 179106 228792 183282 228848
rect 183338 228792 183343 228848
rect 179045 228790 183343 228792
rect 179045 228787 179111 228790
rect 183277 228787 183343 228790
rect 192661 228850 192727 228853
rect 195697 228850 195763 228853
rect 192661 228848 195763 228850
rect 192661 228792 192666 228848
rect 192722 228792 195702 228848
rect 195758 228792 195763 228848
rect 192661 228790 195763 228792
rect 192661 228787 192727 228790
rect 195697 228787 195763 228790
rect 489913 228850 489979 228853
rect 495801 228850 495867 228853
rect 489913 228848 495867 228850
rect 489913 228792 489918 228848
rect 489974 228792 495806 228848
rect 495862 228792 495867 228848
rect 489913 228790 495867 228792
rect 489913 228787 489979 228790
rect 495801 228787 495867 228790
rect 505093 228850 505159 228853
rect 513557 228850 513623 228853
rect 505093 228848 513623 228850
rect 505093 228792 505098 228848
rect 505154 228792 513562 228848
rect 513618 228792 513623 228848
rect 505093 228790 513623 228792
rect 505093 228787 505159 228790
rect 513557 228787 513623 228790
rect 50337 228578 50403 228581
rect 647233 228578 647299 228581
rect 50337 228576 647299 228578
rect 50337 228520 50342 228576
rect 50398 228520 647238 228576
rect 647294 228520 647299 228576
rect 50337 228518 647299 228520
rect 50337 228515 50403 228518
rect 647233 228515 647299 228518
rect 50521 228306 50587 228309
rect 650545 228306 650611 228309
rect 50521 228304 650611 228306
rect 50521 228248 50526 228304
rect 50582 228248 650550 228304
rect 650606 228248 650611 228304
rect 50521 228246 650611 228248
rect 50521 228243 50587 228246
rect 650545 228243 650611 228246
rect 154757 228034 154823 228037
rect 147998 228032 154823 228034
rect 147998 227976 154762 228032
rect 154818 227976 154823 228032
rect 147998 227974 154823 227976
rect 147998 227901 148058 227974
rect 154757 227971 154823 227974
rect 147949 227896 148058 227901
rect 147949 227840 147954 227896
rect 148010 227840 148058 227896
rect 147949 227838 148058 227840
rect 495433 227898 495499 227901
rect 504909 227898 504975 227901
rect 495433 227896 504975 227898
rect 495433 227840 495438 227896
rect 495494 227840 504914 227896
rect 504970 227840 504975 227896
rect 495433 227838 504975 227840
rect 147949 227835 148015 227838
rect 495433 227835 495499 227838
rect 504909 227835 504975 227838
rect 149513 227762 149579 227765
rect 155493 227762 155559 227765
rect 149513 227760 155559 227762
rect 149513 227704 149518 227760
rect 149574 227704 155498 227760
rect 155554 227704 155559 227760
rect 149513 227702 155559 227704
rect 149513 227699 149579 227702
rect 155493 227699 155559 227702
rect 485313 227762 485379 227765
rect 490741 227762 490807 227765
rect 485313 227760 490807 227762
rect 485313 227704 485318 227760
rect 485374 227704 490746 227760
rect 490802 227704 490807 227760
rect 485313 227702 490807 227704
rect 485313 227699 485379 227702
rect 490741 227699 490807 227702
rect 46381 227490 46447 227493
rect 647509 227490 647575 227493
rect 46381 227488 647575 227490
rect 46381 227432 46386 227488
rect 46442 227432 647514 227488
rect 647570 227432 647575 227488
rect 46381 227430 647575 227432
rect 46381 227427 46447 227430
rect 647509 227427 647575 227430
rect 42057 227354 42123 227357
rect 42374 227354 42380 227356
rect 42057 227352 42380 227354
rect 42057 227296 42062 227352
rect 42118 227296 42380 227352
rect 42057 227294 42380 227296
rect 42057 227291 42123 227294
rect 42374 227292 42380 227294
rect 42444 227292 42450 227356
rect 52085 227218 52151 227221
rect 656341 227218 656407 227221
rect 52085 227216 656407 227218
rect 52085 227160 52090 227216
rect 52146 227160 656346 227216
rect 656402 227160 656407 227216
rect 52085 227158 656407 227160
rect 52085 227155 52151 227158
rect 656341 227155 656407 227158
rect 47761 226946 47827 226949
rect 651649 226946 651715 226949
rect 47761 226944 651715 226946
rect 47761 226888 47766 226944
rect 47822 226888 651654 226944
rect 651710 226888 651715 226944
rect 47761 226886 651715 226888
rect 47761 226883 47827 226886
rect 651649 226883 651715 226886
rect 55857 226674 55923 226677
rect 646405 226674 646471 226677
rect 55857 226672 646471 226674
rect 55857 226616 55862 226672
rect 55918 226616 646410 226672
rect 646466 226616 646471 226672
rect 55857 226614 646471 226616
rect 55857 226611 55923 226614
rect 646405 226611 646471 226614
rect 143441 226402 143507 226405
rect 147673 226402 147739 226405
rect 143441 226400 147739 226402
rect 143441 226344 143446 226400
rect 143502 226344 147678 226400
rect 147734 226344 147739 226400
rect 143441 226342 147739 226344
rect 143441 226339 143507 226342
rect 147673 226339 147739 226342
rect 151077 226402 151143 226405
rect 156873 226402 156939 226405
rect 151077 226400 156939 226402
rect 151077 226344 151082 226400
rect 151138 226344 156878 226400
rect 156934 226344 156939 226400
rect 151077 226342 156939 226344
rect 151077 226339 151143 226342
rect 156873 226339 156939 226342
rect 505093 226402 505159 226405
rect 510153 226402 510219 226405
rect 505093 226400 510219 226402
rect 505093 226344 505098 226400
rect 505154 226344 510158 226400
rect 510214 226344 510219 226400
rect 505093 226342 510219 226344
rect 505093 226339 505159 226342
rect 510153 226339 510219 226342
rect 483657 226266 483723 226269
rect 491937 226266 492003 226269
rect 483657 226264 492003 226266
rect 483657 226208 483662 226264
rect 483718 226208 491942 226264
rect 491998 226208 492003 226264
rect 483657 226206 492003 226208
rect 483657 226203 483723 226206
rect 491937 226203 492003 226206
rect 141601 225994 141667 225997
rect 148501 225994 148567 225997
rect 141601 225992 148567 225994
rect 141601 225936 141606 225992
rect 141662 225936 148506 225992
rect 148562 225936 148567 225992
rect 141601 225934 148567 225936
rect 141601 225931 141667 225934
rect 148501 225931 148567 225934
rect 156505 225994 156571 225997
rect 157425 225994 157491 225997
rect 156505 225992 157491 225994
rect 156505 225936 156510 225992
rect 156566 225936 157430 225992
rect 157486 225936 157491 225992
rect 156505 225934 157491 225936
rect 156505 225931 156571 225934
rect 157425 225931 157491 225934
rect 181253 225994 181319 225997
rect 181989 225994 182055 225997
rect 181253 225992 182055 225994
rect 181253 225936 181258 225992
rect 181314 225936 181994 225992
rect 182050 225936 182055 225992
rect 181253 225934 182055 225936
rect 181253 225931 181319 225934
rect 181989 225931 182055 225934
rect 199285 225994 199351 225997
rect 199837 225994 199903 225997
rect 199285 225992 199903 225994
rect 199285 225936 199290 225992
rect 199346 225936 199842 225992
rect 199898 225936 199903 225992
rect 199285 225934 199903 225936
rect 199285 225931 199351 225934
rect 199837 225931 199903 225934
rect 484301 225994 484367 225997
rect 488073 225994 488139 225997
rect 484301 225992 488139 225994
rect 484301 225936 484306 225992
rect 484362 225936 488078 225992
rect 488134 225936 488139 225992
rect 484301 225934 488139 225936
rect 484301 225931 484367 225934
rect 488073 225931 488139 225934
rect 489867 225994 489933 225997
rect 504909 225994 504975 225997
rect 489867 225992 504975 225994
rect 489867 225936 489872 225992
rect 489928 225936 504914 225992
rect 504970 225936 504975 225992
rect 489867 225934 504975 225936
rect 489867 225931 489933 225934
rect 504909 225931 504975 225934
rect 514569 225994 514635 225997
rect 516777 225994 516843 225997
rect 514569 225992 516843 225994
rect 514569 225936 514574 225992
rect 514630 225936 516782 225992
rect 516838 225936 516843 225992
rect 514569 225934 516843 225936
rect 514569 225931 514635 225934
rect 516777 225931 516843 225934
rect 151537 225722 151603 225725
rect 137970 225720 151603 225722
rect 137970 225664 151542 225720
rect 151598 225664 151603 225720
rect 137970 225662 151603 225664
rect 58985 225586 59051 225589
rect 137970 225586 138030 225662
rect 151537 225659 151603 225662
rect 190177 225722 190243 225725
rect 190729 225722 190795 225725
rect 190177 225720 190795 225722
rect 190177 225664 190182 225720
rect 190238 225664 190734 225720
rect 190790 225664 190795 225720
rect 190177 225662 190795 225664
rect 190177 225659 190243 225662
rect 190729 225659 190795 225662
rect 58985 225584 138030 225586
rect 58985 225528 58990 225584
rect 59046 225528 138030 225584
rect 157287 225618 157353 225623
rect 157287 225562 157292 225618
rect 157348 225586 157353 225618
rect 162301 225586 162367 225589
rect 157348 225584 162367 225586
rect 157348 225562 162306 225584
rect 157287 225557 162306 225562
rect 58985 225526 138030 225528
rect 157290 225528 162306 225557
rect 162362 225528 162367 225584
rect 157290 225526 162367 225528
rect 58985 225523 59051 225526
rect 162301 225523 162367 225526
rect 440969 225586 441035 225589
rect 504725 225586 504791 225589
rect 505185 225586 505251 225589
rect 440969 225584 489930 225586
rect 440969 225528 440974 225584
rect 441030 225528 489930 225584
rect 440969 225526 489930 225528
rect 440969 225523 441035 225526
rect 147765 225450 147831 225453
rect 157149 225450 157215 225453
rect 147765 225448 157215 225450
rect 147765 225392 147770 225448
rect 147826 225392 157154 225448
rect 157210 225392 157215 225448
rect 147765 225390 157215 225392
rect 147765 225387 147831 225390
rect 157149 225387 157215 225390
rect 162669 225450 162735 225453
rect 169017 225450 169083 225453
rect 162669 225448 169083 225450
rect 162669 225392 162674 225448
rect 162730 225392 169022 225448
rect 169078 225392 169083 225448
rect 162669 225390 169083 225392
rect 162669 225387 162735 225390
rect 169017 225387 169083 225390
rect 186129 225450 186195 225453
rect 190269 225450 190335 225453
rect 186129 225448 190335 225450
rect 186129 225392 186134 225448
rect 186190 225392 190274 225448
rect 190330 225392 190335 225448
rect 186129 225390 190335 225392
rect 186129 225387 186195 225390
rect 190269 225387 190335 225390
rect 489870 225314 489930 225526
rect 504725 225584 505251 225586
rect 504725 225528 504730 225584
rect 504786 225528 505190 225584
rect 505246 225528 505251 225584
rect 504725 225526 505251 225528
rect 504725 225523 504791 225526
rect 505185 225523 505251 225526
rect 493869 225314 493935 225317
rect 613285 225314 613351 225317
rect 489870 225312 613351 225314
rect 489870 225256 493874 225312
rect 493930 225256 613290 225312
rect 613346 225256 613351 225312
rect 489870 225254 613351 225256
rect 493869 225251 493935 225254
rect 613285 225251 613351 225254
rect 43621 225042 43687 225045
rect 669129 225042 669195 225045
rect 43621 225040 669195 225042
rect 43621 224984 43626 225040
rect 43682 224984 669134 225040
rect 669190 224984 669195 225040
rect 43621 224982 669195 224984
rect 43621 224979 43687 224982
rect 669129 224979 669195 224982
rect 203885 224770 203951 224773
rect 204989 224770 205055 224773
rect 203885 224768 205055 224770
rect 203885 224712 203890 224768
rect 203946 224712 204994 224768
rect 205050 224712 205055 224768
rect 203885 224710 205055 224712
rect 203885 224707 203951 224710
rect 204989 224707 205055 224710
rect 483657 224770 483723 224773
rect 486233 224770 486299 224773
rect 483657 224768 486299 224770
rect 483657 224712 483662 224768
rect 483718 224712 486238 224768
rect 486294 224712 486299 224768
rect 483657 224710 486299 224712
rect 483657 224707 483723 224710
rect 486233 224707 486299 224710
rect 142153 224498 142219 224501
rect 149053 224498 149119 224501
rect 142153 224496 149119 224498
rect 142153 224440 142158 224496
rect 142214 224440 149058 224496
rect 149114 224440 149119 224496
rect 142153 224438 149119 224440
rect 142153 224435 142219 224438
rect 149053 224435 149119 224438
rect 484853 224498 484919 224501
rect 485865 224498 485931 224501
rect 484853 224496 485931 224498
rect 484853 224440 484858 224496
rect 484914 224440 485870 224496
rect 485926 224440 485931 224496
rect 484853 224438 485931 224440
rect 484853 224435 484919 224438
rect 485865 224435 485931 224438
rect 557349 224498 557415 224501
rect 558545 224498 558611 224501
rect 557349 224496 558611 224498
rect 557349 224440 557354 224496
rect 557410 224440 558550 224496
rect 558606 224440 558611 224496
rect 557349 224438 558611 224440
rect 557349 224435 557415 224438
rect 558545 224435 558611 224438
rect 172237 224362 172303 224365
rect 176377 224362 176443 224365
rect 172237 224360 176443 224362
rect 172237 224304 172242 224360
rect 172298 224304 176382 224360
rect 176438 224304 176443 224360
rect 172237 224302 176443 224304
rect 172237 224299 172303 224302
rect 176377 224299 176443 224302
rect 140681 224226 140747 224229
rect 142245 224226 142311 224229
rect 140681 224224 142311 224226
rect 140681 224168 140686 224224
rect 140742 224168 142250 224224
rect 142306 224168 142311 224224
rect 140681 224166 142311 224168
rect 140681 224163 140747 224166
rect 142245 224163 142311 224166
rect 146661 224226 146727 224229
rect 150801 224226 150867 224229
rect 146661 224224 150867 224226
rect 146661 224168 146666 224224
rect 146722 224168 150806 224224
rect 150862 224168 150867 224224
rect 146661 224166 150867 224168
rect 146661 224163 146727 224166
rect 150801 224163 150867 224166
rect 152273 224226 152339 224229
rect 159265 224226 159331 224229
rect 152273 224224 159331 224226
rect 152273 224168 152278 224224
rect 152334 224168 159270 224224
rect 159326 224168 159331 224224
rect 152273 224166 159331 224168
rect 152273 224163 152339 224166
rect 159265 224163 159331 224166
rect 481817 224226 481883 224229
rect 482645 224226 482711 224229
rect 611629 224226 611695 224229
rect 481817 224224 611695 224226
rect 481817 224168 481822 224224
rect 481878 224168 482650 224224
rect 482706 224168 611634 224224
rect 611690 224168 611695 224224
rect 481817 224166 611695 224168
rect 481817 224163 481883 224166
rect 482645 224163 482711 224166
rect 611629 224163 611695 224166
rect 50337 223954 50403 223957
rect 662413 223954 662479 223957
rect 50337 223952 662479 223954
rect 50337 223896 50342 223952
rect 50398 223896 662418 223952
rect 662474 223896 662479 223952
rect 50337 223894 662479 223896
rect 50337 223891 50403 223894
rect 662413 223891 662479 223894
rect 41689 223682 41755 223685
rect 668945 223682 669011 223685
rect 41689 223680 669011 223682
rect 41689 223624 41694 223680
rect 41750 223624 668950 223680
rect 669006 223624 669011 223680
rect 41689 223622 669011 223624
rect 41689 223619 41755 223622
rect 668945 223619 669011 223622
rect 675661 223546 675727 223549
rect 675661 223544 676292 223546
rect 675661 223488 675666 223544
rect 675722 223488 676292 223544
rect 675661 223486 676292 223488
rect 675661 223483 675727 223486
rect 160461 223410 160527 223413
rect 163773 223410 163839 223413
rect 160461 223408 163839 223410
rect 160461 223352 160466 223408
rect 160522 223352 163778 223408
rect 163834 223352 163839 223408
rect 160461 223350 163839 223352
rect 160461 223347 160527 223350
rect 163773 223347 163839 223350
rect 486785 223410 486851 223413
rect 498193 223410 498259 223413
rect 486785 223408 498259 223410
rect 486785 223352 486790 223408
rect 486846 223352 498198 223408
rect 498254 223352 498259 223408
rect 486785 223350 498259 223352
rect 486785 223347 486851 223350
rect 498193 223347 498259 223350
rect 555417 223410 555483 223413
rect 558545 223410 558611 223413
rect 555417 223408 558611 223410
rect 555417 223352 555422 223408
rect 555478 223352 558550 223408
rect 558606 223352 558611 223408
rect 555417 223350 558611 223352
rect 555417 223347 555483 223350
rect 558545 223347 558611 223350
rect 157425 223274 157491 223277
rect 152966 223272 157491 223274
rect 152966 223216 157430 223272
rect 157486 223216 157491 223272
rect 152966 223214 157491 223216
rect 71405 223138 71471 223141
rect 152966 223138 153026 223214
rect 157425 223211 157491 223214
rect 487061 223138 487127 223141
rect 71405 223136 153026 223138
rect 71405 223080 71410 223136
rect 71466 223080 153026 223136
rect 71405 223078 153026 223080
rect 483062 223136 487127 223138
rect 483062 223080 487066 223136
rect 487122 223080 487127 223136
rect 483062 223078 487127 223080
rect 71405 223075 71471 223078
rect 483062 223039 483122 223078
rect 487061 223075 487127 223078
rect 502517 223138 502583 223141
rect 614389 223138 614455 223141
rect 502517 223136 614455 223138
rect 502517 223080 502522 223136
rect 502578 223080 614394 223136
rect 614450 223080 614455 223136
rect 502517 223078 614455 223080
rect 502517 223075 502583 223078
rect 614389 223075 614455 223078
rect 675109 223138 675175 223141
rect 675109 223136 676292 223138
rect 675109 223080 675114 223136
rect 675170 223080 676292 223136
rect 675109 223078 676292 223080
rect 675109 223075 675175 223078
rect 483013 223034 483122 223039
rect 483013 222978 483018 223034
rect 483074 222978 483122 223034
rect 483013 222976 483122 222978
rect 483013 222973 483079 222976
rect 68737 222866 68803 222869
rect 155217 222866 155283 222869
rect 68737 222864 155283 222866
rect 68737 222808 68742 222864
rect 68798 222808 155222 222864
rect 155278 222808 155283 222864
rect 68737 222806 155283 222808
rect 68737 222803 68803 222806
rect 155217 222803 155283 222806
rect 156413 222866 156479 222869
rect 161105 222866 161171 222869
rect 156413 222864 161171 222866
rect 156413 222808 156418 222864
rect 156474 222808 161110 222864
rect 161166 222808 161171 222864
rect 156413 222806 161171 222808
rect 156413 222803 156479 222806
rect 161105 222803 161171 222806
rect 449525 222866 449591 222869
rect 510153 222866 510219 222869
rect 449525 222864 510219 222866
rect 449525 222808 449530 222864
rect 449586 222808 510158 222864
rect 510214 222808 510219 222864
rect 449525 222806 510219 222808
rect 449525 222803 449591 222806
rect 510153 222803 510219 222806
rect 548701 222866 548767 222869
rect 556337 222866 556403 222869
rect 548701 222864 556403 222866
rect 548701 222808 548706 222864
rect 548762 222808 556342 222864
rect 556398 222808 556403 222864
rect 548701 222806 556403 222808
rect 548701 222803 548767 222806
rect 556337 222803 556403 222806
rect 557993 222866 558059 222869
rect 559833 222866 559899 222869
rect 557993 222864 559899 222866
rect 557993 222808 557998 222864
rect 558054 222808 559838 222864
rect 559894 222808 559899 222864
rect 557993 222806 559899 222808
rect 557993 222803 558059 222806
rect 559833 222803 559899 222806
rect 675477 222730 675543 222733
rect 675477 222728 676292 222730
rect 675477 222672 675482 222728
rect 675538 222672 676292 222728
rect 675477 222670 676292 222672
rect 675477 222667 675543 222670
rect 40677 222594 40743 222597
rect 42609 222594 42675 222597
rect 40677 222592 42675 222594
rect 40677 222536 40682 222592
rect 40738 222536 42614 222592
rect 42670 222536 42675 222592
rect 40677 222534 42675 222536
rect 40677 222531 40743 222534
rect 42609 222531 42675 222534
rect 145925 222594 145991 222597
rect 147121 222594 147187 222597
rect 145925 222592 147187 222594
rect 145925 222536 145930 222592
rect 145986 222536 147126 222592
rect 147182 222536 147187 222592
rect 145925 222534 147187 222536
rect 145925 222531 145991 222534
rect 147121 222531 147187 222534
rect 151905 222594 151971 222597
rect 160921 222594 160987 222597
rect 151905 222592 160987 222594
rect 151905 222536 151910 222592
rect 151966 222536 160926 222592
rect 160982 222536 160987 222592
rect 151905 222534 160987 222536
rect 151905 222531 151971 222534
rect 160921 222531 160987 222534
rect 161565 222594 161631 222597
rect 164601 222594 164667 222597
rect 161565 222592 164667 222594
rect 161565 222536 161570 222592
rect 161626 222536 164606 222592
rect 164662 222536 164667 222592
rect 161565 222534 164667 222536
rect 161565 222531 161631 222534
rect 164601 222531 164667 222534
rect 484669 222594 484735 222597
rect 486233 222594 486299 222597
rect 484669 222592 486299 222594
rect 484669 222536 484674 222592
rect 484730 222536 486238 222592
rect 486294 222536 486299 222592
rect 484669 222534 486299 222536
rect 484669 222531 484735 222534
rect 486233 222531 486299 222534
rect 518893 222594 518959 222597
rect 618529 222594 618595 222597
rect 518893 222592 618595 222594
rect 518893 222536 518898 222592
rect 518954 222536 618534 222592
rect 618590 222536 618595 222592
rect 518893 222534 618595 222536
rect 518893 222531 518959 222534
rect 618529 222531 618595 222534
rect 28533 222322 28599 222325
rect 666737 222322 666803 222325
rect 28533 222320 666803 222322
rect 28533 222264 28538 222320
rect 28594 222264 666742 222320
rect 666798 222264 666803 222320
rect 28533 222262 666803 222264
rect 28533 222259 28599 222262
rect 666737 222259 666803 222262
rect 675293 222322 675359 222325
rect 675293 222320 676292 222322
rect 675293 222264 675298 222320
rect 675354 222264 676292 222320
rect 675293 222262 676292 222264
rect 675293 222259 675359 222262
rect 131757 222050 131823 222053
rect 661493 222050 661559 222053
rect 131757 222048 661559 222050
rect 131757 221992 131762 222048
rect 131818 221992 661498 222048
rect 661554 221992 661559 222048
rect 131757 221990 661559 221992
rect 131757 221987 131823 221990
rect 661493 221987 661559 221990
rect 675293 221914 675359 221917
rect 675293 221912 676292 221914
rect 675293 221856 675298 221912
rect 675354 221856 676292 221912
rect 675293 221854 676292 221856
rect 675293 221851 675359 221854
rect 128997 221778 129063 221781
rect 662597 221778 662663 221781
rect 128997 221776 662663 221778
rect 128997 221720 129002 221776
rect 129058 221720 662602 221776
rect 662658 221720 662663 221776
rect 128997 221718 662663 221720
rect 128997 221715 129063 221718
rect 662597 221715 662663 221718
rect 47577 221642 47643 221645
rect 47577 221640 64890 221642
rect 47577 221584 47582 221640
rect 47638 221584 64890 221640
rect 47577 221582 64890 221584
rect 47577 221579 47643 221582
rect 64830 221506 64890 221582
rect 663793 221506 663859 221509
rect 64830 221504 663859 221506
rect 64830 221448 663798 221504
rect 663854 221448 663859 221504
rect 64830 221446 663859 221448
rect 663793 221443 663859 221446
rect 675477 221506 675543 221509
rect 675477 221504 676292 221506
rect 675477 221448 675482 221504
rect 675538 221448 676292 221504
rect 675477 221446 676292 221448
rect 675477 221443 675543 221446
rect 147029 221234 147095 221237
rect 148317 221234 148383 221237
rect 147029 221232 148383 221234
rect 147029 221176 147034 221232
rect 147090 221176 148322 221232
rect 148378 221176 148383 221232
rect 147029 221174 148383 221176
rect 147029 221171 147095 221174
rect 148317 221171 148383 221174
rect 150709 221234 150775 221237
rect 152273 221234 152339 221237
rect 150709 221232 152339 221234
rect 150709 221176 150714 221232
rect 150770 221176 152278 221232
rect 152334 221176 152339 221232
rect 150709 221174 152339 221176
rect 150709 221171 150775 221174
rect 152273 221171 152339 221174
rect 161381 221234 161447 221237
rect 161565 221234 161631 221237
rect 161381 221232 161631 221234
rect 161381 221176 161386 221232
rect 161442 221176 161570 221232
rect 161626 221176 161631 221232
rect 161381 221174 161631 221176
rect 161381 221171 161447 221174
rect 161565 221171 161631 221174
rect 525977 221234 526043 221237
rect 529749 221234 529815 221237
rect 525977 221232 529815 221234
rect 525977 221176 525982 221232
rect 526038 221176 529754 221232
rect 529810 221176 529815 221232
rect 525977 221174 529815 221176
rect 525977 221171 526043 221174
rect 529749 221171 529815 221174
rect 533521 221234 533587 221237
rect 536649 221234 536715 221237
rect 533521 221232 536715 221234
rect 533521 221176 533526 221232
rect 533582 221176 536654 221232
rect 536710 221176 536715 221232
rect 533521 221174 536715 221176
rect 533521 221171 533587 221174
rect 536649 221171 536715 221174
rect 553485 221234 553551 221237
rect 554865 221234 554931 221237
rect 553485 221232 554931 221234
rect 553485 221176 553490 221232
rect 553546 221176 554870 221232
rect 554926 221176 554931 221232
rect 553485 221174 554931 221176
rect 553485 221171 553551 221174
rect 554865 221171 554931 221174
rect 592033 221234 592099 221237
rect 594149 221234 594215 221237
rect 592033 221232 594215 221234
rect 592033 221176 592038 221232
rect 592094 221176 594154 221232
rect 594210 221176 594215 221232
rect 592033 221174 594215 221176
rect 592033 221171 592099 221174
rect 594149 221171 594215 221174
rect 543549 221098 543615 221101
rect 550817 221098 550883 221101
rect 553301 221098 553367 221101
rect 543549 221096 553367 221098
rect 543549 221040 543554 221096
rect 543610 221040 550822 221096
rect 550878 221040 553306 221096
rect 553362 221040 553367 221096
rect 543549 221038 553367 221040
rect 543549 221035 543615 221038
rect 550817 221035 550883 221038
rect 553301 221035 553367 221038
rect 675477 221098 675543 221101
rect 675477 221096 676292 221098
rect 675477 221040 675482 221096
rect 675538 221040 676292 221096
rect 675477 221038 676292 221040
rect 675477 221035 675543 221038
rect 525057 220962 525123 220965
rect 533981 220962 534047 220965
rect 525057 220960 534047 220962
rect 525057 220904 525062 220960
rect 525118 220904 533986 220960
rect 534042 220904 534047 220960
rect 525057 220902 534047 220904
rect 525057 220899 525123 220902
rect 533981 220899 534047 220902
rect 562777 220962 562843 220965
rect 562777 220960 566290 220962
rect 562777 220904 562782 220960
rect 562838 220904 566290 220960
rect 562777 220902 566290 220904
rect 562777 220899 562843 220902
rect 538397 220826 538463 220829
rect 545205 220826 545271 220829
rect 538397 220824 545271 220826
rect 538397 220768 538402 220824
rect 538458 220768 545210 220824
rect 545266 220768 545271 220824
rect 538397 220766 545271 220768
rect 566230 220826 566290 220902
rect 567285 220826 567351 220829
rect 566230 220824 567351 220826
rect 566230 220768 567290 220824
rect 567346 220768 567351 220824
rect 566230 220766 567351 220768
rect 538397 220763 538463 220766
rect 545205 220763 545271 220766
rect 567285 220763 567351 220766
rect 553117 220690 553183 220693
rect 562961 220690 563027 220693
rect 553117 220688 553226 220690
rect 553117 220632 553122 220688
rect 553178 220632 553226 220688
rect 553117 220627 553226 220632
rect 543365 220554 543431 220557
rect 545757 220554 545823 220557
rect 543365 220552 545823 220554
rect 543365 220496 543370 220552
rect 543426 220496 545762 220552
rect 545818 220496 545823 220552
rect 543365 220494 545823 220496
rect 553166 220554 553226 220627
rect 562918 220688 563027 220690
rect 562918 220632 562966 220688
rect 563022 220632 563027 220688
rect 562918 220627 563027 220632
rect 675293 220690 675359 220693
rect 675293 220688 676292 220690
rect 675293 220632 675298 220688
rect 675354 220632 676292 220688
rect 675293 220630 676292 220632
rect 675293 220627 675359 220630
rect 553485 220554 553551 220557
rect 553166 220552 553551 220554
rect 553166 220496 553490 220552
rect 553546 220496 553551 220552
rect 553166 220494 553551 220496
rect 543365 220491 543431 220494
rect 545757 220491 545823 220494
rect 553485 220491 553551 220494
rect 553669 220554 553735 220557
rect 560661 220554 560727 220557
rect 562918 220554 562978 220627
rect 553669 220552 562978 220554
rect 553669 220496 553674 220552
rect 553730 220496 560666 220552
rect 560722 220496 562978 220552
rect 553669 220494 562978 220496
rect 564617 220554 564683 220557
rect 565353 220554 565419 220557
rect 564617 220552 565419 220554
rect 564617 220496 564622 220552
rect 564678 220496 565358 220552
rect 565414 220496 565419 220552
rect 564617 220494 565419 220496
rect 553669 220491 553735 220494
rect 560661 220491 560727 220494
rect 564617 220491 564683 220494
rect 565353 220491 565419 220494
rect 572529 220554 572595 220557
rect 574921 220554 574987 220557
rect 572529 220552 574987 220554
rect 572529 220496 572534 220552
rect 572590 220496 574926 220552
rect 574982 220496 574987 220552
rect 572529 220494 574987 220496
rect 572529 220491 572595 220494
rect 574921 220491 574987 220494
rect 144729 220418 144795 220421
rect 149237 220418 149303 220421
rect 144729 220416 149303 220418
rect 144729 220360 144734 220416
rect 144790 220360 149242 220416
rect 149298 220360 149303 220416
rect 144729 220358 149303 220360
rect 144729 220355 144795 220358
rect 149237 220355 149303 220358
rect 153929 220418 153995 220421
rect 156229 220418 156295 220421
rect 153929 220416 156295 220418
rect 153929 220360 153934 220416
rect 153990 220360 156234 220416
rect 156290 220360 156295 220416
rect 153929 220358 156295 220360
rect 153929 220355 153995 220358
rect 156229 220355 156295 220358
rect 524321 220282 524387 220285
rect 596265 220282 596331 220285
rect 524321 220280 596331 220282
rect 524321 220224 524326 220280
rect 524382 220224 596270 220280
rect 596326 220224 596331 220280
rect 524321 220222 596331 220224
rect 524321 220219 524387 220222
rect 596265 220219 596331 220222
rect 674649 220282 674715 220285
rect 674649 220280 676292 220282
rect 674649 220224 674654 220280
rect 674710 220224 676292 220280
rect 674649 220222 676292 220224
rect 674649 220219 674715 220222
rect 73061 220146 73127 220149
rect 158805 220146 158871 220149
rect 73061 220144 158871 220146
rect 73061 220088 73066 220144
rect 73122 220088 158810 220144
rect 158866 220088 158871 220144
rect 73061 220086 158871 220088
rect 73061 220083 73127 220086
rect 158805 220083 158871 220086
rect 483289 220146 483355 220149
rect 485865 220146 485931 220149
rect 483289 220144 485931 220146
rect 483289 220088 483294 220144
rect 483350 220088 485870 220144
rect 485926 220088 485931 220144
rect 483289 220086 485931 220088
rect 483289 220083 483355 220086
rect 485865 220083 485931 220086
rect 50981 220010 51047 220013
rect 164417 220010 164483 220013
rect 168557 220010 168623 220013
rect 50981 220008 54034 220010
rect 50981 219952 50986 220008
rect 51042 219952 54034 220008
rect 50981 219950 54034 219952
rect 50981 219947 51047 219950
rect 53974 219466 54034 219950
rect 164417 220008 168623 220010
rect 164417 219952 164422 220008
rect 164478 219952 168562 220008
rect 168618 219952 168623 220008
rect 164417 219950 168623 219952
rect 164417 219947 164483 219950
rect 168557 219947 168623 219950
rect 503529 220010 503595 220013
rect 598013 220010 598079 220013
rect 503529 220008 598079 220010
rect 503529 219952 503534 220008
rect 503590 219952 598018 220008
rect 598074 219952 598079 220008
rect 503529 219950 598079 219952
rect 503529 219947 503595 219950
rect 598013 219947 598079 219950
rect 675477 219874 675543 219877
rect 675477 219872 676292 219874
rect 675477 219816 675482 219872
rect 675538 219816 676292 219872
rect 675477 219814 676292 219816
rect 675477 219811 675543 219814
rect 54201 219738 54267 219741
rect 663977 219738 664043 219741
rect 54201 219736 664043 219738
rect 54201 219680 54206 219736
rect 54262 219680 663982 219736
rect 664038 219680 664043 219736
rect 54201 219678 664043 219680
rect 54201 219675 54267 219678
rect 663977 219675 664043 219678
rect 668393 219466 668459 219469
rect 53974 219464 668459 219466
rect 53974 219408 668398 219464
rect 668454 219408 668459 219464
rect 53974 219406 668459 219408
rect 668393 219403 668459 219406
rect 675477 219466 675543 219469
rect 675477 219464 676292 219466
rect 675477 219408 675482 219464
rect 675538 219408 676292 219464
rect 675477 219406 676292 219408
rect 675477 219403 675543 219406
rect 126421 219194 126487 219197
rect 128629 219194 128695 219197
rect 126421 219192 128695 219194
rect 126421 219136 126426 219192
rect 126482 219136 128634 219192
rect 128690 219136 128695 219192
rect 126421 219134 128695 219136
rect 126421 219131 126487 219134
rect 128629 219131 128695 219134
rect 137921 219194 137987 219197
rect 138473 219194 138539 219197
rect 137921 219192 138539 219194
rect 137921 219136 137926 219192
rect 137982 219136 138478 219192
rect 138534 219136 138539 219192
rect 137921 219134 138539 219136
rect 137921 219131 137987 219134
rect 138473 219131 138539 219134
rect 142245 219194 142311 219197
rect 144729 219194 144795 219197
rect 142245 219192 144795 219194
rect 142245 219136 142250 219192
rect 142306 219136 144734 219192
rect 144790 219136 144795 219192
rect 142245 219134 144795 219136
rect 142245 219131 142311 219134
rect 144729 219131 144795 219134
rect 156597 219194 156663 219197
rect 163221 219194 163287 219197
rect 156597 219192 163287 219194
rect 156597 219136 156602 219192
rect 156658 219136 163226 219192
rect 163282 219136 163287 219192
rect 156597 219134 163287 219136
rect 156597 219131 156663 219134
rect 163221 219131 163287 219134
rect 183185 219194 183251 219197
rect 189901 219194 189967 219197
rect 183185 219192 189967 219194
rect 183185 219136 183190 219192
rect 183246 219136 189906 219192
rect 189962 219136 189967 219192
rect 183185 219134 189967 219136
rect 183185 219131 183251 219134
rect 189901 219131 189967 219134
rect 489545 219194 489611 219197
rect 494421 219194 494487 219197
rect 489545 219192 494487 219194
rect 489545 219136 489550 219192
rect 489606 219136 494426 219192
rect 494482 219136 494487 219192
rect 489545 219134 494487 219136
rect 489545 219131 489611 219134
rect 494421 219131 494487 219134
rect 567469 219194 567535 219197
rect 572529 219194 572595 219197
rect 574185 219196 574251 219197
rect 574134 219194 574140 219196
rect 567469 219192 572595 219194
rect 567469 219136 567474 219192
rect 567530 219136 572534 219192
rect 572590 219136 572595 219192
rect 567469 219134 572595 219136
rect 574094 219134 574140 219194
rect 574204 219192 574251 219196
rect 574246 219136 574251 219192
rect 567469 219131 567535 219134
rect 572529 219131 572595 219134
rect 574134 219132 574140 219134
rect 574204 219132 574251 219136
rect 574502 219132 574508 219196
rect 574572 219194 574578 219196
rect 575105 219194 575171 219197
rect 574572 219192 575171 219194
rect 574572 219136 575110 219192
rect 575166 219136 575171 219192
rect 574572 219134 575171 219136
rect 574572 219132 574578 219134
rect 574185 219131 574251 219132
rect 575105 219131 575171 219134
rect 499573 219060 499639 219061
rect 499573 219056 499620 219060
rect 499684 219058 499690 219060
rect 500217 219058 500283 219061
rect 499684 219056 500283 219058
rect 499573 219000 499578 219056
rect 499684 219000 500222 219056
rect 500278 219000 500283 219056
rect 499573 218996 499620 219000
rect 499684 218998 500283 219000
rect 499684 218996 499690 218998
rect 499573 218995 499639 218996
rect 500217 218995 500283 218998
rect 675569 219058 675635 219061
rect 675569 219056 676292 219058
rect 675569 219000 675574 219056
rect 675630 219000 676292 219056
rect 675569 218998 676292 219000
rect 675569 218995 675635 218998
rect 130193 218922 130259 218925
rect 184197 218922 184263 218925
rect 130193 218920 184263 218922
rect 130193 218864 130198 218920
rect 130254 218864 184202 218920
rect 184258 218864 184263 218920
rect 130193 218862 184263 218864
rect 130193 218859 130259 218862
rect 184197 218859 184263 218862
rect 442441 218922 442507 218925
rect 512729 218922 512795 218925
rect 616873 218922 616939 218925
rect 442441 218920 485146 218922
rect 442441 218864 442446 218920
rect 442502 218864 485146 218920
rect 442441 218862 485146 218864
rect 442441 218859 442507 218862
rect 202873 218786 202939 218789
rect 205495 218786 205561 218789
rect 202873 218784 205561 218786
rect 202873 218728 202878 218784
rect 202934 218728 205500 218784
rect 205556 218728 205561 218784
rect 202873 218726 205561 218728
rect 485086 218786 485146 218862
rect 512729 218920 616939 218922
rect 512729 218864 512734 218920
rect 512790 218864 616878 218920
rect 616934 218864 616939 218920
rect 512729 218862 616939 218864
rect 512729 218859 512795 218862
rect 616873 218859 616939 218862
rect 487889 218786 487955 218789
rect 485086 218784 487955 218786
rect 485086 218728 487894 218784
rect 487950 218728 487955 218784
rect 485086 218726 487955 218728
rect 202873 218723 202939 218726
rect 205495 218723 205561 218726
rect 487889 218723 487955 218726
rect 77201 218650 77267 218653
rect 156597 218650 156663 218653
rect 77201 218648 156663 218650
rect 77201 218592 77206 218648
rect 77262 218592 156602 218648
rect 156658 218592 156663 218648
rect 77201 218590 156663 218592
rect 77201 218587 77267 218590
rect 156597 218587 156663 218590
rect 191925 218650 191991 218653
rect 196617 218650 196683 218653
rect 191925 218648 196683 218650
rect 191925 218592 191930 218648
rect 191986 218592 196622 218648
rect 196678 218592 196683 218648
rect 191925 218590 196683 218592
rect 191925 218587 191991 218590
rect 196617 218587 196683 218590
rect 435357 218650 435423 218653
rect 484577 218650 484643 218653
rect 435357 218648 484643 218650
rect 435357 218592 435362 218648
rect 435418 218592 484582 218648
rect 484638 218592 484643 218648
rect 435357 218590 484643 218592
rect 435357 218587 435423 218590
rect 484577 218587 484643 218590
rect 505737 218650 505803 218653
rect 508313 218650 508379 218653
rect 505737 218648 508379 218650
rect 505737 218592 505742 218648
rect 505798 218592 508318 218648
rect 508374 218592 508379 218648
rect 505737 218590 508379 218592
rect 505737 218587 505803 218590
rect 508313 218587 508379 218590
rect 510153 218650 510219 218653
rect 616137 218650 616203 218653
rect 510153 218648 616203 218650
rect 510153 218592 510158 218648
rect 510214 218592 616142 218648
rect 616198 218592 616203 218648
rect 510153 218590 616203 218592
rect 510153 218587 510219 218590
rect 616137 218587 616203 218590
rect 675518 218588 675524 218652
rect 675588 218650 675594 218652
rect 675588 218590 676292 218650
rect 675588 218588 675594 218590
rect 161289 218514 161355 218517
rect 161749 218514 161815 218517
rect 161289 218512 161815 218514
rect 161289 218456 161294 218512
rect 161350 218456 161754 218512
rect 161810 218456 161815 218512
rect 161289 218454 161815 218456
rect 161289 218451 161355 218454
rect 161749 218451 161815 218454
rect 183553 218514 183619 218517
rect 185301 218514 185367 218517
rect 183553 218512 185367 218514
rect 183553 218456 183558 218512
rect 183614 218456 185306 218512
rect 185362 218456 185367 218512
rect 183553 218454 185367 218456
rect 183553 218451 183619 218454
rect 185301 218451 185367 218454
rect 205449 218514 205515 218517
rect 205633 218514 205699 218517
rect 205449 218512 205699 218514
rect 205449 218456 205454 218512
rect 205510 218456 205638 218512
rect 205694 218456 205699 218512
rect 205449 218454 205699 218456
rect 205449 218451 205515 218454
rect 205633 218451 205699 218454
rect 487613 218514 487679 218517
rect 491109 218514 491175 218517
rect 487613 218512 491175 218514
rect 487613 218456 487618 218512
rect 487674 218456 491114 218512
rect 491170 218456 491175 218512
rect 487613 218454 491175 218456
rect 487613 218451 487679 218454
rect 491109 218451 491175 218454
rect 39757 218378 39823 218381
rect 43437 218378 43503 218381
rect 39757 218376 43503 218378
rect 39757 218320 39762 218376
rect 39818 218320 43442 218376
rect 43498 218320 43503 218376
rect 39757 218318 43503 218320
rect 39757 218315 39823 218318
rect 43437 218315 43503 218318
rect 150065 218378 150131 218381
rect 151905 218378 151971 218381
rect 150065 218376 151971 218378
rect 150065 218320 150070 218376
rect 150126 218320 151910 218376
rect 151966 218320 151971 218376
rect 150065 218318 151971 218320
rect 150065 218315 150131 218318
rect 151905 218315 151971 218318
rect 478781 218378 478847 218381
rect 482185 218378 482251 218381
rect 609605 218378 609671 218381
rect 478781 218376 482251 218378
rect 478781 218320 478786 218376
rect 478842 218320 482190 218376
rect 482246 218320 482251 218376
rect 478781 218318 482251 218320
rect 478781 218315 478847 218318
rect 482185 218315 482251 218318
rect 508086 218376 609671 218378
rect 508086 218320 609610 218376
rect 609666 218320 609671 218376
rect 508086 218318 609671 218320
rect 152549 218242 152615 218245
rect 161289 218242 161355 218245
rect 152549 218240 161355 218242
rect 152549 218184 152554 218240
rect 152610 218184 161294 218240
rect 161350 218184 161355 218240
rect 152549 218182 161355 218184
rect 152549 218179 152615 218182
rect 161289 218179 161355 218182
rect 161473 218242 161539 218245
rect 167545 218242 167611 218245
rect 161473 218240 167611 218242
rect 161473 218184 161478 218240
rect 161534 218184 167550 218240
rect 167606 218184 167611 218240
rect 161473 218182 167611 218184
rect 161473 218179 161539 218182
rect 167545 218179 167611 218182
rect 215201 218242 215267 218245
rect 217317 218242 217383 218245
rect 215201 218240 217383 218242
rect 215201 218184 215206 218240
rect 215262 218184 217322 218240
rect 217378 218184 217383 218240
rect 215201 218182 217383 218184
rect 215201 218179 215267 218182
rect 217317 218179 217383 218182
rect 490557 218242 490623 218245
rect 491293 218242 491359 218245
rect 490557 218240 491359 218242
rect 490557 218184 490562 218240
rect 490618 218184 491298 218240
rect 491354 218184 491359 218240
rect 490557 218182 491359 218184
rect 490557 218179 490623 218182
rect 491293 218179 491359 218182
rect 40217 218106 40283 218109
rect 47945 218106 48011 218109
rect 40217 218104 48011 218106
rect 40217 218048 40222 218104
rect 40278 218048 47950 218104
rect 48006 218048 48011 218104
rect 40217 218046 48011 218048
rect 40217 218043 40283 218046
rect 47945 218043 48011 218046
rect 143441 218106 143507 218109
rect 151445 218106 151511 218109
rect 143441 218104 151511 218106
rect 143441 218048 143446 218104
rect 143502 218048 151450 218104
rect 151506 218048 151511 218104
rect 143441 218046 151511 218048
rect 143441 218043 143507 218046
rect 151445 218043 151511 218046
rect 484577 218106 484643 218109
rect 489821 218106 489887 218109
rect 490373 218108 490439 218109
rect 490373 218106 490420 218108
rect 484577 218104 489887 218106
rect 484577 218048 484582 218104
rect 484638 218048 489826 218104
rect 489882 218048 489887 218104
rect 484577 218046 489887 218048
rect 490328 218104 490420 218106
rect 490328 218048 490378 218104
rect 490328 218046 490420 218048
rect 484577 218043 484643 218046
rect 489821 218043 489887 218046
rect 490373 218044 490420 218046
rect 490484 218044 490490 218108
rect 507117 218106 507183 218109
rect 507669 218106 507735 218109
rect 508086 218106 508146 218318
rect 609605 218315 609671 218318
rect 675753 218242 675819 218245
rect 675753 218240 676292 218242
rect 675753 218184 675758 218240
rect 675814 218184 676292 218240
rect 675753 218182 676292 218184
rect 675753 218179 675819 218182
rect 507117 218104 508146 218106
rect 507117 218048 507122 218104
rect 507178 218048 507674 218104
rect 507730 218048 508146 218104
rect 507117 218046 508146 218048
rect 508313 218106 508379 218109
rect 615033 218106 615099 218109
rect 508313 218104 615099 218106
rect 508313 218048 508318 218104
rect 508374 218048 615038 218104
rect 615094 218048 615099 218104
rect 508313 218046 615099 218048
rect 490373 218043 490439 218044
rect 507117 218043 507183 218046
rect 507669 218043 507735 218046
rect 508313 218043 508379 218046
rect 615033 218043 615099 218046
rect 493685 217972 493751 217973
rect 493685 217970 493732 217972
rect 493640 217968 493732 217970
rect 493640 217912 493690 217968
rect 493640 217910 493732 217912
rect 493685 217908 493732 217910
rect 493796 217908 493802 217972
rect 669446 217908 669452 217972
rect 669516 217970 669522 217972
rect 670601 217970 670667 217973
rect 669516 217968 670667 217970
rect 669516 217912 670606 217968
rect 670662 217912 670667 217968
rect 669516 217910 670667 217912
rect 669516 217908 669522 217910
rect 493685 217907 493751 217908
rect 670601 217907 670667 217910
rect 564801 217834 564867 217837
rect 566038 217834 566044 217836
rect 564801 217832 566044 217834
rect 564801 217776 564806 217832
rect 564862 217776 566044 217832
rect 564801 217774 566044 217776
rect 564801 217771 564867 217774
rect 566038 217772 566044 217774
rect 566108 217772 566114 217836
rect 567285 217834 567351 217837
rect 574277 217834 574343 217837
rect 567285 217832 574343 217834
rect 567285 217776 567290 217832
rect 567346 217776 574282 217832
rect 574338 217776 574343 217832
rect 567285 217774 574343 217776
rect 567285 217771 567351 217774
rect 574277 217771 574343 217774
rect 675201 217834 675267 217837
rect 675201 217832 676292 217834
rect 675201 217776 675206 217832
rect 675262 217776 676292 217832
rect 675201 217774 676292 217776
rect 675201 217771 675267 217774
rect 501229 217564 501295 217565
rect 501229 217562 501276 217564
rect 501184 217560 501276 217562
rect 501184 217504 501234 217560
rect 501184 217502 501276 217504
rect 501229 217500 501276 217502
rect 501340 217500 501346 217564
rect 503345 217562 503411 217565
rect 595161 217562 595227 217565
rect 503345 217560 595227 217562
rect 503345 217504 503350 217560
rect 503406 217504 595166 217560
rect 595222 217504 595227 217560
rect 503345 217502 595227 217504
rect 501229 217499 501295 217500
rect 503345 217499 503411 217502
rect 595161 217499 595227 217502
rect 601509 217562 601575 217565
rect 603441 217562 603507 217565
rect 601509 217560 603507 217562
rect 601509 217504 601514 217560
rect 601570 217504 603446 217560
rect 603502 217504 603507 217560
rect 601509 217502 603507 217504
rect 601509 217499 601575 217502
rect 603441 217499 603507 217502
rect 675702 217364 675708 217428
rect 675772 217426 675778 217428
rect 675772 217366 676292 217426
rect 675772 217364 675778 217366
rect 491109 217292 491175 217293
rect 491109 217288 491156 217292
rect 491220 217290 491226 217292
rect 495249 217290 495315 217293
rect 595713 217290 595779 217293
rect 491109 217232 491114 217288
rect 491109 217228 491156 217232
rect 491220 217230 491266 217290
rect 495249 217288 595779 217290
rect 495249 217232 495254 217288
rect 495310 217232 595718 217288
rect 595774 217232 595779 217288
rect 495249 217230 595779 217232
rect 491220 217228 491226 217230
rect 491109 217227 491175 217228
rect 495249 217227 495315 217230
rect 595713 217227 595779 217230
rect 601325 217290 601391 217293
rect 603073 217290 603139 217293
rect 601325 217288 603139 217290
rect 601325 217232 601330 217288
rect 601386 217232 603078 217288
rect 603134 217232 603139 217288
rect 601325 217230 603139 217232
rect 601325 217227 601391 217230
rect 603073 217227 603139 217230
rect 491385 217154 491451 217157
rect 491385 217152 492690 217154
rect 491385 217096 491390 217152
rect 491446 217096 492690 217152
rect 491385 217094 492690 217096
rect 491385 217091 491451 217094
rect 492630 217018 492690 217094
rect 492630 216958 495450 217018
rect 495390 216746 495450 216958
rect 501270 216956 501276 217020
rect 501340 217018 501346 217020
rect 596817 217018 596883 217021
rect 501340 217016 596883 217018
rect 501340 216960 596822 217016
rect 596878 216960 596883 217016
rect 501340 216958 596883 216960
rect 501340 216956 501346 216958
rect 596817 216955 596883 216958
rect 675385 217018 675451 217021
rect 675385 217016 676292 217018
rect 675385 216960 675390 217016
rect 675446 216960 676292 217016
rect 675385 216958 676292 216960
rect 675385 216955 675451 216958
rect 575473 216746 575539 216749
rect 495390 216744 575539 216746
rect 495390 216688 575478 216744
rect 575534 216688 575539 216744
rect 495390 216686 575539 216688
rect 575473 216683 575539 216686
rect 575790 216684 575796 216748
rect 575860 216746 575866 216748
rect 612825 216746 612891 216749
rect 575860 216744 612891 216746
rect 575860 216688 612830 216744
rect 612886 216688 612891 216744
rect 575860 216686 612891 216688
rect 575860 216684 575866 216686
rect 612825 216683 612891 216686
rect 670969 216612 671035 216613
rect 670918 216610 670924 216612
rect 670878 216550 670924 216610
rect 670988 216608 671035 216612
rect 671030 216552 671035 216608
rect 670918 216548 670924 216550
rect 670988 216548 671035 216552
rect 675334 216548 675340 216612
rect 675404 216610 675410 216612
rect 675404 216550 676292 216610
rect 675404 216548 675410 216550
rect 670969 216547 671035 216548
rect 574369 216476 574435 216477
rect 574318 216474 574324 216476
rect 574278 216414 574324 216474
rect 574388 216472 574435 216476
rect 574430 216416 574435 216472
rect 574318 216412 574324 216414
rect 574388 216412 574435 216416
rect 574369 216411 574435 216412
rect 671102 216140 671108 216204
rect 671172 216202 671178 216204
rect 671889 216202 671955 216205
rect 671172 216200 671955 216202
rect 671172 216144 671894 216200
rect 671950 216144 671955 216200
rect 671172 216142 671955 216144
rect 671172 216140 671178 216142
rect 671889 216139 671955 216142
rect 675385 216202 675451 216205
rect 675385 216200 676292 216202
rect 675385 216144 675390 216200
rect 675446 216144 676292 216200
rect 675385 216142 676292 216144
rect 675385 216139 675451 216142
rect 566038 216004 566044 216068
rect 566108 216066 566114 216068
rect 574921 216066 574987 216069
rect 566108 216064 574987 216066
rect 566108 216008 574926 216064
rect 574982 216008 574987 216064
rect 566108 216006 574987 216008
rect 566108 216004 566114 216006
rect 574921 216003 574987 216006
rect 575982 215386 576042 215764
rect 676170 215734 676292 215794
rect 676170 215658 676230 215734
rect 672030 215598 676230 215658
rect 672030 215525 672090 215598
rect 671981 215520 672090 215525
rect 671981 215464 671986 215520
rect 672042 215464 672090 215520
rect 671981 215462 672090 215464
rect 671981 215459 672047 215462
rect 578877 215386 578943 215389
rect 575982 215384 578943 215386
rect 575982 215328 578882 215384
rect 578938 215328 578943 215384
rect 575982 215326 578943 215328
rect 578877 215323 578943 215326
rect 674465 215386 674531 215389
rect 674465 215384 676292 215386
rect 674465 215328 674470 215384
rect 674526 215328 676292 215384
rect 674465 215326 676292 215328
rect 674465 215323 674531 215326
rect 676029 214978 676095 214981
rect 676029 214976 676292 214978
rect 35390 214709 35450 214948
rect 676029 214920 676034 214976
rect 676090 214920 676292 214976
rect 676029 214918 676292 214920
rect 676029 214915 676095 214918
rect 35341 214704 35450 214709
rect 35341 214648 35346 214704
rect 35402 214648 35450 214704
rect 35341 214646 35450 214648
rect 35341 214643 35407 214646
rect 35758 214301 35818 214540
rect 675886 214508 675892 214572
rect 675956 214570 675962 214572
rect 675956 214510 676292 214570
rect 675956 214508 675962 214510
rect 35525 214298 35591 214301
rect 35525 214296 35634 214298
rect 35525 214240 35530 214296
rect 35586 214240 35634 214296
rect 35525 214235 35634 214240
rect 35758 214296 35867 214301
rect 35758 214240 35806 214296
rect 35862 214240 35867 214296
rect 35758 214238 35867 214240
rect 35801 214235 35867 214238
rect 39757 214298 39823 214301
rect 45553 214298 45619 214301
rect 39757 214296 45619 214298
rect 39757 214240 39762 214296
rect 39818 214240 45558 214296
rect 45614 214240 45619 214296
rect 39757 214238 45619 214240
rect 39757 214235 39823 214238
rect 45553 214235 45619 214238
rect 35574 214132 35634 214235
rect 674925 214162 674991 214165
rect 674925 214160 676292 214162
rect 674925 214104 674930 214160
rect 674986 214104 676292 214160
rect 674925 214102 676292 214104
rect 674925 214099 674991 214102
rect 673678 213964 673684 214028
rect 673748 214026 673754 214028
rect 673913 214026 673979 214029
rect 673748 214024 673979 214026
rect 673748 213968 673918 214024
rect 673974 213968 673979 214024
rect 673748 213966 673979 213968
rect 673748 213964 673754 213966
rect 673913 213963 673979 213966
rect 675477 213754 675543 213757
rect 675477 213752 676292 213754
rect 35758 213485 35818 213724
rect 675477 213696 675482 213752
rect 675538 213696 676292 213752
rect 675477 213694 676292 213696
rect 675477 213691 675543 213694
rect 35758 213480 35867 213485
rect 35758 213424 35806 213480
rect 35862 213424 35867 213480
rect 35758 213422 35867 213424
rect 35801 213419 35867 213422
rect 675477 213346 675543 213349
rect 675477 213344 676292 213346
rect 35574 213077 35634 213316
rect 35574 213072 35683 213077
rect 35574 213016 35622 213072
rect 35678 213016 35683 213072
rect 35574 213014 35683 213016
rect 35617 213011 35683 213014
rect 39297 213074 39363 213077
rect 44173 213074 44239 213077
rect 39297 213072 44239 213074
rect 39297 213016 39302 213072
rect 39358 213016 44178 213072
rect 44234 213016 44239 213072
rect 39297 213014 44239 213016
rect 39297 213011 39363 213014
rect 44173 213011 44239 213014
rect 575982 212938 576042 213316
rect 675477 213288 675482 213344
rect 675538 213288 676292 213344
rect 675477 213286 676292 213288
rect 675477 213283 675543 213286
rect 578325 212938 578391 212941
rect 575982 212936 578391 212938
rect 35758 212669 35818 212908
rect 575982 212880 578330 212936
rect 578386 212880 578391 212936
rect 575982 212878 578391 212880
rect 578325 212875 578391 212878
rect 28533 212666 28599 212669
rect 28533 212664 28642 212666
rect 28533 212608 28538 212664
rect 28594 212608 28642 212664
rect 28533 212603 28642 212608
rect 35758 212664 35867 212669
rect 35758 212608 35806 212664
rect 35862 212608 35867 212664
rect 35758 212606 35867 212608
rect 35801 212603 35867 212606
rect 41229 212666 41295 212669
rect 42149 212666 42215 212669
rect 41229 212664 42215 212666
rect 41229 212608 41234 212664
rect 41290 212608 42154 212664
rect 42210 212608 42215 212664
rect 41229 212606 42215 212608
rect 41229 212603 41295 212606
rect 42149 212603 42215 212606
rect 672533 212666 672599 212669
rect 672942 212666 672948 212668
rect 672533 212664 672948 212666
rect 672533 212608 672538 212664
rect 672594 212608 672948 212664
rect 672533 212606 672948 212608
rect 672533 212603 672599 212606
rect 672942 212604 672948 212606
rect 673012 212604 673018 212668
rect 28582 212500 28642 212603
rect 683070 212533 683130 212908
rect 683070 212528 683179 212533
rect 683070 212500 683118 212528
rect 683100 212472 683118 212500
rect 683174 212472 683179 212528
rect 683100 212470 683179 212472
rect 683113 212467 683179 212470
rect 675334 212332 675340 212396
rect 675404 212394 675410 212396
rect 675886 212394 675892 212396
rect 675404 212334 675892 212394
rect 675404 212332 675410 212334
rect 675886 212332 675892 212334
rect 675956 212332 675962 212396
rect 41045 212258 41111 212261
rect 43621 212258 43687 212261
rect 41045 212256 43687 212258
rect 41045 212200 41050 212256
rect 41106 212200 43626 212256
rect 43682 212200 43687 212256
rect 41045 212198 43687 212200
rect 41045 212195 41111 212198
rect 43621 212195 43687 212198
rect 675477 212122 675543 212125
rect 675477 212120 676292 212122
rect 35758 211853 35818 212092
rect 675477 212064 675482 212120
rect 675538 212064 676292 212120
rect 675477 212062 676292 212064
rect 675477 212059 675543 212062
rect 35758 211848 35867 211853
rect 35758 211792 35806 211848
rect 35862 211792 35867 211848
rect 35758 211790 35867 211792
rect 35801 211787 35867 211790
rect 41229 211850 41295 211853
rect 43805 211850 43871 211853
rect 41229 211848 43871 211850
rect 41229 211792 41234 211848
rect 41290 211792 43810 211848
rect 43866 211792 43871 211848
rect 41229 211790 43871 211792
rect 41229 211787 41295 211790
rect 43805 211787 43871 211790
rect 35574 211445 35634 211684
rect 35574 211440 35683 211445
rect 35574 211384 35622 211440
rect 35678 211384 35683 211440
rect 35574 211382 35683 211384
rect 35617 211379 35683 211382
rect 39665 211442 39731 211445
rect 42885 211442 42951 211445
rect 39665 211440 42951 211442
rect 39665 211384 39670 211440
rect 39726 211384 42890 211440
rect 42946 211384 42951 211440
rect 39665 211382 42951 211384
rect 39665 211379 39731 211382
rect 42885 211379 42951 211382
rect 676029 211442 676095 211445
rect 676438 211442 676444 211444
rect 676029 211440 676444 211442
rect 676029 211384 676034 211440
rect 676090 211384 676444 211440
rect 676029 211382 676444 211384
rect 676029 211379 676095 211382
rect 676438 211380 676444 211382
rect 676508 211380 676514 211444
rect 35758 211037 35818 211276
rect 665817 211170 665883 211173
rect 670785 211172 670851 211173
rect 667974 211170 667980 211172
rect 665817 211168 667980 211170
rect 665817 211112 665822 211168
rect 665878 211112 667980 211168
rect 665817 211110 667980 211112
rect 665817 211107 665883 211110
rect 667974 211108 667980 211110
rect 668044 211108 668050 211172
rect 669630 211170 669636 211172
rect 669270 211110 669636 211170
rect 35758 211032 35867 211037
rect 35758 210976 35806 211032
rect 35862 210976 35867 211032
rect 35758 210974 35867 210976
rect 35801 210971 35867 210974
rect 664437 210898 664503 210901
rect 669270 210898 669330 211110
rect 669630 211108 669636 211110
rect 669700 211108 669706 211172
rect 670734 211170 670740 211172
rect 670694 211110 670740 211170
rect 670804 211168 670851 211172
rect 670846 211112 670851 211168
rect 670734 211108 670740 211110
rect 670804 211108 670851 211112
rect 675886 211108 675892 211172
rect 675956 211170 675962 211172
rect 683113 211170 683179 211173
rect 675956 211168 683179 211170
rect 675956 211112 683118 211168
rect 683174 211112 683179 211168
rect 675956 211110 683179 211112
rect 675956 211108 675962 211110
rect 670785 211107 670851 211108
rect 683113 211107 683179 211110
rect 664437 210896 669330 210898
rect 35574 210629 35634 210868
rect 35574 210624 35683 210629
rect 35574 210568 35622 210624
rect 35678 210568 35683 210624
rect 35574 210566 35683 210568
rect 35617 210563 35683 210566
rect 35758 210221 35818 210460
rect 575982 210354 576042 210868
rect 664437 210840 664442 210896
rect 664498 210840 669330 210896
rect 664437 210838 669330 210840
rect 670785 210898 670851 210901
rect 671102 210898 671108 210900
rect 670785 210896 671108 210898
rect 670785 210840 670790 210896
rect 670846 210840 671108 210896
rect 670785 210838 671108 210840
rect 664437 210835 664503 210838
rect 670785 210835 670851 210838
rect 671102 210836 671108 210838
rect 671172 210836 671178 210900
rect 666686 210428 666692 210492
rect 666756 210490 666762 210492
rect 667054 210490 667060 210492
rect 666756 210430 667060 210490
rect 666756 210428 666762 210430
rect 667054 210428 667060 210430
rect 667124 210428 667130 210492
rect 672349 210490 672415 210493
rect 673126 210490 673132 210492
rect 672349 210488 673132 210490
rect 672349 210432 672354 210488
rect 672410 210432 673132 210488
rect 672349 210430 673132 210432
rect 672349 210427 672415 210430
rect 673126 210428 673132 210430
rect 673196 210428 673202 210492
rect 673494 210428 673500 210492
rect 673564 210490 673570 210492
rect 673729 210490 673795 210493
rect 673564 210488 673795 210490
rect 673564 210432 673734 210488
rect 673790 210432 673795 210488
rect 673564 210430 673795 210432
rect 673564 210428 673570 210430
rect 673729 210427 673795 210430
rect 675518 210428 675524 210492
rect 675588 210490 675594 210492
rect 676070 210490 676076 210492
rect 675588 210430 676076 210490
rect 675588 210428 675594 210430
rect 676070 210428 676076 210430
rect 676140 210428 676146 210492
rect 579521 210354 579587 210357
rect 575982 210352 579587 210354
rect 575982 210296 579526 210352
rect 579582 210296 579587 210352
rect 575982 210294 579587 210296
rect 579521 210291 579587 210294
rect 35758 210216 35867 210221
rect 35758 210160 35806 210216
rect 35862 210160 35867 210216
rect 35758 210158 35867 210160
rect 35801 210155 35867 210158
rect 41822 210082 41828 210084
rect 41492 210022 41828 210082
rect 41822 210020 41828 210022
rect 41892 210020 41898 210084
rect 35574 209405 35634 209644
rect 35574 209400 35683 209405
rect 35574 209344 35622 209400
rect 35678 209344 35683 209400
rect 35574 209342 35683 209344
rect 35617 209339 35683 209342
rect 672349 209266 672415 209269
rect 673310 209266 673316 209268
rect 672349 209264 673316 209266
rect 30238 208997 30298 209236
rect 672349 209208 672354 209264
rect 672410 209208 673316 209264
rect 672349 209206 673316 209208
rect 672349 209203 672415 209206
rect 673310 209204 673316 209206
rect 673380 209204 673386 209268
rect 30238 208992 30347 208997
rect 35801 208994 35867 208997
rect 30238 208936 30286 208992
rect 30342 208936 30347 208992
rect 30238 208934 30347 208936
rect 30281 208931 30347 208934
rect 35758 208992 35867 208994
rect 35758 208936 35806 208992
rect 35862 208936 35867 208992
rect 35758 208931 35867 208936
rect 35758 208828 35818 208931
rect 39665 208586 39731 208589
rect 43069 208586 43135 208589
rect 579521 208586 579587 208589
rect 39665 208584 43135 208586
rect 39665 208528 39670 208584
rect 39726 208528 43074 208584
rect 43130 208528 43135 208584
rect 39665 208526 43135 208528
rect 39665 208523 39731 208526
rect 43069 208523 43135 208526
rect 575798 208584 579587 208586
rect 575798 208528 579526 208584
rect 579582 208528 579587 208584
rect 575798 208526 579587 208528
rect 575798 208420 575858 208526
rect 579521 208523 579587 208526
rect 40910 208180 40970 208420
rect 589457 208314 589523 208317
rect 589457 208312 592602 208314
rect 589457 208256 589462 208312
rect 589518 208256 592602 208312
rect 589457 208254 592602 208256
rect 589457 208251 589523 208254
rect 40902 208116 40908 208180
rect 40972 208116 40978 208180
rect 592542 208080 592602 208254
rect 40542 207772 40602 208012
rect 40534 207708 40540 207772
rect 40604 207708 40610 207772
rect 35574 207365 35634 207604
rect 35525 207360 35634 207365
rect 35801 207362 35867 207365
rect 667974 207362 667980 207364
rect 35525 207304 35530 207360
rect 35586 207304 35634 207360
rect 35525 207302 35634 207304
rect 35758 207360 35867 207362
rect 35758 207304 35806 207360
rect 35862 207304 35867 207360
rect 35525 207299 35591 207302
rect 35758 207299 35867 207304
rect 666878 207302 667980 207362
rect 35758 207196 35818 207299
rect 666878 207294 666938 207302
rect 667974 207300 667980 207302
rect 668044 207300 668050 207364
rect 666356 207234 666938 207294
rect 39757 206954 39823 206957
rect 42885 206954 42951 206957
rect 39757 206952 42951 206954
rect 39757 206896 39762 206952
rect 39818 206896 42890 206952
rect 42946 206896 42951 206952
rect 39757 206894 42951 206896
rect 39757 206891 39823 206894
rect 42885 206891 42951 206894
rect 589549 206954 589615 206957
rect 589549 206952 592602 206954
rect 589549 206896 589554 206952
rect 589610 206896 592602 206952
rect 589549 206894 592602 206896
rect 589549 206891 589615 206894
rect 35574 206549 35634 206788
rect 35574 206544 35683 206549
rect 35574 206488 35622 206544
rect 35678 206488 35683 206544
rect 35574 206486 35683 206488
rect 35617 206483 35683 206486
rect 592542 206448 592602 206894
rect 35801 206138 35867 206141
rect 40726 206140 40786 206380
rect 35758 206136 35867 206138
rect 35758 206080 35806 206136
rect 35862 206080 35867 206136
rect 35758 206075 35867 206080
rect 40718 206076 40724 206140
rect 40788 206076 40794 206140
rect 35758 205972 35818 206075
rect 575982 205866 576042 205972
rect 579521 205866 579587 205869
rect 575982 205864 579587 205866
rect 575982 205808 579526 205864
rect 579582 205808 579587 205864
rect 575982 205806 579587 205808
rect 579521 205803 579587 205806
rect 40033 205730 40099 205733
rect 41454 205730 41460 205732
rect 40033 205728 41460 205730
rect 40033 205672 40038 205728
rect 40094 205672 41460 205728
rect 40033 205670 41460 205672
rect 40033 205667 40099 205670
rect 41454 205668 41460 205670
rect 41524 205668 41530 205732
rect 35574 205325 35634 205564
rect 669262 205396 669268 205460
rect 669332 205458 669338 205460
rect 669630 205458 669636 205460
rect 669332 205398 669636 205458
rect 669332 205396 669338 205398
rect 669630 205396 669636 205398
rect 669700 205396 669706 205460
rect 35574 205320 35683 205325
rect 35574 205264 35622 205320
rect 35678 205264 35683 205320
rect 35574 205262 35683 205264
rect 35617 205259 35683 205262
rect 39573 205322 39639 205325
rect 44173 205322 44239 205325
rect 39573 205320 44239 205322
rect 39573 205264 39578 205320
rect 39634 205264 44178 205320
rect 44234 205264 44239 205320
rect 39573 205262 44239 205264
rect 39573 205259 39639 205262
rect 44173 205259 44239 205262
rect 589457 205186 589523 205189
rect 589457 205184 592602 205186
rect 35758 204917 35818 205156
rect 589457 205128 589462 205184
rect 589518 205128 592602 205184
rect 589457 205126 592602 205128
rect 589457 205123 589523 205126
rect 35758 204912 35867 204917
rect 35758 204856 35806 204912
rect 35862 204856 35867 204912
rect 35758 204854 35867 204856
rect 35801 204851 35867 204854
rect 40309 204914 40375 204917
rect 43253 204914 43319 204917
rect 40309 204912 43319 204914
rect 40309 204856 40314 204912
rect 40370 204856 43258 204912
rect 43314 204856 43319 204912
rect 40309 204854 43319 204856
rect 40309 204851 40375 204854
rect 43253 204851 43319 204854
rect 592542 204816 592602 205126
rect 675753 205050 675819 205053
rect 676254 205050 676260 205052
rect 675753 205048 676260 205050
rect 675753 204992 675758 205048
rect 675814 204992 676260 205048
rect 675753 204990 676260 204992
rect 675753 204987 675819 204990
rect 676254 204988 676260 204990
rect 676324 204988 676330 205052
rect 35574 204509 35634 204748
rect 35525 204504 35634 204509
rect 35801 204506 35867 204509
rect 35525 204448 35530 204504
rect 35586 204448 35634 204504
rect 35525 204446 35634 204448
rect 35758 204504 35867 204506
rect 35758 204448 35806 204504
rect 35862 204448 35867 204504
rect 35525 204443 35591 204446
rect 35758 204443 35867 204448
rect 39389 204506 39455 204509
rect 43437 204506 43503 204509
rect 39389 204504 43503 204506
rect 39389 204448 39394 204504
rect 39450 204448 43442 204504
rect 43498 204448 43503 204504
rect 39389 204446 43503 204448
rect 39389 204443 39455 204446
rect 43437 204443 43503 204446
rect 35758 204340 35818 204443
rect 39941 204098 40007 204101
rect 44541 204098 44607 204101
rect 669446 204098 669452 204100
rect 39941 204096 44607 204098
rect 39941 204040 39946 204096
rect 40002 204040 44546 204096
rect 44602 204040 44607 204096
rect 39941 204038 44607 204040
rect 39941 204035 40007 204038
rect 44541 204035 44607 204038
rect 666878 204038 669452 204098
rect 666878 204030 666938 204038
rect 669446 204036 669452 204038
rect 669516 204036 669522 204100
rect 666356 203970 666938 204030
rect 35574 203693 35634 203932
rect 35574 203688 35683 203693
rect 35574 203632 35622 203688
rect 35678 203632 35683 203688
rect 35574 203630 35683 203632
rect 35617 203627 35683 203630
rect 41137 203690 41203 203693
rect 43621 203690 43687 203693
rect 41137 203688 43687 203690
rect 41137 203632 41142 203688
rect 41198 203632 43626 203688
rect 43682 203632 43687 203688
rect 41137 203630 43687 203632
rect 41137 203627 41203 203630
rect 43621 203627 43687 203630
rect 589457 203690 589523 203693
rect 589457 203688 592602 203690
rect 589457 203632 589462 203688
rect 589518 203632 592602 203688
rect 589457 203630 592602 203632
rect 589457 203627 589523 203630
rect 35758 203285 35818 203524
rect 35758 203280 35867 203285
rect 35758 203224 35806 203280
rect 35862 203224 35867 203280
rect 35758 203222 35867 203224
rect 35801 203219 35867 203222
rect 41229 203282 41295 203285
rect 43805 203282 43871 203285
rect 41229 203280 43871 203282
rect 41229 203224 41234 203280
rect 41290 203224 43810 203280
rect 43866 203224 43871 203280
rect 41229 203222 43871 203224
rect 575982 203282 576042 203524
rect 578325 203282 578391 203285
rect 575982 203280 578391 203282
rect 575982 203224 578330 203280
rect 578386 203224 578391 203280
rect 575982 203222 578391 203224
rect 41229 203219 41295 203222
rect 43805 203219 43871 203222
rect 578325 203219 578391 203222
rect 592542 203184 592602 203630
rect 668158 202466 668164 202468
rect 666694 202406 668164 202466
rect 666694 202398 666754 202406
rect 668158 202404 668164 202406
rect 668228 202404 668234 202468
rect 666356 202338 666754 202398
rect 589457 202194 589523 202197
rect 589457 202192 592602 202194
rect 589457 202136 589462 202192
rect 589518 202136 592602 202192
rect 589457 202134 592602 202136
rect 589457 202131 589523 202134
rect 592542 201552 592602 202134
rect 670785 201514 670851 201517
rect 670785 201512 672044 201514
rect 670785 201456 670790 201512
rect 670846 201510 672044 201512
rect 670846 201456 672090 201510
rect 670785 201454 672090 201456
rect 670785 201451 670851 201454
rect 671984 201450 672090 201454
rect 672030 201378 672090 201450
rect 676806 201378 676812 201380
rect 672030 201318 676812 201378
rect 676806 201316 676812 201318
rect 676876 201316 676882 201380
rect 30281 200698 30347 200701
rect 41638 200698 41644 200700
rect 30281 200696 41644 200698
rect 30281 200640 30286 200696
rect 30342 200640 41644 200696
rect 30281 200638 41644 200640
rect 30281 200635 30347 200638
rect 41638 200636 41644 200638
rect 41708 200636 41714 200700
rect 575982 200698 576042 201076
rect 579153 200698 579219 200701
rect 575982 200696 579219 200698
rect 575982 200640 579158 200696
rect 579214 200640 579219 200696
rect 575982 200638 579219 200640
rect 579153 200635 579219 200638
rect 675753 200018 675819 200021
rect 676622 200018 676628 200020
rect 675753 200016 676628 200018
rect 675753 199960 675758 200016
rect 675814 199960 676628 200016
rect 675753 199958 676628 199960
rect 675753 199955 675819 199958
rect 676622 199956 676628 199958
rect 676692 199956 676698 200020
rect 589457 199882 589523 199885
rect 589457 199880 592572 199882
rect 589457 199824 589462 199880
rect 589518 199824 592572 199880
rect 589457 199822 592572 199824
rect 589457 199819 589523 199822
rect 666870 199134 666876 199136
rect 666356 199074 666876 199134
rect 666870 199072 666876 199074
rect 666940 199072 666946 199136
rect 590561 198658 590627 198661
rect 590561 198656 592602 198658
rect 575982 198114 576042 198628
rect 590561 198600 590566 198656
rect 590622 198600 592602 198656
rect 590561 198598 592602 198600
rect 590561 198595 590627 198598
rect 592542 198288 592602 198598
rect 675753 198388 675819 198389
rect 675702 198386 675708 198388
rect 675662 198326 675708 198386
rect 675772 198384 675819 198388
rect 675814 198328 675819 198384
rect 675702 198324 675708 198326
rect 675772 198324 675819 198328
rect 675753 198323 675819 198324
rect 578877 198114 578943 198117
rect 575982 198112 578943 198114
rect 575982 198056 578882 198112
rect 578938 198056 578943 198112
rect 575982 198054 578943 198056
rect 578877 198051 578943 198054
rect 668342 197570 668348 197572
rect 666694 197510 668348 197570
rect 666694 197502 666754 197510
rect 668342 197508 668348 197510
rect 668412 197508 668418 197572
rect 666356 197442 666754 197502
rect 40902 197100 40908 197164
rect 40972 197162 40978 197164
rect 41781 197162 41847 197165
rect 40972 197160 41847 197162
rect 40972 197104 41786 197160
rect 41842 197104 41847 197160
rect 40972 197102 41847 197104
rect 40972 197100 40978 197102
rect 41781 197099 41847 197102
rect 589457 197026 589523 197029
rect 675753 197026 675819 197029
rect 676438 197026 676444 197028
rect 589457 197024 592602 197026
rect 589457 196968 589462 197024
rect 589518 196968 592602 197024
rect 589457 196966 592602 196968
rect 589457 196963 589523 196966
rect 592542 196656 592602 196966
rect 675753 197024 676444 197026
rect 675753 196968 675758 197024
rect 675814 196968 676444 197024
rect 675753 196966 676444 196968
rect 675753 196963 675819 196966
rect 676438 196964 676444 196966
rect 676508 196964 676514 197028
rect 575982 196074 576042 196180
rect 579521 196074 579587 196077
rect 575982 196072 579587 196074
rect 575982 196016 579526 196072
rect 579582 196016 579587 196072
rect 575982 196014 579587 196016
rect 579521 196011 579587 196014
rect 589549 195530 589615 195533
rect 589549 195528 592602 195530
rect 589549 195472 589554 195528
rect 589610 195472 592602 195528
rect 589549 195470 592602 195472
rect 589549 195467 589615 195470
rect 41781 195260 41847 195261
rect 41781 195256 41828 195260
rect 41892 195258 41898 195260
rect 41781 195200 41786 195256
rect 41781 195196 41828 195200
rect 41892 195198 41938 195258
rect 41892 195196 41898 195198
rect 41781 195195 41847 195196
rect 592542 195024 592602 195470
rect 666870 194238 666876 194240
rect 666356 194178 666876 194238
rect 666870 194176 666876 194178
rect 666940 194176 666946 194240
rect 579521 193898 579587 193901
rect 575798 193896 579587 193898
rect 575798 193840 579526 193896
rect 579582 193840 579587 193896
rect 575798 193838 579587 193840
rect 575798 193732 575858 193838
rect 579521 193835 579587 193838
rect 589549 193626 589615 193629
rect 589549 193624 592602 193626
rect 589549 193568 589554 193624
rect 589610 193568 592602 193624
rect 589549 193566 592602 193568
rect 589549 193563 589615 193566
rect 592542 193392 592602 193566
rect 670601 193354 670667 193357
rect 675109 193354 675175 193357
rect 670601 193352 675175 193354
rect 670601 193296 670606 193352
rect 670662 193296 675114 193352
rect 675170 193296 675175 193352
rect 670601 193294 675175 193296
rect 670601 193291 670667 193294
rect 675109 193291 675175 193294
rect 675753 193218 675819 193221
rect 676070 193218 676076 193220
rect 675753 193216 676076 193218
rect 675753 193160 675758 193216
rect 675814 193160 676076 193216
rect 675753 193158 676076 193160
rect 675753 193155 675819 193158
rect 676070 193156 676076 193158
rect 676140 193156 676146 193220
rect 675661 192810 675727 192813
rect 675886 192810 675892 192812
rect 675661 192808 675892 192810
rect 675661 192752 675666 192808
rect 675722 192752 675892 192808
rect 675661 192750 675892 192752
rect 675661 192747 675727 192750
rect 675886 192748 675892 192750
rect 675956 192748 675962 192812
rect 666921 192674 666987 192677
rect 666694 192672 666987 192674
rect 666694 192616 666926 192672
rect 666982 192616 666987 192672
rect 666694 192614 666987 192616
rect 666694 192606 666754 192614
rect 666921 192611 666987 192614
rect 666356 192546 666754 192606
rect 589457 191722 589523 191725
rect 589457 191720 592572 191722
rect 589457 191664 589462 191720
rect 589518 191664 592572 191720
rect 589457 191662 592572 191664
rect 589457 191659 589523 191662
rect 40718 191524 40724 191588
rect 40788 191586 40794 191588
rect 41781 191586 41847 191589
rect 40788 191584 41847 191586
rect 40788 191528 41786 191584
rect 41842 191528 41847 191584
rect 40788 191526 41847 191528
rect 40788 191524 40794 191526
rect 41781 191523 41847 191526
rect 575982 191178 576042 191284
rect 579521 191178 579587 191181
rect 575982 191176 579587 191178
rect 575982 191120 579526 191176
rect 579582 191120 579587 191176
rect 575982 191118 579587 191120
rect 579521 191115 579587 191118
rect 589457 190090 589523 190093
rect 673545 190090 673611 190093
rect 675845 190090 675911 190093
rect 589457 190088 592572 190090
rect 589457 190032 589462 190088
rect 589518 190032 592572 190088
rect 589457 190030 592572 190032
rect 673545 190088 675911 190090
rect 673545 190032 673550 190088
rect 673606 190032 675850 190088
rect 675906 190032 675911 190088
rect 673545 190030 675911 190032
rect 589457 190027 589523 190030
rect 673545 190027 673611 190030
rect 675845 190027 675911 190030
rect 666686 189342 666692 189344
rect 666356 189282 666692 189342
rect 666686 189280 666692 189282
rect 666756 189280 666762 189344
rect 579521 189002 579587 189005
rect 575798 189000 579587 189002
rect 575798 188944 579526 189000
rect 579582 188944 579587 189000
rect 575798 188942 579587 188944
rect 575798 188836 575858 188942
rect 579521 188939 579587 188942
rect 589641 188458 589707 188461
rect 589641 188456 592572 188458
rect 589641 188400 589646 188456
rect 589702 188400 592572 188456
rect 589641 188398 592572 188400
rect 589641 188395 589707 188398
rect 668117 187778 668183 187781
rect 666694 187776 668183 187778
rect 666694 187720 668122 187776
rect 668178 187720 668183 187776
rect 666694 187718 668183 187720
rect 666694 187710 666754 187718
rect 668117 187715 668183 187718
rect 666356 187650 666754 187710
rect 589457 186826 589523 186829
rect 589457 186824 592572 186826
rect 589457 186768 589462 186824
rect 589518 186768 592572 186824
rect 589457 186766 592572 186768
rect 589457 186763 589523 186766
rect 579521 186690 579587 186693
rect 575798 186688 579587 186690
rect 575798 186632 579526 186688
rect 579582 186632 579587 186688
rect 575798 186630 579587 186632
rect 575798 186388 575858 186630
rect 579521 186627 579587 186630
rect 41781 185876 41847 185877
rect 41781 185872 41828 185876
rect 41892 185874 41898 185876
rect 41781 185816 41786 185872
rect 41781 185812 41828 185816
rect 41892 185814 41938 185874
rect 41892 185812 41898 185814
rect 41781 185811 41847 185812
rect 589457 185194 589523 185197
rect 589457 185192 592572 185194
rect 589457 185136 589462 185192
rect 589518 185136 592572 185192
rect 589457 185134 592572 185136
rect 589457 185131 589523 185134
rect 666553 184786 666619 184789
rect 666553 184784 666938 184786
rect 666553 184728 666558 184784
rect 666614 184728 666938 184784
rect 666553 184726 666938 184728
rect 666553 184723 666619 184726
rect 666878 184446 666938 184726
rect 666356 184386 666938 184446
rect 578509 184378 578575 184381
rect 575798 184376 578575 184378
rect 575798 184320 578514 184376
rect 578570 184320 578575 184376
rect 575798 184318 578575 184320
rect 41454 184044 41460 184108
rect 41524 184106 41530 184108
rect 41781 184106 41847 184109
rect 41524 184104 41847 184106
rect 41524 184048 41786 184104
rect 41842 184048 41847 184104
rect 41524 184046 41847 184048
rect 41524 184044 41530 184046
rect 41781 184043 41847 184046
rect 575798 183940 575858 184318
rect 578509 184315 578575 184318
rect 589457 183562 589523 183565
rect 672349 183562 672415 183565
rect 673177 183564 673243 183565
rect 672758 183562 672764 183564
rect 589457 183560 592572 183562
rect 589457 183504 589462 183560
rect 589518 183504 592572 183560
rect 589457 183502 592572 183504
rect 672349 183560 672764 183562
rect 672349 183504 672354 183560
rect 672410 183504 672764 183560
rect 672349 183502 672764 183504
rect 589457 183499 589523 183502
rect 672349 183499 672415 183502
rect 672758 183500 672764 183502
rect 672828 183500 672834 183564
rect 673126 183562 673132 183564
rect 673086 183502 673132 183562
rect 673196 183560 673243 183564
rect 673238 183504 673243 183560
rect 673126 183500 673132 183502
rect 673196 183500 673243 183504
rect 673177 183499 673243 183500
rect 40534 183364 40540 183428
rect 40604 183426 40610 183428
rect 41781 183426 41847 183429
rect 40604 183424 41847 183426
rect 40604 183368 41786 183424
rect 41842 183368 41847 183424
rect 40604 183366 41847 183368
rect 40604 183364 40610 183366
rect 41781 183363 41847 183366
rect 669221 182882 669287 182885
rect 666694 182880 669287 182882
rect 666694 182824 669226 182880
rect 669282 182824 669287 182880
rect 666694 182822 669287 182824
rect 666694 182814 666754 182822
rect 669221 182819 669287 182822
rect 666356 182754 666754 182814
rect 579429 182066 579495 182069
rect 575798 182064 579495 182066
rect 575798 182008 579434 182064
rect 579490 182008 579495 182064
rect 575798 182006 579495 182008
rect 575798 181492 575858 182006
rect 579429 182003 579495 182006
rect 589457 181930 589523 181933
rect 589457 181928 592572 181930
rect 589457 181872 589462 181928
rect 589518 181872 592572 181928
rect 589457 181870 592572 181872
rect 589457 181867 589523 181870
rect 589457 180298 589523 180301
rect 589457 180296 592572 180298
rect 589457 180240 589462 180296
rect 589518 180240 592572 180296
rect 589457 180238 592572 180240
rect 589457 180235 589523 180238
rect 669446 179618 669452 179620
rect 666694 179558 669452 179618
rect 666694 179550 666754 179558
rect 669446 179556 669452 179558
rect 669516 179556 669522 179620
rect 666356 179490 666754 179550
rect 578325 179210 578391 179213
rect 575798 179208 578391 179210
rect 575798 179152 578330 179208
rect 578386 179152 578391 179208
rect 575798 179150 578391 179152
rect 575798 179044 575858 179150
rect 578325 179147 578391 179150
rect 589457 178666 589523 178669
rect 589457 178664 592572 178666
rect 589457 178608 589462 178664
rect 589518 178608 592572 178664
rect 589457 178606 592572 178608
rect 589457 178603 589523 178606
rect 675293 178530 675359 178533
rect 675293 178528 676292 178530
rect 675293 178472 675298 178528
rect 675354 178472 676292 178528
rect 675293 178470 676292 178472
rect 675293 178467 675359 178470
rect 675477 178122 675543 178125
rect 675477 178120 676292 178122
rect 675477 178064 675482 178120
rect 675538 178064 676292 178120
rect 675477 178062 676292 178064
rect 675477 178059 675543 178062
rect 667933 177986 667999 177989
rect 666694 177984 667999 177986
rect 666694 177928 667938 177984
rect 667994 177928 667999 177984
rect 666694 177926 667999 177928
rect 666694 177918 666754 177926
rect 667933 177923 667999 177926
rect 666356 177858 666754 177918
rect 683113 177714 683179 177717
rect 683100 177712 683179 177714
rect 683100 177656 683118 177712
rect 683174 177656 683179 177712
rect 683100 177654 683179 177656
rect 683113 177651 683179 177654
rect 675293 177306 675359 177309
rect 675293 177304 676292 177306
rect 675293 177248 675298 177304
rect 675354 177248 676292 177304
rect 675293 177246 676292 177248
rect 675293 177243 675359 177246
rect 589457 177034 589523 177037
rect 589457 177032 592572 177034
rect 589457 176976 589462 177032
rect 589518 176976 592572 177032
rect 589457 176974 592572 176976
rect 589457 176971 589523 176974
rect 675477 176898 675543 176901
rect 675477 176896 676292 176898
rect 675477 176840 675482 176896
rect 675538 176840 676292 176896
rect 675477 176838 676292 176840
rect 675477 176835 675543 176838
rect 669129 176626 669195 176629
rect 669129 176624 676230 176626
rect 575982 176490 576042 176596
rect 669129 176568 669134 176624
rect 669190 176568 676230 176624
rect 669129 176566 676230 176568
rect 669129 176563 669195 176566
rect 579521 176490 579587 176493
rect 575982 176488 579587 176490
rect 575982 176432 579526 176488
rect 579582 176432 579587 176488
rect 575982 176430 579587 176432
rect 676170 176490 676230 176566
rect 676170 176430 676292 176490
rect 579521 176427 579587 176430
rect 674741 176082 674807 176085
rect 674741 176080 676292 176082
rect 674741 176024 674746 176080
rect 674802 176024 676292 176080
rect 674741 176022 676292 176024
rect 674741 176019 674807 176022
rect 674557 175674 674623 175677
rect 674557 175672 676292 175674
rect 674557 175616 674562 175672
rect 674618 175616 676292 175672
rect 674557 175614 676292 175616
rect 674557 175611 674623 175614
rect 589273 175402 589339 175405
rect 589273 175400 592572 175402
rect 589273 175344 589278 175400
rect 589334 175344 592572 175400
rect 589273 175342 592572 175344
rect 589273 175339 589339 175342
rect 675477 175266 675543 175269
rect 675477 175264 676292 175266
rect 675477 175208 675482 175264
rect 675538 175208 676292 175264
rect 675477 175206 676292 175208
rect 675477 175203 675543 175206
rect 676170 174798 676292 174858
rect 578693 174722 578759 174725
rect 667933 174722 667999 174725
rect 575798 174720 578759 174722
rect 575798 174664 578698 174720
rect 578754 174664 578759 174720
rect 575798 174662 578759 174664
rect 575798 174148 575858 174662
rect 578693 174659 578759 174662
rect 666694 174720 667999 174722
rect 666694 174664 667938 174720
rect 667994 174664 667999 174720
rect 666694 174662 667999 174664
rect 666694 174654 666754 174662
rect 667933 174659 667999 174662
rect 675886 174660 675892 174724
rect 675956 174722 675962 174724
rect 676170 174722 676230 174798
rect 675956 174662 676230 174722
rect 675956 174660 675962 174662
rect 666356 174594 666754 174654
rect 674465 174450 674531 174453
rect 674465 174448 676292 174450
rect 674465 174392 674470 174448
rect 674526 174392 676292 174448
rect 674465 174390 676292 174392
rect 674465 174387 674531 174390
rect 675293 174042 675359 174045
rect 675293 174040 676292 174042
rect 675293 173984 675298 174040
rect 675354 173984 676292 174040
rect 675293 173982 676292 173984
rect 675293 173979 675359 173982
rect 589733 173770 589799 173773
rect 589733 173768 592572 173770
rect 589733 173712 589738 173768
rect 589794 173712 592572 173768
rect 589733 173710 592572 173712
rect 589733 173707 589799 173710
rect 675702 173572 675708 173636
rect 675772 173634 675778 173636
rect 675772 173574 676292 173634
rect 675772 173572 675778 173574
rect 675845 173226 675911 173229
rect 675845 173224 676292 173226
rect 675845 173168 675850 173224
rect 675906 173168 676292 173224
rect 675845 173166 676292 173168
rect 675845 173163 675911 173166
rect 673310 173090 673316 173092
rect 666694 173030 673316 173090
rect 666694 173022 666754 173030
rect 673310 173028 673316 173030
rect 673380 173028 673386 173092
rect 666356 172962 666754 173022
rect 675109 172818 675175 172821
rect 675109 172816 676292 172818
rect 675109 172760 675114 172816
rect 675170 172760 676292 172816
rect 675109 172758 676292 172760
rect 675109 172755 675175 172758
rect 675334 172348 675340 172412
rect 675404 172410 675410 172412
rect 675404 172350 676292 172410
rect 675404 172348 675410 172350
rect 579521 172138 579587 172141
rect 575798 172136 579587 172138
rect 575798 172080 579526 172136
rect 579582 172080 579587 172136
rect 575798 172078 579587 172080
rect 575798 171700 575858 172078
rect 579521 172075 579587 172078
rect 589457 172138 589523 172141
rect 589457 172136 592572 172138
rect 589457 172080 589462 172136
rect 589518 172080 592572 172136
rect 589457 172078 592572 172080
rect 589457 172075 589523 172078
rect 675477 172002 675543 172005
rect 675477 172000 676292 172002
rect 675477 171944 675482 172000
rect 675538 171944 676292 172000
rect 675477 171942 676292 171944
rect 675477 171939 675543 171942
rect 678237 171594 678303 171597
rect 678237 171592 678316 171594
rect 678237 171536 678242 171592
rect 678298 171536 678316 171592
rect 678237 171534 678316 171536
rect 678237 171531 678303 171534
rect 675477 171186 675543 171189
rect 675477 171184 676292 171186
rect 675477 171128 675482 171184
rect 675538 171128 676292 171184
rect 675477 171126 676292 171128
rect 675477 171123 675543 171126
rect 675886 170716 675892 170780
rect 675956 170778 675962 170780
rect 675956 170718 676292 170778
rect 675956 170716 675962 170718
rect 588537 170506 588603 170509
rect 588537 170504 592572 170506
rect 588537 170448 588542 170504
rect 588598 170448 592572 170504
rect 588537 170446 592572 170448
rect 588537 170443 588603 170446
rect 675477 170370 675543 170373
rect 675477 170368 676292 170370
rect 675477 170312 675482 170368
rect 675538 170312 676292 170368
rect 675477 170310 676292 170312
rect 675477 170307 675543 170310
rect 676673 169962 676739 169965
rect 676660 169960 676739 169962
rect 676660 169904 676678 169960
rect 676734 169904 676739 169960
rect 676660 169902 676739 169904
rect 676673 169899 676739 169902
rect 666356 169698 666754 169758
rect 666694 169690 666754 169698
rect 667933 169690 667999 169693
rect 666694 169688 667999 169690
rect 666694 169632 667938 169688
rect 667994 169632 667999 169688
rect 666694 169630 667999 169632
rect 667933 169627 667999 169630
rect 579245 169554 579311 169557
rect 575798 169552 579311 169554
rect 575798 169496 579250 169552
rect 579306 169496 579311 169552
rect 575798 169494 579311 169496
rect 575798 169252 575858 169494
rect 579245 169491 579311 169494
rect 676170 169494 676292 169554
rect 675886 169356 675892 169420
rect 675956 169418 675962 169420
rect 676170 169418 676230 169494
rect 675956 169358 676230 169418
rect 675956 169356 675962 169358
rect 675477 169146 675543 169149
rect 675477 169144 676292 169146
rect 675477 169088 675482 169144
rect 675538 169088 676292 169144
rect 675477 169086 676292 169088
rect 675477 169083 675543 169086
rect 589457 168874 589523 168877
rect 589457 168872 592572 168874
rect 589457 168816 589462 168872
rect 589518 168816 592572 168872
rect 589457 168814 592572 168816
rect 589457 168811 589523 168814
rect 675477 168738 675543 168741
rect 675477 168736 676292 168738
rect 675477 168680 675482 168736
rect 675538 168680 676292 168736
rect 675477 168678 676292 168680
rect 675477 168675 675543 168678
rect 672165 168330 672231 168333
rect 672942 168330 672948 168332
rect 672165 168328 672948 168330
rect 672165 168272 672170 168328
rect 672226 168272 672948 168328
rect 672165 168270 672948 168272
rect 672165 168267 672231 168270
rect 672942 168268 672948 168270
rect 673012 168268 673018 168332
rect 675477 168330 675543 168333
rect 675477 168328 676292 168330
rect 675477 168272 675482 168328
rect 675538 168272 676292 168328
rect 675477 168270 676292 168272
rect 675477 168267 675543 168270
rect 668577 168194 668643 168197
rect 666694 168192 668643 168194
rect 666694 168136 668582 168192
rect 668638 168136 668643 168192
rect 666694 168134 668643 168136
rect 666694 168126 666754 168134
rect 668577 168131 668643 168134
rect 666356 168066 666754 168126
rect 675477 167922 675543 167925
rect 675477 167920 676292 167922
rect 675477 167864 675482 167920
rect 675538 167864 676292 167920
rect 675477 167862 676292 167864
rect 675477 167859 675543 167862
rect 675702 167588 675708 167652
rect 675772 167650 675778 167652
rect 675772 167590 676230 167650
rect 675772 167588 675778 167590
rect 676170 167514 676230 167590
rect 676170 167454 676292 167514
rect 589457 167242 589523 167245
rect 589457 167240 592572 167242
rect 589457 167184 589462 167240
rect 589518 167184 592572 167240
rect 589457 167182 592572 167184
rect 589457 167179 589523 167182
rect 675477 167106 675543 167109
rect 675477 167104 676292 167106
rect 675477 167048 675482 167104
rect 675538 167048 676292 167104
rect 675477 167046 676292 167048
rect 675477 167043 675543 167046
rect 578877 166970 578943 166973
rect 575798 166968 578943 166970
rect 575798 166912 578882 166968
rect 578938 166912 578943 166968
rect 575798 166910 578943 166912
rect 575798 166804 575858 166910
rect 578877 166907 578943 166910
rect 676673 166428 676739 166429
rect 676622 166426 676628 166428
rect 676582 166366 676628 166426
rect 676692 166424 676739 166428
rect 676734 166368 676739 166424
rect 676622 166364 676628 166366
rect 676692 166364 676739 166368
rect 676673 166363 676739 166364
rect 668577 165746 668643 165749
rect 670918 165746 670924 165748
rect 668577 165744 670924 165746
rect 668577 165688 668582 165744
rect 668638 165688 670924 165744
rect 668577 165686 670924 165688
rect 668577 165683 668643 165686
rect 670918 165684 670924 165686
rect 670988 165684 670994 165748
rect 589457 165610 589523 165613
rect 589457 165608 592572 165610
rect 589457 165552 589462 165608
rect 589518 165552 592572 165608
rect 589457 165550 592572 165552
rect 589457 165547 589523 165550
rect 668025 164930 668091 164933
rect 666694 164928 668091 164930
rect 666694 164872 668030 164928
rect 668086 164872 668091 164928
rect 666694 164870 668091 164872
rect 666694 164862 666754 164870
rect 668025 164867 668091 164870
rect 666356 164802 666754 164862
rect 579521 164522 579587 164525
rect 575798 164520 579587 164522
rect 575798 164464 579526 164520
rect 579582 164464 579587 164520
rect 575798 164462 579587 164464
rect 575798 164356 575858 164462
rect 579521 164459 579587 164462
rect 589733 163978 589799 163981
rect 589733 163976 592572 163978
rect 589733 163920 589738 163976
rect 589794 163920 592572 163976
rect 589733 163918 592572 163920
rect 589733 163915 589799 163918
rect 668577 163298 668643 163301
rect 666694 163296 668643 163298
rect 666694 163240 668582 163296
rect 668638 163240 668643 163296
rect 666694 163238 668643 163240
rect 666694 163230 666754 163238
rect 668577 163235 668643 163238
rect 666356 163170 666754 163230
rect 579521 162482 579587 162485
rect 575798 162480 579587 162482
rect 575798 162424 579526 162480
rect 579582 162424 579587 162480
rect 575798 162422 579587 162424
rect 575798 161908 575858 162422
rect 579521 162419 579587 162422
rect 590101 162346 590167 162349
rect 590101 162344 592572 162346
rect 590101 162288 590106 162344
rect 590162 162288 592572 162344
rect 590101 162286 592572 162288
rect 590101 162283 590167 162286
rect 675334 162148 675340 162212
rect 675404 162210 675410 162212
rect 675886 162210 675892 162212
rect 675404 162150 675892 162210
rect 675404 162148 675410 162150
rect 675886 162148 675892 162150
rect 675956 162148 675962 162212
rect 675518 161332 675524 161396
rect 675588 161394 675594 161396
rect 675845 161394 675911 161397
rect 675588 161392 675911 161394
rect 675588 161336 675850 161392
rect 675906 161336 675911 161392
rect 675588 161334 675911 161336
rect 675588 161332 675594 161334
rect 675845 161331 675911 161334
rect 589457 160714 589523 160717
rect 589457 160712 592572 160714
rect 589457 160656 589462 160712
rect 589518 160656 592572 160712
rect 589457 160654 592572 160656
rect 589457 160651 589523 160654
rect 675569 160172 675635 160173
rect 675518 160108 675524 160172
rect 675588 160170 675635 160172
rect 675588 160168 675680 160170
rect 675630 160112 675680 160168
rect 675588 160110 675680 160112
rect 675588 160108 675635 160110
rect 675569 160107 675635 160108
rect 666921 160034 666987 160037
rect 666694 160032 666987 160034
rect 666694 159976 666926 160032
rect 666982 159976 666987 160032
rect 666694 159974 666987 159976
rect 666694 159966 666754 159974
rect 666921 159971 666987 159974
rect 666356 159906 666754 159966
rect 579521 159762 579587 159765
rect 575798 159760 579587 159762
rect 575798 159704 579526 159760
rect 579582 159704 579587 159760
rect 575798 159702 579587 159704
rect 575798 159460 575858 159702
rect 579521 159699 579587 159702
rect 588721 159082 588787 159085
rect 588721 159080 592572 159082
rect 588721 159024 588726 159080
rect 588782 159024 592572 159080
rect 588721 159022 592572 159024
rect 588721 159019 588787 159022
rect 668761 158402 668827 158405
rect 666694 158400 668827 158402
rect 666694 158344 668766 158400
rect 668822 158344 668827 158400
rect 666694 158342 668827 158344
rect 666694 158334 666754 158342
rect 668761 158339 668827 158342
rect 666356 158274 666754 158334
rect 589457 157450 589523 157453
rect 589457 157448 592572 157450
rect 589457 157392 589462 157448
rect 589518 157392 592572 157448
rect 589457 157390 592572 157392
rect 589457 157387 589523 157390
rect 579245 157178 579311 157181
rect 575798 157176 579311 157178
rect 575798 157120 579250 157176
rect 579306 157120 579311 157176
rect 575798 157118 579311 157120
rect 575798 157012 575858 157118
rect 579245 157115 579311 157118
rect 675753 156498 675819 156501
rect 676438 156498 676444 156500
rect 675753 156496 676444 156498
rect 675753 156440 675758 156496
rect 675814 156440 676444 156496
rect 675753 156438 676444 156440
rect 675753 156435 675819 156438
rect 676438 156436 676444 156438
rect 676508 156436 676514 156500
rect 589365 155818 589431 155821
rect 589365 155816 592572 155818
rect 589365 155760 589370 155816
rect 589426 155760 592572 155816
rect 589365 155758 592572 155760
rect 589365 155755 589431 155758
rect 675753 155682 675819 155685
rect 676254 155682 676260 155684
rect 675753 155680 676260 155682
rect 675753 155624 675758 155680
rect 675814 155624 676260 155680
rect 675753 155622 676260 155624
rect 675753 155619 675819 155622
rect 676254 155620 676260 155622
rect 676324 155620 676330 155684
rect 578693 155138 578759 155141
rect 670734 155138 670740 155140
rect 575798 155136 578759 155138
rect 575798 155080 578698 155136
rect 578754 155080 578759 155136
rect 575798 155078 578759 155080
rect 575798 154564 575858 155078
rect 578693 155075 578759 155078
rect 666694 155078 670740 155138
rect 666694 155070 666754 155078
rect 670734 155076 670740 155078
rect 670804 155076 670810 155140
rect 666356 155010 666754 155070
rect 589457 154186 589523 154189
rect 589457 154184 592572 154186
rect 589457 154128 589462 154184
rect 589518 154128 592572 154184
rect 589457 154126 592572 154128
rect 589457 154123 589523 154126
rect 666356 153378 666938 153438
rect 666878 153370 666938 153378
rect 673678 153370 673684 153372
rect 666878 153310 673684 153370
rect 673678 153308 673684 153310
rect 673748 153308 673754 153372
rect 675661 153098 675727 153101
rect 675886 153098 675892 153100
rect 675661 153096 675892 153098
rect 675661 153040 675666 153096
rect 675722 153040 675892 153096
rect 675661 153038 675892 153040
rect 675661 153035 675727 153038
rect 675886 153036 675892 153038
rect 675956 153036 675962 153100
rect 578325 152690 578391 152693
rect 575798 152688 578391 152690
rect 575798 152632 578330 152688
rect 578386 152632 578391 152688
rect 575798 152630 578391 152632
rect 575798 152116 575858 152630
rect 578325 152627 578391 152630
rect 589733 152554 589799 152557
rect 589733 152552 592572 152554
rect 589733 152496 589738 152552
rect 589794 152496 592572 152552
rect 589733 152494 592572 152496
rect 589733 152491 589799 152494
rect 675753 151466 675819 151469
rect 676622 151466 676628 151468
rect 675753 151464 676628 151466
rect 675753 151408 675758 151464
rect 675814 151408 676628 151464
rect 675753 151406 676628 151408
rect 675753 151403 675819 151406
rect 676622 151404 676628 151406
rect 676692 151404 676698 151468
rect 589917 150922 589983 150925
rect 589917 150920 592572 150922
rect 589917 150864 589922 150920
rect 589978 150864 592572 150920
rect 589917 150862 592572 150864
rect 589917 150859 589983 150862
rect 668761 150242 668827 150245
rect 666694 150240 668827 150242
rect 666694 150184 668766 150240
rect 668822 150184 668827 150240
rect 666694 150182 668827 150184
rect 666694 150174 666754 150182
rect 668761 150179 668827 150182
rect 666356 150114 666754 150174
rect 579521 150106 579587 150109
rect 575798 150104 579587 150106
rect 575798 150048 579526 150104
rect 579582 150048 579587 150104
rect 575798 150046 579587 150048
rect 575798 149668 575858 150046
rect 579521 150043 579587 150046
rect 589273 149290 589339 149293
rect 589273 149288 592572 149290
rect 589273 149232 589278 149288
rect 589334 149232 592572 149288
rect 589273 149230 592572 149232
rect 589273 149227 589339 149230
rect 666356 148482 666938 148542
rect 666878 148474 666938 148482
rect 673494 148474 673500 148476
rect 666878 148414 673500 148474
rect 673494 148412 673500 148414
rect 673564 148412 673570 148476
rect 675753 148474 675819 148477
rect 676070 148474 676076 148476
rect 675753 148472 676076 148474
rect 675753 148416 675758 148472
rect 675814 148416 676076 148472
rect 675753 148414 676076 148416
rect 675753 148411 675819 148414
rect 676070 148412 676076 148414
rect 676140 148412 676146 148476
rect 578417 147658 578483 147661
rect 575798 147656 578483 147658
rect 575798 147600 578422 147656
rect 578478 147600 578483 147656
rect 575798 147598 578483 147600
rect 575798 147220 575858 147598
rect 578417 147595 578483 147598
rect 589457 147658 589523 147661
rect 675661 147660 675727 147661
rect 589457 147656 592572 147658
rect 589457 147600 589462 147656
rect 589518 147600 592572 147656
rect 589457 147598 592572 147600
rect 675661 147656 675708 147660
rect 675772 147658 675778 147660
rect 675661 147600 675666 147656
rect 589457 147595 589523 147598
rect 675661 147596 675708 147600
rect 675772 147598 675818 147658
rect 675772 147596 675778 147598
rect 675661 147595 675727 147596
rect 589457 146026 589523 146029
rect 589457 146024 592572 146026
rect 589457 145968 589462 146024
rect 589518 145968 592572 146024
rect 589457 145966 592572 145968
rect 589457 145963 589523 145966
rect 668761 145346 668827 145349
rect 666694 145344 668827 145346
rect 666694 145288 668766 145344
rect 668822 145288 668827 145344
rect 666694 145286 668827 145288
rect 666694 145278 666754 145286
rect 668761 145283 668827 145286
rect 666356 145218 666754 145278
rect 575982 144666 576042 144772
rect 578785 144666 578851 144669
rect 575982 144664 578851 144666
rect 575982 144608 578790 144664
rect 578846 144608 578851 144664
rect 575982 144606 578851 144608
rect 578785 144603 578851 144606
rect 588537 144394 588603 144397
rect 588537 144392 592572 144394
rect 588537 144336 588542 144392
rect 588598 144336 592572 144392
rect 588537 144334 592572 144336
rect 588537 144331 588603 144334
rect 668577 143714 668643 143717
rect 666694 143712 668643 143714
rect 666694 143656 668582 143712
rect 668638 143656 668643 143712
rect 666694 143654 668643 143656
rect 666694 143646 666754 143654
rect 668577 143651 668643 143654
rect 666356 143586 666754 143646
rect 579245 142898 579311 142901
rect 575798 142896 579311 142898
rect 575798 142840 579250 142896
rect 579306 142840 579311 142896
rect 575798 142838 579311 142840
rect 575798 142324 575858 142838
rect 579245 142835 579311 142838
rect 590285 142762 590351 142765
rect 590285 142760 592572 142762
rect 590285 142704 590290 142760
rect 590346 142704 592572 142760
rect 590285 142702 592572 142704
rect 590285 142699 590351 142702
rect 589457 141130 589523 141133
rect 589457 141128 592572 141130
rect 589457 141072 589462 141128
rect 589518 141072 592572 141128
rect 589457 141070 592572 141072
rect 589457 141067 589523 141070
rect 668669 140450 668735 140453
rect 666694 140448 668735 140450
rect 666694 140392 668674 140448
rect 668730 140392 668735 140448
rect 666694 140390 668735 140392
rect 666694 140382 666754 140390
rect 668669 140387 668735 140390
rect 666356 140322 666754 140382
rect 579521 140314 579587 140317
rect 575798 140312 579587 140314
rect 575798 140256 579526 140312
rect 579582 140256 579587 140312
rect 575798 140254 579587 140256
rect 575798 139876 575858 140254
rect 579521 140251 579587 140254
rect 589457 139498 589523 139501
rect 589457 139496 592572 139498
rect 589457 139440 589462 139496
rect 589518 139440 592572 139496
rect 589457 139438 592572 139440
rect 589457 139435 589523 139438
rect 666356 138690 666754 138750
rect 666694 138682 666754 138690
rect 668761 138682 668827 138685
rect 666694 138680 668827 138682
rect 666694 138624 668766 138680
rect 668822 138624 668827 138680
rect 666694 138622 668827 138624
rect 668761 138619 668827 138622
rect 589917 137866 589983 137869
rect 589917 137864 592572 137866
rect 589917 137808 589922 137864
rect 589978 137808 592572 137864
rect 589917 137806 592572 137808
rect 589917 137803 589983 137806
rect 578325 137730 578391 137733
rect 575798 137728 578391 137730
rect 575798 137672 578330 137728
rect 578386 137672 578391 137728
rect 575798 137670 578391 137672
rect 575798 137428 575858 137670
rect 578325 137667 578391 137670
rect 589457 136234 589523 136237
rect 589457 136232 592572 136234
rect 589457 136176 589462 136232
rect 589518 136176 592572 136232
rect 589457 136174 592572 136176
rect 589457 136171 589523 136174
rect 668761 135554 668827 135557
rect 666694 135552 668827 135554
rect 666694 135496 668766 135552
rect 668822 135496 668827 135552
rect 666694 135494 668827 135496
rect 666694 135486 666754 135494
rect 668761 135491 668827 135494
rect 666356 135426 666754 135486
rect 579337 135146 579403 135149
rect 575798 135144 579403 135146
rect 575798 135088 579342 135144
rect 579398 135088 579403 135144
rect 575798 135086 579403 135088
rect 575798 134980 575858 135086
rect 579337 135083 579403 135086
rect 589457 134602 589523 134605
rect 589457 134600 592572 134602
rect 589457 134544 589462 134600
rect 589518 134544 592572 134600
rect 589457 134542 592572 134544
rect 589457 134539 589523 134542
rect 666356 133794 666754 133854
rect 666694 133786 666754 133794
rect 672942 133786 672948 133788
rect 666694 133726 672948 133786
rect 672942 133724 672948 133726
rect 673012 133724 673018 133788
rect 675293 133378 675359 133381
rect 675293 133376 676292 133378
rect 675293 133320 675298 133376
rect 675354 133320 676292 133376
rect 675293 133318 676292 133320
rect 675293 133315 675359 133318
rect 578325 133106 578391 133109
rect 575798 133104 578391 133106
rect 575798 133048 578330 133104
rect 578386 133048 578391 133104
rect 575798 133046 578391 133048
rect 575798 132532 575858 133046
rect 578325 133043 578391 133046
rect 589457 132970 589523 132973
rect 675477 132970 675543 132973
rect 589457 132968 592572 132970
rect 589457 132912 589462 132968
rect 589518 132912 592572 132968
rect 589457 132910 592572 132912
rect 675477 132968 676292 132970
rect 675477 132912 675482 132968
rect 675538 132912 676292 132968
rect 675477 132910 676292 132912
rect 589457 132907 589523 132910
rect 675477 132907 675543 132910
rect 675477 132562 675543 132565
rect 675477 132560 676292 132562
rect 675477 132504 675482 132560
rect 675538 132504 676292 132560
rect 675477 132502 676292 132504
rect 675477 132499 675543 132502
rect 675293 132154 675359 132157
rect 675293 132152 676292 132154
rect 675293 132096 675298 132152
rect 675354 132096 676292 132152
rect 675293 132094 676292 132096
rect 675293 132091 675359 132094
rect 675477 131746 675543 131749
rect 675477 131744 676292 131746
rect 675477 131688 675482 131744
rect 675538 131688 676292 131744
rect 675477 131686 676292 131688
rect 675477 131683 675543 131686
rect 588905 131338 588971 131341
rect 674649 131338 674715 131341
rect 588905 131336 592572 131338
rect 588905 131280 588910 131336
rect 588966 131280 592572 131336
rect 588905 131278 592572 131280
rect 674649 131336 676292 131338
rect 674649 131280 674654 131336
rect 674710 131280 676292 131336
rect 674649 131278 676292 131280
rect 588905 131275 588971 131278
rect 674649 131275 674715 131278
rect 675477 130930 675543 130933
rect 675477 130928 676292 130930
rect 675477 130872 675482 130928
rect 675538 130872 676292 130928
rect 675477 130870 676292 130872
rect 675477 130867 675543 130870
rect 579061 130658 579127 130661
rect 667933 130658 667999 130661
rect 575798 130656 579127 130658
rect 575798 130600 579066 130656
rect 579122 130600 579127 130656
rect 575798 130598 579127 130600
rect 575798 130084 575858 130598
rect 579061 130595 579127 130598
rect 666694 130656 667999 130658
rect 666694 130600 667938 130656
rect 667994 130600 667999 130656
rect 666694 130598 667999 130600
rect 666694 130590 666754 130598
rect 667933 130595 667999 130598
rect 666356 130530 666754 130590
rect 675477 130522 675543 130525
rect 675477 130520 676292 130522
rect 675477 130464 675482 130520
rect 675538 130464 676292 130520
rect 675477 130462 676292 130464
rect 675477 130459 675543 130462
rect 675477 130114 675543 130117
rect 675477 130112 676292 130114
rect 675477 130056 675482 130112
rect 675538 130056 676292 130112
rect 675477 130054 676292 130056
rect 675477 130051 675543 130054
rect 589457 129706 589523 129709
rect 674465 129706 674531 129709
rect 589457 129704 592572 129706
rect 589457 129648 589462 129704
rect 589518 129648 592572 129704
rect 589457 129646 592572 129648
rect 674465 129704 676292 129706
rect 674465 129648 674470 129704
rect 674526 129648 676292 129704
rect 674465 129646 676292 129648
rect 589457 129643 589523 129646
rect 674465 129643 674531 129646
rect 675477 129298 675543 129301
rect 675477 129296 676292 129298
rect 675477 129240 675482 129296
rect 675538 129240 676292 129296
rect 675477 129238 676292 129240
rect 675477 129235 675543 129238
rect 669221 129026 669287 129029
rect 666694 129024 669287 129026
rect 666694 128968 669226 129024
rect 669282 128968 669287 129024
rect 666694 128966 669287 128968
rect 666694 128958 666754 128966
rect 669221 128963 669287 128966
rect 666356 128898 666754 128958
rect 676262 128620 676322 128860
rect 676254 128556 676260 128620
rect 676324 128556 676330 128620
rect 676070 128148 676076 128212
rect 676140 128210 676146 128212
rect 676262 128210 676322 128452
rect 676140 128150 676322 128210
rect 676140 128148 676146 128150
rect 590101 128074 590167 128077
rect 590101 128072 592572 128074
rect 590101 128016 590106 128072
rect 590162 128016 592572 128072
rect 590101 128014 592572 128016
rect 590101 128011 590167 128014
rect 579521 127938 579587 127941
rect 575798 127936 579587 127938
rect 575798 127880 579526 127936
rect 579582 127880 579587 127936
rect 575798 127878 579587 127880
rect 575798 127636 575858 127878
rect 579521 127875 579587 127878
rect 679574 127805 679634 128044
rect 679574 127800 679683 127805
rect 679574 127744 679622 127800
rect 679678 127744 679683 127800
rect 679574 127742 679683 127744
rect 679617 127739 679683 127742
rect 674833 127666 674899 127669
rect 674833 127664 676292 127666
rect 674833 127608 674838 127664
rect 674894 127608 676292 127664
rect 674833 127606 676292 127608
rect 674833 127603 674899 127606
rect 675886 127196 675892 127260
rect 675956 127258 675962 127260
rect 675956 127198 676292 127258
rect 675956 127196 675962 127198
rect 683070 126581 683130 126820
rect 683070 126576 683179 126581
rect 683070 126520 683118 126576
rect 683174 126520 683179 126576
rect 683070 126518 683179 126520
rect 683113 126515 683179 126518
rect 589273 126442 589339 126445
rect 675017 126442 675083 126445
rect 589273 126440 592572 126442
rect 589273 126384 589278 126440
rect 589334 126384 592572 126440
rect 589273 126382 592572 126384
rect 675017 126440 676292 126442
rect 675017 126384 675022 126440
rect 675078 126384 676292 126440
rect 675017 126382 676292 126384
rect 589273 126379 589339 126382
rect 675017 126379 675083 126382
rect 675477 126034 675543 126037
rect 675477 126032 676292 126034
rect 675477 125976 675482 126032
rect 675538 125976 676292 126032
rect 675477 125974 676292 125976
rect 675477 125971 675543 125974
rect 667933 125762 667999 125765
rect 666694 125760 667999 125762
rect 666694 125704 667938 125760
rect 667994 125704 667999 125760
rect 666694 125702 667999 125704
rect 666694 125694 666754 125702
rect 667933 125699 667999 125702
rect 666356 125634 666754 125694
rect 675477 125626 675543 125629
rect 675477 125624 676292 125626
rect 675477 125568 675482 125624
rect 675538 125568 676292 125624
rect 675477 125566 676292 125568
rect 675477 125563 675543 125566
rect 578877 125354 578943 125357
rect 575798 125352 578943 125354
rect 575798 125296 578882 125352
rect 578938 125296 578943 125352
rect 575798 125294 578943 125296
rect 575798 125188 575858 125294
rect 578877 125291 578943 125294
rect 674373 125218 674439 125221
rect 674373 125216 676292 125218
rect 674373 125160 674378 125216
rect 674434 125160 676292 125216
rect 674373 125158 676292 125160
rect 674373 125155 674439 125158
rect 588721 124810 588787 124813
rect 675477 124810 675543 124813
rect 588721 124808 592572 124810
rect 588721 124752 588726 124808
rect 588782 124752 592572 124808
rect 588721 124750 592572 124752
rect 675477 124808 676292 124810
rect 675477 124752 675482 124808
rect 675538 124752 676292 124808
rect 675477 124750 676292 124752
rect 588721 124747 588787 124750
rect 675477 124747 675543 124750
rect 676806 124476 676812 124540
rect 676876 124538 676882 124540
rect 683113 124538 683179 124541
rect 676876 124536 683179 124538
rect 676876 124480 683118 124536
rect 683174 124480 683179 124536
rect 676876 124478 683179 124480
rect 676876 124476 676882 124478
rect 683113 124475 683179 124478
rect 683070 124133 683130 124372
rect 669221 124130 669287 124133
rect 666694 124128 669287 124130
rect 666694 124072 669226 124128
rect 669282 124072 669287 124128
rect 666694 124070 669287 124072
rect 683070 124128 683179 124133
rect 683070 124072 683118 124128
rect 683174 124072 683179 124128
rect 683070 124070 683179 124072
rect 666694 124062 666754 124070
rect 669221 124067 669287 124070
rect 683113 124067 683179 124070
rect 666356 124002 666754 124062
rect 675293 123994 675359 123997
rect 675293 123992 676292 123994
rect 675293 123936 675298 123992
rect 675354 123936 676292 123992
rect 675293 123934 676292 123936
rect 675293 123931 675359 123934
rect 674649 123586 674715 123589
rect 674649 123584 676292 123586
rect 674649 123528 674654 123584
rect 674710 123528 676292 123584
rect 674649 123526 676292 123528
rect 674649 123523 674715 123526
rect 590285 123178 590351 123181
rect 675477 123178 675543 123181
rect 590285 123176 592572 123178
rect 590285 123120 590290 123176
rect 590346 123120 592572 123176
rect 590285 123118 592572 123120
rect 675477 123176 676292 123178
rect 675477 123120 675482 123176
rect 675538 123120 676292 123176
rect 675477 123118 676292 123120
rect 590285 123115 590351 123118
rect 675477 123115 675543 123118
rect 575982 122634 576042 122740
rect 578877 122634 578943 122637
rect 575982 122632 578943 122634
rect 575982 122576 578882 122632
rect 578938 122576 578943 122632
rect 575982 122574 578943 122576
rect 578877 122571 578943 122574
rect 675293 122498 675359 122501
rect 676262 122498 676322 122740
rect 675293 122496 676322 122498
rect 675293 122440 675298 122496
rect 675354 122440 676322 122496
rect 675293 122438 676322 122440
rect 675293 122435 675359 122438
rect 677550 122093 677610 122332
rect 677550 122088 677659 122093
rect 677550 122032 677598 122088
rect 677654 122032 677659 122088
rect 677550 122030 677659 122032
rect 677593 122027 677659 122030
rect 675477 121954 675543 121957
rect 675477 121952 676292 121954
rect 675477 121896 675482 121952
rect 675538 121896 676292 121952
rect 675477 121894 676292 121896
rect 675477 121891 675543 121894
rect 589457 121546 589523 121549
rect 589457 121544 592572 121546
rect 589457 121488 589462 121544
rect 589518 121488 592572 121544
rect 589457 121486 592572 121488
rect 589457 121483 589523 121486
rect 578417 120866 578483 120869
rect 668209 120866 668275 120869
rect 575798 120864 578483 120866
rect 575798 120808 578422 120864
rect 578478 120808 578483 120864
rect 575798 120806 578483 120808
rect 575798 120292 575858 120806
rect 578417 120803 578483 120806
rect 666694 120864 668275 120866
rect 666694 120808 668214 120864
rect 668270 120808 668275 120864
rect 666694 120806 668275 120808
rect 666694 120798 666754 120806
rect 668209 120803 668275 120806
rect 666356 120738 666754 120798
rect 589457 119914 589523 119917
rect 589457 119912 592572 119914
rect 589457 119856 589462 119912
rect 589518 119856 592572 119912
rect 589457 119854 592572 119856
rect 589457 119851 589523 119854
rect 669129 119234 669195 119237
rect 666694 119232 669195 119234
rect 666694 119176 669134 119232
rect 669190 119176 669195 119232
rect 666694 119174 669195 119176
rect 666694 119166 666754 119174
rect 669129 119171 669195 119174
rect 666356 119106 666754 119166
rect 578509 118282 578575 118285
rect 575798 118280 578575 118282
rect 575798 118224 578514 118280
rect 578570 118224 578575 118280
rect 575798 118222 578575 118224
rect 575798 117844 575858 118222
rect 578509 118219 578575 118222
rect 589457 118282 589523 118285
rect 589457 118280 592572 118282
rect 589457 118224 589462 118280
rect 589518 118224 592572 118280
rect 589457 118222 592572 118224
rect 589457 118219 589523 118222
rect 667933 117602 667999 117605
rect 666694 117600 667999 117602
rect 666694 117544 667938 117600
rect 667994 117544 667999 117600
rect 666694 117542 667999 117544
rect 666694 117534 666754 117542
rect 667933 117539 667999 117542
rect 666356 117474 666754 117534
rect 676990 117268 676996 117332
rect 677060 117330 677066 117332
rect 683113 117330 683179 117333
rect 677060 117328 683179 117330
rect 677060 117272 683118 117328
rect 683174 117272 683179 117328
rect 677060 117270 683179 117272
rect 677060 117268 677066 117270
rect 683113 117267 683179 117270
rect 675702 116996 675708 117060
rect 675772 117058 675778 117060
rect 677593 117058 677659 117061
rect 675772 117056 677659 117058
rect 675772 117000 677598 117056
rect 677654 117000 677659 117056
rect 675772 116998 677659 117000
rect 675772 116996 675778 116998
rect 677593 116995 677659 116998
rect 589457 116650 589523 116653
rect 589457 116648 592572 116650
rect 589457 116592 589462 116648
rect 589518 116592 592572 116648
rect 589457 116590 592572 116592
rect 589457 116587 589523 116590
rect 666356 115842 666754 115902
rect 666694 115834 666754 115842
rect 668393 115834 668459 115837
rect 666694 115832 668459 115834
rect 666694 115776 668398 115832
rect 668454 115776 668459 115832
rect 666694 115774 668459 115776
rect 668393 115771 668459 115774
rect 579245 115698 579311 115701
rect 575798 115696 579311 115698
rect 575798 115640 579250 115696
rect 579306 115640 579311 115696
rect 575798 115638 579311 115640
rect 575798 115396 575858 115638
rect 579245 115635 579311 115638
rect 589917 115018 589983 115021
rect 589917 115016 592572 115018
rect 589917 114960 589922 115016
rect 589978 114960 592572 115016
rect 589917 114958 592572 114960
rect 589917 114955 589983 114958
rect 668393 114338 668459 114341
rect 666694 114336 668459 114338
rect 666694 114280 668398 114336
rect 668454 114280 668459 114336
rect 666694 114278 668459 114280
rect 666694 114270 666754 114278
rect 668393 114275 668459 114278
rect 666356 114210 666754 114270
rect 589457 113386 589523 113389
rect 589457 113384 592572 113386
rect 589457 113328 589462 113384
rect 589518 113328 592572 113384
rect 589457 113326 592572 113328
rect 589457 113323 589523 113326
rect 579521 113114 579587 113117
rect 575798 113112 579587 113114
rect 575798 113056 579526 113112
rect 579582 113056 579587 113112
rect 575798 113054 579587 113056
rect 575798 112948 575858 113054
rect 579521 113051 579587 113054
rect 675293 113114 675359 113117
rect 676254 113114 676260 113116
rect 675293 113112 676260 113114
rect 675293 113056 675298 113112
rect 675354 113056 676260 113112
rect 675293 113054 676260 113056
rect 675293 113051 675359 113054
rect 676254 113052 676260 113054
rect 676324 113052 676330 113116
rect 668025 112706 668091 112709
rect 666694 112704 668091 112706
rect 666694 112648 668030 112704
rect 668086 112648 668091 112704
rect 666694 112646 668091 112648
rect 666694 112638 666754 112646
rect 668025 112643 668091 112646
rect 666356 112578 666754 112638
rect 589641 111754 589707 111757
rect 589641 111752 592572 111754
rect 589641 111696 589646 111752
rect 589702 111696 592572 111752
rect 589641 111694 592572 111696
rect 589641 111691 589707 111694
rect 579521 111074 579587 111077
rect 668761 111074 668827 111077
rect 575798 111072 579587 111074
rect 575798 111016 579526 111072
rect 579582 111016 579587 111072
rect 575798 111014 579587 111016
rect 575798 110500 575858 111014
rect 579521 111011 579587 111014
rect 666694 111072 668827 111074
rect 666694 111016 668766 111072
rect 668822 111016 668827 111072
rect 666694 111014 668827 111016
rect 666694 111006 666754 111014
rect 668761 111011 668827 111014
rect 666356 110946 666754 111006
rect 675753 110394 675819 110397
rect 676990 110394 676996 110396
rect 675753 110392 676996 110394
rect 675753 110336 675758 110392
rect 675814 110336 676996 110392
rect 675753 110334 676996 110336
rect 675753 110331 675819 110334
rect 676990 110332 676996 110334
rect 677060 110332 677066 110396
rect 589457 110122 589523 110125
rect 589457 110120 592572 110122
rect 589457 110064 589462 110120
rect 589518 110064 592572 110120
rect 589457 110062 592572 110064
rect 589457 110059 589523 110062
rect 666737 109374 666803 109377
rect 666356 109372 666803 109374
rect 666356 109316 666742 109372
rect 666798 109316 666803 109372
rect 666356 109314 666803 109316
rect 666737 109311 666803 109314
rect 579245 108490 579311 108493
rect 575798 108488 579311 108490
rect 575798 108432 579250 108488
rect 579306 108432 579311 108488
rect 575798 108430 579311 108432
rect 575798 108052 575858 108430
rect 579245 108427 579311 108430
rect 589457 108490 589523 108493
rect 589457 108488 592572 108490
rect 589457 108432 589462 108488
rect 589518 108432 592572 108488
rect 589457 108430 592572 108432
rect 589457 108427 589523 108430
rect 675661 108082 675727 108085
rect 675886 108082 675892 108084
rect 675661 108080 675892 108082
rect 675661 108024 675666 108080
rect 675722 108024 675892 108080
rect 675661 108022 675892 108024
rect 675661 108019 675727 108022
rect 675886 108020 675892 108022
rect 675956 108020 675962 108084
rect 666356 107682 666754 107742
rect 666694 107674 666754 107682
rect 669221 107674 669287 107677
rect 666694 107672 669287 107674
rect 666694 107616 669226 107672
rect 669282 107616 669287 107672
rect 666694 107614 669287 107616
rect 669221 107611 669287 107614
rect 589457 106858 589523 106861
rect 589457 106856 592572 106858
rect 589457 106800 589462 106856
rect 589518 106800 592572 106856
rect 589457 106798 592572 106800
rect 589457 106795 589523 106798
rect 673361 106314 673427 106317
rect 675109 106314 675175 106317
rect 673361 106312 675175 106314
rect 673361 106256 673366 106312
rect 673422 106256 675114 106312
rect 675170 106256 675175 106312
rect 673361 106254 675175 106256
rect 673361 106251 673427 106254
rect 675109 106251 675175 106254
rect 666356 106050 666754 106110
rect 666694 106042 666754 106050
rect 668945 106042 669011 106045
rect 666694 106040 669011 106042
rect 666694 105984 668950 106040
rect 669006 105984 669011 106040
rect 666694 105982 669011 105984
rect 668945 105979 669011 105982
rect 578325 105906 578391 105909
rect 575798 105904 578391 105906
rect 575798 105848 578330 105904
rect 578386 105848 578391 105904
rect 575798 105846 578391 105848
rect 575798 105604 575858 105846
rect 578325 105843 578391 105846
rect 589457 105226 589523 105229
rect 589457 105224 592572 105226
rect 589457 105168 589462 105224
rect 589518 105168 592572 105224
rect 589457 105166 592572 105168
rect 589457 105163 589523 105166
rect 669129 104546 669195 104549
rect 666694 104544 669195 104546
rect 666694 104488 669134 104544
rect 669190 104488 669195 104544
rect 666694 104486 669195 104488
rect 666694 104478 666754 104486
rect 669129 104483 669195 104486
rect 666356 104418 666754 104478
rect 589457 103594 589523 103597
rect 589457 103592 592572 103594
rect 589457 103536 589462 103592
rect 589518 103536 592572 103592
rect 589457 103534 592572 103536
rect 589457 103531 589523 103534
rect 579521 103458 579587 103461
rect 575798 103456 579587 103458
rect 575798 103400 579526 103456
rect 579582 103400 579587 103456
rect 575798 103398 579587 103400
rect 575798 103156 575858 103398
rect 579521 103395 579587 103398
rect 675753 103186 675819 103189
rect 676070 103186 676076 103188
rect 675753 103184 676076 103186
rect 675753 103128 675758 103184
rect 675814 103128 676076 103184
rect 675753 103126 676076 103128
rect 675753 103123 675819 103126
rect 676070 103124 676076 103126
rect 676140 103124 676146 103188
rect 668577 102914 668643 102917
rect 666694 102912 668643 102914
rect 666694 102856 668582 102912
rect 668638 102856 668643 102912
rect 666694 102854 668643 102856
rect 666694 102846 666754 102854
rect 668577 102851 668643 102854
rect 666356 102786 666754 102846
rect 675661 102644 675727 102645
rect 675661 102640 675708 102644
rect 675772 102642 675778 102644
rect 675661 102584 675666 102640
rect 675661 102580 675708 102584
rect 675772 102582 675818 102642
rect 675772 102580 675778 102582
rect 675661 102579 675727 102580
rect 589365 101962 589431 101965
rect 589365 101960 592572 101962
rect 589365 101904 589370 101960
rect 589426 101904 592572 101960
rect 589365 101902 592572 101904
rect 589365 101899 589431 101902
rect 675753 101418 675819 101421
rect 676806 101418 676812 101420
rect 675753 101416 676812 101418
rect 675753 101360 675758 101416
rect 675814 101360 676812 101416
rect 675753 101358 676812 101360
rect 675753 101355 675819 101358
rect 676806 101356 676812 101358
rect 676876 101356 676882 101420
rect 575982 100602 576042 100708
rect 579245 100602 579311 100605
rect 575982 100600 579311 100602
rect 575982 100544 579250 100600
rect 579306 100544 579311 100600
rect 575982 100542 579311 100544
rect 579245 100539 579311 100542
rect 579521 98834 579587 98837
rect 575798 98832 579587 98834
rect 575798 98776 579526 98832
rect 579582 98776 579587 98832
rect 575798 98774 579587 98776
rect 575798 98260 575858 98774
rect 579521 98771 579587 98774
rect 637021 96930 637087 96933
rect 637246 96930 637252 96932
rect 637021 96928 637252 96930
rect 637021 96872 637026 96928
rect 637082 96872 637252 96928
rect 637021 96870 637252 96872
rect 637021 96867 637087 96870
rect 637246 96868 637252 96870
rect 637316 96868 637322 96932
rect 578601 96250 578667 96253
rect 575798 96248 578667 96250
rect 575798 96192 578606 96248
rect 578662 96192 578667 96248
rect 575798 96190 578667 96192
rect 575798 95812 575858 96190
rect 578601 96187 578667 96190
rect 634670 95644 634676 95708
rect 634740 95706 634746 95708
rect 635917 95706 635983 95709
rect 634740 95704 635983 95706
rect 634740 95648 635922 95704
rect 635978 95648 635983 95704
rect 634740 95646 635983 95648
rect 634740 95644 634746 95646
rect 635917 95643 635983 95646
rect 626441 95434 626507 95437
rect 626441 95432 628268 95434
rect 626441 95376 626446 95432
rect 626502 95376 628268 95432
rect 626441 95374 628268 95376
rect 626441 95371 626507 95374
rect 642633 95162 642699 95165
rect 642590 95160 642699 95162
rect 642590 95104 642638 95160
rect 642694 95104 642699 95160
rect 642590 95099 642699 95104
rect 642590 94588 642650 95099
rect 626073 94482 626139 94485
rect 626073 94480 628268 94482
rect 626073 94424 626078 94480
rect 626134 94424 628268 94480
rect 626073 94422 628268 94424
rect 626073 94419 626139 94422
rect 653949 94210 654015 94213
rect 653949 94208 656788 94210
rect 653949 94152 653954 94208
rect 654010 94152 656788 94208
rect 653949 94150 656788 94152
rect 653949 94147 654015 94150
rect 579521 93666 579587 93669
rect 575798 93664 579587 93666
rect 575798 93608 579526 93664
rect 579582 93608 579587 93664
rect 575798 93606 579587 93608
rect 575798 93364 575858 93606
rect 579521 93603 579587 93606
rect 626441 93530 626507 93533
rect 626441 93528 628268 93530
rect 626441 93472 626446 93528
rect 626502 93472 628268 93528
rect 626441 93470 628268 93472
rect 626441 93467 626507 93470
rect 654317 93394 654383 93397
rect 665725 93394 665791 93397
rect 654317 93392 656788 93394
rect 654317 93336 654322 93392
rect 654378 93336 656788 93392
rect 654317 93334 656788 93336
rect 663596 93392 665791 93394
rect 663596 93336 665730 93392
rect 665786 93336 665791 93392
rect 663596 93334 665791 93336
rect 654317 93331 654383 93334
rect 665725 93331 665791 93334
rect 663241 93122 663307 93125
rect 663198 93120 663307 93122
rect 663198 93064 663246 93120
rect 663302 93064 663307 93120
rect 663198 93059 663307 93064
rect 626257 92578 626323 92581
rect 654133 92578 654199 92581
rect 626257 92576 628268 92578
rect 626257 92520 626262 92576
rect 626318 92520 628268 92576
rect 626257 92518 628268 92520
rect 654133 92576 656788 92578
rect 654133 92520 654138 92576
rect 654194 92520 656788 92576
rect 663198 92548 663258 93059
rect 654133 92518 656788 92520
rect 626257 92515 626323 92518
rect 654133 92515 654199 92518
rect 644473 92170 644539 92173
rect 642988 92168 644539 92170
rect 642988 92112 644478 92168
rect 644534 92112 644539 92168
rect 642988 92110 644539 92112
rect 644473 92107 644539 92110
rect 665173 91762 665239 91765
rect 663596 91760 665239 91762
rect 663596 91704 665178 91760
rect 665234 91704 665239 91760
rect 663596 91702 665239 91704
rect 665173 91699 665239 91702
rect 625429 91626 625495 91629
rect 625429 91624 628268 91626
rect 625429 91568 625434 91624
rect 625490 91568 628268 91624
rect 625429 91566 628268 91568
rect 625429 91563 625495 91566
rect 654317 91490 654383 91493
rect 654317 91488 656788 91490
rect 654317 91432 654322 91488
rect 654378 91432 656788 91488
rect 654317 91430 656788 91432
rect 654317 91427 654383 91430
rect 579521 91082 579587 91085
rect 575798 91080 579587 91082
rect 575798 91024 579526 91080
rect 579582 91024 579587 91080
rect 575798 91022 579587 91024
rect 575798 90916 575858 91022
rect 579521 91019 579587 91022
rect 626441 90674 626507 90677
rect 654133 90674 654199 90677
rect 665357 90674 665423 90677
rect 626441 90672 628268 90674
rect 626441 90616 626446 90672
rect 626502 90616 628268 90672
rect 626441 90614 628268 90616
rect 654133 90672 656788 90674
rect 654133 90616 654138 90672
rect 654194 90616 656788 90672
rect 654133 90614 656788 90616
rect 663596 90672 665423 90674
rect 663596 90616 665362 90672
rect 665418 90616 665423 90672
rect 663596 90614 665423 90616
rect 626441 90611 626507 90614
rect 654133 90611 654199 90614
rect 665357 90611 665423 90614
rect 663793 90402 663859 90405
rect 663566 90400 663859 90402
rect 663566 90344 663798 90400
rect 663854 90344 663859 90400
rect 663566 90342 663859 90344
rect 655789 89858 655855 89861
rect 655789 89856 656788 89858
rect 655789 89800 655794 89856
rect 655850 89800 656788 89856
rect 663566 89828 663626 90342
rect 663793 90339 663859 90342
rect 655789 89798 656788 89800
rect 655789 89795 655855 89798
rect 626441 89722 626507 89725
rect 644749 89722 644815 89725
rect 626441 89720 628268 89722
rect 626441 89664 626446 89720
rect 626502 89664 628268 89720
rect 626441 89662 628268 89664
rect 642988 89720 644815 89722
rect 642988 89664 644754 89720
rect 644810 89664 644815 89720
rect 642988 89662 644815 89664
rect 626441 89659 626507 89662
rect 644749 89659 644815 89662
rect 578509 89042 578575 89045
rect 663977 89042 664043 89045
rect 575798 89040 578575 89042
rect 575798 88984 578514 89040
rect 578570 88984 578575 89040
rect 575798 88982 578575 88984
rect 663596 89040 664043 89042
rect 663596 88984 663982 89040
rect 664038 88984 664043 89040
rect 663596 88982 664043 88984
rect 575798 88468 575858 88982
rect 578509 88979 578575 88982
rect 663977 88979 664043 88982
rect 624969 88634 625035 88637
rect 628238 88634 628298 88876
rect 624969 88632 628298 88634
rect 624969 88576 624974 88632
rect 625030 88576 628298 88632
rect 624969 88574 628298 88576
rect 624969 88571 625035 88574
rect 626441 87954 626507 87957
rect 626441 87952 628268 87954
rect 626441 87896 626446 87952
rect 626502 87896 628268 87952
rect 626441 87894 628268 87896
rect 626441 87891 626507 87894
rect 643921 87138 643987 87141
rect 642988 87136 643987 87138
rect 642988 87080 643926 87136
rect 643982 87080 643987 87136
rect 642988 87078 643987 87080
rect 643921 87075 643987 87078
rect 625613 87002 625679 87005
rect 625613 87000 628268 87002
rect 625613 86944 625618 87000
rect 625674 86944 628268 87000
rect 625613 86942 628268 86944
rect 625613 86939 625679 86942
rect 579521 86458 579587 86461
rect 575798 86456 579587 86458
rect 575798 86400 579526 86456
rect 579582 86400 579587 86456
rect 575798 86398 579587 86400
rect 575798 86020 575858 86398
rect 579521 86395 579587 86398
rect 626441 86050 626507 86053
rect 626441 86048 628268 86050
rect 626441 85992 626446 86048
rect 626502 85992 628268 86048
rect 626441 85990 628268 85992
rect 626441 85987 626507 85990
rect 626441 85098 626507 85101
rect 626441 85096 628268 85098
rect 626441 85040 626446 85096
rect 626502 85040 628268 85096
rect 626441 85038 628268 85040
rect 626441 85035 626507 85038
rect 643461 84690 643527 84693
rect 642988 84688 643527 84690
rect 642988 84632 643466 84688
rect 643522 84632 643527 84688
rect 642988 84630 643527 84632
rect 643461 84627 643527 84630
rect 626441 84146 626507 84149
rect 626441 84144 628268 84146
rect 626441 84088 626446 84144
rect 626502 84088 628268 84144
rect 626441 84086 628268 84088
rect 626441 84083 626507 84086
rect 579337 83874 579403 83877
rect 575798 83872 579403 83874
rect 575798 83816 579342 83872
rect 579398 83816 579403 83872
rect 575798 83814 579403 83816
rect 575798 83572 575858 83814
rect 579337 83811 579403 83814
rect 626257 83194 626323 83197
rect 626257 83192 628268 83194
rect 626257 83136 626262 83192
rect 626318 83136 628268 83192
rect 626257 83134 628268 83136
rect 626257 83131 626323 83134
rect 643093 82786 643159 82789
rect 642774 82784 643159 82786
rect 642774 82728 643098 82784
rect 643154 82728 643159 82784
rect 642774 82726 643159 82728
rect 642774 82212 642834 82726
rect 643093 82723 643159 82726
rect 628606 81701 628666 82212
rect 628557 81696 628666 81701
rect 628557 81640 628562 81696
rect 628618 81640 628666 81696
rect 628557 81638 628666 81640
rect 628557 81635 628623 81638
rect 579521 81426 579587 81429
rect 575798 81424 579587 81426
rect 575798 81368 579526 81424
rect 579582 81368 579587 81424
rect 575798 81366 579587 81368
rect 575798 81124 575858 81366
rect 579521 81363 579587 81366
rect 628790 80882 628850 81396
rect 629201 80882 629267 80885
rect 628790 80880 629267 80882
rect 628790 80824 629206 80880
rect 629262 80824 629267 80880
rect 628790 80822 629267 80824
rect 629201 80819 629267 80822
rect 579061 79250 579127 79253
rect 575798 79248 579127 79250
rect 575798 79192 579066 79248
rect 579122 79192 579127 79248
rect 575798 79190 579127 79192
rect 575798 78676 575858 79190
rect 579061 79187 579127 79190
rect 637113 78572 637179 78573
rect 637062 78570 637068 78572
rect 637022 78510 637068 78570
rect 637132 78568 637179 78572
rect 637174 78512 637179 78568
rect 637062 78508 637068 78510
rect 637132 78508 637179 78512
rect 637113 78507 637179 78508
rect 633893 77754 633959 77757
rect 634670 77754 634676 77756
rect 633893 77752 634676 77754
rect 633893 77696 633898 77752
rect 633954 77696 634676 77752
rect 633893 77694 634676 77696
rect 633893 77691 633959 77694
rect 634670 77692 634676 77694
rect 634740 77692 634746 77756
rect 578877 76802 578943 76805
rect 575798 76800 578943 76802
rect 575798 76744 578882 76800
rect 578938 76744 578943 76800
rect 575798 76742 578943 76744
rect 575798 76228 575858 76742
rect 578877 76739 578943 76742
rect 646865 74490 646931 74493
rect 646668 74488 646931 74490
rect 646668 74432 646870 74488
rect 646926 74432 646931 74488
rect 646668 74430 646931 74432
rect 646865 74427 646931 74430
rect 579521 74218 579587 74221
rect 575798 74216 579587 74218
rect 575798 74160 579526 74216
rect 579582 74160 579587 74216
rect 575798 74158 579587 74160
rect 575798 73780 575858 74158
rect 579521 74155 579587 74158
rect 647417 72994 647483 72997
rect 646668 72992 647483 72994
rect 646668 72936 647422 72992
rect 647478 72936 647483 72992
rect 646668 72934 647483 72936
rect 647417 72931 647483 72934
rect 646129 71770 646195 71773
rect 646086 71768 646195 71770
rect 646086 71712 646134 71768
rect 646190 71712 646195 71768
rect 646086 71707 646195 71712
rect 579521 71498 579587 71501
rect 575798 71496 579587 71498
rect 575798 71440 579526 71496
rect 579582 71440 579587 71496
rect 646086 71468 646146 71707
rect 575798 71438 579587 71440
rect 575798 71332 575858 71438
rect 579521 71435 579587 71438
rect 646313 70410 646379 70413
rect 646270 70408 646379 70410
rect 646270 70352 646318 70408
rect 646374 70352 646379 70408
rect 646270 70347 646379 70352
rect 646270 69972 646330 70347
rect 575982 68778 576042 68884
rect 578509 68778 578575 68781
rect 575982 68776 578575 68778
rect 575982 68720 578514 68776
rect 578570 68720 578575 68776
rect 575982 68718 578575 68720
rect 578509 68715 578575 68718
rect 647601 68506 647667 68509
rect 646668 68504 647667 68506
rect 646668 68448 647606 68504
rect 647662 68448 647667 68504
rect 646668 68446 647667 68448
rect 647601 68443 647667 68446
rect 579521 67010 579587 67013
rect 648981 67010 649047 67013
rect 575798 67008 579587 67010
rect 575798 66952 579526 67008
rect 579582 66952 579587 67008
rect 575798 66950 579587 66952
rect 646668 67008 649047 67010
rect 646668 66952 648986 67008
rect 649042 66952 649047 67008
rect 646668 66950 649047 66952
rect 575798 66436 575858 66950
rect 579521 66947 579587 66950
rect 648981 66947 649047 66950
rect 646129 66058 646195 66061
rect 646086 66056 646195 66058
rect 646086 66000 646134 66056
rect 646190 66000 646195 66056
rect 646086 65995 646195 66000
rect 646086 65484 646146 65995
rect 579245 64562 579311 64565
rect 575798 64560 579311 64562
rect 575798 64504 579250 64560
rect 579306 64504 579311 64560
rect 575798 64502 579311 64504
rect 575798 63988 575858 64502
rect 579245 64499 579311 64502
rect 648797 64018 648863 64021
rect 646668 64016 648863 64018
rect 646668 63960 648802 64016
rect 648858 63960 648863 64016
rect 646668 63958 648863 63960
rect 648797 63955 648863 63958
rect 578509 61842 578575 61845
rect 575798 61840 578575 61842
rect 575798 61784 578514 61840
rect 578570 61784 578575 61840
rect 575798 61782 578575 61784
rect 575798 61540 575858 61782
rect 578509 61779 578575 61782
rect 575982 58986 576042 59092
rect 579521 58986 579587 58989
rect 575982 58984 579587 58986
rect 575982 58928 579526 58984
rect 579582 58928 579587 58984
rect 575982 58926 579587 58928
rect 579521 58923 579587 58926
rect 579061 57218 579127 57221
rect 575798 57216 579127 57218
rect 575798 57160 579066 57216
rect 579122 57160 579127 57216
rect 575798 57158 579127 57160
rect 575798 56644 575858 57158
rect 579061 57155 579127 57158
rect 578509 54770 578575 54773
rect 575798 54768 578575 54770
rect 575798 54712 578514 54768
rect 578570 54712 578575 54768
rect 575798 54710 578575 54712
rect 575798 54196 575858 54710
rect 578509 54707 578575 54710
rect 409638 53076 409644 53140
rect 409708 53138 409714 53140
rect 591297 53138 591363 53141
rect 409708 53136 591363 53138
rect 409708 53080 591302 53136
rect 591358 53080 591363 53136
rect 409708 53078 591363 53080
rect 409708 53076 409714 53078
rect 591297 53075 591363 53078
rect 464838 51716 464844 51780
rect 464908 51778 464914 51780
rect 603073 51778 603139 51781
rect 464908 51776 603139 51778
rect 464908 51720 603078 51776
rect 603134 51720 603139 51776
rect 464908 51718 603139 51720
rect 464908 51716 464914 51718
rect 603073 51715 603139 51718
rect 497549 50554 497615 50557
rect 525742 50554 525748 50556
rect 497549 50552 525748 50554
rect 497549 50496 497554 50552
rect 497610 50496 525748 50552
rect 497549 50494 525748 50496
rect 497549 50491 497615 50494
rect 525742 50492 525748 50494
rect 525812 50492 525818 50556
rect 529790 50492 529796 50556
rect 529860 50554 529866 50556
rect 549253 50554 549319 50557
rect 529860 50552 549319 50554
rect 529860 50496 549258 50552
rect 549314 50496 549319 50552
rect 529860 50494 549319 50496
rect 529860 50492 529866 50494
rect 549253 50491 549319 50494
rect 78581 50282 78647 50285
rect 147622 50282 147628 50284
rect 78581 50280 147628 50282
rect 78581 50224 78586 50280
rect 78642 50224 147628 50280
rect 78581 50222 147628 50224
rect 78581 50219 78647 50222
rect 147622 50220 147628 50222
rect 147692 50220 147698 50284
rect 460790 50220 460796 50284
rect 460860 50282 460866 50284
rect 601877 50282 601943 50285
rect 460860 50280 601943 50282
rect 460860 50224 601882 50280
rect 601938 50224 601943 50280
rect 460860 50222 601943 50224
rect 460860 50220 460866 50222
rect 601877 50219 601943 50222
rect 131021 49740 131087 49741
rect 131021 49736 131068 49740
rect 131132 49738 131138 49740
rect 131021 49680 131026 49736
rect 131021 49676 131068 49680
rect 131132 49678 131178 49738
rect 131132 49676 131138 49678
rect 131021 49675 131087 49676
rect 411110 49132 411116 49196
rect 411180 49194 411186 49196
rect 600313 49194 600379 49197
rect 411180 49192 600379 49194
rect 411180 49136 600318 49192
rect 600374 49136 600379 49192
rect 411180 49134 600379 49136
rect 411180 49132 411186 49134
rect 600313 49131 600379 49134
rect 365478 48860 365484 48924
rect 365548 48922 365554 48924
rect 596173 48922 596239 48925
rect 365548 48920 596239 48922
rect 365548 48864 596178 48920
rect 596234 48864 596239 48920
rect 365548 48862 596239 48864
rect 365548 48860 365554 48862
rect 596173 48859 596239 48862
rect 663793 48514 663859 48517
rect 662094 48512 663859 48514
rect 661480 48456 663798 48512
rect 663854 48456 663859 48512
rect 661480 48454 663859 48456
rect 661480 48452 662154 48454
rect 663793 48451 663859 48454
rect 416630 48044 416636 48108
rect 416700 48106 416706 48108
rect 598933 48106 598999 48109
rect 416700 48104 598999 48106
rect 416700 48048 598938 48104
rect 598994 48048 598999 48104
rect 416700 48046 598999 48048
rect 416700 48044 416706 48046
rect 598933 48043 598999 48046
rect 361982 47772 361988 47836
rect 362052 47834 362058 47836
rect 594057 47834 594123 47837
rect 662597 47834 662663 47837
rect 362052 47832 594123 47834
rect 362052 47776 594062 47832
rect 594118 47776 594123 47832
rect 661910 47832 662663 47834
rect 661910 47791 662602 47832
rect 362052 47774 594123 47776
rect 362052 47772 362058 47774
rect 594057 47771 594123 47774
rect 661388 47776 662602 47791
rect 662658 47776 662663 47832
rect 661388 47774 662663 47776
rect 661388 47731 661970 47774
rect 662597 47771 662663 47774
rect 147622 47500 147628 47564
rect 147692 47562 147698 47564
rect 147692 47502 171150 47562
rect 147692 47500 147698 47502
rect 151905 47290 151971 47293
rect 146710 47288 151971 47290
rect 146710 47232 151910 47288
rect 151966 47232 151971 47288
rect 146710 47230 151971 47232
rect 171090 47290 171150 47502
rect 187550 47500 187556 47564
rect 187620 47562 187626 47564
rect 624417 47562 624483 47565
rect 187620 47560 624483 47562
rect 187620 47504 624422 47560
rect 624478 47504 624483 47560
rect 187620 47502 624483 47504
rect 187620 47500 187626 47502
rect 624417 47499 624483 47502
rect 662413 47426 662479 47429
rect 661388 47424 662479 47426
rect 661388 47368 662418 47424
rect 662474 47368 662479 47424
rect 661388 47366 662479 47368
rect 662413 47363 662479 47366
rect 514702 47290 514708 47292
rect 171090 47230 514708 47290
rect 131062 46956 131068 47020
rect 131132 47018 131138 47020
rect 146710 47018 146770 47230
rect 151905 47227 151971 47230
rect 514702 47228 514708 47230
rect 514772 47228 514778 47292
rect 499573 47018 499639 47021
rect 518566 47018 518572 47020
rect 131132 46958 146770 47018
rect 238710 46958 267750 47018
rect 131132 46956 131138 46958
rect 151905 45930 151971 45933
rect 238710 45930 238770 46958
rect 151905 45928 238770 45930
rect 151905 45872 151910 45928
rect 151966 45872 238770 45928
rect 151905 45870 238770 45872
rect 267690 45930 267750 46958
rect 499573 47016 518572 47018
rect 499573 46960 499578 47016
rect 499634 46960 518572 47016
rect 499573 46958 518572 46960
rect 499573 46955 499639 46958
rect 518566 46956 518572 46958
rect 518636 46956 518642 47020
rect 306966 46412 306972 46476
rect 307036 46474 307042 46476
rect 592677 46474 592743 46477
rect 307036 46472 592743 46474
rect 307036 46416 592682 46472
rect 592738 46416 592743 46472
rect 307036 46414 592743 46416
rect 307036 46412 307042 46414
rect 592677 46411 592743 46414
rect 310094 46140 310100 46204
rect 310164 46202 310170 46204
rect 597553 46202 597619 46205
rect 310164 46200 597619 46202
rect 310164 46144 597558 46200
rect 597614 46144 597619 46200
rect 310164 46142 597619 46144
rect 310164 46140 310170 46142
rect 597553 46139 597619 46142
rect 521694 45930 521700 45932
rect 267690 45870 521700 45930
rect 151905 45867 151971 45870
rect 521694 45868 521700 45870
rect 521764 45868 521770 45932
rect 445017 45114 445083 45117
rect 520406 45114 520412 45116
rect 445017 45112 520412 45114
rect 445017 45056 445022 45112
rect 445078 45056 520412 45112
rect 445017 45054 520412 45056
rect 445017 45051 445083 45054
rect 520406 45052 520412 45054
rect 520476 45052 520482 45116
rect 471646 44780 471652 44844
rect 471716 44842 471722 44844
rect 601693 44842 601759 44845
rect 471716 44840 601759 44842
rect 471716 44784 601698 44840
rect 601754 44784 601759 44840
rect 471716 44782 601759 44784
rect 471716 44780 471722 44782
rect 601693 44779 601759 44782
rect 474457 43482 474523 43485
rect 604453 43482 604519 43485
rect 474457 43480 604519 43482
rect 474457 43424 474462 43480
rect 474518 43424 604458 43480
rect 604514 43424 604519 43480
rect 474457 43422 604519 43424
rect 474457 43419 474523 43422
rect 604453 43419 604519 43422
rect 409597 42804 409663 42805
rect 411069 42804 411135 42805
rect 416589 42804 416655 42805
rect 464889 42804 464955 42805
rect 409597 42800 409644 42804
rect 409708 42802 409714 42804
rect 409597 42744 409602 42800
rect 409597 42740 409644 42744
rect 409708 42742 409754 42802
rect 411069 42800 411116 42804
rect 411180 42802 411186 42804
rect 416589 42802 416636 42804
rect 411069 42744 411074 42800
rect 409708 42740 409714 42742
rect 411069 42740 411116 42744
rect 411180 42742 411226 42802
rect 416544 42800 416636 42802
rect 416544 42744 416594 42800
rect 416544 42742 416636 42744
rect 411180 42740 411186 42742
rect 416589 42740 416636 42742
rect 416700 42740 416706 42804
rect 464838 42802 464844 42804
rect 464798 42742 464844 42802
rect 464908 42800 464955 42804
rect 464950 42744 464955 42800
rect 464838 42740 464844 42742
rect 464908 42740 464955 42744
rect 409597 42739 409663 42740
rect 411069 42739 411135 42740
rect 416589 42739 416655 42740
rect 464889 42739 464955 42740
rect 306971 42396 307037 42397
rect 310099 42396 310165 42397
rect 518617 42396 518683 42397
rect 306966 42394 306972 42396
rect 306880 42334 306972 42394
rect 306966 42332 306972 42334
rect 307036 42332 307042 42396
rect 310094 42394 310100 42396
rect 310008 42334 310100 42394
rect 310094 42332 310100 42334
rect 310164 42332 310170 42396
rect 518566 42332 518572 42396
rect 518636 42394 518683 42396
rect 518636 42392 518728 42394
rect 518678 42336 518728 42392
rect 518636 42334 518728 42336
rect 518636 42332 518683 42334
rect 306971 42331 307037 42332
rect 310099 42331 310165 42332
rect 518617 42331 518683 42332
rect 187509 42124 187575 42125
rect 361941 42124 362007 42125
rect 187509 42122 187556 42124
rect 187464 42120 187556 42122
rect 187464 42064 187514 42120
rect 187464 42062 187556 42064
rect 187509 42060 187556 42062
rect 187620 42060 187626 42124
rect 361941 42122 361988 42124
rect 361896 42120 361988 42122
rect 361896 42064 361946 42120
rect 361896 42062 361988 42064
rect 361941 42060 361988 42062
rect 362052 42060 362058 42124
rect 365161 42122 365227 42125
rect 365478 42122 365484 42124
rect 365161 42120 365484 42122
rect 365161 42064 365166 42120
rect 365222 42064 365484 42120
rect 365161 42062 365484 42064
rect 187509 42059 187575 42060
rect 361941 42059 362007 42060
rect 365161 42059 365227 42062
rect 365478 42060 365484 42062
rect 365548 42060 365554 42124
rect 460565 42122 460631 42125
rect 471605 42124 471671 42125
rect 460790 42122 460796 42124
rect 460565 42120 460796 42122
rect 460565 42064 460570 42120
rect 460626 42064 460796 42120
rect 460565 42062 460796 42064
rect 460565 42059 460631 42062
rect 460790 42060 460796 42062
rect 460860 42060 460866 42124
rect 471605 42122 471652 42124
rect 471560 42120 471652 42122
rect 471560 42064 471610 42120
rect 471560 42062 471652 42064
rect 471605 42060 471652 42062
rect 471716 42060 471722 42124
rect 514702 42060 514708 42124
rect 514772 42122 514778 42124
rect 514937 42122 515003 42125
rect 520457 42124 520523 42125
rect 514772 42120 515003 42122
rect 514772 42064 514942 42120
rect 514998 42064 515003 42120
rect 514772 42062 515003 42064
rect 514772 42060 514778 42062
rect 471605 42059 471671 42060
rect 514937 42059 515003 42062
rect 520406 42060 520412 42124
rect 520476 42122 520523 42124
rect 520476 42120 520568 42122
rect 520518 42064 520568 42120
rect 520476 42062 520568 42064
rect 520476 42060 520523 42062
rect 525742 42060 525748 42124
rect 525812 42122 525818 42124
rect 525977 42122 526043 42125
rect 525812 42120 526043 42122
rect 525812 42064 525982 42120
rect 526038 42064 526043 42120
rect 525812 42062 526043 42064
rect 525812 42060 525818 42062
rect 520457 42059 520523 42060
rect 525977 42059 526043 42062
rect 529565 42122 529631 42125
rect 529790 42122 529796 42124
rect 529565 42120 529796 42122
rect 529565 42064 529570 42120
rect 529626 42064 529796 42120
rect 529565 42062 529796 42064
rect 529565 42059 529631 42062
rect 529790 42060 529796 42062
rect 529860 42060 529866 42124
rect 521653 41988 521719 41989
rect 521653 41986 521700 41988
rect 521608 41984 521700 41986
rect 521608 41928 521658 41984
rect 521608 41926 521700 41928
rect 521653 41924 521700 41926
rect 521764 41924 521770 41988
rect 521653 41923 521719 41924
<< via3 >>
rect 195100 997656 195164 997660
rect 195100 997600 195150 997656
rect 195150 997600 195164 997656
rect 195100 997596 195164 997600
rect 87828 997188 87892 997252
rect 180564 997188 180628 997252
rect 183876 997188 183940 997252
rect 292804 996780 292868 996844
rect 527956 996780 528020 996844
rect 192524 996372 192588 996436
rect 183876 995692 183940 995756
rect 189580 995752 189644 995756
rect 189580 995696 189594 995752
rect 189594 995696 189644 995752
rect 189580 995692 189644 995696
rect 186268 995420 186332 995484
rect 192524 995480 192588 995484
rect 192524 995424 192538 995480
rect 192538 995424 192588 995480
rect 192524 995420 192588 995424
rect 194548 995420 194612 995484
rect 87828 995008 87892 995012
rect 87828 994952 87842 995008
rect 87842 994952 87892 995008
rect 87828 994948 87892 994952
rect 293540 996372 293604 996436
rect 293540 995752 293604 995756
rect 293540 995696 293554 995752
rect 293554 995696 293604 995752
rect 293540 995692 293604 995696
rect 298508 995692 298572 995756
rect 474044 996644 474108 996708
rect 627868 996644 627932 996708
rect 474780 996372 474844 996436
rect 528324 996508 528388 996572
rect 506428 995828 506492 995892
rect 485636 995752 485700 995756
rect 485636 995696 485650 995752
rect 485650 995696 485700 995752
rect 485636 995692 485700 995696
rect 527956 995752 528020 995756
rect 527956 995696 528006 995752
rect 528006 995696 528020 995752
rect 527956 995692 528020 995696
rect 528324 995692 528388 995756
rect 536604 995752 536668 995756
rect 536604 995696 536618 995752
rect 536618 995696 536668 995752
rect 536604 995692 536668 995696
rect 556108 995556 556172 995620
rect 286732 995480 286796 995484
rect 286732 995424 286746 995480
rect 286746 995424 286796 995480
rect 286732 995420 286796 995424
rect 292804 995420 292868 995484
rect 474044 995480 474108 995484
rect 474044 995424 474094 995480
rect 474094 995424 474108 995480
rect 474044 995420 474108 995424
rect 474780 995480 474844 995484
rect 474780 995424 474794 995480
rect 474794 995424 474844 995480
rect 474780 995420 474844 995424
rect 480116 995420 480180 995484
rect 627868 995752 627932 995756
rect 627868 995696 627918 995752
rect 627918 995696 627932 995752
rect 627868 995692 627932 995696
rect 242940 995208 243004 995212
rect 242940 995152 242944 995208
rect 242944 995152 243000 995208
rect 243000 995152 243004 995208
rect 242940 995148 243004 995152
rect 180564 994528 180628 994532
rect 180564 994472 180614 994528
rect 180614 994472 180628 994528
rect 180564 994468 180628 994472
rect 480116 994196 480180 994260
rect 242940 992836 243004 992900
rect 41460 968764 41524 968828
rect 42012 967192 42076 967196
rect 42012 967136 42026 967192
rect 42026 967136 42076 967192
rect 42012 967132 42076 967136
rect 675340 966512 675404 966516
rect 675340 966456 675390 966512
rect 675390 966456 675404 966512
rect 675340 966452 675404 966456
rect 676076 965092 676140 965156
rect 675156 963384 675220 963388
rect 675156 963328 675206 963384
rect 675206 963328 675220 963384
rect 675156 963324 675220 963328
rect 41828 962160 41892 962164
rect 41828 962104 41842 962160
rect 41842 962104 41892 962160
rect 41828 962100 41892 962104
rect 676628 961964 676692 962028
rect 675156 959380 675220 959444
rect 41276 959108 41340 959172
rect 676812 958292 676876 958356
rect 40724 956524 40788 956588
rect 676996 956388 677060 956452
rect 40540 955436 40604 955500
rect 675892 953940 675956 954004
rect 41460 952852 41524 952916
rect 41644 952172 41708 952236
rect 41276 951764 41340 951828
rect 42012 951628 42076 951692
rect 676628 951492 676692 951556
rect 676076 949996 676140 950060
rect 675892 949240 675956 949244
rect 675892 949184 675942 949240
rect 675942 949184 675956 949240
rect 675892 949180 675956 949184
rect 675340 948908 675404 948972
rect 41828 938980 41892 939044
rect 41828 936532 41892 936596
rect 676996 931908 677060 931972
rect 676812 930684 676876 930748
rect 676076 877100 676140 877164
rect 676996 876420 677060 876484
rect 675340 874032 675404 874036
rect 675340 873976 675390 874032
rect 675390 873976 675404 874032
rect 675340 873972 675404 873976
rect 676812 872748 676876 872812
rect 673868 872204 673932 872268
rect 675340 869620 675404 869684
rect 675892 869620 675956 869684
rect 674420 854312 674484 854316
rect 674420 854256 674470 854312
rect 674470 854256 674484 854312
rect 674420 854252 674484 854256
rect 42012 813180 42076 813244
rect 40540 810698 40604 810762
rect 40724 810562 40788 810626
rect 41828 809296 41892 809300
rect 41828 809240 41842 809296
rect 41842 809240 41892 809296
rect 41828 809236 41892 809240
rect 40908 805020 40972 805084
rect 41828 803796 41892 803860
rect 40356 800728 40420 800732
rect 40356 800672 40370 800728
rect 40370 800672 40420 800728
rect 40356 800668 40420 800672
rect 41092 800668 41156 800732
rect 41092 796180 41156 796244
rect 40356 794412 40420 794476
rect 40908 793460 40972 793524
rect 41644 791556 41708 791620
rect 40540 790196 40604 790260
rect 40724 789924 40788 789988
rect 41460 788156 41524 788220
rect 41828 787884 41892 787948
rect 674236 784212 674300 784276
rect 674972 780328 675036 780332
rect 674972 780272 674986 780328
rect 674986 780272 675036 780328
rect 674972 780268 675036 780272
rect 675156 779860 675220 779924
rect 675156 775372 675220 775436
rect 674972 773332 675036 773396
rect 676076 772652 676140 772716
rect 673868 772380 673932 772444
rect 674420 771972 674484 772036
rect 675892 771292 675956 771356
rect 41460 769796 41524 769860
rect 40908 765716 40972 765780
rect 40540 765308 40604 765372
rect 40724 764900 40788 764964
rect 676996 761832 677060 761836
rect 676996 761776 677010 761832
rect 677010 761776 677060 761832
rect 676996 761772 677060 761776
rect 41828 759596 41892 759660
rect 41644 757692 41708 757756
rect 675892 753748 675956 753812
rect 42196 751632 42260 751636
rect 42196 751576 42246 751632
rect 42246 751576 42260 751632
rect 42196 751572 42260 751576
rect 40908 751028 40972 751092
rect 676076 751028 676140 751092
rect 42196 750484 42260 750548
rect 40724 750348 40788 750412
rect 40540 749396 40604 749460
rect 41828 745588 41892 745652
rect 41644 745044 41708 745108
rect 41460 743684 41524 743748
rect 675524 743064 675588 743068
rect 675524 743008 675574 743064
rect 675574 743008 675588 743064
rect 675524 743004 675588 743008
rect 674420 738652 674484 738716
rect 674604 738108 674668 738172
rect 675340 735116 675404 735180
rect 676812 733620 676876 733684
rect 674604 725868 674668 725932
rect 41828 725792 41892 725796
rect 41828 725736 41842 725792
rect 41842 725736 41892 725792
rect 41828 725732 41892 725736
rect 40724 721708 40788 721772
rect 40908 721708 40972 721772
rect 41644 721708 41708 721772
rect 676076 721516 676140 721580
rect 40540 718524 40604 718588
rect 41828 716756 41892 716820
rect 42564 714716 42628 714780
rect 40356 714172 40420 714236
rect 42380 714172 42444 714236
rect 42012 713900 42076 713964
rect 677732 713488 677796 713492
rect 677732 713432 677746 713488
rect 677746 713432 677796 713488
rect 677732 713428 677796 713432
rect 40356 712132 40420 712196
rect 42564 711588 42628 711652
rect 42012 710364 42076 710428
rect 40724 709412 40788 709476
rect 674236 709140 674300 709204
rect 40908 708460 40972 708524
rect 40540 707236 40604 707300
rect 42380 706556 42444 706620
rect 41460 702476 41524 702540
rect 41644 701388 41708 701452
rect 41828 701116 41892 701180
rect 675340 696824 675404 696828
rect 675340 696768 675390 696824
rect 675390 696768 675404 696824
rect 675340 696764 675404 696768
rect 674052 694588 674116 694652
rect 676996 694044 677060 694108
rect 674604 692956 674668 693020
rect 675340 685884 675404 685948
rect 41828 682408 41892 682412
rect 41828 682352 41842 682408
rect 41842 682352 41892 682408
rect 41828 682348 41892 682352
rect 676076 681804 676140 681868
rect 41828 680368 41892 680372
rect 41828 680312 41842 680368
rect 41842 680312 41892 680368
rect 41828 680308 41892 680312
rect 40540 678928 40604 678992
rect 40724 678928 40788 678992
rect 674420 674052 674484 674116
rect 41828 672692 41892 672756
rect 41092 671196 41156 671260
rect 40908 670924 40972 670988
rect 40908 667932 40972 667996
rect 41092 667388 41156 667452
rect 676996 666572 677060 666636
rect 40724 666436 40788 666500
rect 42012 666436 42076 666500
rect 676812 665348 676876 665412
rect 42012 664048 42076 664052
rect 42012 663992 42026 664048
rect 42026 663992 42076 664048
rect 42012 663988 42076 663992
rect 40540 662628 40604 662692
rect 41460 659636 41524 659700
rect 41644 658548 41708 658612
rect 41828 658276 41892 658340
rect 675524 652896 675588 652900
rect 675524 652840 675574 652896
rect 675574 652840 675588 652896
rect 675524 652836 675588 652840
rect 675156 650176 675220 650180
rect 675156 650120 675206 650176
rect 675206 650120 675220 650176
rect 675156 650116 675220 650120
rect 674236 648892 674300 648956
rect 675156 647940 675220 648004
rect 674972 643920 675036 643924
rect 674972 643864 674986 643920
rect 674986 643864 675036 643920
rect 674972 643860 675036 643864
rect 41460 640596 41524 640660
rect 676812 640188 676876 640252
rect 674972 638148 675036 638212
rect 675524 637604 675588 637668
rect 41644 637332 41708 637396
rect 40540 636924 40604 636988
rect 674052 636788 674116 636852
rect 40908 636108 40972 636172
rect 40724 635700 40788 635764
rect 41828 635292 41892 635356
rect 675156 631408 675220 631412
rect 675156 631352 675206 631408
rect 675206 631352 675220 631408
rect 675156 631348 675220 631352
rect 676076 631348 676140 631412
rect 42196 626724 42260 626788
rect 40908 625228 40972 625292
rect 42012 625228 42076 625292
rect 674604 623596 674668 623660
rect 42012 621480 42076 621484
rect 42012 621424 42026 621480
rect 42026 621424 42076 621480
rect 42012 621420 42076 621424
rect 42196 620196 42260 620260
rect 40724 619788 40788 619852
rect 40540 618972 40604 619036
rect 41828 618700 41892 618764
rect 671476 616796 671540 616860
rect 41460 615980 41524 616044
rect 41828 612776 41892 612780
rect 41828 612720 41842 612776
rect 41842 612720 41892 612776
rect 41828 612716 41892 612720
rect 671476 608696 671540 608700
rect 671476 608640 671526 608696
rect 671526 608640 671540 608696
rect 671476 608636 671540 608640
rect 674420 604420 674484 604484
rect 674604 602924 674668 602988
rect 42012 596396 42076 596460
rect 41828 596048 41892 596052
rect 41828 595992 41842 596048
rect 41842 595992 41892 596048
rect 41828 595988 41892 595992
rect 676076 592860 676140 592924
rect 675156 592588 675220 592652
rect 40724 589656 40788 589660
rect 40724 589600 40774 589656
rect 40774 589600 40788 589656
rect 40724 589596 40788 589600
rect 40908 589460 40972 589524
rect 40540 589384 40604 589388
rect 40540 589328 40590 589384
rect 40590 589328 40604 589384
rect 40540 589324 40604 589328
rect 41828 587148 41892 587212
rect 676076 586196 676140 586260
rect 41092 584836 41156 584900
rect 42012 584836 42076 584900
rect 40356 584564 40420 584628
rect 42564 584564 42628 584628
rect 42012 582584 42076 582588
rect 42012 582528 42026 582584
rect 42026 582528 42076 582584
rect 42012 582524 42076 582528
rect 41092 580484 41156 580548
rect 40356 580212 40420 580276
rect 40908 579940 40972 580004
rect 42564 576540 42628 576604
rect 676812 576404 676876 576468
rect 40540 575452 40604 575516
rect 40724 574636 40788 574700
rect 41460 573956 41524 574020
rect 674236 573276 674300 573340
rect 41828 572188 41892 572252
rect 41644 571916 41708 571980
rect 676996 571508 677060 571572
rect 675340 561912 675404 561916
rect 675340 561856 675390 561912
rect 675390 561856 675404 561912
rect 675340 561852 675404 561856
rect 675524 559464 675588 559468
rect 675524 559408 675538 559464
rect 675538 559408 675588 559464
rect 675524 559404 675588 559408
rect 676812 558996 676876 559060
rect 42380 553964 42444 554028
rect 42196 552740 42260 552804
rect 41828 550428 41892 550492
rect 675156 550292 675220 550356
rect 675524 547904 675588 547908
rect 675524 547848 675538 547904
rect 675538 547848 675588 547904
rect 675524 547844 675588 547848
rect 675340 547572 675404 547636
rect 41644 546348 41708 546412
rect 41460 546076 41524 546140
rect 42380 546076 42444 546140
rect 40908 545804 40972 545868
rect 41828 545804 41892 545868
rect 675156 545864 675220 545868
rect 675156 545808 675206 545864
rect 675206 545808 675220 545864
rect 675156 545804 675220 545808
rect 40724 545532 40788 545596
rect 40540 545260 40604 545324
rect 676076 545124 676140 545188
rect 40908 538188 40972 538252
rect 40724 536828 40788 536892
rect 40540 533292 40604 533356
rect 41828 532612 41892 532676
rect 676996 531388 677060 531452
rect 41644 529756 41708 529820
rect 674420 528804 674484 528868
rect 41460 527580 41524 527644
rect 674604 527036 674668 527100
rect 673868 525812 673932 525876
rect 676812 500924 676876 500988
rect 41460 431156 41524 431220
rect 41460 428198 41524 428262
rect 41828 426396 41892 426460
rect 41828 425580 41892 425644
rect 40724 422248 40788 422312
rect 42012 421908 42076 421972
rect 40540 418644 40604 418708
rect 42012 418644 42076 418708
rect 41828 418372 41892 418436
rect 40724 407492 40788 407556
rect 40540 403820 40604 403884
rect 41828 401976 41892 401980
rect 41828 401920 41842 401976
rect 41842 401920 41892 401976
rect 41828 401916 41892 401920
rect 41460 400012 41524 400076
rect 41828 398848 41892 398852
rect 41828 398792 41842 398848
rect 41842 398792 41892 398848
rect 41828 398788 41892 398792
rect 676076 398788 676140 398852
rect 676260 396748 676324 396812
rect 676628 395116 676692 395180
rect 676444 394708 676508 394772
rect 672948 394572 673012 394636
rect 675892 389812 675956 389876
rect 675708 388452 675772 388516
rect 676260 384916 676324 384980
rect 41460 382196 41524 382260
rect 676444 380564 676508 380628
rect 41644 380156 41708 380220
rect 40908 379340 40972 379404
rect 41828 378932 41892 378996
rect 675708 378720 675772 378724
rect 675708 378664 675758 378720
rect 675758 378664 675772 378720
rect 675708 378660 675772 378664
rect 40540 378524 40604 378588
rect 40724 378116 40788 378180
rect 674788 377980 674852 378044
rect 676628 377300 676692 377364
rect 676076 374988 676140 375052
rect 675892 372948 675956 373012
rect 674788 372540 674852 372604
rect 40908 365604 40972 365668
rect 40724 363700 40788 363764
rect 40540 360572 40604 360636
rect 41828 358728 41892 358732
rect 41828 358672 41878 358728
rect 41878 358672 41892 358728
rect 41828 358668 41892 358672
rect 41460 356900 41524 356964
rect 42012 355736 42076 355740
rect 42012 355680 42026 355736
rect 42026 355680 42076 355736
rect 42012 355676 42076 355680
rect 675340 354180 675404 354244
rect 675524 352956 675588 353020
rect 675708 352140 675772 352204
rect 675892 351732 675956 351796
rect 675892 350916 675956 350980
rect 675892 350100 675956 350164
rect 675340 345476 675404 345540
rect 675892 345476 675956 345540
rect 671844 345264 671908 345268
rect 671844 345208 671858 345264
rect 671858 345208 671908 345264
rect 671844 345204 671908 345208
rect 671292 344932 671356 344996
rect 671844 340444 671908 340508
rect 676628 340308 676692 340372
rect 41460 339764 41524 339828
rect 41828 339492 41892 339556
rect 675892 339356 675956 339420
rect 41644 338540 41708 338604
rect 675524 337784 675588 337788
rect 675524 337728 675574 337784
rect 675574 337728 675588 337784
rect 675524 337724 675588 337728
rect 40540 337316 40604 337380
rect 676444 336636 676508 336700
rect 40724 336092 40788 336156
rect 676260 332284 676324 332348
rect 676076 326844 676140 326908
rect 41828 324864 41892 324868
rect 41828 324808 41842 324864
rect 41842 324808 41892 324864
rect 41828 324804 41892 324808
rect 40724 322764 40788 322828
rect 41828 315616 41892 315620
rect 41828 315560 41842 315616
rect 41842 315560 41892 315616
rect 41828 315556 41892 315560
rect 41460 313652 41524 313716
rect 40540 312972 40604 313036
rect 675892 308756 675956 308820
rect 676076 304914 676140 304978
rect 676076 302968 676140 302972
rect 676076 302912 676090 302968
rect 676090 302912 676140 302968
rect 676076 302908 676140 302912
rect 676444 301608 676508 301612
rect 676444 301552 676458 301608
rect 676458 301552 676508 301608
rect 676444 301548 676508 301552
rect 675892 299372 675956 299436
rect 675708 297332 675772 297396
rect 41828 296788 41892 296852
rect 675524 296516 675588 296580
rect 42012 296380 42076 296444
rect 675524 295352 675588 295356
rect 675524 295296 675574 295352
rect 675574 295296 675588 295352
rect 675524 295292 675588 295296
rect 40540 292588 40604 292592
rect 40540 292532 40554 292588
rect 40554 292532 40604 292588
rect 40540 292528 40604 292532
rect 40724 292528 40788 292592
rect 40908 292528 40972 292592
rect 41828 292300 41892 292364
rect 676444 291484 676508 291548
rect 676260 290940 676324 291004
rect 676628 286996 676692 287060
rect 676076 283596 676140 283660
rect 675892 282780 675956 282844
rect 675708 281616 675772 281620
rect 675708 281560 675722 281616
rect 675722 281560 675772 281616
rect 675708 281556 675772 281560
rect 42012 281480 42076 281484
rect 42012 281424 42026 281480
rect 42026 281424 42076 281480
rect 42012 281420 42076 281424
rect 671292 278700 671356 278764
rect 672948 278700 673012 278764
rect 673868 278564 673932 278628
rect 40908 277884 40972 277948
rect 673868 277612 673932 277676
rect 40724 277340 40788 277404
rect 40540 273396 40604 273460
rect 41828 272368 41892 272372
rect 41828 272312 41842 272368
rect 41842 272312 41892 272368
rect 41828 272308 41892 272312
rect 41460 270404 41524 270468
rect 674788 264148 674852 264212
rect 676076 263604 676140 263668
rect 676996 261564 677060 261628
rect 676812 260748 676876 260812
rect 40724 249732 40788 249796
rect 673868 249792 673932 249796
rect 673868 249736 673918 249792
rect 673918 249736 673932 249792
rect 673868 249732 673932 249736
rect 674788 249732 674852 249796
rect 676076 249732 676140 249796
rect 40540 249324 40604 249388
rect 676996 248236 677060 248300
rect 676812 246604 676876 246668
rect 666876 246060 666940 246124
rect 666508 245924 666572 245988
rect 668164 245984 668228 245988
rect 668164 245928 668178 245984
rect 668178 245928 668228 245984
rect 668164 245924 668228 245928
rect 666692 245652 666756 245716
rect 668348 245712 668412 245716
rect 668348 245656 668362 245712
rect 668362 245656 668412 245712
rect 668348 245652 668412 245656
rect 675340 243264 675404 243268
rect 675340 243208 675354 243264
rect 675354 243208 675404 243264
rect 675340 243204 675404 243208
rect 675340 238640 675404 238644
rect 675340 238584 675390 238640
rect 675390 238584 675404 238640
rect 675340 238580 675404 238584
rect 42380 237356 42444 237420
rect 40724 236540 40788 236604
rect 40540 234500 40604 234564
rect 147812 230964 147876 231028
rect 147812 230420 147876 230484
rect 42380 227292 42444 227356
rect 574140 219192 574204 219196
rect 574140 219136 574190 219192
rect 574190 219136 574204 219192
rect 574140 219132 574204 219136
rect 574508 219132 574572 219196
rect 499620 219056 499684 219060
rect 499620 219000 499634 219056
rect 499634 219000 499684 219056
rect 499620 218996 499684 219000
rect 675524 218588 675588 218652
rect 490420 218104 490484 218108
rect 490420 218048 490434 218104
rect 490434 218048 490484 218104
rect 490420 218044 490484 218048
rect 493732 217968 493796 217972
rect 493732 217912 493746 217968
rect 493746 217912 493796 217968
rect 493732 217908 493796 217912
rect 669452 217908 669516 217972
rect 566044 217772 566108 217836
rect 501276 217560 501340 217564
rect 501276 217504 501290 217560
rect 501290 217504 501340 217560
rect 501276 217500 501340 217504
rect 675708 217364 675772 217428
rect 491156 217288 491220 217292
rect 491156 217232 491170 217288
rect 491170 217232 491220 217288
rect 491156 217228 491220 217232
rect 501276 216956 501340 217020
rect 575796 216684 575860 216748
rect 670924 216608 670988 216612
rect 670924 216552 670974 216608
rect 670974 216552 670988 216608
rect 670924 216548 670988 216552
rect 675340 216548 675404 216612
rect 574324 216472 574388 216476
rect 574324 216416 574374 216472
rect 574374 216416 574388 216472
rect 574324 216412 574388 216416
rect 671108 216140 671172 216204
rect 566044 216004 566108 216068
rect 675892 214508 675956 214572
rect 673684 213964 673748 214028
rect 672948 212604 673012 212668
rect 675340 212332 675404 212396
rect 675892 212332 675956 212396
rect 676444 211380 676508 211444
rect 667980 211108 668044 211172
rect 669636 211108 669700 211172
rect 670740 211168 670804 211172
rect 670740 211112 670790 211168
rect 670790 211112 670804 211168
rect 670740 211108 670804 211112
rect 675892 211108 675956 211172
rect 671108 210836 671172 210900
rect 666692 210428 666756 210492
rect 667060 210428 667124 210492
rect 673132 210428 673196 210492
rect 673500 210428 673564 210492
rect 675524 210428 675588 210492
rect 676076 210428 676140 210492
rect 41828 210020 41892 210084
rect 673316 209204 673380 209268
rect 40908 208116 40972 208180
rect 40540 207708 40604 207772
rect 667980 207300 668044 207364
rect 40724 206076 40788 206140
rect 41460 205668 41524 205732
rect 669268 205396 669332 205460
rect 669636 205396 669700 205460
rect 676260 204988 676324 205052
rect 669452 204036 669516 204100
rect 668164 202404 668228 202468
rect 676812 201316 676876 201380
rect 41644 200636 41708 200700
rect 676628 199956 676692 200020
rect 666876 199072 666940 199136
rect 675708 198384 675772 198388
rect 675708 198328 675758 198384
rect 675758 198328 675772 198384
rect 675708 198324 675772 198328
rect 668348 197508 668412 197572
rect 40908 197100 40972 197164
rect 676444 196964 676508 197028
rect 41828 195256 41892 195260
rect 41828 195200 41842 195256
rect 41842 195200 41892 195256
rect 41828 195196 41892 195200
rect 666876 194176 666940 194240
rect 676076 193156 676140 193220
rect 675892 192748 675956 192812
rect 40724 191524 40788 191588
rect 666692 189280 666756 189344
rect 41828 185872 41892 185876
rect 41828 185816 41842 185872
rect 41842 185816 41892 185872
rect 41828 185812 41892 185816
rect 41460 184044 41524 184108
rect 672764 183500 672828 183564
rect 673132 183560 673196 183564
rect 673132 183504 673182 183560
rect 673182 183504 673196 183560
rect 673132 183500 673196 183504
rect 40540 183364 40604 183428
rect 669452 179556 669516 179620
rect 675892 174660 675956 174724
rect 675708 173572 675772 173636
rect 673316 173028 673380 173092
rect 675340 172348 675404 172412
rect 675892 170716 675956 170780
rect 675892 169356 675956 169420
rect 672948 168268 673012 168332
rect 675708 167588 675772 167652
rect 676628 166424 676692 166428
rect 676628 166368 676678 166424
rect 676678 166368 676692 166424
rect 676628 166364 676692 166368
rect 670924 165684 670988 165748
rect 675340 162148 675404 162212
rect 675892 162148 675956 162212
rect 675524 161332 675588 161396
rect 675524 160168 675588 160172
rect 675524 160112 675574 160168
rect 675574 160112 675588 160168
rect 675524 160108 675588 160112
rect 676444 156436 676508 156500
rect 676260 155620 676324 155684
rect 670740 155076 670804 155140
rect 673684 153308 673748 153372
rect 675892 153036 675956 153100
rect 676628 151404 676692 151468
rect 673500 148412 673564 148476
rect 676076 148412 676140 148476
rect 675708 147656 675772 147660
rect 675708 147600 675722 147656
rect 675722 147600 675772 147656
rect 675708 147596 675772 147600
rect 672948 133724 673012 133788
rect 676260 128556 676324 128620
rect 676076 128148 676140 128212
rect 675892 127196 675956 127260
rect 676812 124476 676876 124540
rect 676996 117268 677060 117332
rect 675708 116996 675772 117060
rect 676260 113052 676324 113116
rect 676996 110332 677060 110396
rect 675892 108020 675956 108084
rect 676076 103124 676140 103188
rect 675708 102640 675772 102644
rect 675708 102584 675722 102640
rect 675722 102584 675772 102640
rect 675708 102580 675772 102584
rect 676812 101356 676876 101420
rect 637252 96868 637316 96932
rect 634676 95644 634740 95708
rect 637068 78568 637132 78572
rect 637068 78512 637118 78568
rect 637118 78512 637132 78568
rect 637068 78508 637132 78512
rect 634676 77692 634740 77756
rect 409644 53076 409708 53140
rect 464844 51716 464908 51780
rect 525748 50492 525812 50556
rect 529796 50492 529860 50556
rect 147628 50220 147692 50284
rect 460796 50220 460860 50284
rect 131068 49736 131132 49740
rect 131068 49680 131082 49736
rect 131082 49680 131132 49736
rect 131068 49676 131132 49680
rect 411116 49132 411180 49196
rect 365484 48860 365548 48924
rect 416636 48044 416700 48108
rect 361988 47772 362052 47836
rect 147628 47500 147692 47564
rect 187556 47500 187620 47564
rect 131068 46956 131132 47020
rect 514708 47228 514772 47292
rect 518572 46956 518636 47020
rect 306972 46412 307036 46476
rect 310100 46140 310164 46204
rect 521700 45868 521764 45932
rect 520412 45052 520476 45116
rect 471652 44780 471716 44844
rect 409644 42800 409708 42804
rect 409644 42744 409658 42800
rect 409658 42744 409708 42800
rect 409644 42740 409708 42744
rect 411116 42800 411180 42804
rect 411116 42744 411130 42800
rect 411130 42744 411180 42800
rect 411116 42740 411180 42744
rect 416636 42800 416700 42804
rect 416636 42744 416650 42800
rect 416650 42744 416700 42800
rect 416636 42740 416700 42744
rect 464844 42800 464908 42804
rect 464844 42744 464894 42800
rect 464894 42744 464908 42800
rect 464844 42740 464908 42744
rect 306972 42392 307036 42396
rect 306972 42336 306976 42392
rect 306976 42336 307032 42392
rect 307032 42336 307036 42392
rect 306972 42332 307036 42336
rect 310100 42392 310164 42396
rect 310100 42336 310104 42392
rect 310104 42336 310160 42392
rect 310160 42336 310164 42392
rect 310100 42332 310164 42336
rect 518572 42392 518636 42396
rect 518572 42336 518622 42392
rect 518622 42336 518636 42392
rect 518572 42332 518636 42336
rect 187556 42120 187620 42124
rect 187556 42064 187570 42120
rect 187570 42064 187620 42120
rect 187556 42060 187620 42064
rect 361988 42120 362052 42124
rect 361988 42064 362002 42120
rect 362002 42064 362052 42120
rect 361988 42060 362052 42064
rect 365484 42060 365548 42124
rect 460796 42060 460860 42124
rect 471652 42120 471716 42124
rect 471652 42064 471666 42120
rect 471666 42064 471716 42120
rect 471652 42060 471716 42064
rect 514708 42060 514772 42124
rect 520412 42120 520476 42124
rect 520412 42064 520462 42120
rect 520462 42064 520476 42120
rect 520412 42060 520476 42064
rect 525748 42060 525812 42124
rect 529796 42060 529860 42124
rect 521700 41984 521764 41988
rect 521700 41928 521714 41984
rect 521714 41928 521764 41984
rect 521700 41924 521764 41928
<< metal4 >>
rect 195099 997660 195165 997661
rect 195099 997596 195100 997660
rect 195164 997596 195165 997660
rect 195099 997595 195165 997596
rect 195102 997338 195162 997595
rect 87827 997252 87893 997253
rect 87827 997188 87828 997252
rect 87892 997188 87893 997252
rect 87827 997187 87893 997188
rect 180563 997252 180629 997253
rect 180563 997188 180564 997252
rect 180628 997188 180629 997252
rect 180563 997187 180629 997188
rect 183875 997252 183941 997253
rect 183875 997188 183876 997252
rect 183940 997188 183941 997252
rect 183875 997187 183941 997188
rect 87830 995013 87890 997187
rect 87827 995012 87893 995013
rect 87827 994948 87828 995012
rect 87892 994948 87893 995012
rect 87827 994947 87893 994948
rect 180566 994533 180626 997187
rect 183878 995757 183938 997187
rect 189582 995757 189642 997102
rect 292803 996844 292869 996845
rect 292803 996780 292804 996844
rect 292868 996780 292869 996844
rect 292803 996779 292869 996780
rect 192523 996436 192589 996437
rect 192523 996372 192524 996436
rect 192588 996372 192589 996436
rect 192523 996371 192589 996372
rect 183875 995756 183941 995757
rect 183875 995692 183876 995756
rect 183940 995692 183941 995756
rect 183875 995691 183941 995692
rect 189579 995756 189645 995757
rect 189579 995692 189580 995756
rect 189644 995692 189645 995756
rect 189579 995691 189645 995692
rect 192526 995485 192586 996371
rect 292806 995485 292866 996779
rect 474043 996708 474109 996709
rect 474043 996644 474044 996708
rect 474108 996644 474109 996708
rect 474043 996643 474109 996644
rect 293539 996436 293605 996437
rect 293539 996372 293540 996436
rect 293604 996372 293605 996436
rect 293539 996371 293605 996372
rect 293542 995757 293602 996371
rect 293539 995756 293605 995757
rect 293539 995692 293540 995756
rect 293604 995692 293605 995756
rect 293539 995691 293605 995692
rect 298507 995756 298573 995757
rect 298507 995692 298508 995756
rect 298572 995692 298573 995756
rect 298507 995691 298573 995692
rect 186267 995484 186333 995485
rect 186267 995420 186268 995484
rect 186332 995420 186333 995484
rect 186267 995419 186333 995420
rect 192523 995484 192589 995485
rect 192523 995420 192524 995484
rect 192588 995420 192589 995484
rect 192523 995419 192589 995420
rect 194547 995484 194613 995485
rect 194547 995420 194548 995484
rect 194612 995420 194613 995484
rect 194547 995419 194613 995420
rect 286731 995484 286797 995485
rect 286731 995420 286732 995484
rect 286796 995420 286797 995484
rect 286731 995419 286797 995420
rect 292803 995484 292869 995485
rect 292803 995420 292804 995484
rect 292868 995420 292869 995484
rect 292803 995419 292869 995420
rect 180563 994532 180629 994533
rect 180563 994468 180564 994532
rect 180628 994468 180629 994532
rect 180563 994467 180629 994468
rect 186270 993258 186330 995419
rect 194550 993258 194610 995419
rect 242939 995212 243005 995213
rect 242939 995148 242940 995212
rect 243004 995148 243005 995212
rect 242939 995147 243005 995148
rect 242942 992901 243002 995147
rect 286734 993258 286794 995419
rect 298510 993258 298570 995691
rect 474046 995485 474106 996643
rect 474779 996436 474845 996437
rect 474779 996372 474780 996436
rect 474844 996372 474845 996436
rect 474779 996371 474845 996372
rect 474782 995485 474842 996371
rect 485638 995757 485698 997102
rect 506430 995893 506490 997102
rect 527955 996844 528021 996845
rect 527955 996780 527956 996844
rect 528020 996780 528021 996844
rect 527955 996779 528021 996780
rect 506427 995892 506493 995893
rect 506427 995828 506428 995892
rect 506492 995828 506493 995892
rect 506427 995827 506493 995828
rect 527958 995757 528018 996779
rect 528323 996572 528389 996573
rect 528323 996508 528324 996572
rect 528388 996508 528389 996572
rect 528323 996507 528389 996508
rect 528326 995757 528386 996507
rect 536606 995757 536666 997102
rect 485635 995756 485701 995757
rect 485635 995692 485636 995756
rect 485700 995692 485701 995756
rect 485635 995691 485701 995692
rect 527955 995756 528021 995757
rect 527955 995692 527956 995756
rect 528020 995692 528021 995756
rect 527955 995691 528021 995692
rect 528323 995756 528389 995757
rect 528323 995692 528324 995756
rect 528388 995692 528389 995756
rect 528323 995691 528389 995692
rect 536603 995756 536669 995757
rect 536603 995692 536604 995756
rect 536668 995692 536669 995756
rect 536603 995691 536669 995692
rect 556110 995621 556170 997102
rect 627867 996708 627933 996709
rect 627867 996644 627868 996708
rect 627932 996644 627933 996708
rect 627867 996643 627933 996644
rect 627870 995757 627930 996643
rect 627867 995756 627933 995757
rect 627867 995692 627868 995756
rect 627932 995692 627933 995756
rect 627867 995691 627933 995692
rect 556107 995620 556173 995621
rect 556107 995556 556108 995620
rect 556172 995556 556173 995620
rect 556107 995555 556173 995556
rect 474043 995484 474109 995485
rect 474043 995420 474044 995484
rect 474108 995420 474109 995484
rect 474043 995419 474109 995420
rect 474779 995484 474845 995485
rect 474779 995420 474780 995484
rect 474844 995420 474845 995484
rect 474779 995419 474845 995420
rect 480115 995484 480181 995485
rect 480115 995420 480116 995484
rect 480180 995420 480181 995484
rect 480115 995419 480181 995420
rect 480118 994261 480178 995419
rect 480115 994260 480181 994261
rect 480115 994196 480116 994260
rect 480180 994196 480181 994260
rect 480115 994195 480181 994196
rect 242939 992900 243005 992901
rect 242939 992836 242940 992900
rect 243004 992836 243005 992900
rect 242939 992835 243005 992836
rect 41459 968828 41525 968829
rect 41459 968764 41460 968828
rect 41524 968764 41525 968828
rect 41459 968763 41525 968764
rect 41275 959172 41341 959173
rect 41275 959108 41276 959172
rect 41340 959108 41341 959172
rect 41275 959107 41341 959108
rect 40723 956588 40789 956589
rect 40723 956524 40724 956588
rect 40788 956524 40789 956588
rect 40723 956523 40789 956524
rect 40539 955500 40605 955501
rect 40539 955436 40540 955500
rect 40604 955436 40605 955500
rect 40539 955435 40605 955436
rect 40542 937050 40602 955435
rect 40726 939450 40786 956523
rect 41278 951829 41338 959107
rect 41462 952917 41522 968763
rect 42011 967196 42077 967197
rect 42011 967132 42012 967196
rect 42076 967132 42077 967196
rect 42011 967131 42077 967132
rect 41827 962164 41893 962165
rect 41827 962100 41828 962164
rect 41892 962100 41893 962164
rect 41827 962099 41893 962100
rect 41830 953610 41890 962099
rect 41646 953550 41890 953610
rect 41459 952916 41525 952917
rect 41459 952852 41460 952916
rect 41524 952852 41525 952916
rect 41459 952851 41525 952852
rect 41646 952237 41706 953550
rect 41643 952236 41709 952237
rect 41643 952172 41644 952236
rect 41708 952172 41709 952236
rect 41643 952171 41709 952172
rect 41275 951828 41341 951829
rect 41275 951764 41276 951828
rect 41340 951764 41341 951828
rect 41275 951763 41341 951764
rect 42014 951693 42074 967131
rect 675339 966516 675405 966517
rect 675339 966452 675340 966516
rect 675404 966452 675405 966516
rect 675339 966451 675405 966452
rect 675155 963388 675221 963389
rect 675155 963324 675156 963388
rect 675220 963324 675221 963388
rect 675155 963323 675221 963324
rect 675158 959445 675218 963323
rect 675155 959444 675221 959445
rect 675155 959380 675156 959444
rect 675220 959380 675221 959444
rect 675155 959379 675221 959380
rect 42011 951692 42077 951693
rect 42011 951628 42012 951692
rect 42076 951628 42077 951692
rect 42011 951627 42077 951628
rect 675342 948973 675402 966451
rect 676075 965156 676141 965157
rect 676075 965092 676076 965156
rect 676140 965092 676141 965156
rect 676075 965091 676141 965092
rect 675891 954004 675957 954005
rect 675891 953940 675892 954004
rect 675956 953940 675957 954004
rect 675891 953939 675957 953940
rect 675894 949245 675954 953939
rect 676078 950061 676138 965091
rect 676627 962028 676693 962029
rect 676627 961964 676628 962028
rect 676692 961964 676693 962028
rect 676627 961963 676693 961964
rect 676630 951557 676690 961963
rect 676811 958356 676877 958357
rect 676811 958292 676812 958356
rect 676876 958292 676877 958356
rect 676811 958291 676877 958292
rect 676627 951556 676693 951557
rect 676627 951492 676628 951556
rect 676692 951492 676693 951556
rect 676627 951491 676693 951492
rect 676075 950060 676141 950061
rect 676075 949996 676076 950060
rect 676140 949996 676141 950060
rect 676075 949995 676141 949996
rect 675891 949244 675957 949245
rect 675891 949180 675892 949244
rect 675956 949180 675957 949244
rect 675891 949179 675957 949180
rect 675339 948972 675405 948973
rect 675339 948908 675340 948972
rect 675404 948908 675405 948972
rect 675339 948907 675405 948908
rect 40726 939390 41890 939450
rect 41830 939045 41890 939390
rect 41827 939044 41893 939045
rect 41827 938980 41828 939044
rect 41892 938980 41893 939044
rect 41827 938979 41893 938980
rect 40542 936990 41890 937050
rect 41830 936597 41890 936990
rect 41827 936596 41893 936597
rect 41827 936532 41828 936596
rect 41892 936532 41893 936596
rect 41827 936531 41893 936532
rect 676814 930749 676874 958291
rect 676995 956452 677061 956453
rect 676995 956388 676996 956452
rect 677060 956388 677061 956452
rect 676995 956387 677061 956388
rect 676998 931973 677058 956387
rect 676995 931972 677061 931973
rect 676995 931908 676996 931972
rect 677060 931908 677061 931972
rect 676995 931907 677061 931908
rect 676811 930748 676877 930749
rect 676811 930684 676812 930748
rect 676876 930684 676877 930748
rect 676811 930683 676877 930684
rect 676075 877164 676141 877165
rect 676075 877100 676076 877164
rect 676140 877100 676141 877164
rect 676075 877099 676141 877100
rect 675339 874036 675405 874037
rect 675339 873972 675340 874036
rect 675404 873972 675405 874036
rect 675339 873971 675405 873972
rect 673867 872268 673933 872269
rect 673867 872204 673868 872268
rect 673932 872204 673933 872268
rect 673867 872203 673933 872204
rect 42011 813244 42077 813245
rect 42011 813180 42012 813244
rect 42076 813180 42077 813244
rect 42011 813179 42077 813180
rect 40539 810762 40605 810763
rect 40539 810698 40540 810762
rect 40604 810698 40605 810762
rect 40539 810697 40605 810698
rect 40355 800732 40421 800733
rect 40355 800668 40356 800732
rect 40420 800668 40421 800732
rect 40355 800667 40421 800668
rect 40358 794477 40418 800667
rect 40355 794476 40421 794477
rect 40355 794412 40356 794476
rect 40420 794412 40421 794476
rect 40355 794411 40421 794412
rect 40542 790261 40602 810697
rect 40723 810626 40789 810627
rect 40723 810562 40724 810626
rect 40788 810562 40789 810626
rect 40723 810561 40789 810562
rect 40539 790260 40605 790261
rect 40539 790196 40540 790260
rect 40604 790196 40605 790260
rect 40539 790195 40605 790196
rect 40726 789989 40786 810561
rect 42014 809570 42074 813179
rect 41462 809510 42074 809570
rect 40907 805084 40973 805085
rect 40907 805020 40908 805084
rect 40972 805020 40973 805084
rect 40907 805019 40973 805020
rect 40910 793525 40970 805019
rect 41091 800732 41157 800733
rect 41091 800668 41092 800732
rect 41156 800668 41157 800732
rect 41091 800667 41157 800668
rect 41094 796245 41154 800667
rect 41091 796244 41157 796245
rect 41091 796180 41092 796244
rect 41156 796180 41157 796244
rect 41091 796179 41157 796180
rect 40907 793524 40973 793525
rect 40907 793460 40908 793524
rect 40972 793460 40973 793524
rect 40907 793459 40973 793460
rect 40723 789988 40789 789989
rect 40723 789924 40724 789988
rect 40788 789924 40789 789988
rect 40723 789923 40789 789924
rect 41462 788221 41522 809510
rect 41827 809300 41893 809301
rect 41827 809236 41828 809300
rect 41892 809236 41893 809300
rect 41827 809235 41893 809236
rect 41830 804570 41890 809235
rect 41646 804510 41890 804570
rect 41646 791621 41706 804510
rect 41827 803860 41893 803861
rect 41827 803796 41828 803860
rect 41892 803796 41893 803860
rect 41827 803795 41893 803796
rect 41643 791620 41709 791621
rect 41643 791556 41644 791620
rect 41708 791556 41709 791620
rect 41643 791555 41709 791556
rect 41459 788220 41525 788221
rect 41459 788156 41460 788220
rect 41524 788156 41525 788220
rect 41459 788155 41525 788156
rect 41830 787949 41890 803795
rect 41827 787948 41893 787949
rect 41827 787884 41828 787948
rect 41892 787884 41893 787948
rect 41827 787883 41893 787884
rect 673870 772445 673930 872203
rect 675342 869685 675402 873971
rect 675339 869684 675405 869685
rect 675339 869620 675340 869684
rect 675404 869620 675405 869684
rect 675339 869619 675405 869620
rect 675891 869684 675957 869685
rect 675891 869620 675892 869684
rect 675956 869620 675957 869684
rect 675891 869619 675957 869620
rect 674419 854316 674485 854317
rect 674419 854252 674420 854316
rect 674484 854252 674485 854316
rect 674419 854251 674485 854252
rect 674235 784276 674301 784277
rect 674235 784212 674236 784276
rect 674300 784212 674301 784276
rect 674235 784211 674301 784212
rect 673867 772444 673933 772445
rect 673867 772380 673868 772444
rect 673932 772380 673933 772444
rect 673867 772379 673933 772380
rect 41459 769860 41525 769861
rect 41459 769796 41460 769860
rect 41524 769796 41525 769860
rect 41459 769795 41525 769796
rect 40907 765780 40973 765781
rect 40907 765716 40908 765780
rect 40972 765716 40973 765780
rect 40907 765715 40973 765716
rect 40539 765372 40605 765373
rect 40539 765308 40540 765372
rect 40604 765308 40605 765372
rect 40539 765307 40605 765308
rect 40542 749461 40602 765307
rect 40723 764964 40789 764965
rect 40723 764900 40724 764964
rect 40788 764900 40789 764964
rect 40723 764899 40789 764900
rect 40726 750413 40786 764899
rect 40910 751093 40970 765715
rect 40907 751092 40973 751093
rect 40907 751028 40908 751092
rect 40972 751028 40973 751092
rect 40907 751027 40973 751028
rect 40723 750412 40789 750413
rect 40723 750348 40724 750412
rect 40788 750348 40789 750412
rect 40723 750347 40789 750348
rect 40539 749460 40605 749461
rect 40539 749396 40540 749460
rect 40604 749396 40605 749460
rect 40539 749395 40605 749396
rect 41462 743749 41522 769795
rect 41827 759660 41893 759661
rect 41827 759596 41828 759660
rect 41892 759596 41893 759660
rect 41827 759595 41893 759596
rect 41643 757756 41709 757757
rect 41643 757692 41644 757756
rect 41708 757692 41709 757756
rect 41643 757691 41709 757692
rect 41646 745109 41706 757691
rect 41830 745653 41890 759595
rect 42195 751636 42261 751637
rect 42195 751572 42196 751636
rect 42260 751572 42261 751636
rect 42195 751571 42261 751572
rect 42198 750549 42258 751571
rect 42195 750548 42261 750549
rect 42195 750484 42196 750548
rect 42260 750484 42261 750548
rect 42195 750483 42261 750484
rect 41827 745652 41893 745653
rect 41827 745588 41828 745652
rect 41892 745588 41893 745652
rect 41827 745587 41893 745588
rect 41643 745108 41709 745109
rect 41643 745044 41644 745108
rect 41708 745044 41709 745108
rect 41643 745043 41709 745044
rect 41459 743748 41525 743749
rect 41459 743684 41460 743748
rect 41524 743684 41525 743748
rect 41459 743683 41525 743684
rect 41827 725796 41893 725797
rect 41827 725732 41828 725796
rect 41892 725732 41893 725796
rect 41827 725731 41893 725732
rect 41830 725250 41890 725731
rect 41462 725190 41890 725250
rect 40723 721772 40789 721773
rect 40723 721708 40724 721772
rect 40788 721708 40789 721772
rect 40723 721707 40789 721708
rect 40907 721772 40973 721773
rect 40907 721708 40908 721772
rect 40972 721708 40973 721772
rect 40907 721707 40973 721708
rect 40539 718588 40605 718589
rect 40539 718524 40540 718588
rect 40604 718524 40605 718588
rect 40539 718523 40605 718524
rect 40355 714236 40421 714237
rect 40355 714172 40356 714236
rect 40420 714172 40421 714236
rect 40355 714171 40421 714172
rect 40358 712197 40418 714171
rect 40355 712196 40421 712197
rect 40355 712132 40356 712196
rect 40420 712132 40421 712196
rect 40355 712131 40421 712132
rect 40542 707301 40602 718523
rect 40726 709477 40786 721707
rect 40723 709476 40789 709477
rect 40723 709412 40724 709476
rect 40788 709412 40789 709476
rect 40723 709411 40789 709412
rect 40910 708525 40970 721707
rect 40907 708524 40973 708525
rect 40907 708460 40908 708524
rect 40972 708460 40973 708524
rect 40907 708459 40973 708460
rect 40539 707300 40605 707301
rect 40539 707236 40540 707300
rect 40604 707236 40605 707300
rect 40539 707235 40605 707236
rect 41462 702541 41522 725190
rect 41643 721772 41709 721773
rect 41643 721708 41644 721772
rect 41708 721708 41709 721772
rect 41643 721707 41709 721708
rect 41459 702540 41525 702541
rect 41459 702476 41460 702540
rect 41524 702476 41525 702540
rect 41459 702475 41525 702476
rect 41646 701453 41706 721707
rect 41827 716820 41893 716821
rect 41827 716756 41828 716820
rect 41892 716756 41893 716820
rect 41827 716755 41893 716756
rect 41643 701452 41709 701453
rect 41643 701388 41644 701452
rect 41708 701388 41709 701452
rect 41643 701387 41709 701388
rect 41830 701181 41890 716755
rect 42563 714780 42629 714781
rect 42563 714716 42564 714780
rect 42628 714716 42629 714780
rect 42563 714715 42629 714716
rect 42379 714236 42445 714237
rect 42379 714172 42380 714236
rect 42444 714172 42445 714236
rect 42379 714171 42445 714172
rect 42011 713964 42077 713965
rect 42011 713900 42012 713964
rect 42076 713900 42077 713964
rect 42011 713899 42077 713900
rect 42014 710429 42074 713899
rect 42011 710428 42077 710429
rect 42011 710364 42012 710428
rect 42076 710364 42077 710428
rect 42011 710363 42077 710364
rect 42382 706621 42442 714171
rect 42566 711653 42626 714715
rect 42563 711652 42629 711653
rect 42563 711588 42564 711652
rect 42628 711588 42629 711652
rect 42563 711587 42629 711588
rect 674238 709205 674298 784211
rect 674422 772037 674482 854251
rect 674971 780332 675037 780333
rect 674971 780268 674972 780332
rect 675036 780268 675037 780332
rect 674971 780267 675037 780268
rect 674974 773397 675034 780267
rect 675155 779924 675221 779925
rect 675155 779860 675156 779924
rect 675220 779860 675221 779924
rect 675155 779859 675221 779860
rect 675158 775437 675218 779859
rect 675155 775436 675221 775437
rect 675155 775372 675156 775436
rect 675220 775372 675221 775436
rect 675155 775371 675221 775372
rect 674971 773396 675037 773397
rect 674971 773332 674972 773396
rect 675036 773332 675037 773396
rect 674971 773331 675037 773332
rect 674419 772036 674485 772037
rect 674419 771972 674420 772036
rect 674484 771972 674485 772036
rect 674419 771971 674485 771972
rect 675894 771357 675954 869619
rect 676078 772717 676138 877099
rect 676995 876484 677061 876485
rect 676995 876420 676996 876484
rect 677060 876420 677061 876484
rect 676995 876419 677061 876420
rect 676811 872812 676877 872813
rect 676811 872748 676812 872812
rect 676876 872748 676877 872812
rect 676811 872747 676877 872748
rect 676075 772716 676141 772717
rect 676075 772652 676076 772716
rect 676140 772652 676141 772716
rect 676075 772651 676141 772652
rect 675891 771356 675957 771357
rect 675891 771292 675892 771356
rect 675956 771292 675957 771356
rect 675891 771291 675957 771292
rect 676814 756270 676874 872747
rect 676998 761837 677058 876419
rect 676995 761836 677061 761837
rect 676995 761772 676996 761836
rect 677060 761772 677061 761836
rect 676995 761771 677061 761772
rect 676630 756210 676874 756270
rect 675891 753812 675957 753813
rect 675891 753748 675892 753812
rect 675956 753810 675957 753812
rect 676630 753810 676690 756210
rect 675956 753750 676690 753810
rect 675956 753748 675957 753750
rect 675891 753747 675957 753748
rect 676075 751092 676141 751093
rect 676075 751028 676076 751092
rect 676140 751090 676141 751092
rect 676140 751030 676322 751090
rect 676140 751028 676141 751030
rect 676075 751027 676141 751028
rect 676262 746610 676322 751030
rect 676262 746550 677058 746610
rect 675523 743068 675589 743069
rect 675523 743004 675524 743068
rect 675588 743004 675589 743068
rect 675523 743003 675589 743004
rect 674419 738716 674485 738717
rect 674419 738652 674420 738716
rect 674484 738652 674485 738716
rect 674419 738651 674485 738652
rect 674235 709204 674301 709205
rect 674235 709140 674236 709204
rect 674300 709140 674301 709204
rect 674235 709139 674301 709140
rect 42379 706620 42445 706621
rect 42379 706556 42380 706620
rect 42444 706556 42445 706620
rect 42379 706555 42445 706556
rect 41827 701180 41893 701181
rect 41827 701116 41828 701180
rect 41892 701116 41893 701180
rect 41827 701115 41893 701116
rect 674051 694652 674117 694653
rect 674051 694588 674052 694652
rect 674116 694588 674117 694652
rect 674051 694587 674117 694588
rect 41827 682412 41893 682413
rect 41827 682410 41828 682412
rect 41462 682350 41828 682410
rect 40539 678992 40605 678993
rect 40539 678928 40540 678992
rect 40604 678928 40605 678992
rect 40539 678927 40605 678928
rect 40723 678992 40789 678993
rect 40723 678928 40724 678992
rect 40788 678928 40789 678992
rect 40723 678927 40789 678928
rect 40542 662693 40602 678927
rect 40726 666501 40786 678927
rect 41091 671260 41157 671261
rect 41091 671196 41092 671260
rect 41156 671196 41157 671260
rect 41091 671195 41157 671196
rect 40907 670988 40973 670989
rect 40907 670924 40908 670988
rect 40972 670924 40973 670988
rect 40907 670923 40973 670924
rect 40910 667997 40970 670923
rect 40907 667996 40973 667997
rect 40907 667932 40908 667996
rect 40972 667932 40973 667996
rect 40907 667931 40973 667932
rect 41094 667453 41154 671195
rect 41091 667452 41157 667453
rect 41091 667388 41092 667452
rect 41156 667388 41157 667452
rect 41091 667387 41157 667388
rect 40723 666500 40789 666501
rect 40723 666436 40724 666500
rect 40788 666436 40789 666500
rect 40723 666435 40789 666436
rect 40539 662692 40605 662693
rect 40539 662628 40540 662692
rect 40604 662628 40605 662692
rect 40539 662627 40605 662628
rect 41462 659701 41522 682350
rect 41827 682348 41828 682350
rect 41892 682348 41893 682412
rect 41827 682347 41893 682348
rect 41827 680372 41893 680373
rect 41827 680370 41828 680372
rect 41646 680310 41828 680370
rect 41459 659700 41525 659701
rect 41459 659636 41460 659700
rect 41524 659636 41525 659700
rect 41459 659635 41525 659636
rect 41646 658613 41706 680310
rect 41827 680308 41828 680310
rect 41892 680308 41893 680372
rect 41827 680307 41893 680308
rect 41827 672756 41893 672757
rect 41827 672692 41828 672756
rect 41892 672692 41893 672756
rect 41827 672691 41893 672692
rect 41643 658612 41709 658613
rect 41643 658548 41644 658612
rect 41708 658548 41709 658612
rect 41643 658547 41709 658548
rect 41830 658341 41890 672691
rect 42011 666500 42077 666501
rect 42011 666436 42012 666500
rect 42076 666436 42077 666500
rect 42011 666435 42077 666436
rect 42014 664053 42074 666435
rect 42011 664052 42077 664053
rect 42011 663988 42012 664052
rect 42076 663988 42077 664052
rect 42011 663987 42077 663988
rect 41827 658340 41893 658341
rect 41827 658276 41828 658340
rect 41892 658276 41893 658340
rect 41827 658275 41893 658276
rect 41459 640660 41525 640661
rect 41459 640596 41460 640660
rect 41524 640596 41525 640660
rect 41459 640595 41525 640596
rect 40539 636988 40605 636989
rect 40539 636924 40540 636988
rect 40604 636924 40605 636988
rect 40539 636923 40605 636924
rect 40542 619037 40602 636923
rect 40907 636172 40973 636173
rect 40907 636108 40908 636172
rect 40972 636108 40973 636172
rect 40907 636107 40973 636108
rect 40723 635764 40789 635765
rect 40723 635700 40724 635764
rect 40788 635700 40789 635764
rect 40723 635699 40789 635700
rect 40726 619853 40786 635699
rect 40910 625293 40970 636107
rect 40907 625292 40973 625293
rect 40907 625228 40908 625292
rect 40972 625228 40973 625292
rect 40907 625227 40973 625228
rect 40723 619852 40789 619853
rect 40723 619788 40724 619852
rect 40788 619788 40789 619852
rect 40723 619787 40789 619788
rect 40539 619036 40605 619037
rect 40539 618972 40540 619036
rect 40604 618972 40605 619036
rect 40539 618971 40605 618972
rect 41462 616045 41522 640595
rect 41643 637396 41709 637397
rect 41643 637332 41644 637396
rect 41708 637332 41709 637396
rect 41643 637331 41709 637332
rect 41646 618270 41706 637331
rect 674054 636853 674114 694587
rect 674422 674117 674482 738651
rect 674603 738172 674669 738173
rect 674603 738108 674604 738172
rect 674668 738108 674669 738172
rect 674603 738107 674669 738108
rect 674606 725933 674666 738107
rect 675526 736950 675586 743003
rect 675342 736890 675586 736950
rect 675342 735181 675402 736890
rect 675339 735180 675405 735181
rect 675339 735116 675340 735180
rect 675404 735116 675405 735180
rect 675339 735115 675405 735116
rect 676811 733684 676877 733685
rect 676811 733620 676812 733684
rect 676876 733620 676877 733684
rect 676811 733619 676877 733620
rect 674603 725932 674669 725933
rect 674603 725868 674604 725932
rect 674668 725868 674669 725932
rect 674603 725867 674669 725868
rect 676075 721580 676141 721581
rect 676075 721516 676076 721580
rect 676140 721516 676141 721580
rect 676075 721515 676141 721516
rect 675339 696828 675405 696829
rect 675339 696764 675340 696828
rect 675404 696764 675405 696828
rect 675339 696763 675405 696764
rect 674603 693020 674669 693021
rect 674603 692956 674604 693020
rect 674668 692956 674669 693020
rect 674603 692955 674669 692956
rect 674419 674116 674485 674117
rect 674419 674052 674420 674116
rect 674484 674052 674485 674116
rect 674419 674051 674485 674052
rect 674235 648956 674301 648957
rect 674235 648892 674236 648956
rect 674300 648892 674301 648956
rect 674235 648891 674301 648892
rect 674051 636852 674117 636853
rect 674051 636788 674052 636852
rect 674116 636788 674117 636852
rect 674051 636787 674117 636788
rect 41827 635356 41893 635357
rect 41827 635292 41828 635356
rect 41892 635292 41893 635356
rect 41827 635291 41893 635292
rect 41830 618765 41890 635291
rect 42195 626788 42261 626789
rect 42195 626724 42196 626788
rect 42260 626724 42261 626788
rect 42195 626723 42261 626724
rect 42011 625292 42077 625293
rect 42011 625228 42012 625292
rect 42076 625228 42077 625292
rect 42011 625227 42077 625228
rect 42014 621485 42074 625227
rect 42011 621484 42077 621485
rect 42011 621420 42012 621484
rect 42076 621420 42077 621484
rect 42011 621419 42077 621420
rect 42198 620261 42258 626723
rect 42195 620260 42261 620261
rect 42195 620196 42196 620260
rect 42260 620196 42261 620260
rect 42195 620195 42261 620196
rect 41827 618764 41893 618765
rect 41827 618700 41828 618764
rect 41892 618700 41893 618764
rect 41827 618699 41893 618700
rect 41646 618210 41890 618270
rect 41459 616044 41525 616045
rect 41459 615980 41460 616044
rect 41524 615980 41525 616044
rect 41459 615979 41525 615980
rect 41830 612781 41890 618210
rect 671475 616860 671541 616861
rect 671475 616796 671476 616860
rect 671540 616796 671541 616860
rect 671475 616795 671541 616796
rect 41827 612780 41893 612781
rect 41827 612716 41828 612780
rect 41892 612716 41893 612780
rect 41827 612715 41893 612716
rect 671478 608701 671538 616795
rect 671475 608700 671541 608701
rect 671475 608636 671476 608700
rect 671540 608636 671541 608700
rect 671475 608635 671541 608636
rect 42011 596460 42077 596461
rect 42011 596396 42012 596460
rect 42076 596396 42077 596460
rect 42011 596395 42077 596396
rect 41827 596052 41893 596053
rect 41827 596050 41828 596052
rect 41462 595990 41828 596050
rect 40723 589660 40789 589661
rect 40723 589596 40724 589660
rect 40788 589596 40789 589660
rect 40723 589595 40789 589596
rect 40539 589388 40605 589389
rect 40539 589324 40540 589388
rect 40604 589324 40605 589388
rect 40539 589323 40605 589324
rect 40355 584628 40421 584629
rect 40355 584564 40356 584628
rect 40420 584564 40421 584628
rect 40355 584563 40421 584564
rect 40358 580277 40418 584563
rect 40355 580276 40421 580277
rect 40355 580212 40356 580276
rect 40420 580212 40421 580276
rect 40355 580211 40421 580212
rect 40542 575517 40602 589323
rect 40539 575516 40605 575517
rect 40539 575452 40540 575516
rect 40604 575452 40605 575516
rect 40539 575451 40605 575452
rect 40726 574701 40786 589595
rect 40907 589524 40973 589525
rect 40907 589460 40908 589524
rect 40972 589460 40973 589524
rect 40907 589459 40973 589460
rect 40910 580005 40970 589459
rect 41091 584900 41157 584901
rect 41091 584836 41092 584900
rect 41156 584836 41157 584900
rect 41091 584835 41157 584836
rect 41094 580549 41154 584835
rect 41091 580548 41157 580549
rect 41091 580484 41092 580548
rect 41156 580484 41157 580548
rect 41091 580483 41157 580484
rect 40907 580004 40973 580005
rect 40907 579940 40908 580004
rect 40972 579940 40973 580004
rect 40907 579939 40973 579940
rect 40723 574700 40789 574701
rect 40723 574636 40724 574700
rect 40788 574636 40789 574700
rect 40723 574635 40789 574636
rect 41462 574021 41522 595990
rect 41827 595988 41828 595990
rect 41892 595988 41893 596052
rect 41827 595987 41893 595988
rect 42014 589290 42074 596395
rect 41646 589230 42074 589290
rect 41459 574020 41525 574021
rect 41459 573956 41460 574020
rect 41524 573956 41525 574020
rect 41459 573955 41525 573956
rect 41646 571981 41706 589230
rect 41827 587212 41893 587213
rect 41827 587148 41828 587212
rect 41892 587148 41893 587212
rect 41827 587147 41893 587148
rect 41830 572253 41890 587147
rect 42011 584900 42077 584901
rect 42011 584836 42012 584900
rect 42076 584836 42077 584900
rect 42011 584835 42077 584836
rect 42014 582589 42074 584835
rect 42563 584628 42629 584629
rect 42563 584564 42564 584628
rect 42628 584564 42629 584628
rect 42563 584563 42629 584564
rect 42011 582588 42077 582589
rect 42011 582524 42012 582588
rect 42076 582524 42077 582588
rect 42011 582523 42077 582524
rect 42566 576605 42626 584563
rect 42563 576604 42629 576605
rect 42563 576540 42564 576604
rect 42628 576540 42629 576604
rect 42563 576539 42629 576540
rect 674238 573341 674298 648891
rect 674606 623661 674666 692955
rect 675342 685949 675402 696763
rect 675339 685948 675405 685949
rect 675339 685884 675340 685948
rect 675404 685884 675405 685948
rect 675339 685883 675405 685884
rect 676078 681869 676138 721515
rect 676075 681868 676141 681869
rect 676075 681804 676076 681868
rect 676140 681804 676141 681868
rect 676075 681803 676141 681804
rect 676814 665413 676874 733619
rect 676998 714870 677058 746550
rect 676998 714810 677794 714870
rect 677734 713493 677794 714810
rect 677731 713492 677797 713493
rect 677731 713428 677732 713492
rect 677796 713428 677797 713492
rect 677731 713427 677797 713428
rect 676995 694108 677061 694109
rect 676995 694044 676996 694108
rect 677060 694044 677061 694108
rect 676995 694043 677061 694044
rect 676998 666637 677058 694043
rect 676995 666636 677061 666637
rect 676995 666572 676996 666636
rect 677060 666572 677061 666636
rect 676995 666571 677061 666572
rect 676811 665412 676877 665413
rect 676811 665348 676812 665412
rect 676876 665348 676877 665412
rect 676811 665347 676877 665348
rect 675523 652900 675589 652901
rect 675523 652836 675524 652900
rect 675588 652836 675589 652900
rect 675523 652835 675589 652836
rect 675155 650180 675221 650181
rect 675155 650116 675156 650180
rect 675220 650116 675221 650180
rect 675155 650115 675221 650116
rect 675158 648005 675218 650115
rect 675155 648004 675221 648005
rect 675155 647940 675156 648004
rect 675220 647940 675221 648004
rect 675155 647939 675221 647940
rect 674971 643924 675037 643925
rect 674971 643860 674972 643924
rect 675036 643860 675037 643924
rect 674971 643859 675037 643860
rect 674974 638213 675034 643859
rect 674971 638212 675037 638213
rect 674971 638148 674972 638212
rect 675036 638148 675037 638212
rect 674971 638147 675037 638148
rect 675526 637669 675586 652835
rect 676811 640252 676877 640253
rect 676811 640188 676812 640252
rect 676876 640188 676877 640252
rect 676811 640187 676877 640188
rect 675523 637668 675589 637669
rect 675523 637604 675524 637668
rect 675588 637604 675589 637668
rect 675523 637603 675589 637604
rect 675155 631412 675221 631413
rect 675155 631348 675156 631412
rect 675220 631348 675221 631412
rect 675155 631347 675221 631348
rect 676075 631412 676141 631413
rect 676075 631348 676076 631412
rect 676140 631348 676141 631412
rect 676075 631347 676141 631348
rect 674603 623660 674669 623661
rect 674603 623596 674604 623660
rect 674668 623596 674669 623660
rect 674603 623595 674669 623596
rect 674419 604484 674485 604485
rect 674419 604420 674420 604484
rect 674484 604420 674485 604484
rect 674419 604419 674485 604420
rect 674235 573340 674301 573341
rect 674235 573276 674236 573340
rect 674300 573276 674301 573340
rect 674235 573275 674301 573276
rect 41827 572252 41893 572253
rect 41827 572188 41828 572252
rect 41892 572188 41893 572252
rect 41827 572187 41893 572188
rect 41643 571980 41709 571981
rect 41643 571916 41644 571980
rect 41708 571916 41709 571980
rect 41643 571915 41709 571916
rect 42379 554028 42445 554029
rect 42379 553964 42380 554028
rect 42444 553964 42445 554028
rect 42379 553963 42445 553964
rect 42195 552804 42261 552805
rect 42195 552740 42196 552804
rect 42260 552740 42261 552804
rect 42195 552739 42261 552740
rect 41827 550492 41893 550493
rect 41827 550428 41828 550492
rect 41892 550428 41893 550492
rect 41827 550427 41893 550428
rect 41643 546412 41709 546413
rect 41643 546348 41644 546412
rect 41708 546348 41709 546412
rect 41643 546347 41709 546348
rect 41459 546140 41525 546141
rect 41459 546076 41460 546140
rect 41524 546076 41525 546140
rect 41459 546075 41525 546076
rect 40907 545868 40973 545869
rect 40907 545804 40908 545868
rect 40972 545804 40973 545868
rect 40907 545803 40973 545804
rect 40723 545596 40789 545597
rect 40723 545532 40724 545596
rect 40788 545532 40789 545596
rect 40723 545531 40789 545532
rect 40539 545324 40605 545325
rect 40539 545260 40540 545324
rect 40604 545260 40605 545324
rect 40539 545259 40605 545260
rect 40542 533357 40602 545259
rect 40726 536893 40786 545531
rect 40910 538253 40970 545803
rect 40907 538252 40973 538253
rect 40907 538188 40908 538252
rect 40972 538188 40973 538252
rect 40907 538187 40973 538188
rect 40723 536892 40789 536893
rect 40723 536828 40724 536892
rect 40788 536828 40789 536892
rect 40723 536827 40789 536828
rect 40539 533356 40605 533357
rect 40539 533292 40540 533356
rect 40604 533292 40605 533356
rect 40539 533291 40605 533292
rect 41462 527645 41522 546075
rect 41646 529821 41706 546347
rect 41830 545869 41890 550427
rect 41827 545868 41893 545869
rect 41827 545804 41828 545868
rect 41892 545804 41893 545868
rect 41827 545803 41893 545804
rect 42198 543750 42258 552739
rect 42382 546141 42442 553963
rect 42379 546140 42445 546141
rect 42379 546076 42380 546140
rect 42444 546076 42445 546140
rect 42379 546075 42445 546076
rect 41830 543690 42258 543750
rect 41830 532677 41890 543690
rect 41827 532676 41893 532677
rect 41827 532612 41828 532676
rect 41892 532612 41893 532676
rect 41827 532611 41893 532612
rect 41643 529820 41709 529821
rect 41643 529756 41644 529820
rect 41708 529756 41709 529820
rect 41643 529755 41709 529756
rect 674422 528869 674482 604419
rect 674603 602988 674669 602989
rect 674603 602924 674604 602988
rect 674668 602924 674669 602988
rect 674603 602923 674669 602924
rect 674419 528868 674485 528869
rect 674419 528804 674420 528868
rect 674484 528804 674485 528868
rect 674419 528803 674485 528804
rect 41459 527644 41525 527645
rect 41459 527580 41460 527644
rect 41524 527580 41525 527644
rect 41459 527579 41525 527580
rect 674606 527101 674666 602923
rect 675158 592653 675218 631347
rect 676078 592925 676138 631347
rect 676075 592924 676141 592925
rect 676075 592860 676076 592924
rect 676140 592860 676141 592924
rect 676075 592859 676141 592860
rect 675155 592652 675221 592653
rect 675155 592588 675156 592652
rect 675220 592588 675221 592652
rect 675155 592587 675221 592588
rect 676075 586260 676141 586261
rect 676075 586196 676076 586260
rect 676140 586196 676141 586260
rect 676075 586195 676141 586196
rect 675339 561916 675405 561917
rect 675339 561852 675340 561916
rect 675404 561852 675405 561916
rect 675339 561851 675405 561852
rect 675155 550356 675221 550357
rect 675155 550292 675156 550356
rect 675220 550292 675221 550356
rect 675155 550291 675221 550292
rect 675158 545869 675218 550291
rect 675342 547637 675402 561851
rect 675523 559468 675589 559469
rect 675523 559404 675524 559468
rect 675588 559404 675589 559468
rect 675523 559403 675589 559404
rect 675526 547909 675586 559403
rect 675523 547908 675589 547909
rect 675523 547844 675524 547908
rect 675588 547844 675589 547908
rect 675523 547843 675589 547844
rect 675339 547636 675405 547637
rect 675339 547572 675340 547636
rect 675404 547572 675405 547636
rect 675339 547571 675405 547572
rect 675155 545868 675221 545869
rect 675155 545804 675156 545868
rect 675220 545804 675221 545868
rect 675155 545803 675221 545804
rect 676078 545189 676138 586195
rect 676814 576469 676874 640187
rect 676811 576468 676877 576469
rect 676811 576404 676812 576468
rect 676876 576404 676877 576468
rect 676811 576403 676877 576404
rect 676995 571572 677061 571573
rect 676995 571508 676996 571572
rect 677060 571508 677061 571572
rect 676995 571507 677061 571508
rect 676811 559060 676877 559061
rect 676811 558996 676812 559060
rect 676876 558996 676877 559060
rect 676811 558995 676877 558996
rect 676075 545188 676141 545189
rect 676075 545124 676076 545188
rect 676140 545124 676141 545188
rect 676075 545123 676141 545124
rect 674603 527100 674669 527101
rect 674603 527036 674604 527100
rect 674668 527036 674669 527100
rect 674603 527035 674669 527036
rect 673867 525876 673933 525877
rect 673867 525812 673868 525876
rect 673932 525812 673933 525876
rect 673867 525811 673933 525812
rect 41459 431220 41525 431221
rect 41459 431156 41460 431220
rect 41524 431156 41525 431220
rect 41459 431155 41525 431156
rect 41462 428263 41522 431155
rect 41459 428262 41525 428263
rect 41459 428198 41460 428262
rect 41524 428198 41525 428262
rect 41459 428197 41525 428198
rect 41827 426460 41893 426461
rect 41827 426396 41828 426460
rect 41892 426396 41893 426460
rect 41827 426395 41893 426396
rect 41830 426050 41890 426395
rect 41462 425990 41890 426050
rect 40723 422312 40789 422313
rect 40723 422248 40724 422312
rect 40788 422248 40789 422312
rect 40723 422247 40789 422248
rect 40539 418708 40605 418709
rect 40539 418644 40540 418708
rect 40604 418644 40605 418708
rect 40539 418643 40605 418644
rect 40542 403885 40602 418643
rect 40726 407557 40786 422247
rect 40723 407556 40789 407557
rect 40723 407492 40724 407556
rect 40788 407492 40789 407556
rect 40723 407491 40789 407492
rect 40539 403884 40605 403885
rect 40539 403820 40540 403884
rect 40604 403820 40605 403884
rect 40539 403819 40605 403820
rect 41462 400077 41522 425990
rect 41827 425644 41893 425645
rect 41827 425580 41828 425644
rect 41892 425580 41893 425644
rect 41827 425579 41893 425580
rect 41830 425370 41890 425579
rect 41646 425310 41890 425370
rect 41459 400076 41525 400077
rect 41459 400012 41460 400076
rect 41524 400012 41525 400076
rect 41459 400011 41525 400012
rect 41646 398850 41706 425310
rect 42011 421972 42077 421973
rect 42011 421908 42012 421972
rect 42076 421908 42077 421972
rect 42011 421907 42077 421908
rect 42014 418709 42074 421907
rect 42011 418708 42077 418709
rect 42011 418644 42012 418708
rect 42076 418644 42077 418708
rect 42011 418643 42077 418644
rect 41827 418436 41893 418437
rect 41827 418372 41828 418436
rect 41892 418372 41893 418436
rect 41827 418371 41893 418372
rect 41830 401981 41890 418371
rect 41827 401980 41893 401981
rect 41827 401916 41828 401980
rect 41892 401916 41893 401980
rect 41827 401915 41893 401916
rect 41827 398852 41893 398853
rect 41827 398850 41828 398852
rect 41646 398790 41828 398850
rect 41827 398788 41828 398790
rect 41892 398788 41893 398852
rect 41827 398787 41893 398788
rect 672947 394636 673013 394637
rect 672947 394572 672948 394636
rect 673012 394572 673013 394636
rect 672947 394571 673013 394572
rect 41459 382260 41525 382261
rect 41459 382196 41460 382260
rect 41524 382196 41525 382260
rect 41459 382195 41525 382196
rect 40907 379404 40973 379405
rect 40907 379340 40908 379404
rect 40972 379340 40973 379404
rect 40907 379339 40973 379340
rect 40539 378588 40605 378589
rect 40539 378524 40540 378588
rect 40604 378524 40605 378588
rect 40539 378523 40605 378524
rect 40542 360637 40602 378523
rect 40723 378180 40789 378181
rect 40723 378116 40724 378180
rect 40788 378116 40789 378180
rect 40723 378115 40789 378116
rect 40726 363765 40786 378115
rect 40910 365669 40970 379339
rect 40907 365668 40973 365669
rect 40907 365604 40908 365668
rect 40972 365604 40973 365668
rect 40907 365603 40973 365604
rect 40723 363764 40789 363765
rect 40723 363700 40724 363764
rect 40788 363700 40789 363764
rect 40723 363699 40789 363700
rect 40539 360636 40605 360637
rect 40539 360572 40540 360636
rect 40604 360572 40605 360636
rect 40539 360571 40605 360572
rect 41462 356965 41522 382195
rect 41643 380220 41709 380221
rect 41643 380156 41644 380220
rect 41708 380156 41709 380220
rect 41643 380155 41709 380156
rect 41646 358730 41706 380155
rect 41827 378996 41893 378997
rect 41827 378932 41828 378996
rect 41892 378932 41893 378996
rect 41827 378931 41893 378932
rect 41830 364350 41890 378931
rect 41830 364290 42074 364350
rect 41827 358732 41893 358733
rect 41827 358730 41828 358732
rect 41646 358670 41828 358730
rect 41827 358668 41828 358670
rect 41892 358668 41893 358732
rect 41827 358667 41893 358668
rect 41459 356964 41525 356965
rect 41459 356900 41460 356964
rect 41524 356900 41525 356964
rect 41459 356899 41525 356900
rect 42014 355741 42074 364290
rect 42011 355740 42077 355741
rect 42011 355676 42012 355740
rect 42076 355676 42077 355740
rect 42011 355675 42077 355676
rect 671843 345268 671909 345269
rect 671843 345204 671844 345268
rect 671908 345204 671909 345268
rect 671843 345203 671909 345204
rect 671291 344996 671357 344997
rect 671291 344932 671292 344996
rect 671356 344932 671357 344996
rect 671291 344931 671357 344932
rect 41459 339828 41525 339829
rect 41459 339764 41460 339828
rect 41524 339764 41525 339828
rect 41459 339763 41525 339764
rect 40539 337380 40605 337381
rect 40539 337316 40540 337380
rect 40604 337316 40605 337380
rect 40539 337315 40605 337316
rect 40542 313037 40602 337315
rect 40723 336156 40789 336157
rect 40723 336092 40724 336156
rect 40788 336092 40789 336156
rect 40723 336091 40789 336092
rect 40726 322829 40786 336091
rect 40723 322828 40789 322829
rect 40723 322764 40724 322828
rect 40788 322764 40789 322828
rect 40723 322763 40789 322764
rect 41462 313717 41522 339763
rect 41827 339556 41893 339557
rect 41827 339492 41828 339556
rect 41892 339492 41893 339556
rect 41827 339491 41893 339492
rect 41643 338604 41709 338605
rect 41643 338540 41644 338604
rect 41708 338540 41709 338604
rect 41643 338539 41709 338540
rect 41646 316050 41706 338539
rect 41830 324869 41890 339491
rect 41827 324868 41893 324869
rect 41827 324804 41828 324868
rect 41892 324804 41893 324868
rect 41827 324803 41893 324804
rect 41646 315990 41890 316050
rect 41830 315621 41890 315990
rect 41827 315620 41893 315621
rect 41827 315556 41828 315620
rect 41892 315556 41893 315620
rect 41827 315555 41893 315556
rect 41459 313716 41525 313717
rect 41459 313652 41460 313716
rect 41524 313652 41525 313716
rect 41459 313651 41525 313652
rect 40539 313036 40605 313037
rect 40539 312972 40540 313036
rect 40604 312972 40605 313036
rect 40539 312971 40605 312972
rect 41827 296852 41893 296853
rect 41827 296788 41828 296852
rect 41892 296788 41893 296852
rect 41827 296787 41893 296788
rect 40539 292592 40605 292593
rect 40539 292528 40540 292592
rect 40604 292528 40605 292592
rect 40539 292527 40605 292528
rect 40723 292592 40789 292593
rect 40723 292528 40724 292592
rect 40788 292528 40789 292592
rect 40723 292527 40789 292528
rect 40907 292592 40973 292593
rect 40907 292528 40908 292592
rect 40972 292528 40973 292592
rect 41830 292590 41890 296787
rect 42011 296444 42077 296445
rect 42011 296380 42012 296444
rect 42076 296380 42077 296444
rect 42011 296379 42077 296380
rect 40907 292527 40973 292528
rect 41462 292530 41890 292590
rect 40542 273461 40602 292527
rect 40726 277405 40786 292527
rect 40910 277949 40970 292527
rect 40907 277948 40973 277949
rect 40907 277884 40908 277948
rect 40972 277884 40973 277948
rect 40907 277883 40973 277884
rect 40723 277404 40789 277405
rect 40723 277340 40724 277404
rect 40788 277340 40789 277404
rect 40723 277339 40789 277340
rect 40539 273460 40605 273461
rect 40539 273396 40540 273460
rect 40604 273396 40605 273460
rect 40539 273395 40605 273396
rect 41462 270469 41522 292530
rect 41827 292364 41893 292365
rect 41827 292300 41828 292364
rect 41892 292300 41893 292364
rect 41827 292299 41893 292300
rect 41830 272373 41890 292299
rect 42014 281485 42074 296379
rect 42011 281484 42077 281485
rect 42011 281420 42012 281484
rect 42076 281420 42077 281484
rect 42011 281419 42077 281420
rect 671294 278765 671354 344931
rect 671846 340509 671906 345203
rect 671843 340508 671909 340509
rect 671843 340444 671844 340508
rect 671908 340444 671909 340508
rect 671843 340443 671909 340444
rect 672950 278765 673010 394571
rect 671291 278764 671357 278765
rect 671291 278700 671292 278764
rect 671356 278700 671357 278764
rect 671291 278699 671357 278700
rect 672947 278764 673013 278765
rect 672947 278700 672948 278764
rect 673012 278700 673013 278764
rect 672947 278699 673013 278700
rect 673870 278629 673930 525811
rect 676814 500989 676874 558995
rect 676998 531453 677058 571507
rect 676995 531452 677061 531453
rect 676995 531388 676996 531452
rect 677060 531388 677061 531452
rect 676995 531387 677061 531388
rect 676811 500988 676877 500989
rect 676811 500924 676812 500988
rect 676876 500924 676877 500988
rect 676811 500923 676877 500924
rect 676075 398852 676141 398853
rect 676075 398788 676076 398852
rect 676140 398788 676141 398852
rect 676075 398787 676141 398788
rect 675891 389876 675957 389877
rect 675891 389812 675892 389876
rect 675956 389812 675957 389876
rect 675891 389811 675957 389812
rect 675707 388516 675773 388517
rect 675707 388452 675708 388516
rect 675772 388452 675773 388516
rect 675707 388451 675773 388452
rect 675710 378725 675770 388451
rect 675707 378724 675773 378725
rect 675707 378660 675708 378724
rect 675772 378660 675773 378724
rect 675707 378659 675773 378660
rect 674787 378044 674853 378045
rect 674787 377980 674788 378044
rect 674852 377980 674853 378044
rect 674787 377979 674853 377980
rect 674790 372605 674850 377979
rect 675894 373013 675954 389811
rect 676078 375053 676138 398787
rect 676259 396812 676325 396813
rect 676259 396748 676260 396812
rect 676324 396748 676325 396812
rect 676259 396747 676325 396748
rect 676262 384981 676322 396747
rect 676627 395180 676693 395181
rect 676627 395116 676628 395180
rect 676692 395116 676693 395180
rect 676627 395115 676693 395116
rect 676443 394772 676509 394773
rect 676443 394708 676444 394772
rect 676508 394708 676509 394772
rect 676443 394707 676509 394708
rect 676259 384980 676325 384981
rect 676259 384916 676260 384980
rect 676324 384916 676325 384980
rect 676259 384915 676325 384916
rect 676446 380629 676506 394707
rect 676443 380628 676509 380629
rect 676443 380564 676444 380628
rect 676508 380564 676509 380628
rect 676443 380563 676509 380564
rect 676630 377365 676690 395115
rect 676627 377364 676693 377365
rect 676627 377300 676628 377364
rect 676692 377300 676693 377364
rect 676627 377299 676693 377300
rect 676075 375052 676141 375053
rect 676075 374988 676076 375052
rect 676140 374988 676141 375052
rect 676075 374987 676141 374988
rect 675891 373012 675957 373013
rect 675891 372948 675892 373012
rect 675956 372948 675957 373012
rect 675891 372947 675957 372948
rect 674787 372604 674853 372605
rect 674787 372540 674788 372604
rect 674852 372540 674853 372604
rect 674787 372539 674853 372540
rect 675339 354244 675405 354245
rect 675339 354180 675340 354244
rect 675404 354180 675405 354244
rect 675339 354179 675405 354180
rect 675342 345541 675402 354179
rect 675523 353020 675589 353021
rect 675523 352956 675524 353020
rect 675588 352956 675589 353020
rect 675523 352955 675589 352956
rect 675339 345540 675405 345541
rect 675339 345476 675340 345540
rect 675404 345476 675405 345540
rect 675339 345475 675405 345476
rect 675526 337789 675586 352955
rect 675707 352204 675773 352205
rect 675707 352140 675708 352204
rect 675772 352140 675773 352204
rect 675707 352139 675773 352140
rect 675710 345810 675770 352139
rect 675891 351796 675957 351797
rect 675891 351732 675892 351796
rect 675956 351732 675957 351796
rect 675891 351731 675957 351732
rect 675894 351250 675954 351731
rect 675894 351190 676690 351250
rect 675891 350980 675957 350981
rect 675891 350916 675892 350980
rect 675956 350916 675957 350980
rect 675891 350915 675957 350916
rect 675894 350570 675954 350915
rect 675894 350510 676506 350570
rect 675891 350164 675957 350165
rect 675891 350100 675892 350164
rect 675956 350100 675957 350164
rect 675891 350099 675957 350100
rect 675894 349890 675954 350099
rect 675894 349830 676322 349890
rect 675710 345750 676138 345810
rect 675891 345540 675957 345541
rect 675891 345476 675892 345540
rect 675956 345476 675957 345540
rect 675891 345475 675957 345476
rect 675894 339421 675954 345475
rect 675891 339420 675957 339421
rect 675891 339356 675892 339420
rect 675956 339356 675957 339420
rect 675891 339355 675957 339356
rect 675523 337788 675589 337789
rect 675523 337724 675524 337788
rect 675588 337724 675589 337788
rect 675523 337723 675589 337724
rect 676078 326909 676138 345750
rect 676262 332349 676322 349830
rect 676446 336701 676506 350510
rect 676630 340373 676690 351190
rect 676627 340372 676693 340373
rect 676627 340308 676628 340372
rect 676692 340308 676693 340372
rect 676627 340307 676693 340308
rect 676443 336700 676509 336701
rect 676443 336636 676444 336700
rect 676508 336636 676509 336700
rect 676443 336635 676509 336636
rect 676259 332348 676325 332349
rect 676259 332284 676260 332348
rect 676324 332284 676325 332348
rect 676259 332283 676325 332284
rect 676075 326908 676141 326909
rect 676075 326844 676076 326908
rect 676140 326844 676141 326908
rect 676075 326843 676141 326844
rect 675891 308820 675957 308821
rect 675891 308756 675892 308820
rect 675956 308756 675957 308820
rect 675891 308755 675957 308756
rect 675894 302250 675954 308755
rect 676078 304979 676322 305010
rect 676075 304978 676322 304979
rect 676075 304914 676076 304978
rect 676140 304950 676322 304978
rect 676140 304914 676141 304950
rect 676075 304913 676141 304914
rect 676262 304330 676322 304950
rect 676262 304270 676690 304330
rect 676075 302972 676141 302973
rect 676075 302908 676076 302972
rect 676140 302970 676141 302972
rect 676140 302910 676322 302970
rect 676140 302908 676141 302910
rect 676075 302907 676141 302908
rect 675894 302190 676138 302250
rect 675891 299436 675957 299437
rect 675891 299372 675892 299436
rect 675956 299372 675957 299436
rect 675891 299371 675957 299372
rect 675707 297396 675773 297397
rect 675707 297332 675708 297396
rect 675772 297332 675773 297396
rect 675707 297331 675773 297332
rect 675523 296580 675589 296581
rect 675523 296516 675524 296580
rect 675588 296516 675589 296580
rect 675523 296515 675589 296516
rect 675526 295357 675586 296515
rect 675523 295356 675589 295357
rect 675523 295292 675524 295356
rect 675588 295292 675589 295356
rect 675523 295291 675589 295292
rect 675710 281621 675770 297331
rect 675894 282845 675954 299371
rect 676078 283661 676138 302190
rect 676262 291005 676322 302910
rect 676443 301612 676509 301613
rect 676443 301548 676444 301612
rect 676508 301548 676509 301612
rect 676443 301547 676509 301548
rect 676446 291549 676506 301547
rect 676443 291548 676509 291549
rect 676443 291484 676444 291548
rect 676508 291484 676509 291548
rect 676443 291483 676509 291484
rect 676259 291004 676325 291005
rect 676259 290940 676260 291004
rect 676324 290940 676325 291004
rect 676259 290939 676325 290940
rect 676630 287061 676690 304270
rect 676627 287060 676693 287061
rect 676627 286996 676628 287060
rect 676692 286996 676693 287060
rect 676627 286995 676693 286996
rect 676075 283660 676141 283661
rect 676075 283596 676076 283660
rect 676140 283596 676141 283660
rect 676075 283595 676141 283596
rect 675891 282844 675957 282845
rect 675891 282780 675892 282844
rect 675956 282780 675957 282844
rect 675891 282779 675957 282780
rect 675707 281620 675773 281621
rect 675707 281556 675708 281620
rect 675772 281556 675773 281620
rect 675707 281555 675773 281556
rect 673867 278628 673933 278629
rect 673867 278564 673868 278628
rect 673932 278564 673933 278628
rect 673867 278563 673933 278564
rect 673867 277676 673933 277677
rect 673867 277612 673868 277676
rect 673932 277612 673933 277676
rect 673867 277611 673933 277612
rect 41827 272372 41893 272373
rect 41827 272308 41828 272372
rect 41892 272308 41893 272372
rect 41827 272307 41893 272308
rect 41459 270468 41525 270469
rect 41459 270404 41460 270468
rect 41524 270404 41525 270468
rect 41459 270403 41525 270404
rect 673870 249797 673930 277611
rect 674787 264212 674853 264213
rect 674787 264148 674788 264212
rect 674852 264148 674853 264212
rect 674787 264147 674853 264148
rect 674790 249797 674850 264147
rect 676075 263668 676141 263669
rect 676075 263604 676076 263668
rect 676140 263604 676141 263668
rect 676075 263603 676141 263604
rect 676078 249797 676138 263603
rect 676995 261628 677061 261629
rect 676995 261564 676996 261628
rect 677060 261564 677061 261628
rect 676995 261563 677061 261564
rect 676811 260812 676877 260813
rect 676811 260748 676812 260812
rect 676876 260748 676877 260812
rect 676811 260747 676877 260748
rect 40723 249796 40789 249797
rect 40723 249732 40724 249796
rect 40788 249732 40789 249796
rect 40723 249731 40789 249732
rect 673867 249796 673933 249797
rect 673867 249732 673868 249796
rect 673932 249732 673933 249796
rect 673867 249731 673933 249732
rect 674787 249796 674853 249797
rect 674787 249732 674788 249796
rect 674852 249732 674853 249796
rect 674787 249731 674853 249732
rect 676075 249796 676141 249797
rect 676075 249732 676076 249796
rect 676140 249732 676141 249796
rect 676075 249731 676141 249732
rect 40539 249388 40605 249389
rect 40539 249324 40540 249388
rect 40604 249324 40605 249388
rect 40539 249323 40605 249324
rect 40542 234565 40602 249323
rect 40726 236605 40786 249731
rect 676814 246669 676874 260747
rect 676998 248301 677058 261563
rect 676995 248300 677061 248301
rect 676995 248236 676996 248300
rect 677060 248236 677061 248300
rect 676995 248235 677061 248236
rect 676811 246668 676877 246669
rect 676811 246604 676812 246668
rect 676876 246604 676877 246668
rect 676811 246603 676877 246604
rect 666875 246124 666941 246125
rect 666875 246060 666876 246124
rect 666940 246060 666941 246124
rect 666875 246059 666941 246060
rect 666507 245988 666573 245989
rect 666507 245924 666508 245988
rect 666572 245924 666573 245988
rect 666507 245923 666573 245924
rect 42379 237420 42445 237421
rect 42379 237356 42380 237420
rect 42444 237356 42445 237420
rect 42379 237355 42445 237356
rect 40723 236604 40789 236605
rect 40723 236540 40724 236604
rect 40788 236540 40789 236604
rect 40723 236539 40789 236540
rect 40539 234564 40605 234565
rect 40539 234500 40540 234564
rect 40604 234500 40605 234564
rect 40539 234499 40605 234500
rect 42382 227357 42442 237355
rect 147811 231028 147877 231029
rect 147811 230964 147812 231028
rect 147876 230964 147877 231028
rect 147811 230963 147877 230964
rect 147814 230485 147874 230963
rect 147811 230484 147877 230485
rect 147811 230420 147812 230484
rect 147876 230420 147877 230484
rect 147811 230419 147877 230420
rect 42379 227356 42445 227357
rect 42379 227292 42380 227356
rect 42444 227292 42445 227356
rect 42379 227291 42445 227292
rect 574507 219196 574573 219197
rect 499622 219061 499682 219182
rect 574139 219132 574140 219182
rect 574204 219132 574205 219182
rect 574139 219131 574205 219132
rect 574507 219132 574508 219196
rect 574572 219132 574573 219196
rect 574507 219131 574573 219132
rect 499619 219060 499685 219061
rect 499619 218996 499620 219060
rect 499684 218996 499685 219060
rect 499619 218995 499685 218996
rect 574510 218738 574570 219131
rect 490422 218109 490482 218502
rect 490419 218108 490485 218109
rect 490419 218044 490420 218108
rect 490484 218044 490485 218108
rect 490419 218043 490485 218044
rect 566043 217836 566109 217837
rect 566043 217772 566044 217836
rect 566108 217772 566109 217836
rect 566043 217771 566109 217772
rect 501275 217564 501341 217565
rect 501275 217500 501276 217564
rect 501340 217500 501341 217564
rect 501275 217499 501341 217500
rect 501278 217021 501338 217499
rect 501275 217020 501341 217021
rect 501275 216956 501276 217020
rect 501340 216956 501341 217020
rect 501275 216955 501341 216956
rect 566046 216069 566106 217771
rect 574326 216477 574386 217142
rect 575798 216749 575858 217822
rect 575795 216748 575861 216749
rect 575795 216684 575796 216748
rect 575860 216684 575861 216748
rect 575795 216683 575861 216684
rect 574323 216476 574389 216477
rect 574323 216412 574324 216476
rect 574388 216412 574389 216476
rect 574323 216411 574389 216412
rect 566043 216068 566109 216069
rect 566043 216004 566044 216068
rect 566108 216004 566109 216068
rect 566043 216003 566109 216004
rect 41827 210084 41893 210085
rect 41827 210020 41828 210084
rect 41892 210020 41893 210084
rect 41827 210019 41893 210020
rect 40907 208180 40973 208181
rect 40907 208116 40908 208180
rect 40972 208116 40973 208180
rect 40907 208115 40973 208116
rect 40539 207772 40605 207773
rect 40539 207708 40540 207772
rect 40604 207708 40605 207772
rect 40539 207707 40605 207708
rect 40542 183429 40602 207707
rect 40723 206140 40789 206141
rect 40723 206076 40724 206140
rect 40788 206076 40789 206140
rect 40723 206075 40789 206076
rect 40726 191589 40786 206075
rect 40910 197165 40970 208115
rect 41459 205732 41525 205733
rect 41459 205668 41460 205732
rect 41524 205668 41525 205732
rect 41459 205667 41525 205668
rect 40907 197164 40973 197165
rect 40907 197100 40908 197164
rect 40972 197100 40973 197164
rect 40907 197099 40973 197100
rect 40723 191588 40789 191589
rect 40723 191524 40724 191588
rect 40788 191524 40789 191588
rect 40723 191523 40789 191524
rect 41462 184109 41522 205667
rect 41643 200700 41709 200701
rect 41643 200636 41644 200700
rect 41708 200636 41709 200700
rect 41643 200635 41709 200636
rect 41646 186330 41706 200635
rect 41830 195261 41890 210019
rect 666510 205650 666570 245923
rect 666691 245716 666757 245717
rect 666691 245652 666692 245716
rect 666756 245652 666757 245716
rect 666691 245651 666757 245652
rect 666694 210493 666754 245651
rect 666691 210492 666757 210493
rect 666691 210428 666692 210492
rect 666756 210428 666757 210492
rect 666691 210427 666757 210428
rect 666510 205590 666754 205650
rect 41827 195260 41893 195261
rect 41827 195196 41828 195260
rect 41892 195196 41893 195260
rect 41827 195195 41893 195196
rect 666694 189345 666754 205590
rect 666878 199137 666938 246059
rect 668163 245988 668229 245989
rect 668163 245924 668164 245988
rect 668228 245924 668229 245988
rect 668163 245923 668229 245924
rect 667979 211172 668045 211173
rect 667979 211108 667980 211172
rect 668044 211108 668045 211172
rect 667979 211107 668045 211108
rect 667059 210492 667125 210493
rect 667059 210428 667060 210492
rect 667124 210428 667125 210492
rect 667059 210427 667125 210428
rect 666875 199136 666941 199137
rect 666875 199072 666876 199136
rect 666940 199072 666941 199136
rect 666875 199071 666941 199072
rect 667062 194850 667122 210427
rect 667982 207365 668042 211107
rect 667979 207364 668045 207365
rect 667979 207300 667980 207364
rect 668044 207300 668045 207364
rect 667979 207299 668045 207300
rect 668166 202469 668226 245923
rect 668347 245716 668413 245717
rect 668347 245652 668348 245716
rect 668412 245652 668413 245716
rect 668347 245651 668413 245652
rect 668163 202468 668229 202469
rect 668163 202404 668164 202468
rect 668228 202404 668229 202468
rect 668163 202403 668229 202404
rect 668350 197573 668410 245651
rect 675339 243268 675405 243269
rect 675339 243204 675340 243268
rect 675404 243204 675405 243268
rect 675339 243203 675405 243204
rect 675342 238645 675402 243203
rect 675339 238644 675405 238645
rect 675339 238580 675340 238644
rect 675404 238580 675405 238644
rect 675339 238579 675405 238580
rect 675523 218652 675589 218653
rect 675523 218588 675524 218652
rect 675588 218588 675589 218652
rect 675523 218587 675589 218588
rect 669451 217972 669517 217973
rect 669451 217908 669452 217972
rect 669516 217908 669517 217972
rect 669451 217907 669517 217908
rect 669454 206410 669514 217907
rect 670923 216612 670989 216613
rect 670923 216548 670924 216612
rect 670988 216548 670989 216612
rect 670923 216547 670989 216548
rect 675339 216612 675405 216613
rect 675339 216548 675340 216612
rect 675404 216548 675405 216612
rect 675339 216547 675405 216548
rect 669635 211172 669701 211173
rect 669635 211108 669636 211172
rect 669700 211108 669701 211172
rect 669635 211107 669701 211108
rect 670739 211172 670805 211173
rect 670739 211108 670740 211172
rect 670804 211108 670805 211172
rect 670739 211107 670805 211108
rect 669270 206350 669514 206410
rect 669270 205461 669330 206350
rect 669638 205730 669698 211107
rect 669454 205670 669698 205730
rect 669267 205460 669333 205461
rect 669267 205396 669268 205460
rect 669332 205396 669333 205460
rect 669267 205395 669333 205396
rect 669454 204101 669514 205670
rect 669635 205460 669701 205461
rect 669635 205396 669636 205460
rect 669700 205396 669701 205460
rect 669635 205395 669701 205396
rect 669451 204100 669517 204101
rect 669451 204036 669452 204100
rect 669516 204036 669517 204100
rect 669451 204035 669517 204036
rect 668347 197572 668413 197573
rect 668347 197508 668348 197572
rect 668412 197508 668413 197572
rect 668347 197507 668413 197508
rect 669638 195990 669698 205395
rect 666878 194790 667122 194850
rect 669454 195930 669698 195990
rect 666878 194241 666938 194790
rect 666875 194240 666941 194241
rect 666875 194176 666876 194240
rect 666940 194176 666941 194240
rect 666875 194175 666941 194176
rect 666691 189344 666757 189345
rect 666691 189280 666692 189344
rect 666756 189280 666757 189344
rect 666691 189279 666757 189280
rect 41646 186270 41890 186330
rect 41830 185877 41890 186270
rect 41827 185876 41893 185877
rect 41827 185812 41828 185876
rect 41892 185812 41893 185876
rect 41827 185811 41893 185812
rect 41459 184108 41525 184109
rect 41459 184044 41460 184108
rect 41524 184044 41525 184108
rect 41459 184043 41525 184044
rect 40539 183428 40605 183429
rect 40539 183364 40540 183428
rect 40604 183364 40605 183428
rect 40539 183363 40605 183364
rect 669454 179621 669514 195930
rect 669451 179620 669517 179621
rect 669451 179556 669452 179620
rect 669516 179556 669517 179620
rect 669451 179555 669517 179556
rect 670742 155141 670802 211107
rect 670926 165749 670986 216547
rect 671107 216204 671173 216205
rect 671107 216140 671108 216204
rect 671172 216140 671173 216204
rect 671107 216139 671173 216140
rect 671110 210901 671170 216139
rect 673683 214028 673749 214029
rect 673683 213964 673684 214028
rect 673748 213964 673749 214028
rect 673683 213963 673749 213964
rect 672947 212668 673013 212669
rect 672947 212604 672948 212668
rect 673012 212604 673013 212668
rect 672947 212603 673013 212604
rect 671107 210900 671173 210901
rect 671107 210836 671108 210900
rect 671172 210836 671173 210900
rect 671107 210835 671173 210836
rect 672950 186330 673010 212603
rect 673131 210492 673197 210493
rect 673131 210428 673132 210492
rect 673196 210428 673197 210492
rect 673131 210427 673197 210428
rect 673499 210492 673565 210493
rect 673499 210428 673500 210492
rect 673564 210428 673565 210492
rect 673499 210427 673565 210428
rect 672766 186270 673010 186330
rect 672766 183565 672826 186270
rect 673134 183565 673194 210427
rect 673315 209268 673381 209269
rect 673315 209204 673316 209268
rect 673380 209204 673381 209268
rect 673315 209203 673381 209204
rect 672763 183564 672829 183565
rect 672763 183500 672764 183564
rect 672828 183500 672829 183564
rect 672763 183499 672829 183500
rect 673131 183564 673197 183565
rect 673131 183500 673132 183564
rect 673196 183500 673197 183564
rect 673131 183499 673197 183500
rect 673318 173093 673378 209203
rect 673315 173092 673381 173093
rect 673315 173028 673316 173092
rect 673380 173028 673381 173092
rect 673315 173027 673381 173028
rect 672947 168332 673013 168333
rect 672947 168268 672948 168332
rect 673012 168268 673013 168332
rect 672947 168267 673013 168268
rect 670923 165748 670989 165749
rect 670923 165684 670924 165748
rect 670988 165684 670989 165748
rect 670923 165683 670989 165684
rect 670739 155140 670805 155141
rect 670739 155076 670740 155140
rect 670804 155076 670805 155140
rect 670739 155075 670805 155076
rect 672950 133789 673010 168267
rect 673502 148477 673562 210427
rect 673686 153373 673746 213963
rect 675342 212397 675402 216547
rect 675339 212396 675405 212397
rect 675339 212332 675340 212396
rect 675404 212332 675405 212396
rect 675339 212331 675405 212332
rect 675526 210493 675586 218587
rect 675707 217428 675773 217429
rect 675707 217364 675708 217428
rect 675772 217364 675773 217428
rect 675707 217363 675773 217364
rect 675523 210492 675589 210493
rect 675523 210428 675524 210492
rect 675588 210428 675589 210492
rect 675523 210427 675589 210428
rect 675710 198389 675770 217363
rect 675891 214572 675957 214573
rect 675891 214508 675892 214572
rect 675956 214508 675957 214572
rect 675891 214507 675957 214508
rect 675894 213210 675954 214507
rect 675894 213150 676690 213210
rect 675891 212396 675957 212397
rect 675891 212332 675892 212396
rect 675956 212332 675957 212396
rect 675891 212331 675957 212332
rect 675894 211850 675954 212331
rect 675894 211790 676322 211850
rect 675891 211172 675957 211173
rect 675891 211108 675892 211172
rect 675956 211108 675957 211172
rect 675891 211107 675957 211108
rect 675707 198388 675773 198389
rect 675707 198324 675708 198388
rect 675772 198324 675773 198388
rect 675707 198323 675773 198324
rect 675894 192813 675954 211107
rect 676075 210492 676141 210493
rect 676075 210428 676076 210492
rect 676140 210428 676141 210492
rect 676075 210427 676141 210428
rect 676078 193221 676138 210427
rect 676262 205053 676322 211790
rect 676443 211444 676509 211445
rect 676443 211380 676444 211444
rect 676508 211380 676509 211444
rect 676443 211379 676509 211380
rect 676259 205052 676325 205053
rect 676259 204988 676260 205052
rect 676324 204988 676325 205052
rect 676259 204987 676325 204988
rect 676446 197029 676506 211379
rect 676630 200021 676690 213150
rect 676811 201380 676877 201381
rect 676811 201316 676812 201380
rect 676876 201316 676877 201380
rect 676811 201315 676877 201316
rect 676627 200020 676693 200021
rect 676627 199956 676628 200020
rect 676692 199956 676693 200020
rect 676627 199955 676693 199956
rect 676443 197028 676509 197029
rect 676443 196964 676444 197028
rect 676508 196964 676509 197028
rect 676443 196963 676509 196964
rect 676075 193220 676141 193221
rect 676075 193156 676076 193220
rect 676140 193156 676141 193220
rect 676075 193155 676141 193156
rect 675891 192812 675957 192813
rect 675891 192748 675892 192812
rect 675956 192748 675957 192812
rect 675891 192747 675957 192748
rect 676814 183570 676874 201315
rect 676262 183510 676874 183570
rect 675891 174724 675957 174725
rect 675891 174660 675892 174724
rect 675956 174660 675957 174724
rect 675891 174659 675957 174660
rect 675894 174450 675954 174659
rect 676262 174450 676322 183510
rect 675894 174390 676322 174450
rect 675707 173636 675773 173637
rect 675707 173572 675708 173636
rect 675772 173572 675773 173636
rect 675707 173571 675773 173572
rect 675339 172412 675405 172413
rect 675339 172348 675340 172412
rect 675404 172348 675405 172412
rect 675339 172347 675405 172348
rect 675342 162213 675402 172347
rect 675710 169010 675770 173571
rect 675891 170780 675957 170781
rect 675891 170716 675892 170780
rect 675956 170716 675957 170780
rect 675891 170715 675957 170716
rect 675894 170370 675954 170715
rect 675894 170310 676506 170370
rect 675894 169630 676322 169690
rect 675894 169421 675954 169630
rect 675891 169420 675957 169421
rect 675891 169356 675892 169420
rect 675956 169356 675957 169420
rect 675891 169355 675957 169356
rect 675710 168950 676138 169010
rect 675707 167652 675773 167653
rect 675707 167588 675708 167652
rect 675772 167588 675773 167652
rect 675707 167587 675773 167588
rect 675339 162212 675405 162213
rect 675339 162148 675340 162212
rect 675404 162148 675405 162212
rect 675339 162147 675405 162148
rect 675523 161396 675589 161397
rect 675523 161332 675524 161396
rect 675588 161332 675589 161396
rect 675523 161331 675589 161332
rect 675526 160173 675586 161331
rect 675523 160172 675589 160173
rect 675523 160108 675524 160172
rect 675588 160108 675589 160172
rect 675523 160107 675589 160108
rect 673683 153372 673749 153373
rect 673683 153308 673684 153372
rect 673748 153308 673749 153372
rect 673683 153307 673749 153308
rect 673499 148476 673565 148477
rect 673499 148412 673500 148476
rect 673564 148412 673565 148476
rect 673499 148411 673565 148412
rect 675710 147661 675770 167587
rect 675891 162212 675957 162213
rect 675891 162148 675892 162212
rect 675956 162148 675957 162212
rect 675891 162147 675957 162148
rect 675894 153101 675954 162147
rect 675891 153100 675957 153101
rect 675891 153036 675892 153100
rect 675956 153036 675957 153100
rect 675891 153035 675957 153036
rect 676078 148477 676138 168950
rect 676262 155685 676322 169630
rect 676446 156501 676506 170310
rect 676627 166428 676693 166429
rect 676627 166364 676628 166428
rect 676692 166364 676693 166428
rect 676627 166363 676693 166364
rect 676443 156500 676509 156501
rect 676443 156436 676444 156500
rect 676508 156436 676509 156500
rect 676443 156435 676509 156436
rect 676259 155684 676325 155685
rect 676259 155620 676260 155684
rect 676324 155620 676325 155684
rect 676259 155619 676325 155620
rect 676630 151469 676690 166363
rect 676627 151468 676693 151469
rect 676627 151404 676628 151468
rect 676692 151404 676693 151468
rect 676627 151403 676693 151404
rect 676075 148476 676141 148477
rect 676075 148412 676076 148476
rect 676140 148412 676141 148476
rect 676075 148411 676141 148412
rect 675707 147660 675773 147661
rect 675707 147596 675708 147660
rect 675772 147596 675773 147660
rect 675707 147595 675773 147596
rect 672947 133788 673013 133789
rect 672947 133724 672948 133788
rect 673012 133724 673013 133788
rect 672947 133723 673013 133724
rect 676259 128620 676325 128621
rect 676259 128556 676260 128620
rect 676324 128556 676325 128620
rect 676259 128555 676325 128556
rect 676075 128212 676141 128213
rect 676075 128148 676076 128212
rect 676140 128148 676141 128212
rect 676075 128147 676141 128148
rect 675891 127260 675957 127261
rect 675891 127196 675892 127260
rect 675956 127196 675957 127260
rect 675891 127195 675957 127196
rect 675707 117060 675773 117061
rect 675707 116996 675708 117060
rect 675772 116996 675773 117060
rect 675707 116995 675773 116996
rect 675710 102645 675770 116995
rect 675894 108085 675954 127195
rect 675891 108084 675957 108085
rect 675891 108020 675892 108084
rect 675956 108020 675957 108084
rect 675891 108019 675957 108020
rect 676078 103189 676138 128147
rect 676262 113117 676322 128555
rect 676811 124540 676877 124541
rect 676811 124476 676812 124540
rect 676876 124476 676877 124540
rect 676811 124475 676877 124476
rect 676259 113116 676325 113117
rect 676259 113052 676260 113116
rect 676324 113052 676325 113116
rect 676259 113051 676325 113052
rect 676075 103188 676141 103189
rect 676075 103124 676076 103188
rect 676140 103124 676141 103188
rect 676075 103123 676141 103124
rect 675707 102644 675773 102645
rect 675707 102580 675708 102644
rect 675772 102580 675773 102644
rect 675707 102579 675773 102580
rect 676814 101421 676874 124475
rect 676995 117332 677061 117333
rect 676995 117268 676996 117332
rect 677060 117268 677061 117332
rect 676995 117267 677061 117268
rect 676998 110397 677058 117267
rect 676995 110396 677061 110397
rect 676995 110332 676996 110396
rect 677060 110332 677061 110396
rect 676995 110331 677061 110332
rect 676811 101420 676877 101421
rect 676811 101356 676812 101420
rect 676876 101356 676877 101420
rect 676811 101355 676877 101356
rect 637251 96932 637317 96933
rect 637251 96868 637252 96932
rect 637316 96868 637317 96932
rect 637251 96867 637317 96868
rect 634675 95708 634741 95709
rect 634675 95644 634676 95708
rect 634740 95644 634741 95708
rect 634675 95643 634741 95644
rect 634678 77757 634738 95643
rect 637254 84210 637314 96867
rect 637070 84150 637314 84210
rect 637070 78573 637130 84150
rect 637067 78572 637133 78573
rect 637067 78508 637068 78572
rect 637132 78508 637133 78572
rect 637067 78507 637133 78508
rect 634675 77756 634741 77757
rect 634675 77692 634676 77756
rect 634740 77692 634741 77756
rect 634675 77691 634741 77692
rect 409643 53140 409709 53141
rect 409643 53076 409644 53140
rect 409708 53076 409709 53140
rect 409643 53075 409709 53076
rect 147627 50284 147693 50285
rect 147627 50220 147628 50284
rect 147692 50220 147693 50284
rect 147627 50219 147693 50220
rect 131067 49740 131133 49741
rect 131067 49676 131068 49740
rect 131132 49676 131133 49740
rect 131067 49675 131133 49676
rect 131070 47021 131130 49675
rect 147630 47565 147690 50219
rect 365483 48924 365549 48925
rect 365483 48860 365484 48924
rect 365548 48860 365549 48924
rect 365483 48859 365549 48860
rect 361987 47836 362053 47837
rect 361987 47772 361988 47836
rect 362052 47772 362053 47836
rect 361987 47771 362053 47772
rect 147627 47564 147693 47565
rect 147627 47500 147628 47564
rect 147692 47500 147693 47564
rect 147627 47499 147693 47500
rect 187555 47564 187621 47565
rect 187555 47500 187556 47564
rect 187620 47500 187621 47564
rect 187555 47499 187621 47500
rect 131067 47020 131133 47021
rect 131067 46956 131068 47020
rect 131132 46956 131133 47020
rect 131067 46955 131133 46956
rect 187558 42125 187618 47499
rect 306971 46476 307037 46477
rect 306971 46412 306972 46476
rect 307036 46412 307037 46476
rect 306971 46411 307037 46412
rect 306974 42397 307034 46411
rect 310099 46204 310165 46205
rect 310099 46140 310100 46204
rect 310164 46140 310165 46204
rect 310099 46139 310165 46140
rect 310102 42397 310162 46139
rect 306971 42396 307037 42397
rect 306971 42332 306972 42396
rect 307036 42332 307037 42396
rect 306971 42331 307037 42332
rect 310099 42396 310165 42397
rect 310099 42332 310100 42396
rect 310164 42332 310165 42396
rect 310099 42331 310165 42332
rect 361990 42125 362050 47771
rect 365486 42125 365546 48859
rect 409646 42805 409706 53075
rect 464843 51780 464909 51781
rect 464843 51716 464844 51780
rect 464908 51716 464909 51780
rect 464843 51715 464909 51716
rect 460795 50284 460861 50285
rect 460795 50220 460796 50284
rect 460860 50220 460861 50284
rect 460795 50219 460861 50220
rect 411115 49196 411181 49197
rect 411115 49132 411116 49196
rect 411180 49132 411181 49196
rect 411115 49131 411181 49132
rect 411118 42805 411178 49131
rect 416635 48108 416701 48109
rect 416635 48044 416636 48108
rect 416700 48044 416701 48108
rect 416635 48043 416701 48044
rect 416638 42805 416698 48043
rect 409643 42804 409709 42805
rect 409643 42740 409644 42804
rect 409708 42740 409709 42804
rect 409643 42739 409709 42740
rect 411115 42804 411181 42805
rect 411115 42740 411116 42804
rect 411180 42740 411181 42804
rect 411115 42739 411181 42740
rect 416635 42804 416701 42805
rect 416635 42740 416636 42804
rect 416700 42740 416701 42804
rect 416635 42739 416701 42740
rect 460798 42125 460858 50219
rect 464846 42805 464906 51715
rect 525747 50556 525813 50557
rect 525747 50492 525748 50556
rect 525812 50492 525813 50556
rect 525747 50491 525813 50492
rect 529795 50556 529861 50557
rect 529795 50492 529796 50556
rect 529860 50492 529861 50556
rect 529795 50491 529861 50492
rect 514707 47292 514773 47293
rect 514707 47228 514708 47292
rect 514772 47228 514773 47292
rect 514707 47227 514773 47228
rect 471651 44844 471717 44845
rect 471651 44780 471652 44844
rect 471716 44780 471717 44844
rect 471651 44779 471717 44780
rect 464843 42804 464909 42805
rect 464843 42740 464844 42804
rect 464908 42740 464909 42804
rect 464843 42739 464909 42740
rect 471654 42125 471714 44779
rect 514710 42125 514770 47227
rect 518571 47020 518637 47021
rect 518571 46956 518572 47020
rect 518636 46956 518637 47020
rect 518571 46955 518637 46956
rect 518574 42397 518634 46955
rect 521699 45932 521765 45933
rect 521699 45868 521700 45932
rect 521764 45868 521765 45932
rect 521699 45867 521765 45868
rect 520411 45116 520477 45117
rect 520411 45052 520412 45116
rect 520476 45052 520477 45116
rect 520411 45051 520477 45052
rect 518571 42396 518637 42397
rect 518571 42332 518572 42396
rect 518636 42332 518637 42396
rect 518571 42331 518637 42332
rect 520414 42125 520474 45051
rect 187555 42124 187621 42125
rect 187555 42060 187556 42124
rect 187620 42060 187621 42124
rect 187555 42059 187621 42060
rect 361987 42124 362053 42125
rect 361987 42060 361988 42124
rect 362052 42060 362053 42124
rect 361987 42059 362053 42060
rect 365483 42124 365549 42125
rect 365483 42060 365484 42124
rect 365548 42060 365549 42124
rect 365483 42059 365549 42060
rect 460795 42124 460861 42125
rect 460795 42060 460796 42124
rect 460860 42060 460861 42124
rect 460795 42059 460861 42060
rect 471651 42124 471717 42125
rect 471651 42060 471652 42124
rect 471716 42060 471717 42124
rect 471651 42059 471717 42060
rect 514707 42124 514773 42125
rect 514707 42060 514708 42124
rect 514772 42060 514773 42124
rect 514707 42059 514773 42060
rect 520411 42124 520477 42125
rect 520411 42060 520412 42124
rect 520476 42060 520477 42124
rect 520411 42059 520477 42060
rect 521702 41989 521762 45867
rect 525750 42125 525810 50491
rect 529798 42125 529858 50491
rect 525747 42124 525813 42125
rect 525747 42060 525748 42124
rect 525812 42060 525813 42124
rect 525747 42059 525813 42060
rect 529795 42124 529861 42125
rect 529795 42060 529796 42124
rect 529860 42060 529861 42124
rect 529795 42059 529861 42060
rect 521699 41988 521765 41989
rect 521699 41924 521700 41988
rect 521764 41924 521765 41988
rect 521699 41923 521765 41924
<< via4 >>
rect 189494 997102 189730 997338
rect 195014 997102 195250 997338
rect 485550 997102 485786 997338
rect 506342 997102 506578 997338
rect 536518 997102 536754 997338
rect 556022 997102 556258 997338
rect 186182 993022 186418 993258
rect 194462 993022 194698 993258
rect 286646 993022 286882 993258
rect 298422 993022 298658 993258
rect 499534 219182 499770 219418
rect 574054 219196 574290 219418
rect 574054 219182 574140 219196
rect 574140 219182 574204 219196
rect 574204 219182 574290 219196
rect 490334 218502 490570 218738
rect 574422 218502 574658 218738
rect 493646 217972 493882 218058
rect 493646 217908 493732 217972
rect 493732 217908 493796 217972
rect 493796 217908 493882 217972
rect 493646 217822 493882 217908
rect 575710 217822 575946 218058
rect 491070 217292 491306 217378
rect 491070 217228 491156 217292
rect 491156 217228 491220 217292
rect 491220 217228 491306 217292
rect 491070 217142 491306 217228
rect 574238 217142 574474 217378
<< metal5 >>
rect 189452 997338 195292 997380
rect 189452 997102 189494 997338
rect 189730 997102 195014 997338
rect 195250 997102 195292 997338
rect 189452 997060 195292 997102
rect 485508 997338 506620 997380
rect 485508 997102 485550 997338
rect 485786 997102 506342 997338
rect 506578 997102 506620 997338
rect 485508 997060 506620 997102
rect 536476 997338 556300 997380
rect 536476 997102 536518 997338
rect 536754 997102 556022 997338
rect 556258 997102 556300 997338
rect 536476 997060 556300 997102
rect 186140 993258 194740 993300
rect 186140 993022 186182 993258
rect 186418 993022 194462 993258
rect 194698 993022 194740 993258
rect 186140 992980 194740 993022
rect 286604 993258 298700 993300
rect 286604 993022 286646 993258
rect 286882 993022 298422 993258
rect 298658 993022 298700 993258
rect 286604 992980 298700 993022
rect 499492 219418 574332 219460
rect 499492 219182 499534 219418
rect 499770 219182 574054 219418
rect 574290 219182 574332 219418
rect 499492 219140 574332 219182
rect 490292 218738 574700 218780
rect 490292 218502 490334 218738
rect 490570 218502 574422 218738
rect 574658 218502 574700 218738
rect 490292 218460 574700 218502
rect 493604 218058 575988 218100
rect 493604 217822 493646 218058
rect 493882 217822 575710 218058
rect 575946 217822 575988 218058
rect 493604 217780 575988 217822
rect 491028 217378 574516 217420
rect 491028 217142 491070 217378
rect 491306 217142 574238 217378
rect 574474 217142 574516 217378
rect 491028 217100 574516 217142
use user_id_programming  user_id_value
timestamp 1665478365
transform 1 0 656624 0 1 88126
box 0 0 7109 7077
use mgmt_core_wrapper  soc
timestamp 1665478365
transform 1 0 52034 0 1 53002
box -156 0 524096 164000
use xres_buf  rstb_level
timestamp 1665478365
transform -1 0 145710 0 -1 50488
box 414 -400 3522 3800
use simple_por  por
timestamp 1665478365
transform 1 0 650146 0 -1 55282
box -14 11 11344 8684
use digital_pll  pll
timestamp 1665478365
transform 1 0 628146 0 1 80944
box 0 0 15000 15000
use housekeeping  housekeeping
timestamp 1665478365
transform 1 0 592434 0 1 100002
box 0 0 74046 110190
use gpio_defaults_block  gpio_defaults_block_0
timestamp 1665478365
transform -1 0 709467 0 1 134000
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_1\[0\]
timestamp 1665478365
transform -1 0 710203 0 1 121000
box 872 416 34000 13000
use caravel_clocking  clock_ctrl
timestamp 1665478365
transform 1 0 626764 0 1 63284
box -38 -48 20000 12000
use gpio_control_block  gpio_control_bidir_1\[1\]
timestamp 1665478365
transform -1 0 710203 0 1 166200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_1
timestamp 1665478365
transform -1 0 709467 0 1 179200
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_2\[2\]
timestamp 1665478365
transform 1 0 7631 0 1 202600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[0\]
timestamp 1665478365
transform -1 0 710203 0 1 211200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_2
timestamp 1665478365
transform -1 0 709467 0 1 224200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_37
timestamp 1665478365
transform 1 0 8367 0 1 215600
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_2\[1\]
timestamp 1665478365
transform 1 0 7631 0 1 245800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[1\]
timestamp 1665478365
transform -1 0 710203 0 1 256400
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_36
timestamp 1665478365
transform 1 0 8367 0 1 258800
box -38 0 6018 2224
use mgmt_protect  mgmt_buffers
timestamp 1665478365
transform 1 0 128180 0 1 232036
box 1066 -400 380400 32400
use spare_logic_block  spare_logic\[0\]
timestamp 1665478365
transform 1 0 88632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[1\]
timestamp 1665478365
transform 1 0 89351 0 1 248673
box 0 0 9000 9000
use spare_logic_block  spare_logic\[2\]
timestamp 1665478365
transform 1 0 575145 0 1 246987
box 0 0 9000 9000
use spare_logic_block  spare_logic\[3\]
timestamp 1665478365
transform 1 0 613558 0 1 245856
box 0 0 9000 9000
use gpio_control_block  gpio_control_bidir_2\[0\]
timestamp 1665478365
transform 1 0 7631 0 1 289000
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_3
timestamp 1665478365
transform -1 0 709467 0 1 269400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[2\]
timestamp 1665478365
transform -1 0 710203 0 1 301400
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_35
timestamp 1665478365
transform 1 0 8367 0 1 302000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_4
timestamp 1665478365
transform -1 0 709467 0 1 314400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[13\]
timestamp 1665478365
transform 1 0 7631 0 1 418600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[14\]
timestamp 1665478365
transform 1 0 7631 0 1 375400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[15\]
timestamp 1665478365
transform 1 0 7631 0 1 332200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_32
timestamp 1665478365
transform 1 0 8367 0 1 431600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_33
timestamp 1665478365
transform 1 0 8367 0 1 388400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_34
timestamp 1665478365
transform 1 0 8367 0 1 345200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[3\]
timestamp 1665478365
transform -1 0 710203 0 1 346400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[4\]
timestamp 1665478365
transform -1 0 710203 0 1 391600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[5\]
timestamp 1665478365
transform -1 0 710203 0 1 479800
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_5
timestamp 1665478365
transform -1 0 709467 0 1 359400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_6
timestamp 1665478365
transform -1 0 709467 0 1 404600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_7
timestamp 1665478365
transform -1 0 709467 0 1 492800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_31
timestamp 1665478365
transform 1 0 8367 0 1 559200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_30
timestamp 1665478365
transform 1 0 8367 0 1 602400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[12\]
timestamp 1665478365
transform 1 0 7631 0 1 546200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[11\]
timestamp 1665478365
transform 1 0 7631 0 1 589400
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_9
timestamp 1665478365
transform -1 0 709467 0 1 581800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_8
timestamp 1665478365
transform -1 0 709467 0 1 536800
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[1\]
timestamp 1665478365
transform -1 0 710203 0 1 568800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[0\]
timestamp 1665478365
transform -1 0 710203 0 1 523800
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_29
timestamp 1665478365
transform 1 0 8367 0 1 645600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_28
timestamp 1665478365
transform 1 0 8367 0 1 688800
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[9\]
timestamp 1665478365
transform 1 0 7631 0 1 675800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[10\]
timestamp 1665478365
transform 1 0 7631 0 1 632600
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_11
timestamp 1665478365
transform -1 0 709467 0 1 672000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_10
timestamp 1665478365
transform -1 0 709467 0 1 627000
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[3\]
timestamp 1665478365
transform -1 0 710203 0 1 659000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[2\]
timestamp 1665478365
transform -1 0 710203 0 1 614000
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_27
timestamp 1665478365
transform 1 0 8367 0 1 732000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_26
timestamp 1665478365
transform 1 0 8367 0 1 775200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[8\]
timestamp 1665478365
transform 1 0 7631 0 1 719000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[7\]
timestamp 1665478365
transform 1 0 7631 0 1 762200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_13
timestamp 1665478365
transform -1 0 709467 0 1 762200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_12
timestamp 1665478365
transform -1 0 709467 0 1 717200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[5\]
timestamp 1665478365
transform -1 0 710203 0 1 749200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[4\]
timestamp 1665478365
transform -1 0 710203 0 1 704200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_25
timestamp 1665478365
transform 1 0 8367 0 1 818400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[6\]
timestamp 1665478365
transform 1 0 7631 0 1 805400
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_24
timestamp 1665478365
transform 1 0 8367 0 1 944200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[5\]
timestamp 1665478365
transform 1 0 7631 0 1 931200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_14
timestamp 1665478365
transform -1 0 709467 0 1 940600
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[6\]
timestamp 1665478365
transform -1 0 710203 0 1 927600
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_23
timestamp 1665478365
transform 0 1 110194 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_22
timestamp 1665478365
transform 0 1 161594 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[4\]
timestamp 1665478365
transform 0 1 97200 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[3\]
timestamp 1665478365
transform 0 1 148600 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_21
timestamp 1665478365
transform 0 1 212994 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[2\]
timestamp 1665478365
transform 0 1 200000 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[1\]
timestamp 1665478365
transform 0 1 251400 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_20
timestamp 1665478365
transform 0 1 264394 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_19
timestamp 1665478365
transform 0 1 315994 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[0\]
timestamp 1665478365
transform 0 1 303000 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_18
timestamp 1665478365
transform 0 1 366394 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_17
timestamp 1665478365
transform 0 1 433794 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[9\]
timestamp 1665478365
transform 0 1 420800 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[10\]
timestamp 1665478365
transform 0 1 353400 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_16
timestamp 1665478365
transform 0 1 510794 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[8\]
timestamp 1665478365
transform 0 1 497800 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_15
timestamp 1665478365
transform 0 1 562194 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[7\]
timestamp 1665478365
transform 0 1 549200 -1 0 1030077
box 872 416 34000 13000
use caravel_power_routing  caravel_power_routing
timestamp 1665478365
transform 1 0 6022 0 1 33900
box 0 0 705792 997796
use user_project_wrapper  mprj
timestamp 1665478365
transform 1 0 65308 0 1 278718
box -8726 -7654 592650 711590
use chip_io  padframe
timestamp 1665478365
transform 1 0 0 0 1 0
box 0 0 717600 1037600
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
