* NGSPICE file created from housekeeping.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_1 abstract view
.subckt sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4bb_1 abstract view
.subckt sky130_fd_sc_hd__nand4bb_1 A_N B_N C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4bb_4 abstract view
.subckt sky130_fd_sc_hd__nand4bb_4 A_N B_N C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtn_1 abstract view
.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4bb_2 abstract view
.subckt sky130_fd_sc_hd__nand4bb_2 A_N B_N C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_1 abstract view
.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_1 abstract view
.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_2 abstract view
.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_2 abstract view
.subckt sky130_fd_sc_hd__a41oi_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_2 abstract view
.subckt sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_1 abstract view
.subckt sky130_fd_sc_hd__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

.subckt housekeeping VGND VPWR debug_in debug_mode debug_oeb debug_out irq[0] irq[1]
+ irq[2] mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13]
+ mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18]
+ mask_rev_in[19] mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23]
+ mask_rev_in[24] mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4]
+ mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14]
+ mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19]
+ mgmt_gpio_in[1] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23]
+ mgmt_gpio_in[24] mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28]
+ mgmt_gpio_in[29] mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32]
+ mgmt_gpio_in[33] mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37]
+ mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7]
+ mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16]
+ mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20]
+ mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2]
+ mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[35] mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4]
+ mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18]
+ mgmt_gpio_out[19] mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22]
+ mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27]
+ mgmt_gpio_out[28] mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31]
+ mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36]
+ mgmt_gpio_out[37] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oeb
+ pad_flash_csb pad_flash_csb_oeb pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ieb
+ pad_flash_io0_oeb pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ieb pad_flash_io1_oeb
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1]
+ pll_div[2] pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0]
+ pll_trim[10] pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16]
+ pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22]
+ pll_trim[23] pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5]
+ pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out[0] pwr_ctrl_out[1]
+ pwr_ctrl_out[2] pwr_ctrl_out[3] qspi_enabled reset ser_rx ser_tx serial_clock serial_data_1
+ serial_data_2 serial_load serial_resetn spi_csb spi_enabled spi_sck spi_sdi spi_sdo
+ spi_sdoenb spimemio_flash_clk spimemio_flash_csb spimemio_flash_io0_di spimemio_flash_io0_do
+ spimemio_flash_io0_oeb spimemio_flash_io1_di spimemio_flash_io1_do spimemio_flash_io1_oeb
+ spimemio_flash_io2_di spimemio_flash_io2_do spimemio_flash_io2_oeb spimemio_flash_io3_di
+ spimemio_flash_io3_do spimemio_flash_io3_oeb trap uart_enabled user_clock usr1_vcc_pwrgood
+ usr1_vdd_pwrgood usr2_vcc_pwrgood usr2_vdd_pwrgood wb_ack_o wb_adr_i[0] wb_adr_i[10]
+ wb_adr_i[11] wb_adr_i[12] wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17]
+ wb_adr_i[18] wb_adr_i[19] wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23]
+ wb_adr_i[24] wb_adr_i[25] wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2]
+ wb_adr_i[30] wb_adr_i[31] wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7]
+ wb_adr_i[8] wb_adr_i[9] wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11]
+ wb_dat_i[12] wb_dat_i[13] wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18]
+ wb_dat_i[19] wb_dat_i[1] wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24]
+ wb_dat_i[25] wb_dat_i[26] wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30]
+ wb_dat_i[31] wb_dat_i[3] wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8]
+ wb_dat_i[9] wb_dat_o[0] wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14]
+ wb_dat_o[15] wb_dat_o[16] wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20]
+ wb_dat_o[21] wb_dat_o[22] wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27]
+ wb_dat_o[28] wb_dat_o[29] wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4]
+ wb_dat_o[5] wb_dat_o[6] wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0]
+ wb_sel_i[1] wb_sel_i[2] wb_sel_i[3] wb_stb_i wb_we_i
XFILLER_140_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6914_ _7258_/CLK _6957_/Q _6869_/X VGND VGND VPWR VPWR _6914_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6845_ _6969_/Q _6845_/A2 _6845_/B1 _6970_/Q VGND VGND VPWR VPWR _6845_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6776_ _7232_/Q _6720_/C _6562_/C _6457_/X _7197_/Q VGND VGND VPWR VPWR _6776_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_168_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3988_ _7174_/Q _6038_/B hold98/A input4/X _3544_/X VGND VGND VPWR VPWR _3988_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_22_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5727_ _5727_/A0 _6006_/A1 _5731_/S VGND VGND VPWR VPWR _5727_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5658_ _6028_/A1 hold532/X _5658_/S VGND VGND VPWR VPWR _5658_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4609_ _5189_/A _5316_/A _5094_/A _5109_/A VGND VGND VPWR VPWR _4760_/B sky130_fd_sc_hd__nand4_4
XFILLER_190_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5589_ _5553_/B _5589_/B _5589_/C VGND VGND VPWR VPWR _5589_/Y sky130_fd_sc_hd__nand3b_1
Xhold340 _5986_/X VGND VGND VPWR VPWR _7563_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7328_ _7557_/CLK _7328_/D fanout623/X VGND VGND VPWR VPWR _7328_/Q sky130_fd_sc_hd__dfrtp_1
Xhold351 _7571_/Q VGND VGND VPWR VPWR hold351/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 _4472_/X VGND VGND VPWR VPWR _7166_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold373 _7510_/Q VGND VGND VPWR VPWR hold373/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold384 _5942_/X VGND VGND VPWR VPWR _7524_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7259_ _7293_/CLK _7259_/D _6886_/A VGND VGND VPWR VPWR _7259_/Q sky130_fd_sc_hd__dfrtp_4
Xhold395 _7165_/Q VGND VGND VPWR VPWR hold395/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1040 _7194_/Q VGND VGND VPWR VPWR _4506_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1051 _4518_/X VGND VGND VPWR VPWR _7204_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1062 _4353_/X VGND VGND VPWR VPWR _7061_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1073 _4299_/X VGND VGND VPWR VPWR _7015_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1084 _5799_/X VGND VGND VPWR VPWR _7397_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1095 _4554_/X VGND VGND VPWR VPWR _7234_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_202 _7422_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_213 _7114_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_224 _7356_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_235 _7657_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_246 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_257 _4199_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_268 _4171_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_279 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4960_ _5146_/A _5112_/B VGND VGND VPWR VPWR _4960_/Y sky130_fd_sc_hd__nand2_8
XFILLER_83_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3911_ _7122_/Q _5903_/A _4535_/B _3843_/X _7296_/Q VGND VGND VPWR VPWR _3911_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_189_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4891_ _4953_/B _4950_/C _4901_/B _5401_/A VGND VGND VPWR VPWR _4891_/Y sky130_fd_sc_hd__nand4b_1
XFILLER_60_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6630_ _7479_/Q _6441_/X _6485_/X _7551_/Q _6629_/X VGND VGND VPWR VPWR _6630_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_60_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3842_ _7191_/Q _3543_/X _4511_/C _3696_/X _7201_/Q VGND VGND VPWR VPWR _3842_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6561_ _7605_/Q _6791_/B _6791_/C _6562_/B VGND VGND VPWR VPWR _6561_/X sky130_fd_sc_hd__and4_1
X_3773_ _7060_/Q _4346_/A _3769_/X _3771_/X _3772_/X VGND VGND VPWR VPWR _3774_/D
+ sky130_fd_sc_hd__a2111o_1
X_5512_ _4992_/D _5512_/B _5512_/C _5512_/D VGND VGND VPWR VPWR _5514_/D sky130_fd_sc_hd__nand4b_1
XFILLER_158_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6492_ _7610_/Q _6451_/X _6453_/X _7554_/Q _6491_/X VGND VGND VPWR VPWR _6492_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5443_ _5018_/Y _5440_/Y _5261_/Y _4879_/X _5392_/D VGND VGND VPWR VPWR _5447_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_172_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5374_ _5476_/A _4813_/B _5322_/A _4806_/X _4814_/A VGND VGND VPWR VPWR _5376_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_99_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7113_ _7233_/CLK _7113_/D fanout599/X VGND VGND VPWR VPWR _7113_/Q sky130_fd_sc_hd__dfstp_1
X_4325_ _4325_/A0 _6864_/A1 _4327_/S VGND VGND VPWR VPWR _4325_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7044_ _7227_/CLK _7044_/D fanout619/X VGND VGND VPWR VPWR _7044_/Q sky130_fd_sc_hd__dfstp_1
X_4256_ hold968/X _4255_/X _4258_/S VGND VGND VPWR VPWR _4256_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4187_ _6951_/Q _4187_/B VGND VGND VPWR VPWR _4188_/A sky130_fd_sc_hd__nor2_2
XFILLER_67_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6828_ _6827_/Y _6971_/Q _6969_/Q _6825_/Y VGND VGND VPWR VPWR _6828_/X sky130_fd_sc_hd__a22o_1
XFILLER_10_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6759_ _6742_/X _6749_/X _6759_/C _6759_/D VGND VGND VPWR VPWR _6759_/X sky130_fd_sc_hd__and4bb_1
XFILLER_183_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold170 _7494_/Q VGND VGND VPWR VPWR hold170/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 _5856_/X VGND VGND VPWR VPWR _7448_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold192 _4441_/X VGND VGND VPWR VPWR _7135_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_120_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4110_ input118/X input119/X _4110_/C _4110_/D VGND VGND VPWR VPWR _4116_/C sky130_fd_sc_hd__and4bb_1
XFILLER_68_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5090_ _5316_/A _5090_/B VGND VGND VPWR VPWR _5090_/Y sky130_fd_sc_hd__nand2_1
XFILLER_1_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4041_ _6914_/Q _7256_/Q _7257_/Q _7258_/Q VGND VGND VPWR VPWR _4174_/B sky130_fd_sc_hd__and4b_1
XFILLER_56_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5992_ hold825/X _6028_/A1 hold63/X VGND VGND VPWR VPWR _5992_/X sky130_fd_sc_hd__mux2_1
X_4943_ _4943_/A _4943_/B VGND VGND VPWR VPWR _4943_/Y sky130_fd_sc_hd__nand2_1
XFILLER_178_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7662_ _7662_/CLK _7662_/D fanout596/X VGND VGND VPWR VPWR _7662_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_177_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4874_ _4943_/A _5261_/D _5389_/B _5389_/C VGND VGND VPWR VPWR _4874_/Y sky130_fd_sc_hd__nand4_1
XFILLER_60_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6613_ _7567_/Q _6099_/B _6720_/D _6454_/X _7359_/Q VGND VGND VPWR VPWR _6613_/X
+ sky130_fd_sc_hd__a32o_1
X_3825_ _7187_/Q _5984_/A _5680_/A _3554_/X _7565_/Q VGND VGND VPWR VPWR _3825_/X
+ sky130_fd_sc_hd__a32o_1
X_7593_ _7607_/CLK _7593_/D fanout624/X VGND VGND VPWR VPWR _7593_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_193_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6544_ _7516_/Q _6645_/B _6562_/C _6458_/X _7420_/Q VGND VGND VPWR VPWR _6544_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_192_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3756_ _7582_/Q _6002_/A _5680_/B _3755_/X VGND VGND VPWR VPWR _3756_/X sky130_fd_sc_hd__a31o_1
XFILLER_118_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_5_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR _7202_/CLK sky130_fd_sc_hd__clkbuf_8
X_6475_ _7629_/Q _6485_/B _6443_/Y _4126_/B VGND VGND VPWR VPWR _6476_/D sky130_fd_sc_hd__a211o_1
XFILLER_165_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3687_ _4195_/A _4505_/B _4481_/A _3565_/X _7327_/Q VGND VGND VPWR VPWR _3687_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_173_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5426_ _5418_/X _5425_/Y _5413_/X _5414_/X VGND VGND VPWR VPWR _5428_/B sky130_fd_sc_hd__o211a_1
Xoutput220 _7698_/X VGND VGND VPWR VPWR mgmt_gpio_out[18] sky130_fd_sc_hd__buf_12
Xoutput231 _7708_/X VGND VGND VPWR VPWR mgmt_gpio_out[28] sky130_fd_sc_hd__buf_12
Xoutput242 _7690_/X VGND VGND VPWR VPWR mgmt_gpio_out[3] sky130_fd_sc_hd__buf_12
Xoutput253 _4186_/Y VGND VGND VPWR VPWR pad_flash_io0_oeb sky130_fd_sc_hd__buf_12
Xoutput264 _7263_/Q VGND VGND VPWR VPWR pll_div[2] sky130_fd_sc_hd__buf_12
XFILLER_102_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5357_ _5551_/A1 _5233_/A _5181_/C _4738_/A _4738_/B VGND VGND VPWR VPWR _5357_/X
+ sky130_fd_sc_hd__o311a_1
Xoutput275 _7136_/Q VGND VGND VPWR VPWR pll_trim[13] sky130_fd_sc_hd__buf_12
XFILLER_87_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput286 _7279_/Q VGND VGND VPWR VPWR pll_trim[23] sky130_fd_sc_hd__buf_12
XFILLER_87_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput297 _7281_/Q VGND VGND VPWR VPWR pwr_ctrl_out[0] sky130_fd_sc_hd__buf_12
X_4308_ _6006_/A1 _4308_/A1 _4312_/S VGND VGND VPWR VPWR _4308_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5288_ _5011_/C _5604_/B1 _4998_/Y _5001_/Y _5088_/Y VGND VGND VPWR VPWR _5288_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_75_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7027_ _7421_/CLK _7027_/D fanout630/X VGND VGND VPWR VPWR _7027_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_75_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4239_ _3618_/Y _4239_/A1 _4239_/S VGND VGND VPWR VPWR _6987_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire347 _3995_/Y VGND VGND VPWR VPWR _4037_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire358 _3667_/Y VGND VGND VPWR VPWR _3692_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_183_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3610_ _7457_/Q _3516_/X _6002_/A _6011_/A _7593_/Q VGND VGND VPWR VPWR _3610_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_175_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4590_ _4706_/D _4590_/B VGND VGND VPWR VPWR _4592_/D sky130_fd_sc_hd__nor2_1
XFILLER_128_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3541_ hold69/X _3622_/A _3622_/B hold96/X VGND VGND VPWR VPWR _4487_/A sky130_fd_sc_hd__and4bb_4
XFILLER_155_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold906 _7505_/Q VGND VGND VPWR VPWR hold906/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold917 _5749_/X VGND VGND VPWR VPWR _7353_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold928 hold928/A VGND VGND VPWR VPWR hold928/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold939 _7476_/Q VGND VGND VPWR VPWR hold939/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6260_ _7559_/Q _6131_/B _6432_/A3 _6160_/X _7375_/Q VGND VGND VPWR VPWR _6260_/X
+ sky130_fd_sc_hd__a32o_1
X_3472_ _7294_/Q _4171_/C _4171_/D VGND VGND VPWR VPWR _3472_/Y sky130_fd_sc_hd__nor3_1
XFILLER_182_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5211_ _5042_/A _5038_/B _5195_/X _5005_/C VGND VGND VPWR VPWR _5215_/B sky130_fd_sc_hd__a22oi_1
X_6191_ _7396_/Q _6114_/X _6119_/X _7412_/Q _6190_/X VGND VGND VPWR VPWR _6191_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_97_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5142_ _4992_/D _5404_/C _4805_/Y _5141_/Y VGND VGND VPWR VPWR _5142_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_96_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1606 _6920_/Q VGND VGND VPWR VPWR _4096_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1617 _4078_/X VGND VGND VPWR VPWR _6928_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1628 _7155_/Q VGND VGND VPWR VPWR _4459_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5073_ _5073_/A _5073_/B _5073_/C VGND VGND VPWR VPWR _5076_/B sky130_fd_sc_hd__nor3_1
Xhold1639 hold68/A VGND VGND VPWR VPWR _5520_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4024_ _7116_/Q _4541_/A _3535_/X _3545_/X _7402_/Q VGND VGND VPWR VPWR _4024_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_65_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5975_ _5993_/A _5975_/B _6038_/C VGND VGND VPWR VPWR _5983_/S sky130_fd_sc_hd__and3_4
XFILLER_52_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4926_ _5375_/C _4926_/B _4934_/C VGND VGND VPWR VPWR _4927_/B sky130_fd_sc_hd__and3_1
X_7714_ _7714_/A VGND VGND VPWR VPWR _7714_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7645_ _7662_/CLK _7645_/D fanout597/X VGND VGND VPWR VPWR _7645_/Q sky130_fd_sc_hd__dfrtp_1
X_4857_ _4633_/Y _4785_/Y _4783_/X _4950_/D VGND VGND VPWR VPWR _4953_/D sky130_fd_sc_hd__o211ai_4
XFILLER_138_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3808_ _7605_/Q _6029_/A _3583_/X input55/X _3807_/X VGND VGND VPWR VPWR _3815_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_165_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7576_ _7601_/CLK _7576_/D fanout611/X VGND VGND VPWR VPWR _7576_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4788_ _5143_/B _4595_/B _4779_/X _4781_/C _4781_/B VGND VGND VPWR VPWR _4788_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_118_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6527_ _7363_/Q _6445_/X _6471_/X _7323_/Q _6526_/X VGND VGND VPWR VPWR _6532_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_181_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3739_ _7462_/Q _4559_/B _5939_/B _3738_/X VGND VGND VPWR VPWR _3739_/X sky130_fd_sc_hd__a31o_1
XFILLER_109_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6458_ _7631_/Q _6485_/B _6645_/B _6771_/C VGND VGND VPWR VPWR _6458_/X sky130_fd_sc_hd__and4_4
XFILLER_134_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5409_ _5407_/A _5189_/D _4972_/C _4848_/Y _4972_/X VGND VGND VPWR VPWR _5409_/X
+ sky130_fd_sc_hd__a311o_1
X_6389_ _6387_/X _6379_/X _6388_/X VGND VGND VPWR VPWR _6389_/X sky130_fd_sc_hd__o21a_1
XFILLER_161_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5760_ _5760_/A0 hold44/A _5767_/S VGND VGND VPWR VPWR hold16/A sky130_fd_sc_hd__mux2_1
XFILLER_61_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4711_ _5186_/C _4946_/A _5186_/B VGND VGND VPWR VPWR _4711_/X sky130_fd_sc_hd__and3_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5691_ _5761_/A1 hold610/X _5695_/S VGND VGND VPWR VPWR _5691_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7430_ _7430_/CLK _7430_/D fanout627/X VGND VGND VPWR VPWR _7430_/Q sky130_fd_sc_hd__dfrtp_4
X_4642_ _4573_/A _4573_/B _5476_/D VGND VGND VPWR VPWR _5046_/B sky130_fd_sc_hd__a21oi_1
X_7361_ _7553_/CLK _7361_/D fanout624/X VGND VGND VPWR VPWR _7361_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_163_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4573_ _4573_/A _4573_/B VGND VGND VPWR VPWR _4950_/D sky130_fd_sc_hd__nand2_4
XFILLER_116_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold703 _5636_/X VGND VGND VPWR VPWR _7260_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold714 hold714/A VGND VGND VPWR VPWR hold714/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap422 _3568_/C VGND VGND VPWR VPWR _5768_/B sky130_fd_sc_hd__buf_6
X_6312_ _7449_/Q _6159_/B _6416_/C _6166_/C VGND VGND VPWR VPWR _6312_/X sky130_fd_sc_hd__o211a_1
X_3524_ hold73/X hold53/X _5686_/B VGND VGND VPWR VPWR _3550_/B sky130_fd_sc_hd__and3_4
X_7292_ _7293_/CLK _7292_/D fanout596/X VGND VGND VPWR VPWR _7292_/Q sky130_fd_sc_hd__dfrtp_4
Xhold725 hold725/A VGND VGND VPWR VPWR hold725/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold736 _7307_/Q VGND VGND VPWR VPWR hold736/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 _5708_/X VGND VGND VPWR VPWR _7316_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold758 _4426_/X VGND VGND VPWR VPWR _7122_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap466 _4215_/B VGND VGND VPWR VPWR _6855_/B1 sky130_fd_sc_hd__clkbuf_1
Xhold769 _7540_/Q VGND VGND VPWR VPWR hold769/X sky130_fd_sc_hd__dlygate4sd3_1
X_6243_ _7470_/Q _6130_/X _6241_/X _6242_/X VGND VGND VPWR VPWR _6243_/X sky130_fd_sc_hd__a211o_1
XFILLER_89_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3455_ _7349_/Q VGND VGND VPWR VPWR _3455_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_143_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6174_ _7547_/Q _6151_/X _6161_/X _7347_/Q _6173_/X VGND VGND VPWR VPWR _6174_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5125_ _5011_/C _4816_/Y _5611_/A2 _4991_/Y VGND VGND VPWR VPWR _5125_/X sky130_fd_sc_hd__a211o_1
Xhold1403 _7314_/Q VGND VGND VPWR VPWR hold277/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1414 _6985_/Q VGND VGND VPWR VPWR _4237_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1425 _7231_/Q VGND VGND VPWR VPWR hold1425/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1436 _5787_/X VGND VGND VPWR VPWR _7386_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1447 _7222_/Q VGND VGND VPWR VPWR hold472/A sky130_fd_sc_hd__dlygate4sd3_1
X_5056_ _5056_/A _5056_/B _5056_/C _5056_/D VGND VGND VPWR VPWR _5056_/Y sky130_fd_sc_hd__nor4_1
Xhold1458 _6636_/X VGND VGND VPWR VPWR _7655_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1469 _7378_/Q VGND VGND VPWR VPWR hold427/A sky130_fd_sc_hd__dlygate4sd3_1
X_4007_ _7346_/Q _5741_/A _4346_/A _7056_/Q _4006_/X VGND VGND VPWR VPWR _4007_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_609 _6039_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5958_ hold555/X _6039_/A1 _5965_/S VGND VGND VPWR VPWR _7538_/D sky130_fd_sc_hd__mux2_1
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4909_ _5000_/C _4836_/A _4777_/Y _4837_/Y _5007_/D VGND VGND VPWR VPWR _4934_/C
+ sky130_fd_sc_hd__o311a_4
XFILLER_166_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5889_ _5889_/A0 _6042_/A1 _5893_/S VGND VGND VPWR VPWR _5889_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7628_ _4167_/A1 _7628_/D fanout620/X VGND VGND VPWR VPWR _7628_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_193_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7559_ _7559_/CLK _7559_/D fanout613/X VGND VGND VPWR VPWR _7559_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_107_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold30 hold30/A VGND VGND VPWR VPWR hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A VGND VGND VPWR VPWR hold41/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold52 hold52/A VGND VGND VPWR VPWR hold52/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A VGND VGND VPWR VPWR hold63/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 hold74/A VGND VGND VPWR VPWR hold74/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold85 hold85/A VGND VGND VPWR VPWR hold85/X sky130_fd_sc_hd__clkbuf_16
XFILLER_76_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold96 hold96/A VGND VGND VPWR VPWR hold96/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_7__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _4167_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_43_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_5 _7244_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_746 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6930_ _7258_/CLK _6930_/D _6885_/X VGND VGND VPWR VPWR _6930_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_82_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6861_ _6861_/A hold98/X _6861_/C VGND VGND VPWR VPWR _6866_/S sky130_fd_sc_hd__and3_4
Xclkbuf_leaf_6_csclk _7236_/CLK VGND VGND VPWR VPWR _7682_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_62_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5812_ hold873/X _6046_/A1 _5812_/S VGND VGND VPWR VPWR _5812_/X sky130_fd_sc_hd__mux2_1
X_6792_ _7045_/Q _6451_/X _6483_/X _7070_/Q VGND VGND VPWR VPWR _6792_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5743_ _6040_/A1 hold984/X _5749_/S VGND VGND VPWR VPWR _7347_/D sky130_fd_sc_hd__mux2_1
XFILLER_148_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5674_ _5674_/A0 _6864_/A1 _5677_/S VGND VGND VPWR VPWR _5674_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4625_ _4948_/A _5074_/A _5189_/D VGND VGND VPWR VPWR _4625_/Y sky130_fd_sc_hd__nand3_2
XFILLER_148_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7413_ _7421_/CLK _7413_/D fanout628/X VGND VGND VPWR VPWR _7413_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_175_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold500 _7275_/Q VGND VGND VPWR VPWR hold500/X sky130_fd_sc_hd__dlygate4sd3_1
X_7344_ _7445_/CLK _7344_/D fanout622/X VGND VGND VPWR VPWR _7344_/Q sky130_fd_sc_hd__dfrtp_1
Xhold511 _7489_/Q VGND VGND VPWR VPWR hold511/X sky130_fd_sc_hd__dlygate4sd3_1
X_4556_ _4556_/A0 _4556_/A1 _4558_/S VGND VGND VPWR VPWR _4556_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold522 _5929_/X VGND VGND VPWR VPWR _7513_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 _5658_/X VGND VGND VPWR VPWR _7279_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3507_ hold188/X hold104/X _4229_/S VGND VGND VPWR VPWR _3673_/C sky130_fd_sc_hd__mux2_8
Xhold544 _4411_/X VGND VGND VPWR VPWR _7110_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7275_ _7462_/CLK _7275_/D fanout604/X VGND VGND VPWR VPWR _7275_/Q sky130_fd_sc_hd__dfstp_4
Xhold555 hold555/A VGND VGND VPWR VPWR hold555/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold566 _7497_/Q VGND VGND VPWR VPWR hold566/X sky130_fd_sc_hd__dlygate4sd3_1
X_4487_ _4487_/A _4487_/B _6861_/C VGND VGND VPWR VPWR _4492_/S sky130_fd_sc_hd__and3_2
XFILLER_143_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold577 _7321_/Q VGND VGND VPWR VPWR hold577/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold588 _5884_/X VGND VGND VPWR VPWR _7473_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6226_ _6159_/B _6212_/X _6225_/X VGND VGND VPWR VPWR _6226_/X sky130_fd_sc_hd__a21o_2
X_3438_ _7485_/Q VGND VGND VPWR VPWR _3438_/Y sky130_fd_sc_hd__inv_2
Xhold599 _4564_/X VGND VGND VPWR VPWR _7243_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6157_ _7626_/Q _6416_/B _6157_/C _6158_/D VGND VGND VPWR VPWR _6157_/X sky130_fd_sc_hd__and4b_4
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1200 _7004_/Q VGND VGND VPWR VPWR _4280_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1211 _4455_/A1 VGND VGND VPWR VPWR hold661/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1222 _4462_/A1 VGND VGND VPWR VPWR hold710/A sky130_fd_sc_hd__dlygate4sd3_1
X_5108_ _5109_/A _5108_/B _5291_/C _5452_/B VGND VGND VPWR VPWR _5108_/Y sky130_fd_sc_hd__nand4_1
Xhold1233 _6816_/A1 VGND VGND VPWR VPWR hold790/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1244 _7080_/Q VGND VGND VPWR VPWR hold570/A sky130_fd_sc_hd__dlygate4sd3_1
X_6088_ _7629_/Q _7628_/Q VGND VGND VPWR VPWR _6455_/C sky130_fd_sc_hd__and2b_4
Xhold1255 _4342_/X VGND VGND VPWR VPWR hold136/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1266 _7215_/Q VGND VGND VPWR VPWR hold967/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5039_ _5313_/B _5093_/C VGND VGND VPWR VPWR _5039_/Y sky130_fd_sc_hd__nand2_1
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1277 _6024_/X VGND VGND VPWR VPWR _7597_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1288 _4552_/X VGND VGND VPWR VPWR _7233_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_406 _4522_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1299 _5797_/X VGND VGND VPWR VPWR _7395_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_417 _6516_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_428 _6192_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_439 _6444_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_607 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput120 wb_adr_i[29] VGND VGND VPWR VPWR _4110_/C sky130_fd_sc_hd__clkbuf_1
Xinput131 wb_cyc_i VGND VGND VPWR VPWR _4116_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput142 wb_dat_i[19] VGND VGND VPWR VPWR _6840_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_163_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput153 wb_dat_i[29] VGND VGND VPWR VPWR _6846_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput164 wb_rstn_i VGND VGND VPWR VPWR input164/X sky130_fd_sc_hd__buf_2
XFILLER_76_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4410_ _4410_/A0 _6865_/A1 _4411_/S VGND VGND VPWR VPWR _4410_/X sky130_fd_sc_hd__mux2_1
X_5390_ _4769_/Y _4953_/C _4862_/Y _4871_/X VGND VGND VPWR VPWR _5390_/X sky130_fd_sc_hd__a211o_1
X_4341_ _5697_/A0 hold456/X _4345_/S VGND VGND VPWR VPWR _4341_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7060_ _7192_/CLK _7060_/D fanout617/X VGND VGND VPWR VPWR _7060_/Q sky130_fd_sc_hd__dfrtp_4
X_4272_ _4271_/X hold999/X _4276_/S VGND VGND VPWR VPWR _4272_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6011_ _6011_/A _6029_/B VGND VGND VPWR VPWR _6019_/S sky130_fd_sc_hd__nand2_8
XFILLER_100_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6913_ _4183_/A1 _6956_/Q _6868_/X VGND VGND VPWR VPWR _6913_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6844_ _6844_/A0 _6843_/X _6853_/S VGND VGND VPWR VPWR _7676_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3987_ _5669_/B _5666_/B _3970_/Y _3974_/X VGND VGND VPWR VPWR _3987_/X sky130_fd_sc_hd__a31o_1
X_6775_ _6775_/A _6775_/B _6775_/C _6775_/D VGND VGND VPWR VPWR _6775_/Y sky130_fd_sc_hd__nor4_1
X_5726_ hold329/X _5843_/A1 _5731_/S VGND VGND VPWR VPWR _5726_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5657_ hold50/X _5657_/A1 _5658_/S VGND VGND VPWR VPWR hold67/A sky130_fd_sc_hd__mux2_1
XFILLER_163_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4608_ _5014_/D _4990_/A VGND VGND VPWR VPWR _4608_/Y sky130_fd_sc_hd__nand2b_2
X_5588_ _5318_/B _5021_/B _5376_/A _4813_/X _5376_/B VGND VGND VPWR VPWR _5589_/C
+ sky130_fd_sc_hd__a2111oi_1
Xhold330 _5726_/X VGND VGND VPWR VPWR _7332_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 _7555_/Q VGND VGND VPWR VPWR hold341/X sky130_fd_sc_hd__dlygate4sd3_1
X_4539_ hold472/X _5673_/A1 _4540_/S VGND VGND VPWR VPWR _7222_/D sky130_fd_sc_hd__mux2_1
XFILLER_104_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7327_ _7435_/CLK _7327_/D fanout623/X VGND VGND VPWR VPWR _7327_/Q sky130_fd_sc_hd__dfrtp_1
Xhold352 _5995_/X VGND VGND VPWR VPWR _7571_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold363 _7032_/Q VGND VGND VPWR VPWR hold363/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 _5926_/X VGND VGND VPWR VPWR _7510_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold385 _7057_/Q VGND VGND VPWR VPWR hold385/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7258_ _7258_/CLK _7258_/D _6911_/X VGND VGND VPWR VPWR _7258_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_117_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold396 _4471_/X VGND VGND VPWR VPWR _7165_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6209_ _7389_/Q _6115_/X _6119_/X _7413_/Q _6208_/X VGND VGND VPWR VPWR _6209_/X
+ sky130_fd_sc_hd__a221o_1
X_7189_ _7207_/CLK _7189_/D fanout633/X VGND VGND VPWR VPWR _7189_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_98_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1030 _4294_/X VGND VGND VPWR VPWR _7011_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1041 _4506_/X VGND VGND VPWR VPWR _7194_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_133_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_727 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1052 _7697_/A VGND VGND VPWR VPWR _4246_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1063 hold1370/X VGND VGND VPWR VPWR _5934_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1074 hold1270/X VGND VGND VPWR VPWR _5889_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1085 hold1540/X VGND VGND VPWR VPWR _4562_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_203 _7430_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1096 _7116_/Q VGND VGND VPWR VPWR _4419_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_214 _7485_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_225 _7356_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_236 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_247 wb_clk_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_258 input41/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_269 _4195_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_71_csclk _7095_/CLK VGND VGND VPWR VPWR _7459_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3910_ _7132_/Q hold56/A hold75/A _7507_/Q _3909_/X VGND VGND VPWR VPWR _3910_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4890_ _4953_/C _4859_/Y _4878_/X _4900_/A VGND VGND VPWR VPWR _4890_/X sky130_fd_sc_hd__o31a_1
X_3841_ _5661_/A _5659_/C _5669_/B _4340_/A VGND VGND VPWR VPWR _3841_/X sky130_fd_sc_hd__o211a_1
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6560_ _6559_/X _6560_/A1 _6611_/S VGND VGND VPWR VPWR _7652_/D sky130_fd_sc_hd__mux2_1
X_3772_ _7342_/Q _6020_/A _4487_/B _3552_/X _7390_/Q VGND VGND VPWR VPWR _3772_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_192_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5511_ _5418_/X _5425_/A _5510_/X _5503_/X _5414_/X VGND VGND VPWR VPWR _5515_/B
+ sky130_fd_sc_hd__o311a_1
X_6491_ _7602_/Q _6456_/X _6460_/X _7442_/Q VGND VGND VPWR VPWR _6491_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5442_ _5245_/X _5442_/B _5442_/C VGND VGND VPWR VPWR _5621_/A sky130_fd_sc_hd__and3b_1
XFILLER_173_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5373_ _5429_/A _5313_/C _5322_/A _5372_/X _5371_/Y VGND VGND VPWR VPWR _5376_/C
+ sky130_fd_sc_hd__a311o_1
XFILLER_172_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_24_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7254_/CLK sky130_fd_sc_hd__clkbuf_16
X_7112_ _7233_/CLK _7112_/D fanout599/X VGND VGND VPWR VPWR _7112_/Q sky130_fd_sc_hd__dfrtp_2
X_4324_ hold738/X _6863_/A1 _4327_/S VGND VGND VPWR VPWR _4324_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7043_ _7558_/CLK _7043_/D fanout615/X VGND VGND VPWR VPWR _7043_/Q sky130_fd_sc_hd__dfrtp_1
X_4255_ hold604/X _5991_/A1 _4257_/S VGND VGND VPWR VPWR _4255_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4186_ _4186_/A VGND VGND VPWR VPWR _4186_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_39_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7408_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_55_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_1_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR _7236_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_94_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6827_ _6827_/A _6827_/B VGND VGND VPWR VPWR _6827_/Y sky130_fd_sc_hd__nand2_1
XFILLER_11_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6758_ _6758_/A _6758_/B _6758_/C _6758_/D VGND VGND VPWR VPWR _6759_/C sky130_fd_sc_hd__nor4_1
XFILLER_10_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5709_ hold9/X _5709_/A1 hold38/X VGND VGND VPWR VPWR hold39/A sky130_fd_sc_hd__mux2_1
X_6689_ _7121_/Q _6441_/X _6456_/X _7159_/Q _6688_/X VGND VGND VPWR VPWR _6689_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_164_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold160 _7579_/Q VGND VGND VPWR VPWR hold160/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 _5908_/X VGND VGND VPWR VPWR _7494_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold182 _7686_/Q VGND VGND VPWR VPWR hold182/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_616 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold193 _7273_/Q VGND VGND VPWR VPWR hold193/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout640 _5008_/C VGND VGND VPWR VPWR _5017_/B sky130_fd_sc_hd__buf_12
XFILLER_120_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4040_ _7258_/Q _7257_/Q _7256_/Q VGND VGND VPWR VPWR _4192_/C sky130_fd_sc_hd__and3_2
XFILLER_49_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5991_ hold726/X _5991_/A1 hold63/X VGND VGND VPWR VPWR _7568_/D sky130_fd_sc_hd__mux2_1
X_4942_ _5375_/C _4957_/B _5261_/D _5389_/C VGND VGND VPWR VPWR _5268_/A sky130_fd_sc_hd__and4_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7661_ _7662_/CLK _7661_/D fanout596/X VGND VGND VPWR VPWR _7661_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4873_ _5452_/A _5389_/C VGND VGND VPWR VPWR _4873_/Y sky130_fd_sc_hd__nand2_2
XFILLER_178_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6612_ _7439_/Q _6097_/X _6445_/C _6483_/X _7391_/Q VGND VGND VPWR VPWR _6612_/X
+ sky130_fd_sc_hd__a32o_1
X_3824_ _7517_/Q _3555_/X _3701_/X _7242_/Q _3823_/X VGND VGND VPWR VPWR _3824_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_178_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7592_ _7601_/CLK _7592_/D fanout611/X VGND VGND VPWR VPWR _7592_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_165_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3755_ _7040_/Q _5678_/C _4505_/B _3695_/X _7050_/Q VGND VGND VPWR VPWR _3755_/X
+ sky130_fd_sc_hd__a32o_1
X_6543_ _7412_/Q _6450_/X _6483_/X _7388_/Q VGND VGND VPWR VPWR _6543_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3686_ _7407_/Q _3545_/X _3684_/X _3685_/X VGND VGND VPWR VPWR _3691_/B sky130_fd_sc_hd__a211o_1
X_6474_ _6474_/A _6474_/B _6474_/C _6474_/D VGND VGND VPWR VPWR _6476_/C sky130_fd_sc_hd__nor4_1
XFILLER_118_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput210 _3452_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[7] sky130_fd_sc_hd__buf_12
X_5425_ _5425_/A _5425_/B _5425_/C _5424_/X VGND VGND VPWR VPWR _5425_/Y sky130_fd_sc_hd__nor4b_1
XFILLER_161_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput221 _7699_/X VGND VGND VPWR VPWR mgmt_gpio_out[19] sky130_fd_sc_hd__buf_12
XFILLER_173_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput232 _7709_/X VGND VGND VPWR VPWR mgmt_gpio_out[29] sky130_fd_sc_hd__buf_12
Xoutput243 _7691_/X VGND VGND VPWR VPWR mgmt_gpio_out[4] sky130_fd_sc_hd__buf_12
Xoutput254 _7713_/X VGND VGND VPWR VPWR pad_flash_io1_do sky130_fd_sc_hd__buf_12
X_5356_ _5551_/A1 _5233_/A _5181_/C _4747_/B VGND VGND VPWR VPWR _5490_/A sky130_fd_sc_hd__o31a_1
Xoutput265 _7264_/Q VGND VGND VPWR VPWR pll_div[3] sky130_fd_sc_hd__buf_12
Xoutput276 _7137_/Q VGND VGND VPWR VPWR pll_trim[14] sky130_fd_sc_hd__buf_12
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput287 _6958_/Q VGND VGND VPWR VPWR pll_trim[24] sky130_fd_sc_hd__buf_12
XFILLER_102_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4307_ _5789_/A1 hold139/X _4312_/S VGND VGND VPWR VPWR _4307_/X sky130_fd_sc_hd__mux2_1
Xoutput298 _7282_/Q VGND VGND VPWR VPWR pwr_ctrl_out[1] sky130_fd_sc_hd__buf_12
XFILLER_87_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5287_ _5011_/C _5604_/B1 _4991_/Y _4998_/Y _5088_/Y VGND VGND VPWR VPWR _5287_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_141_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4238_ _3655_/Y _4238_/A1 _4239_/S VGND VGND VPWR VPWR _6986_/D sky130_fd_sc_hd__mux2_1
X_7026_ _7583_/CLK _7026_/D fanout630/X VGND VGND VPWR VPWR _7026_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4169_ _7634_/Q _7289_/Q _7292_/Q VGND VGND VPWR VPWR _4169_/X sky130_fd_sc_hd__mux2_2
XFILLER_83_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire348 _3883_/Y VGND VGND VPWR VPWR _3902_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire359 _3597_/Y VGND VGND VPWR VPWR _3618_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_191_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout470 _6445_/C VGND VGND VPWR VPWR _6771_/C sky130_fd_sc_hd__buf_6
XFILLER_65_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3540_ _3673_/B _3622_/A VGND VGND VPWR VPWR _5659_/C sky130_fd_sc_hd__nor2_8
Xhold907 _5920_/X VGND VGND VPWR VPWR _7505_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold918 _7593_/Q VGND VGND VPWR VPWR hold918/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_127_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3471_ _3474_/A1 _3470_/B hold1641/X VGND VGND VPWR VPWR _6954_/D sky130_fd_sc_hd__o21bai_1
XFILLER_143_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold929 _7343_/Q VGND VGND VPWR VPWR hold929/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5210_ _5196_/A _5061_/A _5005_/C _4985_/B _5110_/C VGND VGND VPWR VPWR _5616_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6190_ _7324_/Q _6067_/X _6145_/C _6077_/X _7380_/Q VGND VGND VPWR VPWR _6190_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_170_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5141_ _5551_/A1 _5322_/A _5071_/C _5140_/X _5139_/Y VGND VGND VPWR VPWR _5141_/Y
+ sky130_fd_sc_hd__a311oi_1
Xhold1607 _7257_/Q VGND VGND VPWR VPWR _3468_/B1 sky130_fd_sc_hd__dlygate4sd3_1
X_5072_ _4673_/X _5322_/A _5068_/C _5318_/B _5551_/A1 VGND VGND VPWR VPWR _5579_/A
+ sky130_fd_sc_hd__a32o_1
Xhold1618 _6929_/Q VGND VGND VPWR VPWR _4070_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1629 _7657_/Q VGND VGND VPWR VPWR _6687_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_4023_ _7434_/Q _4541_/A _5984_/B _3585_/X _7330_/Q VGND VGND VPWR VPWR _4023_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5974_ hold851/X _6046_/A1 _5974_/S VGND VGND VPWR VPWR _5974_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7713_ _7713_/A VGND VGND VPWR VPWR _7713_/X sky130_fd_sc_hd__clkbuf_2
X_4925_ _5452_/A _4957_/C _4925_/C VGND VGND VPWR VPWR _4927_/A sky130_fd_sc_hd__and3_1
X_7644_ _7657_/CLK _7644_/D fanout606/X VGND VGND VPWR VPWR _7644_/Q sky130_fd_sc_hd__dfrtp_1
X_4856_ _5476_/A _4966_/A _4946_/B VGND VGND VPWR VPWR _4955_/A sky130_fd_sc_hd__and3_1
XFILLER_193_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3807_ _7685_/Q _6861_/A hold98/A _3779_/X VGND VGND VPWR VPWR _3807_/X sky130_fd_sc_hd__a31o_1
X_7575_ _7601_/CLK _7575_/D fanout611/X VGND VGND VPWR VPWR _7575_/Q sky130_fd_sc_hd__dfrtp_1
X_4787_ _4633_/Y _4785_/Y _4782_/Y _5096_/A VGND VGND VPWR VPWR _4787_/Y sky130_fd_sc_hd__a2bb2oi_2
XFILLER_20_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6526_ _7515_/Q _6645_/B _6562_/C _6474_/C _7371_/Q VGND VGND VPWR VPWR _6526_/X
+ sky130_fd_sc_hd__a32o_1
X_3738_ _7265_/Q _5939_/B _5678_/C _3710_/X _7075_/Q VGND VGND VPWR VPWR _3738_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_118_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6457_ _6791_/B _6791_/D _6645_/C VGND VGND VPWR VPWR _6457_/X sky130_fd_sc_hd__and3_4
XFILLER_173_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3669_ _7551_/Q _3514_/X _3558_/X _7559_/Q _3668_/X VGND VGND VPWR VPWR _3678_/A
+ sky130_fd_sc_hd__a221o_1
X_5408_ _5042_/A _4972_/C _4850_/X _5280_/X _5406_/X VGND VGND VPWR VPWR _5408_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_134_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6388_ _7038_/Q _6082_/Y _6811_/S VGND VGND VPWR VPWR _6388_/X sky130_fd_sc_hd__o21ba_1
XFILLER_161_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5339_ _4629_/Y _4657_/Y _4750_/Y _4821_/Y _5011_/C VGND VGND VPWR VPWR _5339_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7009_ _7584_/CLK _7009_/D fanout613/X VGND VGND VPWR VPWR _7692_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_75_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_6__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _7679_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4710_ _4760_/D _4760_/C _4760_/B _4946_/A VGND VGND VPWR VPWR _4710_/Y sky130_fd_sc_hd__nand4_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5690_ _6012_/A0 _5690_/A1 _5695_/S VGND VGND VPWR VPWR _5690_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4641_ _5096_/A _4637_/A _4639_/Y _4584_/Y VGND VGND VPWR VPWR _5476_/D sky130_fd_sc_hd__o2bb2ai_4
XFILLER_175_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4572_ _4573_/A _4573_/B VGND VGND VPWR VPWR _4572_/X sky130_fd_sc_hd__and2_4
X_7360_ _7568_/CLK _7360_/D fanout622/X VGND VGND VPWR VPWR _7360_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_162_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap412 _3546_/C VGND VGND VPWR VPWR _6020_/A sky130_fd_sc_hd__clkbuf_16
Xhold704 hold704/A VGND VGND VPWR VPWR hold704/X sky130_fd_sc_hd__dlygate4sd3_1
X_6311_ _7361_/Q _6159_/B _6137_/X _6157_/X _7505_/Q VGND VGND VPWR VPWR _6311_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_116_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3523_ hold53/X _5686_/B VGND VGND VPWR VPWR _5768_/C sky130_fd_sc_hd__and2_4
Xhold715 hold715/A VGND VGND VPWR VPWR wb_dat_o[9] sky130_fd_sc_hd__buf_12
XFILLER_116_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7291_ _7291_/CLK hold51/X fanout596/X VGND VGND VPWR VPWR _7291_/Q sky130_fd_sc_hd__dfrtp_1
Xhold726 hold726/A VGND VGND VPWR VPWR hold726/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold737 _5698_/X VGND VGND VPWR VPWR _7307_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap456 _6113_/Y VGND VGND VPWR VPWR wire455/A sky130_fd_sc_hd__clkbuf_2
Xhold748 _7696_/A VGND VGND VPWR VPWR hold748/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold759 _7495_/Q VGND VGND VPWR VPWR hold759/X sky130_fd_sc_hd__dlygate4sd3_1
X_6242_ _7526_/Q _6309_/B _6334_/C _6157_/X _7502_/Q VGND VGND VPWR VPWR _6242_/X
+ sky130_fd_sc_hd__a32o_1
X_3454_ _7357_/Q VGND VGND VPWR VPWR _3454_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_170_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6173_ _7491_/Q _6309_/B _6407_/A3 _6144_/X _7539_/Q VGND VGND VPWR VPWR _6173_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_130_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5124_ _4948_/A _4704_/A _5611_/A2 _4991_/Y _5123_/X VGND VGND VPWR VPWR _5124_/Y
+ sky130_fd_sc_hd__o41ai_1
Xhold1404 _7295_/Q VGND VGND VPWR VPWR _5683_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1415 _7514_/Q VGND VGND VPWR VPWR hold297/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1426 _4550_/X VGND VGND VPWR VPWR _7231_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1437 _7123_/Q VGND VGND VPWR VPWR hold1437/X sky130_fd_sc_hd__dlygate4sd3_1
X_5055_ _5036_/X _5055_/B _5055_/C _5055_/D VGND VGND VPWR VPWR _5056_/D sky130_fd_sc_hd__nand4b_1
Xhold1448 _7659_/Q VGND VGND VPWR VPWR _6761_/B1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1459 _7482_/Q VGND VGND VPWR VPWR hold365/A sky130_fd_sc_hd__dlygate4sd3_1
X_4006_ _7209_/Q hold70/A _4511_/C _3696_/X _7199_/Q VGND VGND VPWR VPWR _4006_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_65_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5957_ _5993_/A _5957_/B _6038_/C VGND VGND VPWR VPWR _5965_/S sky130_fd_sc_hd__and3_4
XFILLER_111_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4908_ _4908_/A _4908_/B _4908_/C VGND VGND VPWR VPWR _4915_/C sky130_fd_sc_hd__nand3_1
XFILLER_139_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5888_ hold939/X _6041_/A1 _5893_/S VGND VGND VPWR VPWR _5888_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7627_ _4167_/A1 _7627_/D fanout619/X VGND VGND VPWR VPWR _7627_/Q sky130_fd_sc_hd__dfstp_2
X_4839_ _4907_/A VGND VGND VPWR VPWR _4935_/B sky130_fd_sc_hd__clkinv_2
XFILLER_138_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7558_ _7558_/CLK _7558_/D fanout615/X VGND VGND VPWR VPWR _7558_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_107_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6509_ _7314_/Q _6759_/D _6109_/X VGND VGND VPWR VPWR _6509_/X sky130_fd_sc_hd__o21a_1
XFILLER_134_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7489_ _7616_/CLK _7489_/D fanout610/X VGND VGND VPWR VPWR _7489_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold20 hold20/A VGND VGND VPWR VPWR hold20/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 hold31/A VGND VGND VPWR VPWR hold31/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold42 hold42/A VGND VGND VPWR VPWR hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hold53/A VGND VGND VPWR VPWR hold53/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 hold64/A VGND VGND VPWR VPWR hold64/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A VGND VGND VPWR VPWR hold75/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 hold86/A VGND VGND VPWR VPWR hold86/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 hold97/A VGND VGND VPWR VPWR hold97/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_6 _5631_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6860_ _6827_/A _6857_/X _6859_/X VGND VGND VPWR VPWR _7681_/D sky130_fd_sc_hd__a21o_1
XFILLER_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5811_ hold694/X _5991_/A1 _5812_/S VGND VGND VPWR VPWR _5811_/X sky130_fd_sc_hd__mux2_1
X_6791_ _7163_/Q _6791_/B _6791_/C _6791_/D VGND VGND VPWR VPWR _6791_/X sky130_fd_sc_hd__and4_1
XFILLER_15_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5742_ _6003_/A1 hold417/X _5749_/S VGND VGND VPWR VPWR _7346_/D sky130_fd_sc_hd__mux2_1
X_5673_ hold444/X _5673_/A1 _5677_/S VGND VGND VPWR VPWR _5673_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7412_ _7430_/CLK _7412_/D fanout627/X VGND VGND VPWR VPWR _7412_/Q sky130_fd_sc_hd__dfrtp_1
X_4624_ _5189_/A _5074_/A _5189_/D VGND VGND VPWR VPWR _5196_/A sky130_fd_sc_hd__and3_4
XFILLER_163_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold501 _7067_/Q VGND VGND VPWR VPWR hold501/X sky130_fd_sc_hd__dlygate4sd3_1
X_7343_ _7408_/CLK _7343_/D fanout628/X VGND VGND VPWR VPWR _7343_/Q sky130_fd_sc_hd__dfrtp_1
X_4555_ hold438/X _5761_/A1 _4558_/S VGND VGND VPWR VPWR _4555_/X sky130_fd_sc_hd__mux2_1
Xhold512 _5902_/X VGND VGND VPWR VPWR _7489_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 _7320_/Q VGND VGND VPWR VPWR hold523/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 hold534/A VGND VGND VPWR VPWR hold534/X sky130_fd_sc_hd__dlygate4sd3_1
X_3506_ hold21/X _3478_/X hold187/X VGND VGND VPWR VPWR _3506_/X sky130_fd_sc_hd__a21bo_1
Xhold545 _7520_/Q VGND VGND VPWR VPWR hold545/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold556 hold556/A VGND VGND VPWR VPWR hold556/X sky130_fd_sc_hd__dlygate4sd3_1
X_7274_ _7286_/CLK _7274_/D fanout598/X VGND VGND VPWR VPWR _7274_/Q sky130_fd_sc_hd__dfstp_1
X_4486_ hold596/X _4564_/A1 _4486_/S VGND VGND VPWR VPWR _4486_/X sky130_fd_sc_hd__mux2_1
Xhold567 _5911_/X VGND VGND VPWR VPWR _7497_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold578 _5713_/X VGND VGND VPWR VPWR _7321_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold589 _7344_/Q VGND VGND VPWR VPWR hold589/X sky130_fd_sc_hd__dlygate4sd3_1
X_6225_ _7421_/Q _6150_/X _6213_/X _6215_/X _6224_/X VGND VGND VPWR VPWR _6225_/X
+ sky130_fd_sc_hd__a2111o_1
X_3437_ hold40/A VGND VGND VPWR VPWR _3437_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6156_ _6131_/B _6143_/X _6148_/X _6155_/X _6140_/X VGND VGND VPWR VPWR _6156_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_106_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1201 _4280_/X VGND VGND VPWR VPWR _7004_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1212 _4452_/A1 VGND VGND VPWR VPWR hold657/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1223 _4447_/A1 VGND VGND VPWR VPWR hold704/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5107_ _5452_/B _5107_/B VGND VGND VPWR VPWR _5127_/B sky130_fd_sc_hd__nand2_1
Xhold1234 _6814_/B2 VGND VGND VPWR VPWR hold941/A sky130_fd_sc_hd__dlygate4sd3_1
X_6087_ _6109_/B _6086_/C _6086_/Y VGND VGND VPWR VPWR _7628_/D sky130_fd_sc_hd__a21oi_1
Xhold1245 _4375_/X VGND VGND VPWR VPWR _7080_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_181_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1256 _7682_/Q VGND VGND VPWR VPWR hold1256/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1267 _4531_/X VGND VGND VPWR VPWR _7215_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1278 _7399_/Q VGND VGND VPWR VPWR hold934/A sky130_fd_sc_hd__dlygate4sd3_1
X_5038_ _5042_/A _5038_/B VGND VGND VPWR VPWR _5051_/C sky130_fd_sc_hd__nand2_1
Xhold1289 _7516_/Q VGND VGND VPWR VPWR hold957/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_407 _5233_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_418 _6131_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_429 _6192_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6989_ _7421_/CLK _6989_/D fanout630/X VGND VGND VPWR VPWR _7697_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_53_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput110 wb_adr_i[1] VGND VGND VPWR VPWR _4992_/A sky130_fd_sc_hd__buf_2
XFILLER_163_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput121 wb_adr_i[2] VGND VGND VPWR VPWR _5462_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput132 wb_dat_i[0] VGND VGND VPWR VPWR _6831_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput143 wb_dat_i[1] VGND VGND VPWR VPWR _6834_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput154 wb_dat_i[2] VGND VGND VPWR VPWR _6837_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput165 wb_sel_i[0] VGND VGND VPWR VPWR _6826_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_64_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4340_ _4340_/A _4493_/C _5680_/B _5686_/D VGND VGND VPWR VPWR _4340_/Y sky130_fd_sc_hd__nand4_4
XFILLER_98_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4271_ hold798/X _5999_/A1 _4275_/S VGND VGND VPWR VPWR _4271_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6010_ hold912/X _6046_/A1 _6010_/S VGND VGND VPWR VPWR _6010_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6912_ _7258_/CLK _6955_/Q _6867_/X VGND VGND VPWR VPWR _6912_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_47_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6843_ _6971_/Q _6843_/A2 _6843_/B1 wire537/X _6842_/X VGND VGND VPWR VPWR _6843_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_23_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6774_ _7049_/Q _6471_/X _6770_/X _6771_/X _6773_/X VGND VGND VPWR VPWR _6775_/D
+ sky130_fd_sc_hd__a2111o_1
X_3986_ _7514_/Q _3555_/X _4388_/A _7091_/Q _3985_/X VGND VGND VPWR VPWR _3986_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5725_ hold980/X _6040_/A1 _5731_/S VGND VGND VPWR VPWR _5725_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5656_ hold85/X _5656_/A1 _5658_/S VGND VGND VPWR VPWR hold86/A sky130_fd_sc_hd__mux2_1
XFILLER_163_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4607_ _5014_/D _4990_/A VGND VGND VPWR VPWR _5109_/A sky130_fd_sc_hd__and2b_4
XFILLER_117_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5587_ _5587_/A _5618_/B VGND VGND VPWR VPWR _5587_/Y sky130_fd_sc_hd__nand2_1
Xhold320 _5744_/X VGND VGND VPWR VPWR _7348_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold331 _7603_/Q VGND VGND VPWR VPWR hold331/X sky130_fd_sc_hd__dlygate4sd3_1
X_7326_ _7430_/CLK _7326_/D fanout627/X VGND VGND VPWR VPWR _7326_/Q sky130_fd_sc_hd__dfrtp_2
X_4538_ _4538_/A0 _6864_/A1 _4540_/S VGND VGND VPWR VPWR _7221_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold342 _5977_/X VGND VGND VPWR VPWR _7555_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 _7595_/Q VGND VGND VPWR VPWR hold353/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold364 _4318_/X VGND VGND VPWR VPWR _7032_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold375 _7042_/Q VGND VGND VPWR VPWR hold375/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7257_ _4183_/A1 _7257_/D _6910_/X VGND VGND VPWR VPWR _7257_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_171_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold386 _4348_/X VGND VGND VPWR VPWR _7057_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4469_ _4487_/B _4469_/B _6861_/C VGND VGND VPWR VPWR _4474_/S sky130_fd_sc_hd__and3_2
XFILLER_89_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold397 _7253_/Q VGND VGND VPWR VPWR hold397/X sky130_fd_sc_hd__dlygate4sd3_1
X_6208_ _4171_/C _6157_/C _6145_/C _6077_/X _7381_/Q VGND VGND VPWR VPWR _6208_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_58_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7188_ _7236_/CLK _7188_/D fanout603/X VGND VGND VPWR VPWR _7188_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6139_ _7506_/Q _6136_/X _6138_/X _7354_/Q _6135_/X VGND VGND VPWR VPWR _6139_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1020 hold1485/X VGND VGND VPWR VPWR _4520_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1031 hold1320/X VGND VGND VPWR VPWR _5763_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1042 _7041_/Q VGND VGND VPWR VPWR _4329_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1053 _4246_/X VGND VGND VPWR VPWR _6989_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1064 _7509_/Q VGND VGND VPWR VPWR _5925_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1075 _7023_/Q VGND VGND VPWR VPWR _4308_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1086 _7389_/Q VGND VGND VPWR VPWR _5790_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1097 _4419_/X VGND VGND VPWR VPWR _7116_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_204 _7445_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_215 hold40/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_226 _7060_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_237 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_248 hold52/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_259 input58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_5_csclk _7236_/CLK VGND VGND VPWR VPWR _7238_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_150_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3840_ _3903_/A1 _3839_/X _3904_/S VGND VGND VPWR VPWR _3840_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3771_ _7350_/Q _5957_/B _4511_/C _3770_/X VGND VGND VPWR VPWR _3771_/X sky130_fd_sc_hd__a31o_1
XFILLER_192_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5510_ _5625_/B _5610_/C _5560_/D _5560_/A VGND VGND VPWR VPWR _5510_/X sky130_fd_sc_hd__and4bb_1
XFILLER_9_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6490_ _7394_/Q _6463_/X _6483_/X _7386_/Q _6455_/X VGND VGND VPWR VPWR _6490_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5441_ _4859_/Y _4960_/Y _5004_/Y _4873_/Y _4912_/Y VGND VGND VPWR VPWR _5442_/C
+ sky130_fd_sc_hd__o32a_1
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5372_ _5551_/A1 _5181_/C _5595_/B _5186_/C _5375_/A VGND VGND VPWR VPWR _5372_/X
+ sky130_fd_sc_hd__o2111a_1
X_7111_ _7233_/CLK _7111_/D fanout599/X VGND VGND VPWR VPWR _7111_/Q sky130_fd_sc_hd__dfrtp_4
X_4323_ _4323_/A0 _5697_/A0 _4327_/S VGND VGND VPWR VPWR _4323_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7042_ _7498_/CLK _7042_/D fanout615/X VGND VGND VPWR VPWR _7042_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_86_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4254_ hold537/X _4253_/X _4258_/S VGND VGND VPWR VPWR _4254_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4185_ _6923_/Q _4185_/B VGND VGND VPWR VPWR _4186_/A sky130_fd_sc_hd__nand2b_2
XFILLER_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6826_ _6827_/A _6826_/A2 _6967_/Q VGND VGND VPWR VPWR _6858_/D sky130_fd_sc_hd__a21bo_1
XFILLER_23_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6757_ _7098_/Q _6444_/X _6459_/X _7118_/Q _6756_/X VGND VGND VPWR VPWR _6758_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_149_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3969_ _6923_/Q _6920_/Q _7285_/Q VGND VGND VPWR VPWR _3970_/A sky130_fd_sc_hd__nor3_1
XFILLER_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5708_ _6041_/A1 hold746/X hold38/X VGND VGND VPWR VPWR _5708_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6688_ _7204_/Q _6099_/B _6720_/D _6454_/X _7189_/Q VGND VGND VPWR VPWR _6688_/X
+ sky130_fd_sc_hd__a32o_1
X_5639_ hold802/X _6863_/A1 _5642_/S VGND VGND VPWR VPWR _5639_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold150 _5923_/X VGND VGND VPWR VPWR _7507_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7309_ _7616_/CLK hold10/X fanout608/X VGND VGND VPWR VPWR _7309_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_105_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold161 _6004_/X VGND VGND VPWR VPWR _7579_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 _7475_/Q VGND VGND VPWR VPWR hold172/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 _6866_/X VGND VGND VPWR VPWR _7686_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 _5652_/X VGND VGND VPWR VPWR _7273_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout630 fanout631/X VGND VGND VPWR VPWR fanout630/X sky130_fd_sc_hd__buf_8
Xfanout641 _4822_/A VGND VGND VPWR VPWR _4948_/B sky130_fd_sc_hd__buf_12
XFILLER_77_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5990_ hold943/X _5999_/A1 hold63/X VGND VGND VPWR VPWR _5990_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4941_ _4941_/A _4941_/B VGND VGND VPWR VPWR _4941_/Y sky130_fd_sc_hd__nor2_1
X_7660_ _7662_/CLK _7660_/D fanout597/X VGND VGND VPWR VPWR _7660_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_178_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4872_ _5146_/B _4836_/B _5017_/A _4865_/C VGND VGND VPWR VPWR _5389_/C sky130_fd_sc_hd__o211a_4
XANTENNA_590 _4116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6611_ _6610_/X _6611_/A1 _6611_/S VGND VGND VPWR VPWR _7654_/D sky130_fd_sc_hd__mux2_1
X_3823_ _7094_/Q _6861_/A _4505_/B _3822_/X VGND VGND VPWR VPWR _3823_/X sky130_fd_sc_hd__a31o_1
X_7591_ _7599_/CLK _7591_/D fanout629/X VGND VGND VPWR VPWR _7591_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_177_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6542_ _7524_/Q _6447_/X _6474_/C _7372_/Q _6538_/X VGND VGND VPWR VPWR _6542_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_186_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3754_ _7233_/Q _5984_/A _5678_/B _3514_/X _7550_/Q VGND VGND VPWR VPWR _3754_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_146_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6473_ _6694_/B _6771_/C _6451_/X _6467_/X _6563_/C VGND VGND VPWR VPWR _6474_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_118_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3685_ input49/X _4481_/A _5666_/B _3571_/X _7359_/Q VGND VGND VPWR VPWR _3685_/X
+ sky130_fd_sc_hd__a32o_1
X_5424_ _5611_/A2 _5013_/Y _5412_/X _5299_/X _5560_/C VGND VGND VPWR VPWR _5424_/X
+ sky130_fd_sc_hd__o311a_1
Xoutput200 _3427_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[32] sky130_fd_sc_hd__buf_12
XFILLER_145_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput211 _3451_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[8] sky130_fd_sc_hd__buf_12
Xoutput222 _4160_/X VGND VGND VPWR VPWR mgmt_gpio_out[1] sky130_fd_sc_hd__buf_12
Xoutput233 _7689_/X VGND VGND VPWR VPWR mgmt_gpio_out[2] sky130_fd_sc_hd__buf_12
XFILLER_160_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput244 _7692_/X VGND VGND VPWR VPWR mgmt_gpio_out[5] sky130_fd_sc_hd__buf_12
X_5355_ _5189_/A _5189_/D _5614_/C _5551_/A1 VGND VGND VPWR VPWR _5595_/C sky130_fd_sc_hd__a211o_2
Xoutput255 _4188_/A VGND VGND VPWR VPWR pad_flash_io1_ieb sky130_fd_sc_hd__buf_12
Xoutput266 _7265_/Q VGND VGND VPWR VPWR pll_div[4] sky130_fd_sc_hd__buf_12
Xoutput277 _7138_/Q VGND VGND VPWR VPWR pll_trim[15] sky130_fd_sc_hd__buf_12
Xoutput288 _6959_/Q VGND VGND VPWR VPWR pll_trim[25] sky130_fd_sc_hd__buf_12
X_4306_ _5761_/A1 hold214/X _4311_/S VGND VGND VPWR VPWR _4306_/X sky130_fd_sc_hd__mux2_1
Xoutput299 _7283_/Q VGND VGND VPWR VPWR pwr_ctrl_out[2] sky130_fd_sc_hd__buf_12
XFILLER_114_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5286_ _5146_/A _5146_/B _5112_/B _5404_/A VGND VGND VPWR VPWR _5313_/A sky130_fd_sc_hd__a22o_2
XFILLER_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7025_ _7583_/CLK _7025_/D fanout629/X VGND VGND VPWR VPWR _7025_/Q sky130_fd_sc_hd__dfrtp_1
X_4237_ _3692_/Y _4237_/A1 _4239_/S VGND VGND VPWR VPWR _6985_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4168_ _7001_/Q input93/X _7297_/Q VGND VGND VPWR VPWR _4168_/X sky130_fd_sc_hd__mux2_4
XFILLER_55_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_5__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _7672_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_67_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4099_ _4099_/A0 input58/X _4099_/S VGND VGND VPWR VPWR _6918_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6809_ _6809_/A _6809_/B _6809_/C _6809_/D VGND VGND VPWR VPWR _6809_/Y sky130_fd_sc_hd__nor4_1
XFILLER_23_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire349 _3774_/Y VGND VGND VPWR VPWR _3775_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_136_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout460 _6427_/A3 VGND VGND VPWR VPWR _6146_/C sky130_fd_sc_hd__clkbuf_16
Xfanout471 _6694_/C VGND VGND VPWR VPWR _6445_/C sky130_fd_sc_hd__buf_4
XFILLER_93_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_23_csclk _7202_/CLK VGND VGND VPWR VPWR _7212_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_38_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7445_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_127_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold908 _7545_/Q VGND VGND VPWR VPWR hold908/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold919 _6019_/X VGND VGND VPWR VPWR _7593_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3470_ _3470_/A _3470_/B VGND VGND VPWR VPWR _7256_/D sky130_fd_sc_hd__xor2_1
XFILLER_170_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5140_ _5313_/C _5071_/B _5517_/A2 _4814_/A VGND VGND VPWR VPWR _5140_/X sky130_fd_sc_hd__a31o_1
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1608 _6977_/Q VGND VGND VPWR VPWR hold117/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5071_ _5429_/A _5071_/B _5071_/C VGND VGND VPWR VPWR _5074_/B sky130_fd_sc_hd__and3_1
Xhold1619 _7246_/Q VGND VGND VPWR VPWR _5439_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4022_ _7224_/Q _4541_/A hold98/A _3552_/X _7386_/Q VGND VGND VPWR VPWR _4022_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_49_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5973_ hold488/X _6045_/A1 _5974_/S VGND VGND VPWR VPWR _5973_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7712_ _7712_/A VGND VGND VPWR VPWR _7712_/X sky130_fd_sc_hd__clkbuf_2
X_4924_ _4924_/A _4924_/B _4924_/C VGND VGND VPWR VPWR _4927_/C sky130_fd_sc_hd__nand3_1
XFILLER_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7643_ _7657_/CLK _7643_/D fanout609/X VGND VGND VPWR VPWR _7643_/Q sky130_fd_sc_hd__dfrtp_1
X_4855_ _4966_/A _4957_/B _4923_/B VGND VGND VPWR VPWR _4961_/A sky130_fd_sc_hd__and3_1
XFILLER_178_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3806_ _7172_/Q _3700_/X _3715_/X _7109_/Q _3805_/X VGND VGND VPWR VPWR _3816_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_166_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7574_ _7606_/CLK _7574_/D fanout606/X VGND VGND VPWR VPWR _7574_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_159_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4786_ _4786_/A _4786_/B VGND VGND VPWR VPWR _4786_/Y sky130_fd_sc_hd__nand2_2
XFILLER_193_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6525_ _7339_/Q _6474_/A _6465_/X _7347_/Q _6524_/X VGND VGND VPWR VPWR _6532_/A
+ sky130_fd_sc_hd__a221o_1
X_3737_ _7470_/Q _3528_/X _3733_/X _3735_/X _3736_/X VGND VGND VPWR VPWR _3753_/A
+ sky130_fd_sc_hd__a2111o_1
X_6456_ _6791_/B _6791_/C _6791_/D VGND VGND VPWR VPWR _6456_/X sky130_fd_sc_hd__and3_4
X_3668_ _7567_/Q _5993_/A _5984_/B _3546_/X _7535_/Q VGND VGND VPWR VPWR _3668_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5407_ _5407_/A _5407_/B _5407_/C _5407_/D VGND VGND VPWR VPWR _5407_/Y sky130_fd_sc_hd__nor4_1
X_6387_ _7241_/Q _6158_/X _6382_/X _6383_/X _6386_/X VGND VGND VPWR VPWR _6387_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_88_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3599_ _7433_/Q _3556_/X _5741_/A _7353_/Q _3598_/X VGND VGND VPWR VPWR _3617_/A
+ sky130_fd_sc_hd__a221o_1
X_5338_ _4660_/C _5585_/A1 _5193_/Y _5015_/Y _4982_/Y VGND VGND VPWR VPWR _5463_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_87_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5269_ _4854_/X _5604_/B1 _4949_/Y _4945_/Y _4811_/Y VGND VGND VPWR VPWR _5273_/B
+ sky130_fd_sc_hd__o32a_1
X_7008_ _7616_/CLK _7008_/D fanout610/X VGND VGND VPWR VPWR _7691_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_56_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4640_ _4584_/Y _4639_/Y _4637_/A _5096_/A VGND VGND VPWR VPWR _5195_/B sky130_fd_sc_hd__a2bb2oi_4
XFILLER_190_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4571_ _4884_/A _5096_/A _5096_/B _5096_/C VGND VGND VPWR VPWR _4573_/B sky130_fd_sc_hd__nand4_4
XFILLER_162_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap402 _3551_/Y VGND VGND VPWR VPWR wire401/A sky130_fd_sc_hd__clkbuf_2
X_6310_ _7521_/Q _6131_/B _6115_/X _6151_/X _7553_/Q VGND VGND VPWR VPWR _6310_/X
+ sky130_fd_sc_hd__a32o_1
X_3522_ hold34/X hold61/X VGND VGND VPWR VPWR _5686_/B sky130_fd_sc_hd__nor2_4
Xhold705 hold705/A VGND VGND VPWR VPWR wb_dat_o[17] sky130_fd_sc_hd__buf_12
X_7290_ _7293_/CLK hold93/X fanout596/X VGND VGND VPWR VPWR hold92/A sky130_fd_sc_hd__dfrtp_1
Xhold716 hold716/A VGND VGND VPWR VPWR hold716/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold727 _7308_/Q VGND VGND VPWR VPWR hold727/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold738 _7037_/Q VGND VGND VPWR VPWR hold738/X sky130_fd_sc_hd__dlygate4sd3_1
X_6241_ _7374_/Q _6082_/B _6127_/X _6151_/X _7550_/Q VGND VGND VPWR VPWR _6241_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_116_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold749 _4244_/X VGND VGND VPWR VPWR _6988_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3453_ _7365_/Q VGND VGND VPWR VPWR _3453_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_131_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6172_ _7355_/Q _6138_/X _6152_/X _7363_/Q _6171_/X VGND VGND VPWR VPWR _6172_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5123_ _4998_/Y _5088_/Y _5108_/Y _5122_/Y VGND VGND VPWR VPWR _5123_/X sky130_fd_sc_hd__o211a_1
Xhold1405 _5683_/X VGND VGND VPWR VPWR hold122/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1416 _7671_/Q VGND VGND VPWR VPWR _6823_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1427 _7176_/Q VGND VGND VPWR VPWR hold1427/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1438 _4427_/X VGND VGND VPWR VPWR _7123_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5054_ _5195_/B _5476_/B _5322_/C _5092_/B VGND VGND VPWR VPWR _5055_/D sky130_fd_sc_hd__nand4_1
Xhold1449 _6737_/X VGND VGND VPWR VPWR _7659_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4005_ _4197_/A _4293_/S _3996_/X _3999_/X _4004_/X VGND VGND VPWR VPWR _4005_/Y
+ sky130_fd_sc_hd__a2111oi_2
XFILLER_72_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5956_ hold853/X _6028_/A1 _5956_/S VGND VGND VPWR VPWR _5956_/X sky130_fd_sc_hd__mux2_1
X_4907_ _4907_/A _4935_/C _4907_/C _4943_/A VGND VGND VPWR VPWR _4908_/B sky130_fd_sc_hd__nand4_1
X_5887_ hold172/X _6031_/A0 _5893_/S VGND VGND VPWR VPWR _5887_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4838_ _4836_/A _4865_/B _4837_/Y VGND VGND VPWR VPWR _4907_/A sky130_fd_sc_hd__o21ai_4
X_7626_ _4167_/A1 _7626_/D fanout620/X VGND VGND VPWR VPWR _7626_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7557_ _7557_/CLK _7557_/D fanout627/X VGND VGND VPWR VPWR _7557_/Q sky130_fd_sc_hd__dfrtp_4
X_4769_ _5407_/A _5189_/D _5429_/D VGND VGND VPWR VPWR _4769_/Y sky130_fd_sc_hd__nand3_4
XFILLER_107_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6508_ _7538_/Q _6479_/X _6493_/X _6507_/X VGND VGND VPWR VPWR _6508_/X sky130_fd_sc_hd__a211o_1
X_7488_ _7616_/CLK _7488_/D fanout610/X VGND VGND VPWR VPWR _7488_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6439_ _6438_/X _6439_/A1 _6812_/S VGND VGND VPWR VPWR _7649_/D sky130_fd_sc_hd__mux2_1
XFILLER_107_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold10 hold10/A VGND VGND VPWR VPWR hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A VGND VGND VPWR VPWR hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A VGND VGND VPWR VPWR hold32/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold43 hold43/A VGND VGND VPWR VPWR hold43/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A VGND VGND VPWR VPWR hold54/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold65 hold65/A VGND VGND VPWR VPWR hold65/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_188_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold76 hold76/A VGND VGND VPWR VPWR hold76/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold87 hold87/A VGND VGND VPWR VPWR hold87/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold98 hold98/A VGND VGND VPWR VPWR hold98/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_7 _5663_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5810_ hold881/X _6044_/A1 _5812_/S VGND VGND VPWR VPWR _5810_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6790_ _7173_/Q _6474_/A _6487_/X _7130_/Q _6789_/X VGND VGND VPWR VPWR _6800_/A
+ sky130_fd_sc_hd__a221o_1
X_5741_ _5741_/A _6029_/B VGND VGND VPWR VPWR _5749_/S sky130_fd_sc_hd__nand2_8
X_5672_ hold260/X _6866_/A1 _5677_/S VGND VGND VPWR VPWR _5672_/X sky130_fd_sc_hd__mux2_1
X_7411_ _7515_/CLK _7411_/D fanout623/X VGND VGND VPWR VPWR _7411_/Q sky130_fd_sc_hd__dfstp_2
X_4623_ _4822_/A _4959_/C VGND VGND VPWR VPWR _5189_/D sky130_fd_sc_hd__nor2_8
XFILLER_129_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7342_ _7518_/CLK _7342_/D fanout627/X VGND VGND VPWR VPWR _7342_/Q sky130_fd_sc_hd__dfrtp_1
X_4554_ _4554_/A0 _6012_/A0 _4558_/S VGND VGND VPWR VPWR _4554_/X sky130_fd_sc_hd__mux2_1
Xhold502 _4360_/X VGND VGND VPWR VPWR _7067_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 hold513/A VGND VGND VPWR VPWR hold513/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold524 _5712_/X VGND VGND VPWR VPWR _7320_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3505_ _3508_/S _3505_/B VGND VGND VPWR VPWR _3505_/Y sky130_fd_sc_hd__nand2_1
X_7273_ _7462_/CLK _7273_/D fanout604/X VGND VGND VPWR VPWR _7273_/Q sky130_fd_sc_hd__dfstp_1
Xhold535 _7201_/Q VGND VGND VPWR VPWR hold535/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 _5937_/X VGND VGND VPWR VPWR _7520_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4485_ hold723/X _5673_/A1 _4486_/S VGND VGND VPWR VPWR _4485_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold557 _7100_/Q VGND VGND VPWR VPWR hold557/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold568 _7065_/Q VGND VGND VPWR VPWR hold568/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold579 _7480_/Q VGND VGND VPWR VPWR hold579/X sky130_fd_sc_hd__dlygate4sd3_1
X_6224_ _6221_/X _6213_/B _6217_/X _6223_/X _6219_/X VGND VGND VPWR VPWR _6224_/X
+ sky130_fd_sc_hd__a2111o_1
X_3436_ _7501_/Q VGND VGND VPWR VPWR _3436_/Y sky130_fd_sc_hd__inv_2
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6155_ _7418_/Q _6150_/X _6151_/X _7546_/Q _6154_/X VGND VGND VPWR VPWR _6155_/X
+ sky130_fd_sc_hd__a221o_2
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1202 _6943_/Q VGND VGND VPWR VPWR _3904_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5106_ _4953_/C _5039_/Y _5064_/Y _4949_/Y _5104_/Y VGND VGND VPWR VPWR _5116_/A
+ sky130_fd_sc_hd__o221a_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1213 _4457_/A1 VGND VGND VPWR VPWR hold674/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1224 _4453_/A1 VGND VGND VPWR VPWR hold721/A sky130_fd_sc_hd__dlygate4sd3_1
X_6086_ _7139_/Q _6109_/B _6086_/C VGND VGND VPWR VPWR _6086_/Y sky130_fd_sc_hd__nor3_1
Xhold1235 _6820_/A1 VGND VGND VPWR VPWR hold833/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1246 _7096_/Q VGND VGND VPWR VPWR hold1246/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1257 _6862_/X VGND VGND VPWR VPWR _7682_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5037_ _5094_/A _5109_/A _5311_/C VGND VGND VPWR VPWR _5038_/B sky130_fd_sc_hd__and3_4
XFILLER_73_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1268 _7424_/Q VGND VGND VPWR VPWR hold78/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1279 _5801_/X VGND VGND VPWR VPWR _7399_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_408 _4769_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_419 _6131_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6988_ _7421_/CLK _6988_/D fanout630/X VGND VGND VPWR VPWR _7696_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5939_ _5984_/A _5939_/B _6038_/C VGND VGND VPWR VPWR _5947_/S sky130_fd_sc_hd__and3_4
XFILLER_21_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7609_ _7609_/CLK _7609_/D fanout614/X VGND VGND VPWR VPWR _7609_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput100 wb_adr_i[10] VGND VGND VPWR VPWR _4586_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput111 wb_adr_i[20] VGND VGND VPWR VPWR _5096_/A sky130_fd_sc_hd__buf_6
Xinput122 wb_adr_i[30] VGND VGND VPWR VPWR input122/X sky130_fd_sc_hd__clkbuf_1
Xinput133 wb_dat_i[10] VGND VGND VPWR VPWR _6836_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput144 wb_dat_i[20] VGND VGND VPWR VPWR _6842_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput155 wb_dat_i[30] VGND VGND VPWR VPWR _6848_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput166 wb_sel_i[1] VGND VGND VPWR VPWR _6857_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4270_ _4269_/X hold636/X _4274_/S VGND VGND VPWR VPWR _4270_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6911_ _6911_/A _6911_/B VGND VGND VPWR VPWR _6911_/X sky130_fd_sc_hd__and2_1
XFILLER_54_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6842_ _6969_/Q _6842_/A2 _6842_/B1 _6970_/Q VGND VGND VPWR VPWR _6842_/X sky130_fd_sc_hd__a22o_1
XFILLER_23_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6773_ _7044_/Q _6451_/X _6485_/X _7217_/Q _6772_/X VGND VGND VPWR VPWR _6773_/X
+ sky130_fd_sc_hd__a221o_1
X_3985_ _7081_/Q _4559_/B _5680_/A _3562_/X _7498_/Q VGND VGND VPWR VPWR _3985_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5724_ _5724_/A0 _6012_/A0 _5731_/S VGND VGND VPWR VPWR _5724_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5655_ _6866_/A1 hold273/X _5658_/S VGND VGND VPWR VPWR _5655_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4606_ _4706_/D _4836_/A _5014_/D VGND VGND VPWR VPWR _4760_/C sky130_fd_sc_hd__o21ai_4
X_5586_ _5586_/A _5586_/B _5586_/C _5586_/D VGND VGND VPWR VPWR _5618_/B sky130_fd_sc_hd__and4_1
XFILLER_117_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold310 _4300_/X VGND VGND VPWR VPWR _7016_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7325_ _7599_/CLK _7325_/D fanout629/X VGND VGND VPWR VPWR _7325_/Q sky130_fd_sc_hd__dfrtp_4
X_4537_ hold750/X _6863_/A1 _4540_/S VGND VGND VPWR VPWR _4537_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold321 _7356_/Q VGND VGND VPWR VPWR hold321/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 _6031_/X VGND VGND VPWR VPWR _7603_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold343 _7211_/Q VGND VGND VPWR VPWR hold343/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold354 _6022_/X VGND VGND VPWR VPWR _7595_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7256_ _4183_/A1 _7256_/D _6909_/X VGND VGND VPWR VPWR _7256_/Q sky130_fd_sc_hd__dfrtp_4
Xhold365 hold365/A VGND VGND VPWR VPWR hold365/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4468_ _4564_/A1 hold563/X _4468_/S VGND VGND VPWR VPWR _7163_/D sky130_fd_sc_hd__mux2_1
Xhold376 _4330_/X VGND VGND VPWR VPWR _7042_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold387 _7168_/Q VGND VGND VPWR VPWR hold387/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold398 _5631_/X VGND VGND VPWR VPWR _7253_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6207_ _6206_/X _6228_/A2 _6812_/S VGND VGND VPWR VPWR _7639_/D sky130_fd_sc_hd__mux2_1
X_3419_ _6939_/Q VGND VGND VPWR VPWR _3419_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7187_ _7255_/CLK _7187_/D fanout616/X VGND VGND VPWR VPWR _7187_/Q sky130_fd_sc_hd__dfrtp_2
X_4399_ hold557/X _4564_/A1 _4399_/S VGND VGND VPWR VPWR _4399_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6138_ _6158_/D _6151_/B _6392_/B _6231_/D VGND VGND VPWR VPWR _6138_/X sky130_fd_sc_hd__and4bb_4
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1010 _7091_/Q VGND VGND VPWR VPWR _4389_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1021 hold1262/X VGND VGND VPWR VPWR _5629_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1032 _7121_/Q VGND VGND VPWR VPWR _4425_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_133_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1043 _4329_/X VGND VGND VPWR VPWR _7041_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1054 _7164_/Q VGND VGND VPWR VPWR _4470_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_6069_ _7624_/Q _7623_/Q VGND VGND VPWR VPWR _6161_/D sky130_fd_sc_hd__nor2_8
Xhold1065 _5925_/X VGND VGND VPWR VPWR _7509_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1076 _4308_/X VGND VGND VPWR VPWR _7023_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1087 _5790_/X VGND VGND VPWR VPWR _7389_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1098 hold1573/X VGND VGND VPWR VPWR _4355_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_205 _7446_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_216 _7083_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_227 _7381_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_238 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_249 input21/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3770_ _7183_/Q _4535_/B _4487_/B _4358_/A _7070_/Q VGND VGND VPWR VPWR _3770_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_158_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5440_ _5452_/A _5452_/B VGND VGND VPWR VPWR _5440_/Y sky130_fd_sc_hd__nand2_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5371_ _5367_/X _5371_/B _5552_/B VGND VGND VPWR VPWR _5371_/Y sky130_fd_sc_hd__nand3b_1
X_7110_ _7130_/CLK _7110_/D fanout602/X VGND VGND VPWR VPWR _7110_/Q sky130_fd_sc_hd__dfrtp_1
X_4322_ _5678_/C _4505_/B _5680_/C VGND VGND VPWR VPWR _4327_/S sky130_fd_sc_hd__and3_2
XFILLER_126_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7041_ _7194_/CLK _7041_/D fanout602/X VGND VGND VPWR VPWR _7041_/Q sky130_fd_sc_hd__dfrtp_1
X_4253_ hold845/X hold85/X _4257_/S VGND VGND VPWR VPWR _4253_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4184_ _6951_/Q _6911_/A VGND VGND VPWR VPWR _4184_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_3_4__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _7676_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_95_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6825_ _6825_/A _6827_/A VGND VGND VPWR VPWR _6825_/Y sky130_fd_sc_hd__nand2_1
XFILLER_23_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3968_ _4038_/B1 _3967_/X _3968_/S VGND VGND VPWR VPWR _3968_/X sky130_fd_sc_hd__mux2_1
X_6756_ _7231_/Q _6720_/C _6536_/C _6755_/X VGND VGND VPWR VPWR _6756_/X sky130_fd_sc_hd__a31o_1
XFILLER_149_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5707_ _6031_/A0 hold141/X hold38/X VGND VGND VPWR VPWR _5707_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6687_ _6686_/X _6687_/A1 _6812_/S VGND VGND VPWR VPWR _7657_/D sky130_fd_sc_hd__mux2_1
XFILLER_164_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3899_ _7420_/Q _3602_/X _3895_/X _3898_/X VGND VGND VPWR VPWR _3899_/X sky130_fd_sc_hd__a211o_1
XFILLER_148_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5638_ _5638_/A0 _5697_/A0 _5642_/S VGND VGND VPWR VPWR _7261_/D sky130_fd_sc_hd__mux2_1
XFILLER_164_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5569_ _5569_/A1 wire535/X _5501_/Y _5568_/X _5558_/Y VGND VGND VPWR VPWR _7248_/D
+ sky130_fd_sc_hd__a221o_1
Xhold140 _4307_/X VGND VGND VPWR VPWR _7022_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_163_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7308_ _7512_/CLK _7308_/D fanout608/X VGND VGND VPWR VPWR _7308_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold151 _7296_/Q VGND VGND VPWR VPWR hold151/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold162 _7614_/Q VGND VGND VPWR VPWR hold162/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 _5887_/X VGND VGND VPWR VPWR _7475_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold184 _7075_/Q VGND VGND VPWR VPWR hold184/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 _7208_/Q VGND VGND VPWR VPWR hold195/X sky130_fd_sc_hd__dlygate4sd3_1
X_7239_ _7682_/CLK _7239_/D fanout603/X VGND VGND VPWR VPWR _7239_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout620 fanout633/X VGND VGND VPWR VPWR fanout620/X sky130_fd_sc_hd__buf_6
Xfanout631 fanout632/X VGND VGND VPWR VPWR fanout631/X sky130_fd_sc_hd__clkbuf_8
Xfanout642 _4992_/C VGND VGND VPWR VPWR _4822_/A sky130_fd_sc_hd__buf_12
XFILLER_92_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4940_ _4946_/A _4957_/B _5452_/A _5389_/C VGND VGND VPWR VPWR _4941_/A sky130_fd_sc_hd__and4_1
X_4871_ _4865_/B _4865_/C _4859_/Y _4860_/B VGND VGND VPWR VPWR _4871_/X sky130_fd_sc_hd__a211o_4
XANTENNA_580 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_591 _4116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6610_ _6610_/A1 _6109_/X _6609_/X _6686_/S VGND VGND VPWR VPWR _6610_/X sky130_fd_sc_hd__o22a_1
X_3822_ _7177_/Q _4481_/A hold98/A _4293_/S _4171_/D VGND VGND VPWR VPWR _3822_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_177_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7590_ _7590_/CLK _7590_/D fanout612/X VGND VGND VPWR VPWR _7590_/Q sky130_fd_sc_hd__dfrtp_1
X_6541_ _7324_/Q _6471_/X _6501_/X _7564_/Q _6536_/X VGND VGND VPWR VPWR _6541_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_193_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3753_ _3753_/A _3753_/B _3753_/C _3753_/D VGND VGND VPWR VPWR _3775_/A sky130_fd_sc_hd__nor4_2
XFILLER_146_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6472_ _6099_/B _6771_/C _6452_/X _6469_/X _6471_/X VGND VGND VPWR VPWR _6478_/C
+ sky130_fd_sc_hd__a2111oi_4
X_3684_ _7599_/Q _3569_/X _5689_/A _7715_/A _3682_/X VGND VGND VPWR VPWR _3684_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_145_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5423_ _5452_/B _5040_/C _5095_/C _5291_/C VGND VGND VPWR VPWR _5423_/X sky130_fd_sc_hd__o211a_1
XFILLER_145_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput201 _3426_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[33] sky130_fd_sc_hd__buf_12
Xoutput212 _3450_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[9] sky130_fd_sc_hd__buf_12
XFILLER_145_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput223 _7700_/X VGND VGND VPWR VPWR mgmt_gpio_out[20] sky130_fd_sc_hd__buf_12
XFILLER_161_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput234 _7710_/X VGND VGND VPWR VPWR mgmt_gpio_out[30] sky130_fd_sc_hd__buf_12
X_5354_ _5236_/Y _5352_/X _5353_/X _5544_/C VGND VGND VPWR VPWR _5354_/X sky130_fd_sc_hd__o31a_1
XFILLER_160_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput245 _4157_/X VGND VGND VPWR VPWR mgmt_gpio_out[6] sky130_fd_sc_hd__buf_12
XFILLER_114_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput256 _4188_/Y VGND VGND VPWR VPWR pad_flash_io1_oeb sky130_fd_sc_hd__buf_12
Xoutput267 _7259_/Q VGND VGND VPWR VPWR pll_ena sky130_fd_sc_hd__buf_12
XFILLER_99_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4305_ _6003_/A1 hold405/X _4311_/S VGND VGND VPWR VPWR _4305_/X sky130_fd_sc_hd__mux2_1
Xoutput278 _7272_/Q VGND VGND VPWR VPWR pll_trim[16] sky130_fd_sc_hd__buf_12
Xoutput289 _6974_/Q VGND VGND VPWR VPWR pll_trim[2] sky130_fd_sc_hd__buf_12
X_5285_ _5407_/A _5429_/D _5407_/B _4825_/Y VGND VGND VPWR VPWR _5285_/X sky130_fd_sc_hd__o31a_4
X_7024_ _7583_/CLK _7024_/D fanout630/X VGND VGND VPWR VPWR _7024_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4236_ _4459_/A0 _4236_/A1 _4239_/S VGND VGND VPWR VPWR _6984_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4167_ _7002_/Q _4167_/A1 _7295_/Q VGND VGND VPWR VPWR _4167_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4098_ _7258_/Q _7256_/Q _4104_/D _7257_/Q VGND VGND VPWR VPWR _4099_/S sky130_fd_sc_hd__and4bb_1
XFILLER_82_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_4_csclk _7236_/CLK VGND VGND VPWR VPWR _7130_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6808_ _7100_/Q _6444_/X _6805_/X _6807_/X VGND VGND VPWR VPWR _6809_/C sky130_fd_sc_hd__a211o_1
XFILLER_23_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6739_ _7161_/Q _6456_/X _6457_/X _7196_/Q VGND VGND VPWR VPWR _6739_/X sky130_fd_sc_hd__a22o_1
XFILLER_149_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout461 _6076_/X VGND VGND VPWR VPWR _6427_/A3 sky130_fd_sc_hd__buf_12
XFILLER_171_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout472 _6442_/Y VGND VGND VPWR VPWR _6694_/C sky130_fd_sc_hd__buf_8
XFILLER_59_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold909 _5965_/X VGND VGND VPWR VPWR _7545_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5070_ _5375_/A _5476_/A _5233_/C _5069_/X VGND VGND VPWR VPWR _5073_/B sky130_fd_sc_hd__a31o_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1609 _6975_/Q VGND VGND VPWR VPWR hold455/A sky130_fd_sc_hd__dlygate4sd3_1
X_4021_ _7538_/Q _5993_/A _5957_/B _4016_/X _4020_/X VGND VGND VPWR VPWR _4036_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_96_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5972_ hold947/X _5999_/A1 _5974_/S VGND VGND VPWR VPWR _5972_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7711_ _7711_/A VGND VGND VPWR VPWR _7711_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4923_ _4943_/A _4923_/B _5452_/A _4934_/C VGND VGND VPWR VPWR _4924_/C sky130_fd_sc_hd__nand4_1
XFILLER_80_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7642_ _7657_/CLK _7642_/D fanout607/X VGND VGND VPWR VPWR _7642_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_100_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4854_ _4865_/B _4865_/C _4907_/C _4860_/B _4935_/B VGND VGND VPWR VPWR _4854_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_138_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3805_ _7237_/Q _5628_/A _4553_/B _3713_/X _7099_/Q VGND VGND VPWR VPWR _3805_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_178_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7573_ _7613_/CLK _7573_/D fanout626/X VGND VGND VPWR VPWR _7573_/Q sky130_fd_sc_hd__dfrtp_4
X_4785_ _4785_/A _4794_/D _4785_/C _5231_/B VGND VGND VPWR VPWR _4785_/Y sky130_fd_sc_hd__nand4_4
X_3736_ _7115_/Q _5903_/A _4529_/B _3583_/X input56/X VGND VGND VPWR VPWR _3736_/X
+ sky130_fd_sc_hd__a32o_1
X_6524_ _7443_/Q _6460_/X _6482_/X _7483_/Q VGND VGND VPWR VPWR _6524_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3667_ _3667_/A _3667_/B _3667_/C _3667_/D VGND VGND VPWR VPWR _3667_/Y sky130_fd_sc_hd__nor4_1
X_6455_ _7354_/Q _6791_/C _6455_/C _6771_/C VGND VGND VPWR VPWR _6455_/X sky130_fd_sc_hd__and4_1
X_5406_ _4961_/A _5452_/B _5404_/X _5572_/B _5403_/Y VGND VGND VPWR VPWR _5406_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_161_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6386_ _7123_/Q _6133_/X _6146_/X _7083_/Q _6385_/X VGND VGND VPWR VPWR _6386_/X
+ sky130_fd_sc_hd__a221o_1
X_3598_ _6979_/Q _3573_/C _4505_/B _3525_/X _7401_/Q VGND VGND VPWR VPWR _3598_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_133_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5337_ _5011_/B _4976_/Y _4982_/Y _5009_/Y _5206_/B VGND VGND VPWR VPWR _5534_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5268_ _5268_/A _5268_/B _5575_/D VGND VGND VPWR VPWR _5273_/A sky130_fd_sc_hd__nor3b_1
XFILLER_125_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7007_ _7616_/CLK _7007_/D fanout610/X VGND VGND VPWR VPWR _7690_/A sky130_fd_sc_hd__dfrtp_1
X_4219_ hold79/X _6838_/A0 _4229_/S VGND VGND VPWR VPWR hold80/A sky130_fd_sc_hd__mux2_4
XFILLER_102_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5199_ _4816_/Y _5611_/A2 _5015_/Y _5193_/Y _5196_/Y VGND VGND VPWR VPWR _5463_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_28_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4570_ _5429_/D _4948_/B _4959_/C _4948_/A VGND VGND VPWR VPWR _4570_/Y sky130_fd_sc_hd__nand4_4
X_3521_ _3622_/A _4340_/A hold23/X VGND VGND VPWR VPWR _5723_/A sky130_fd_sc_hd__and3_4
Xhold706 hold706/A VGND VGND VPWR VPWR hold706/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold717 hold717/A VGND VGND VPWR VPWR hold717/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold728 _5699_/X VGND VGND VPWR VPWR _7308_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap436 _7341_/Q VGND VGND VPWR VPWR _4171_/C sky130_fd_sc_hd__buf_12
X_6240_ _7518_/Q _6131_/B _6115_/X _6159_/X _7438_/Q VGND VGND VPWR VPWR _6240_/X
+ sky130_fd_sc_hd__a32o_1
Xmax_cap447 _6466_/X VGND VGND VPWR VPWR _6807_/A2 sky130_fd_sc_hd__buf_6
Xhold739 _4324_/X VGND VGND VPWR VPWR _7037_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3452_ _7373_/Q VGND VGND VPWR VPWR _3452_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6171_ _7523_/Q _6131_/B _6334_/C _6145_/X _7459_/Q VGND VGND VPWR VPWR _6171_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_69_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5122_ _4948_/B _5090_/B _5034_/C _5121_/Y VGND VGND VPWR VPWR _5122_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1406 _7349_/Q VGND VGND VPWR VPWR hold1406/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1417 _7602_/Q VGND VGND VPWR VPWR hold503/A sky130_fd_sc_hd__dlygate4sd3_1
X_5053_ _5109_/A _5311_/A _5131_/B _5311_/C VGND VGND VPWR VPWR _5055_/C sky130_fd_sc_hd__nand4_1
Xhold1428 _4484_/X VGND VGND VPWR VPWR _7176_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1439 _7346_/Q VGND VGND VPWR VPWR hold417/A sky130_fd_sc_hd__dlygate4sd3_1
X_4004_ _7219_/Q _4547_/A _4535_/B _4001_/X _4003_/X VGND VGND VPWR VPWR _4004_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_37_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5955_ hold469/X _6045_/A1 _5956_/S VGND VGND VPWR VPWR _5955_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4906_ _4906_/A _4906_/B _4906_/C _4906_/D VGND VGND VPWR VPWR _4908_/A sky130_fd_sc_hd__nor4_1
X_5886_ hold280/X _6039_/A1 _5893_/S VGND VGND VPWR VPWR _7474_/D sky130_fd_sc_hd__mux2_1
XFILLER_139_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7625_ _4167_/A1 _7625_/D fanout620/X VGND VGND VPWR VPWR _7625_/Q sky130_fd_sc_hd__dfrtp_1
X_4837_ _4599_/Y _4777_/Y _4990_/A VGND VGND VPWR VPWR _4837_/Y sky130_fd_sc_hd__o21bai_2
XFILLER_138_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7556_ _7603_/CLK _7556_/D fanout611/X VGND VGND VPWR VPWR _7556_/Q sky130_fd_sc_hd__dfrtp_1
X_4768_ _5407_/A _5189_/D _5429_/D VGND VGND VPWR VPWR _5181_/C sky130_fd_sc_hd__and3_4
XFILLER_146_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6507_ _7346_/Q _6465_/X _6809_/D _6497_/X _6506_/X VGND VGND VPWR VPWR _6507_/X
+ sky130_fd_sc_hd__a2111o_2
X_3719_ _7255_/Q _5628_/A _4505_/B _5849_/A _7446_/Q VGND VGND VPWR VPWR _3719_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_147_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7487_ _7512_/CLK _7487_/D fanout608/X VGND VGND VPWR VPWR _7487_/Q sky130_fd_sc_hd__dfrtp_4
X_4699_ _5407_/A _4704_/A VGND VGND VPWR VPWR _5429_/A sky130_fd_sc_hd__nor2_8
XFILLER_134_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6438_ _6438_/A1 _6109_/X _6437_/X _6811_/S VGND VGND VPWR VPWR _6438_/X sky130_fd_sc_hd__o22a_1
XFILLER_136_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6369_ _7181_/Q wire455/A _6141_/X _7201_/Q _6368_/X VGND VGND VPWR VPWR _6369_/X
+ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_22_csclk _7202_/CLK VGND VGND VPWR VPWR _7398_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_102_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold11 hold11/A VGND VGND VPWR VPWR hold11/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold22 hold22/A VGND VGND VPWR VPWR hold22/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 hold33/A VGND VGND VPWR VPWR hold33/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold44 hold44/A VGND VGND VPWR VPWR hold44/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A VGND VGND VPWR VPWR hold55/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold66 hold66/A VGND VGND VPWR VPWR hold66/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold77 hold77/A VGND VGND VPWR VPWR hold77/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 hold88/A VGND VGND VPWR VPWR hold88/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold99 hold99/A VGND VGND VPWR VPWR hold99/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_37_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7421_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_56_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_mgmt_gpio_in[4] mgmt_gpio_in[4] VGND VGND VPWR VPWR clkbuf_0_mgmt_gpio_in[4]/X
+ sky130_fd_sc_hd__clkbuf_16
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_8 _5734_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5740_ hold900/X _6046_/A1 _5740_/S VGND VGND VPWR VPWR _5740_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5671_ _5678_/C _5678_/B _5680_/C VGND VGND VPWR VPWR _5677_/S sky130_fd_sc_hd__and3_2
XFILLER_30_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7410_ _7586_/CLK _7410_/D fanout625/X VGND VGND VPWR VPWR _7410_/Q sky130_fd_sc_hd__dfstp_1
X_4622_ _4822_/A _5074_/A _5189_/A VGND VGND VPWR VPWR _4622_/Y sky130_fd_sc_hd__nand3b_1
X_4553_ _5628_/A _4553_/B _6861_/C VGND VGND VPWR VPWR _4558_/S sky130_fd_sc_hd__and3_2
X_7341_ _7445_/CLK _7341_/D fanout628/X VGND VGND VPWR VPWR _7341_/Q sky130_fd_sc_hd__dfrtp_4
Xhold503 hold503/A VGND VGND VPWR VPWR hold503/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold514 _7138_/Q VGND VGND VPWR VPWR hold514/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3504_ _4229_/S hold95/X hold119/X hold69/X VGND VGND VPWR VPWR _3713_/A sky130_fd_sc_hd__o211a_4
Xhold525 _7053_/Q VGND VGND VPWR VPWR hold525/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7272_ _7286_/CLK _7272_/D fanout598/X VGND VGND VPWR VPWR _7272_/Q sky130_fd_sc_hd__dfstp_1
X_4484_ _4484_/A0 _4556_/A1 _4486_/S VGND VGND VPWR VPWR _4484_/X sky130_fd_sc_hd__mux2_1
Xhold536 _4514_/X VGND VGND VPWR VPWR _7201_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 _7700_/A VGND VGND VPWR VPWR hold547/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold558 _4399_/X VGND VGND VPWR VPWR _7100_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3435_ _7509_/Q VGND VGND VPWR VPWR _3435_/Y sky130_fd_sc_hd__inv_2
Xhold569 _4357_/X VGND VGND VPWR VPWR _7065_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6223_ _7549_/Q _6151_/X _6159_/X _7437_/Q _6222_/X VGND VGND VPWR VPWR _6223_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6154_ _7362_/Q _6159_/B _6141_/X _6153_/X _7562_/Q VGND VGND VPWR VPWR _6154_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1203 _4238_/A1 VGND VGND VPWR VPWR hold594/A sky130_fd_sc_hd__dlygate4sd3_1
X_5105_ _4953_/C _5039_/Y _5064_/Y _4949_/Y VGND VGND VPWR VPWR _5105_/Y sky130_fd_sc_hd__o22ai_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1214 _4458_/A1 VGND VGND VPWR VPWR hold684/A sky130_fd_sc_hd__dlygate4sd3_1
X_6085_ _6159_/B _6084_/X _6083_/X VGND VGND VPWR VPWR _7627_/D sky130_fd_sc_hd__o21ai_1
Xhold1225 _6822_/A1 VGND VGND VPWR VPWR hold632/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1236 _7027_/Q VGND VGND VPWR VPWR _4312_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1247 _4395_/X VGND VGND VPWR VPWR _7096_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5036_ _5061_/A _5042_/A _5092_/B VGND VGND VPWR VPWR _5036_/X sky130_fd_sc_hd__and3_1
Xhold1258 _7526_/Q VGND VGND VPWR VPWR hold421/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1269 _5829_/X VGND VGND VPWR VPWR _7424_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_409 _5401_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6987_ _7672_/CLK _6987_/D VGND VGND VPWR VPWR _6987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5938_ hold885/X _6028_/A1 _5938_/S VGND VGND VPWR VPWR _5938_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5869_ hold203/X _5869_/A1 _5875_/S VGND VGND VPWR VPWR _5869_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7608_ _7608_/CLK _7608_/D fanout611/X VGND VGND VPWR VPWR _7608_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_181_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7539_ _7541_/CLK _7539_/D fanout609/X VGND VGND VPWR VPWR _7539_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_119_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput101 wb_adr_i[11] VGND VGND VPWR VPWR _4586_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput112 wb_adr_i[21] VGND VGND VPWR VPWR _4884_/A sky130_fd_sc_hd__buf_8
XFILLER_103_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput123 wb_adr_i[31] VGND VGND VPWR VPWR input123/X sky130_fd_sc_hd__clkbuf_1
Xinput134 wb_dat_i[11] VGND VGND VPWR VPWR _6839_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput145 wb_dat_i[21] VGND VGND VPWR VPWR _6845_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput156 wb_dat_i[31] VGND VGND VPWR VPWR _6851_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput167 wb_sel_i[2] VGND VGND VPWR VPWR _6825_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_29_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__1128_ clkbuf_0__1128_/X VGND VGND VPWR VPWR _6820_/A0 sky130_fd_sc_hd__clkbuf_16
XFILLER_153_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_3__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _7662_/CLK sky130_fd_sc_hd__clkbuf_16
X_7634__648 VGND VGND VPWR VPWR _7634_/D _7634__648/LO sky130_fd_sc_hd__conb_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6910_ _6911_/A _6911_/B VGND VGND VPWR VPWR _6910_/X sky130_fd_sc_hd__and2_1
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6841_ _6841_/A0 _6840_/X _6853_/S VGND VGND VPWR VPWR _7675_/D sky130_fd_sc_hd__mux2_1
XFILLER_90_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6772_ _7182_/Q _6465_/X _6483_/X _7069_/Q VGND VGND VPWR VPWR _6772_/X sky130_fd_sc_hd__a22o_1
X_3984_ _7506_/Q _6861_/A _5993_/B _3972_/X _3983_/X VGND VGND VPWR VPWR _3995_/C
+ sky130_fd_sc_hd__a311o_1
XFILLER_167_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5723_ _5723_/A _5759_/B _6029_/B VGND VGND VPWR VPWR _5731_/S sky130_fd_sc_hd__and3_4
XFILLER_148_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5654_ _5673_/A1 hold500/X _5658_/S VGND VGND VPWR VPWR _5654_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4605_ _4706_/D _4836_/A _4604_/Y VGND VGND VPWR VPWR _4760_/D sky130_fd_sc_hd__o21ai_4
XFILLER_117_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5585_ _5585_/A1 _4993_/Y _5018_/Y _5047_/C _5340_/X VGND VGND VPWR VPWR _5586_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_163_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold300 _5947_/X VGND VGND VPWR VPWR _7529_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold311 _7444_/Q VGND VGND VPWR VPWR hold311/X sky130_fd_sc_hd__dlygate4sd3_1
X_7324_ _7430_/CLK _7324_/D fanout627/X VGND VGND VPWR VPWR _7324_/Q sky130_fd_sc_hd__dfrtp_4
X_4536_ _4536_/A0 _5697_/A0 _4540_/S VGND VGND VPWR VPWR _7219_/D sky130_fd_sc_hd__mux2_1
Xhold322 _5753_/X VGND VGND VPWR VPWR _7356_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 _7083_/Q VGND VGND VPWR VPWR hold333/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold344 _4526_/X VGND VGND VPWR VPWR _7211_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 _7372_/Q VGND VGND VPWR VPWR hold355/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 _7030_/Q VGND VGND VPWR VPWR hold366/X sky130_fd_sc_hd__dlygate4sd3_1
X_7255_ _7255_/CLK _7255_/D fanout618/X VGND VGND VPWR VPWR _7255_/Q sky130_fd_sc_hd__dfrtp_2
X_4467_ _5673_/A1 hold725/X _4468_/S VGND VGND VPWR VPWR _7162_/D sky130_fd_sc_hd__mux2_1
Xhold377 _7043_/Q VGND VGND VPWR VPWR hold377/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold388 _4474_/X VGND VGND VPWR VPWR _7168_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold399 hold399/A VGND VGND VPWR VPWR hold399/X sky130_fd_sc_hd__dlygate4sd3_1
X_6206_ _6206_/A1 _6109_/X _6205_/X _6686_/S VGND VGND VPWR VPWR _6206_/X sky130_fd_sc_hd__o22a_1
XFILLER_132_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7186_ _7231_/CLK _7186_/D fanout600/X VGND VGND VPWR VPWR _7186_/Q sky130_fd_sc_hd__dfstp_1
X_4398_ _4398_/A0 _6865_/A1 _4399_/S VGND VGND VPWR VPWR _4398_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1000 _4272_/X VGND VGND VPWR VPWR _7001_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6137_ _7624_/Q _6151_/B _6392_/B _7623_/Q VGND VGND VPWR VPWR _6137_/X sky130_fd_sc_hd__and4bb_4
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1011 _4389_/X VGND VGND VPWR VPWR _7091_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1022 hold1444/X VGND VGND VPWR VPWR _4409_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1033 _4425_/X VGND VGND VPWR VPWR _7121_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1044 _7086_/Q VGND VGND VPWR VPWR _4383_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6068_ _7623_/Q _7624_/Q VGND VGND VPWR VPWR _6166_/B sky130_fd_sc_hd__and2b_4
XFILLER_73_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1055 _4470_/X VGND VGND VPWR VPWR _7164_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1066 hold1374/X VGND VGND VPWR VPWR _6042_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1077 hold1284/X VGND VGND VPWR VPWR _5970_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5019_ _4992_/C _4992_/D _5189_/A _4992_/B _5015_/Y VGND VGND VPWR VPWR _5019_/X
+ sky130_fd_sc_hd__a2111o_1
Xhold1088 hold1361/X VGND VGND VPWR VPWR _5916_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1099 _7303_/Q VGND VGND VPWR VPWR _5693_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_206 _7252_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_217 _7082_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_228 _7382_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_239 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_740 _6809_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5370_ _4763_/X _5153_/C _5369_/X VGND VGND VPWR VPWR _5552_/B sky130_fd_sc_hd__a21oi_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4321_ hold571/X _6028_/A1 _4321_/S VGND VGND VPWR VPWR _4321_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4252_ hold547/X _4251_/X _4258_/S VGND VGND VPWR VPWR _4252_/X sky130_fd_sc_hd__mux2_1
X_7040_ _7291_/CLK _7040_/D fanout596/X VGND VGND VPWR VPWR _7040_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_101_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4183_ input83/X _4183_/A1 _6951_/Q VGND VGND VPWR VPWR _4183_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6824_ _6827_/A _6857_/A2 _6970_/Q VGND VGND VPWR VPWR _6829_/C sky130_fd_sc_hd__a21bo_1
XFILLER_23_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6755_ _7186_/Q _6452_/X _6464_/X _7684_/Q _6754_/X VGND VGND VPWR VPWR _6755_/X
+ sky130_fd_sc_hd__a221o_1
X_3967_ _3966_/X _6943_/Q _3967_/S VGND VGND VPWR VPWR _3967_/X sky130_fd_sc_hd__mux2_1
X_5706_ _6039_/A1 hold277/X hold38/X VGND VGND VPWR VPWR _7314_/D sky130_fd_sc_hd__mux2_1
X_6686_ _6685_/X _6686_/A1 _6686_/S VGND VGND VPWR VPWR _6686_/X sky130_fd_sc_hd__mux2_1
X_3898_ _7356_/Q hold24/A _4511_/C _3897_/X VGND VGND VPWR VPWR _3898_/X sky130_fd_sc_hd__a31o_1
XFILLER_164_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5637_ _5939_/B _5678_/C _5680_/C VGND VGND VPWR VPWR _5642_/S sky130_fd_sc_hd__and3_2
XFILLER_136_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5568_ _5297_/A _5322_/A _5071_/C _5567_/Y VGND VGND VPWR VPWR _5568_/X sky130_fd_sc_hd__a31o_1
XFILLER_151_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold130 _4493_/Y VGND VGND VPWR VPWR _4498_/S sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7307_ _7307_/CLK _7307_/D _6911_/A VGND VGND VPWR VPWR _7307_/Q sky130_fd_sc_hd__dfrtp_1
Xhold141 _7315_/Q VGND VGND VPWR VPWR hold141/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4519_ hold440/X _5869_/A1 _4522_/S VGND VGND VPWR VPWR _4519_/X sky130_fd_sc_hd__mux2_1
Xhold152 _5684_/X VGND VGND VPWR VPWR _7296_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 _6043_/X VGND VGND VPWR VPWR _7614_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5499_ _5478_/X _5544_/C _5498_/X VGND VGND VPWR VPWR _5499_/Y sky130_fd_sc_hd__a21oi_2
Xhold174 _7502_/Q VGND VGND VPWR VPWR hold174/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 _4369_/X VGND VGND VPWR VPWR _7075_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7238_ _7238_/CLK _7238_/D fanout603/X VGND VGND VPWR VPWR _7238_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_132_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout610 fanout611/X VGND VGND VPWR VPWR fanout610/X sky130_fd_sc_hd__buf_8
Xhold196 _4522_/X VGND VGND VPWR VPWR _7208_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout621 fanout632/X VGND VGND VPWR VPWR fanout621/X sky130_fd_sc_hd__buf_8
XFILLER_132_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout632 fanout633/X VGND VGND VPWR VPWR fanout632/X sky130_fd_sc_hd__buf_8
Xfanout643 _4992_/D VGND VGND VPWR VPWR _4959_/C sky130_fd_sc_hd__buf_12
XFILLER_86_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7169_ _7242_/CLK _7169_/D fanout616/X VGND VGND VPWR VPWR _7169_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_37_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4870_ _4946_/A _5452_/A _5389_/B _4957_/C VGND VGND VPWR VPWR _4904_/D sky130_fd_sc_hd__nand4_1
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_570 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_581 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_592 _4116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3821_ _7275_/Q _3573_/C _5680_/A _3817_/X _3820_/X VGND VGND VPWR VPWR _3821_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_20_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6540_ _7604_/Q _6456_/X _6468_/X _7588_/Q _6539_/X VGND VGND VPWR VPWR _6540_/X
+ sky130_fd_sc_hd__a221o_1
X_3752_ input7/X _3573_/X _3749_/X _3750_/X _3751_/X VGND VGND VPWR VPWR _3753_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_192_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6471_ _6645_/B _6771_/C _6645_/C VGND VGND VPWR VPWR _6471_/X sky130_fd_sc_hd__and3_4
X_3683_ _5682_/A _5659_/C _4481_/A VGND VGND VPWR VPWR _5689_/A sky130_fd_sc_hd__and3_4
X_5422_ _4823_/Y _5103_/X _5009_/Y _5611_/A2 VGND VGND VPWR VPWR _5560_/C sky130_fd_sc_hd__a211o_1
XFILLER_146_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput202 _3425_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[34] sky130_fd_sc_hd__buf_12
Xoutput213 _4161_/X VGND VGND VPWR VPWR mgmt_gpio_out[0] sky130_fd_sc_hd__buf_12
XFILLER_161_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput224 _7701_/X VGND VGND VPWR VPWR mgmt_gpio_out[21] sky130_fd_sc_hd__buf_12
Xoutput235 _7711_/X VGND VGND VPWR VPWR mgmt_gpio_out[31] sky130_fd_sc_hd__buf_12
X_5353_ _4946_/A _5401_/A _5512_/B _5322_/A VGND VGND VPWR VPWR _5353_/X sky130_fd_sc_hd__o211a_1
Xoutput246 _7693_/X VGND VGND VPWR VPWR mgmt_gpio_out[7] sky130_fd_sc_hd__buf_12
Xoutput257 _7269_/Q VGND VGND VPWR VPWR pll90_sel[0] sky130_fd_sc_hd__buf_12
Xoutput268 _7266_/Q VGND VGND VPWR VPWR pll_sel[0] sky130_fd_sc_hd__buf_12
X_4304_ _7294_/Q _4171_/C _4171_/D _4257_/S _6029_/B VGND VGND VPWR VPWR _4304_/Y
+ sky130_fd_sc_hd__o311ai_4
Xoutput279 _7273_/Q VGND VGND VPWR VPWR pll_trim[17] sky130_fd_sc_hd__buf_12
X_5284_ _5011_/C _5604_/B1 _4987_/Y _5127_/C VGND VGND VPWR VPWR _5310_/A sky130_fd_sc_hd__o31a_1
XFILLER_4_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7023_ _7421_/CLK _7023_/D fanout630/X VGND VGND VPWR VPWR _7023_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4235_ _3838_/Y _4235_/A1 _4239_/S VGND VGND VPWR VPWR _6983_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4166_ _7003_/Q user_clock _7296_/Q VGND VGND VPWR VPWR _4166_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4097_ _4097_/A0 input58/X _4097_/S VGND VGND VPWR VPWR _6919_/D sky130_fd_sc_hd__mux2_1
XFILLER_82_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6807_ _7238_/Q _6807_/A2 _6471_/X _7050_/Q _6806_/X VGND VGND VPWR VPWR _6807_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_23_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4999_ _5614_/A _4999_/B _5311_/A VGND VGND VPWR VPWR _5056_/A sky130_fd_sc_hd__and3_1
XFILLER_23_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6738_ _7043_/Q _6451_/X _6468_/X _7176_/Q VGND VGND VPWR VPWR _6738_/X sky130_fd_sc_hd__a22o_1
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6669_ _7457_/Q _6459_/X _6482_/X _7489_/Q _6668_/X VGND VGND VPWR VPWR _6675_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_109_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout473 _6562_/B VGND VGND VPWR VPWR _6791_/D sky130_fd_sc_hd__buf_12
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4020_ _7298_/Q _5682_/C _5984_/B _4017_/X _4019_/X VGND VGND VPWR VPWR _4020_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_96_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5971_ hold176/X _6043_/A1 _5974_/S VGND VGND VPWR VPWR _5971_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7710_ _7710_/A VGND VGND VPWR VPWR _7710_/X sky130_fd_sc_hd__clkbuf_1
X_4922_ _5181_/C _4923_/B _5452_/A _4934_/C VGND VGND VPWR VPWR _4924_/B sky130_fd_sc_hd__nand4_1
X_7641_ _7657_/CLK _7641_/D fanout609/X VGND VGND VPWR VPWR _7641_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4853_ _4923_/B _4907_/A _4853_/C VGND VGND VPWR VPWR _4946_/B sky130_fd_sc_hd__and3_1
XFILLER_20_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3804_ _7461_/Q _3549_/X _3716_/X _7264_/Q _3803_/X VGND VGND VPWR VPWR _3816_/B
+ sky130_fd_sc_hd__a221o_2
X_7572_ _7602_/CLK _7572_/D fanout615/X VGND VGND VPWR VPWR _7572_/Q sky130_fd_sc_hd__dfrtp_1
X_4784_ _4785_/A _4794_/D _4785_/C _5231_/B VGND VGND VPWR VPWR _4786_/B sky130_fd_sc_hd__and4_1
XFILLER_119_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6523_ _6523_/A _6523_/B _6523_/C _6523_/D VGND VGND VPWR VPWR _6523_/Y sky130_fd_sc_hd__nor4_1
X_3735_ _7606_/Q _5957_/B _5680_/B _3734_/X VGND VGND VPWR VPWR _3735_/X sky130_fd_sc_hd__a31o_1
XFILLER_146_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6454_ _6791_/C _6455_/C _6771_/C VGND VGND VPWR VPWR _6454_/X sky130_fd_sc_hd__and3_4
X_3666_ _7399_/Q _3525_/X _3663_/X _3665_/X VGND VGND VPWR VPWR _3667_/D sky130_fd_sc_hd__a211o_1
XFILLER_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5405_ _5407_/C _4937_/Y _5270_/X _5274_/X VGND VGND VPWR VPWR _5572_/B sky130_fd_sc_hd__o31ai_1
X_6385_ _7191_/Q _6159_/B _6427_/B1 _6384_/X VGND VGND VPWR VPWR _6385_/X sky130_fd_sc_hd__a31o_1
X_3597_ _7529_/Q _3561_/X _3593_/X _3594_/X _3596_/X VGND VGND VPWR VPWR _3597_/Y
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_133_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5336_ _5109_/A _4977_/X _4981_/X _5007_/Y _5209_/B VGND VGND VPWR VPWR _5617_/A
+ sky130_fd_sc_hd__a221oi_2
X_5267_ _4570_/Y _4859_/Y _4937_/Y _4888_/Y _4854_/X VGND VGND VPWR VPWR _5575_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_102_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7006_ _7616_/CLK _7006_/D fanout610/X VGND VGND VPWR VPWR _7689_/A sky130_fd_sc_hd__dfrtp_1
X_4218_ hold740/X _6863_/A1 _4230_/S VGND VGND VPWR VPWR _4218_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5198_ _4984_/Y _5018_/Y _5196_/Y _5197_/Y VGND VGND VPWR VPWR _5586_/A sky130_fd_sc_hd__o22a_1
XFILLER_55_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4149_ _4149_/A _4196_/B VGND VGND VPWR VPWR _4149_/Y sky130_fd_sc_hd__nand2_8
XFILLER_55_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3520_ hold69/X _3559_/B VGND VGND VPWR VPWR _4340_/A sky130_fd_sc_hd__nor2_8
XFILLER_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold707 hold707/A VGND VGND VPWR VPWR wb_dat_o[6] sky130_fd_sc_hd__buf_12
XFILLER_128_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold718 hold718/A VGND VGND VPWR VPWR hold718/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold729 _7092_/Q VGND VGND VPWR VPWR hold729/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap437 _4966_/B VGND VGND VPWR VPWR _4899_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_115_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3451_ _7381_/Q VGND VGND VPWR VPWR _3451_/Y sky130_fd_sc_hd__clkinv_2
Xmax_cap448 _6119_/X VGND VGND VPWR VPWR _6428_/B1 sky130_fd_sc_hd__buf_12
Xmax_cap459 _6077_/X VGND VGND VPWR VPWR _6428_/A2 sky130_fd_sc_hd__buf_12
XFILLER_131_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6170_ _7451_/Q _6213_/B _6170_/C VGND VGND VPWR VPWR _6170_/X sky130_fd_sc_hd__and3_1
XFILLER_130_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_3_csclk _7236_/CLK VGND VGND VPWR VPWR _7215_/CLK sky130_fd_sc_hd__clkbuf_16
X_5121_ _5120_/Y _5121_/B _5121_/C _5121_/D VGND VGND VPWR VPWR _5121_/Y sky130_fd_sc_hd__nand4b_1
Xhold1407 _6962_/Q VGND VGND VPWR VPWR _6968_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1418 _6983_/Q VGND VGND VPWR VPWR _4235_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5052_ _5512_/C _5038_/B _5051_/Y VGND VGND VPWR VPWR _5055_/B sky130_fd_sc_hd__a21oi_1
Xhold1429 _6986_/Q VGND VGND VPWR VPWR _4238_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4003_ _7281_/Q _5993_/B _5680_/B _3976_/X _4002_/X VGND VGND VPWR VPWR _4003_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_93_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5954_ hold963/X _5999_/A1 _5956_/S VGND VGND VPWR VPWR _5954_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4905_ _5375_/C _4935_/C _5389_/B VGND VGND VPWR VPWR _4906_/C sky130_fd_sc_hd__and3_1
XFILLER_21_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5885_ _5903_/A _5957_/B _6038_/C VGND VGND VPWR VPWR _5893_/S sky130_fd_sc_hd__and3_4
XFILLER_21_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7624_ _4167_/A1 _7624_/D fanout619/X VGND VGND VPWR VPWR _7624_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_21_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4836_ _4836_/A _4836_/B _5146_/B VGND VGND VPWR VPWR _4836_/Y sky130_fd_sc_hd__nor3_2
XFILLER_178_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7555_ _7603_/CLK _7555_/D fanout606/X VGND VGND VPWR VPWR _7555_/Q sky130_fd_sc_hd__dfstp_2
X_4767_ _5407_/A _4810_/C VGND VGND VPWR VPWR _4767_/Y sky130_fd_sc_hd__nand2_2
X_6506_ _7466_/Q _6487_/X _6498_/X _6499_/X _6505_/X VGND VGND VPWR VPWR _6506_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_146_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3718_ _7334_/Q _5939_/B _4487_/B _3571_/X _7358_/Q VGND VGND VPWR VPWR _3718_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7486_ _7512_/CLK _7486_/D fanout608/X VGND VGND VPWR VPWR _7486_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_147_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4698_ _4738_/A _5297_/A _4740_/D _5358_/B VGND VGND VPWR VPWR _4722_/A sky130_fd_sc_hd__and4_1
X_6437_ _7040_/Q _6082_/Y _6423_/X _6436_/X VGND VGND VPWR VPWR _6437_/X sky130_fd_sc_hd__o22a_1
XFILLER_146_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3649_ _7464_/Q _3549_/X _3561_/X _7528_/Q _3648_/X VGND VGND VPWR VPWR _3649_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_106_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6368_ _7068_/Q _6231_/D _6146_/C _6149_/X _7088_/Q VGND VGND VPWR VPWR _6368_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5319_ _5319_/A _5602_/B _5319_/C VGND VGND VPWR VPWR _5319_/Y sky130_fd_sc_hd__nor3_1
XFILLER_102_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6299_ _7337_/Q _6166_/B _6145_/C _6149_/X _7425_/Q VGND VGND VPWR VPWR _6299_/X
+ sky130_fd_sc_hd__a32o_1
Xhold12 hold12/A VGND VGND VPWR VPWR hold8/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 hold23/A VGND VGND VPWR VPWR hold23/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_728 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold34 hold34/A VGND VGND VPWR VPWR hold34/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold45 hold45/A VGND VGND VPWR VPWR hold45/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A VGND VGND VPWR VPWR hold56/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold67 hold67/A VGND VGND VPWR VPWR hold67/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold78 hold78/A VGND VGND VPWR VPWR hold78/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 hold89/A VGND VGND VPWR VPWR hold89/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_9 hold24/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_2__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _7657_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_86_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5670_ _5697_/A0 _5669_/Y _5686_/D _5668_/X VGND VGND VPWR VPWR _5670_/X sky130_fd_sc_hd__o211a_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4621_ _4948_/B _5316_/C VGND VGND VPWR VPWR _5233_/A sky130_fd_sc_hd__nor2_4
XFILLER_190_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7340_ _7562_/CLK _7340_/D fanout621/X VGND VGND VPWR VPWR _7340_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_129_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4552_ hold247/X _6866_/A1 _4552_/S VGND VGND VPWR VPWR _4552_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold504 hold504/A VGND VGND VPWR VPWR hold504/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3503_ _4229_/S hold95/X _3502_/Y VGND VGND VPWR VPWR hold96/A sky130_fd_sc_hd__o21ai_2
Xhold515 _4444_/X VGND VGND VPWR VPWR _7138_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7271_ _7291_/CLK hold99/X fanout596/X VGND VGND VPWR VPWR _7271_/Q sky130_fd_sc_hd__dfrtp_4
Xhold526 _4343_/X VGND VGND VPWR VPWR _7053_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4483_ hold463/X _5869_/A1 _4486_/S VGND VGND VPWR VPWR _4483_/X sky130_fd_sc_hd__mux2_1
Xhold537 _7701_/A VGND VGND VPWR VPWR hold537/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold548 _4252_/X VGND VGND VPWR VPWR _6992_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold559 _7576_/Q VGND VGND VPWR VPWR hold559/X sky130_fd_sc_hd__dlygate4sd3_1
X_6222_ _7365_/Q _6159_/B _6141_/X _6132_/X _7453_/Q VGND VGND VPWR VPWR _6222_/X
+ sky130_fd_sc_hd__a32o_1
X_3434_ _7517_/Q VGND VGND VPWR VPWR _3434_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6153_ _6158_/D _6392_/B _6159_/A VGND VGND VPWR VPWR _6153_/X sky130_fd_sc_hd__and3_4
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5104_ _5318_/C _5111_/D _5311_/C _5112_/B VGND VGND VPWR VPWR _5104_/Y sky130_fd_sc_hd__nand4_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1204 _4449_/A1 VGND VGND VPWR VPWR hold612/A sky130_fd_sc_hd__dlygate4sd3_1
X_6084_ _7139_/Q _6109_/B _6416_/C _6166_/C VGND VGND VPWR VPWR _6084_/X sky130_fd_sc_hd__o211a_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1215 _4459_/A1 VGND VGND VPWR VPWR hold686/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1226 _6821_/A1 VGND VGND VPWR VPWR hold634/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1237 _7291_/Q VGND VGND VPWR VPWR _5676_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1248 _7454_/Q VGND VGND VPWR VPWR hold251/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5035_ _5614_/A _5191_/C _5092_/B VGND VGND VPWR VPWR _5056_/C sky130_fd_sc_hd__and3_1
Xhold1259 _5944_/X VGND VGND VPWR VPWR _7526_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6986_ _7672_/CLK _6986_/D VGND VGND VPWR VPWR _6986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5937_ hold545/X _6045_/A1 _5938_/S VGND VGND VPWR VPWR _5937_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5868_ hold296/X _6039_/A1 _5875_/S VGND VGND VPWR VPWR _5868_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7607_ _7607_/CLK _7607_/D fanout624/X VGND VGND VPWR VPWR _7607_/Q sky130_fd_sc_hd__dfrtp_1
X_4819_ _5017_/A _5017_/B VGND VGND VPWR VPWR _5040_/A sky130_fd_sc_hd__nor2_4
XFILLER_193_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5799_ _5799_/A0 _6006_/A1 _5803_/S VGND VGND VPWR VPWR _5799_/X sky130_fd_sc_hd__mux2_1
X_7538_ _7558_/CLK _7538_/D fanout615/X VGND VGND VPWR VPWR _7538_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7469_ _7583_/CLK _7469_/D fanout631/X VGND VGND VPWR VPWR _7469_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_1_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput102 wb_adr_i[12] VGND VGND VPWR VPWR _4585_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput113 wb_adr_i[22] VGND VGND VPWR VPWR _5096_/C sky130_fd_sc_hd__buf_2
XFILLER_49_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput124 wb_adr_i[3] VGND VGND VPWR VPWR _4992_/C sky130_fd_sc_hd__buf_2
XFILLER_193_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput135 wb_dat_i[12] VGND VGND VPWR VPWR _6842_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput146 wb_dat_i[22] VGND VGND VPWR VPWR _6849_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput157 wb_dat_i[3] VGND VGND VPWR VPWR _6840_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput168 wb_sel_i[3] VGND VGND VPWR VPWR _6827_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_102_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6840_ _6969_/Q _6840_/A2 _6840_/B1 wire537/X _6839_/X VGND VGND VPWR VPWR _6840_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_23_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6771_ _7202_/Q _6771_/B _6771_/C VGND VGND VPWR VPWR _6771_/X sky130_fd_sc_hd__and3_1
XFILLER_16_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3983_ input34/X _5957_/B _3573_/C _3982_/X VGND VGND VPWR VPWR _3983_/X sky130_fd_sc_hd__a31o_1
XFILLER_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5722_ hold894/X _6046_/A1 _5722_/S VGND VGND VPWR VPWR _5722_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_21_csclk _7202_/CLK VGND VGND VPWR VPWR _7586_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_176_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5653_ _6864_/A1 _5653_/A1 _5658_/S VGND VGND VPWR VPWR _5653_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4604_ _4568_/Y _4599_/Y _4990_/A VGND VGND VPWR VPWR _4604_/Y sky130_fd_sc_hd__o21bai_4
X_5584_ _4629_/Y _4674_/Y _5193_/Y _5011_/A VGND VGND VPWR VPWR _5586_/C sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_36_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7583_/CLK sky130_fd_sc_hd__clkbuf_16
X_7323_ _7515_/CLK _7323_/D fanout621/X VGND VGND VPWR VPWR _7323_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_163_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4535_ _4547_/A _4535_/B _5680_/C VGND VGND VPWR VPWR _4540_/S sky130_fd_sc_hd__and3_2
Xhold301 _7406_/Q VGND VGND VPWR VPWR hold301/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 _5852_/X VGND VGND VPWR VPWR _7444_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 _7404_/Q VGND VGND VPWR VPWR hold323/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 _4379_/X VGND VGND VPWR VPWR _7083_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold345 _7564_/Q VGND VGND VPWR VPWR hold345/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7254_ _7254_/CLK _7254_/D fanout618/X VGND VGND VPWR VPWR _7254_/Q sky130_fd_sc_hd__dfrtp_2
X_4466_ _4556_/A1 _4466_/A1 _4468_/S VGND VGND VPWR VPWR _4466_/X sky130_fd_sc_hd__mux2_1
Xhold356 _5771_/X VGND VGND VPWR VPWR _7372_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 _4316_/X VGND VGND VPWR VPWR _7030_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold378 _4331_/X VGND VGND VPWR VPWR _7043_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6205_ wire377/X _6192_/Y _6082_/Y _7316_/Q VGND VGND VPWR VPWR _6205_/X sky130_fd_sc_hd__o2bb2a_1
Xhold389 _7183_/Q VGND VGND VPWR VPWR hold389/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7185_ _7286_/CLK _7185_/D fanout600/X VGND VGND VPWR VPWR _7185_/Q sky130_fd_sc_hd__dfrtp_1
X_4397_ _4397_/A0 _4556_/A1 _4399_/S VGND VGND VPWR VPWR _4397_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6136_ _6158_/D _6161_/D _6146_/C VGND VGND VPWR VPWR _6136_/X sky130_fd_sc_hd__and3_4
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1001 _7199_/Q VGND VGND VPWR VPWR _4512_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1012 hold1491/X VGND VGND VPWR VPWR _4397_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1023 hold1340/X VGND VGND VPWR VPWR _4401_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1034 hold1310/X VGND VGND VPWR VPWR _5844_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_6067_ _7624_/Q _7623_/Q VGND VGND VPWR VPWR _6067_/X sky130_fd_sc_hd__and2b_4
Xhold1045 _4383_/X VGND VGND VPWR VPWR _7086_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1056 _7179_/Q VGND VGND VPWR VPWR _4488_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 hold1264/X VGND VGND VPWR VPWR _6033_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5018_ _5094_/A _5094_/D VGND VGND VPWR VPWR _5018_/Y sky130_fd_sc_hd__nand2_4
Xhold1078 _7239_/Q VGND VGND VPWR VPWR _4560_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1089 _7533_/Q VGND VGND VPWR VPWR _5952_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_207 _7450_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_218 hold87/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_229 _6954_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6969_ _7668_/CLK _6969_/D _6815_/A VGND VGND VPWR VPWR _6969_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_186_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold890 _7186_/Q VGND VGND VPWR VPWR hold890/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1590 _7278_/Q VGND VGND VPWR VPWR _5657_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_730 _6002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_741 _6809_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4320_ hold734/X _5991_/A1 _4321_/S VGND VGND VPWR VPWR _4320_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4251_ hold241/X _5935_/A1 _4257_/S VGND VGND VPWR VPWR _4251_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4182_ _6923_/Q _6911_/A VGND VGND VPWR VPWR _4182_/Y sky130_fd_sc_hd__nor2_1
XFILLER_95_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6823_ _3618_/Y _6823_/A1 _6823_/S VGND VGND VPWR VPWR _7671_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6754_ _7253_/Q _6460_/X _6481_/X _7211_/Q VGND VGND VPWR VPWR _6754_/X sky130_fd_sc_hd__a22o_1
X_3966_ _7112_/Q _3703_/X _3913_/X _3921_/X _3965_/Y VGND VGND VPWR VPWR _3966_/X
+ sky130_fd_sc_hd__a2111o_4
X_5705_ hold37/X hold29/X VGND VGND VPWR VPWR hold38/A sky130_fd_sc_hd__nand2_4
X_6685_ _6675_/Y wire366/X _7321_/Q _6759_/D VGND VGND VPWR VPWR _6685_/X sky130_fd_sc_hd__o2bb2a_1
X_3897_ _7436_/Q _3579_/X _4346_/A _7058_/Q _3896_/X VGND VGND VPWR VPWR _3897_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_176_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5636_ hold702/X _6863_/A1 _5636_/S VGND VGND VPWR VPWR _5636_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5567_ _5567_/A _5567_/B VGND VGND VPWR VPWR _5567_/Y sky130_fd_sc_hd__nand2_1
Xhold120 _3713_/A VGND VGND VPWR VPWR _4511_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7306_ _7307_/CLK _7306_/D _6911_/A VGND VGND VPWR VPWR _7306_/Q sky130_fd_sc_hd__dfrtp_1
Xhold131 _4495_/X VGND VGND VPWR VPWR _7185_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4518_ _4518_/A0 _6012_/A0 _4522_/S VGND VGND VPWR VPWR _4518_/X sky130_fd_sc_hd__mux2_1
Xhold142 _5707_/X VGND VGND VPWR VPWR _7315_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold153 _6928_/Q VGND VGND VPWR VPWR hold153/X sky130_fd_sc_hd__dlygate4sd3_1
X_5498_ _4813_/X _5376_/A _5496_/X _5495_/X _5497_/X VGND VGND VPWR VPWR _5498_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_132_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold164 _7364_/Q VGND VGND VPWR VPWR hold164/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 _5917_/X VGND VGND VPWR VPWR _7502_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7237_ _7242_/CLK _7237_/D fanout616/X VGND VGND VPWR VPWR _7237_/Q sky130_fd_sc_hd__dfrtp_2
Xhold186 _6925_/Q VGND VGND VPWR VPWR _3505_/B sky130_fd_sc_hd__dlygate4sd3_1
X_4449_ _3838_/Y _4449_/A1 _4453_/S VGND VGND VPWR VPWR _7146_/D sky130_fd_sc_hd__mux2_1
Xhold197 _7539_/Q VGND VGND VPWR VPWR hold197/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout600 fanout603/X VGND VGND VPWR VPWR fanout600/X sky130_fd_sc_hd__buf_6
XFILLER_104_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout611 fanout612/X VGND VGND VPWR VPWR fanout611/X sky130_fd_sc_hd__buf_8
XFILLER_104_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout622 fanout623/X VGND VGND VPWR VPWR fanout622/X sky130_fd_sc_hd__buf_8
Xfanout633 input75/X VGND VGND VPWR VPWR fanout633/X sky130_fd_sc_hd__buf_12
Xfanout644 _5462_/A1 VGND VGND VPWR VPWR _4992_/D sky130_fd_sc_hd__buf_12
X_7168_ _7254_/CLK _7168_/D fanout617/X VGND VGND VPWR VPWR _7168_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_98_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6119_ _6151_/B _6392_/B _6416_/C VGND VGND VPWR VPWR _6119_/X sky130_fd_sc_hd__and3_4
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7099_ _7242_/CLK _7099_/D fanout616/X VGND VGND VPWR VPWR _7099_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_560 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_571 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_582 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3820_ _7453_/Q _6861_/A _6002_/A _3819_/X VGND VGND VPWR VPWR _3820_/X sky130_fd_sc_hd__a31o_1
XANTENNA_593 _4116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3751_ _7598_/Q _6020_/A _5680_/B _3714_/X _7223_/Q VGND VGND VPWR VPWR _3751_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_185_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6470_ _6791_/C _6487_/A _6771_/C VGND VGND VPWR VPWR _6474_/C sky130_fd_sc_hd__and3_4
X_3682_ _7351_/Q _5957_/B _5759_/B _3585_/X _7335_/Q VGND VGND VPWR VPWR _3682_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_145_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5421_ _5429_/A _5512_/B _5313_/B _5295_/X VGND VGND VPWR VPWR _5425_/C sky130_fd_sc_hd__a31o_1
XFILLER_161_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput203 _4150_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[35] sky130_fd_sc_hd__buf_12
Xoutput214 _4154_/X VGND VGND VPWR VPWR mgmt_gpio_out[10] sky130_fd_sc_hd__buf_12
X_5352_ _5614_/C _5322_/A _5068_/C _5350_/Y _5579_/B VGND VGND VPWR VPWR _5352_/X
+ sky130_fd_sc_hd__a311o_1
Xoutput225 _7702_/X VGND VGND VPWR VPWR mgmt_gpio_out[22] sky130_fd_sc_hd__buf_12
Xoutput236 _4151_/X VGND VGND VPWR VPWR mgmt_gpio_out[32] sky130_fd_sc_hd__buf_12
XFILLER_99_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput247 _4156_/X VGND VGND VPWR VPWR mgmt_gpio_out[8] sky130_fd_sc_hd__buf_12
XFILLER_114_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4303_ hold125/X hold102/X _4303_/S VGND VGND VPWR VPWR _4303_/X sky130_fd_sc_hd__mux2_1
Xoutput258 _7270_/Q VGND VGND VPWR VPWR pll90_sel[1] sky130_fd_sc_hd__buf_12
XFILLER_114_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput269 _7267_/Q VGND VGND VPWR VPWR pll_sel[1] sky130_fd_sc_hd__buf_12
X_5283_ _5512_/B _5512_/C _5512_/D _5138_/A VGND VGND VPWR VPWR _5565_/A sky130_fd_sc_hd__a31o_1
XFILLER_99_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7022_ _7421_/CLK _7022_/D fanout630/X VGND VGND VPWR VPWR _7022_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4234_ _3902_/Y _4234_/A1 _4239_/S VGND VGND VPWR VPWR _6982_/D sky130_fd_sc_hd__mux2_1
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4165_ _7317_/Q input1/X _4164_/Y VGND VGND VPWR VPWR _4165_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_114_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4096_ _4096_/A0 input58/X _4096_/S VGND VGND VPWR VPWR _6920_/D sky130_fd_sc_hd__mux2_1
XFILLER_70_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6806_ _7243_/Q _6694_/B _6720_/D _6452_/X _7188_/Q VGND VGND VPWR VPWR _6806_/X
+ sky130_fd_sc_hd__a32o_1
X_4998_ _5109_/A _5108_/B VGND VGND VPWR VPWR _4998_/Y sky130_fd_sc_hd__nand2_8
XFILLER_149_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6737_ _6736_/X _6761_/B1 _6812_/S VGND VGND VPWR VPWR _6737_/X sky130_fd_sc_hd__mux2_1
X_3949_ _6959_/Q _5678_/C _6002_/A _3674_/X _7267_/Q VGND VGND VPWR VPWR _3949_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_139_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6668_ _7497_/Q _6694_/B _6720_/D _6485_/X _7553_/Q VGND VGND VPWR VPWR _6668_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_139_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5619_ _4859_/Y _4960_/Y _5001_/Y _4871_/X _4912_/Y VGND VGND VPWR VPWR _5619_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_137_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6599_ _7614_/Q _6451_/X _6457_/X _7574_/Q _6598_/X VGND VGND VPWR VPWR _6599_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_164_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout430 _5061_/A VGND VGND VPWR VPWR _5614_/A sky130_fd_sc_hd__buf_4
XFILLER_120_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout485 _6080_/Y VGND VGND VPWR VPWR _6166_/C sky130_fd_sc_hd__buf_12
XFILLER_101_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5970_ _5970_/A0 _6042_/A1 _5974_/S VGND VGND VPWR VPWR _7549_/D sky130_fd_sc_hd__mux2_1
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4921_ _4921_/A _4921_/B _4921_/C VGND VGND VPWR VPWR _4924_/A sky130_fd_sc_hd__nor3_1
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7640_ _7657_/CLK _7640_/D fanout607/X VGND VGND VPWR VPWR _7640_/Q sky130_fd_sc_hd__dfrtp_1
X_4852_ _4599_/Y _4777_/Y _4779_/X _4833_/X _4830_/Y VGND VGND VPWR VPWR _4923_/B
+ sky130_fd_sc_hd__o221a_2
XANTENNA_390 _3584_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3803_ hold87/A _4547_/A _5939_/B _3710_/X _7074_/Q VGND VGND VPWR VPWR _3803_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_20_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7571_ _7603_/CLK _7571_/D fanout606/X VGND VGND VPWR VPWR _7571_/Q sky130_fd_sc_hd__dfstp_1
X_4783_ _4785_/C _4785_/A _4786_/A _5231_/B _4794_/D VGND VGND VPWR VPWR _4783_/X
+ sky130_fd_sc_hd__a41o_2
XFILLER_165_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6522_ _7475_/Q _6441_/X _6453_/X _7555_/Q _6521_/X VGND VGND VPWR VPWR _6523_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3734_ input48/X _5680_/B _5666_/B _7135_/Q hold56/A VGND VGND VPWR VPWR _3734_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_119_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6453_ _7631_/Q _6485_/B _6469_/A _6563_/C VGND VGND VPWR VPWR _6453_/X sky130_fd_sc_hd__and4_4
XFILLER_9_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3665_ _7471_/Q _3528_/X hold56/A _7136_/Q _3664_/X VGND VGND VPWR VPWR _3665_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5404_ _5404_/A _5404_/B _5404_/C VGND VGND VPWR VPWR _5404_/X sky130_fd_sc_hd__and3_1
XFILLER_174_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6384_ _7253_/Q _6159_/B _6161_/D _6166_/C VGND VGND VPWR VPWR _6384_/X sky130_fd_sc_hd__o211a_1
XFILLER_161_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3596_ _7601_/Q _3569_/X _3574_/X input28/X _3595_/X VGND VGND VPWR VPWR _3596_/X
+ sky130_fd_sc_hd__a221o_1
X_5335_ _5046_/A _5061_/A _5005_/C _4981_/X _5110_/C VGND VGND VPWR VPWR _5616_/C
+ sky130_fd_sc_hd__a32o_1
XFILLER_102_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5266_ _4937_/Y _5088_/Y _5263_/Y _5264_/Y VGND VGND VPWR VPWR _5268_/B sky130_fd_sc_hd__o211ai_1
XFILLER_87_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7005_ _7307_/CLK _7005_/D _6886_/A VGND VGND VPWR VPWR _7005_/Q sky130_fd_sc_hd__dfrtp_1
X_4217_ _4217_/A0 _5697_/A0 _4230_/S VGND VGND VPWR VPWR _6972_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5197_ _5197_/A _5197_/B VGND VGND VPWR VPWR _5197_/Y sky130_fd_sc_hd__nand2_1
X_4148_ _7605_/Q _4147_/A _4147_/Y VGND VGND VPWR VPWR _4148_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_56_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4079_ hold94/A _6925_/Q hold21/A _4079_/B1 VGND VGND VPWR VPWR _4079_/X sky130_fd_sc_hd__a31o_1
XFILLER_71_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_1__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _7668_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_59_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold708 _7376_/Q VGND VGND VPWR VPWR hold708/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_156_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold719 _7112_/Q VGND VGND VPWR VPWR hold719/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3450_ _7389_/Q VGND VGND VPWR VPWR _3450_/Y sky130_fd_sc_hd__clkinv_2
Xmax_cap438 _4953_/B VGND VGND VPWR VPWR _5407_/D sky130_fd_sc_hd__buf_4
XFILLER_143_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap449 _6114_/X VGND VGND VPWR VPWR _6334_/C sky130_fd_sc_hd__buf_12
XFILLER_171_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5120_ _5004_/Y _5088_/Y _5090_/Y _5001_/Y _5119_/Y VGND VGND VPWR VPWR _5120_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5051_ _5051_/A _5051_/B _5051_/C _5466_/B VGND VGND VPWR VPWR _5051_/Y sky130_fd_sc_hd__nand4_1
Xhold1408 hold83/A VGND VGND VPWR VPWR _4057_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1419 _7610_/Q VGND VGND VPWR VPWR hold293/A sky130_fd_sc_hd__dlygate4sd3_1
X_4002_ _7294_/Q _5680_/A _6038_/B _3843_/X _7297_/Q VGND VGND VPWR VPWR _4002_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_38_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5953_ hold415/X _6043_/A1 _5956_/S VGND VGND VPWR VPWR _5953_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4904_ _4904_/A _4904_/B _4904_/C _4904_/D VGND VGND VPWR VPWR _4906_/D sky130_fd_sc_hd__nand4_1
X_5884_ hold587/X _6028_/A1 _5884_/S VGND VGND VPWR VPWR _5884_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7623_ _4167_/A1 _7623_/D fanout620/X VGND VGND VPWR VPWR _7623_/Q sky130_fd_sc_hd__dfrtp_4
X_4835_ _5146_/B _4836_/B _4865_/C VGND VGND VPWR VPWR _4877_/C sky130_fd_sc_hd__o21ai_2
XFILLER_178_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7554_ _7566_/CLK _7554_/D fanout615/X VGND VGND VPWR VPWR _7554_/Q sky130_fd_sc_hd__dfstp_1
X_4766_ _4822_/A _5189_/A _5429_/D VGND VGND VPWR VPWR _4813_/C sky130_fd_sc_hd__and3b_2
X_6505_ _7570_/Q _6457_/X _6500_/X _6503_/X _6504_/X VGND VGND VPWR VPWR _6505_/X
+ sky130_fd_sc_hd__a2111o_1
X_3717_ _4541_/A _3717_/B _4493_/C VGND VGND VPWR VPWR _4382_/A sky130_fd_sc_hd__and3_2
X_7485_ _7497_/CLK hold26/X fanout607/X VGND VGND VPWR VPWR _7485_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_162_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4697_ _4747_/B _5476_/A _5364_/B _5358_/B VGND VGND VPWR VPWR _5203_/C sky130_fd_sc_hd__nand4_2
XFILLER_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6436_ _7218_/Q _6151_/X _6429_/X _6432_/X _6435_/X VGND VGND VPWR VPWR _6436_/X
+ sky130_fd_sc_hd__a2111o_1
X_3648_ _7472_/Q _3528_/X _3574_/X input27/X _3647_/X VGND VGND VPWR VPWR _3648_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_136_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6367_ _6366_/X _6390_/A2 _6812_/S VGND VGND VPWR VPWR _7646_/D sky130_fd_sc_hd__mux2_1
X_3579_ _3905_/B _5628_/A _5661_/B VGND VGND VPWR VPWR _3579_/X sky130_fd_sc_hd__and3_2
X_5318_ _5318_/A _5318_/B _5318_/C VGND VGND VPWR VPWR _5319_/A sky130_fd_sc_hd__and3_1
XFILLER_114_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6298_ _6297_/X _6320_/A2 _6611_/S VGND VGND VPWR VPWR _7643_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold13 hold13/A VGND VGND VPWR VPWR hold13/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold24 hold24/A VGND VGND VPWR VPWR hold24/X sky130_fd_sc_hd__dlygate4sd3_1
X_5249_ _5401_/A _5313_/B _5249_/C VGND VGND VPWR VPWR _5249_/X sky130_fd_sc_hd__and3_1
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold35 hold35/A VGND VGND VPWR VPWR hold35/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold46 hold46/A VGND VGND VPWR VPWR hold46/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 hold57/A VGND VGND VPWR VPWR hold57/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold68 hold68/A VGND VGND VPWR VPWR hold68/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A VGND VGND VPWR VPWR hold79/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4620_ _4948_/A _5074_/A VGND VGND VPWR VPWR _5316_/C sky130_fd_sc_hd__nand2_4
XFILLER_187_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4551_ hold471/X _5673_/A1 _4552_/S VGND VGND VPWR VPWR _7232_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3502_ _4229_/S _3502_/B VGND VGND VPWR VPWR _3502_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold505 hold505/A VGND VGND VPWR VPWR hold505/X sky130_fd_sc_hd__dlygate4sd3_1
X_7270_ _7291_/CLK _7270_/D fanout596/X VGND VGND VPWR VPWR _7270_/Q sky130_fd_sc_hd__dfstp_2
Xhold516 _7496_/Q VGND VGND VPWR VPWR hold516/X sky130_fd_sc_hd__dlygate4sd3_1
X_4482_ _4482_/A0 _6862_/A1 _4486_/S VGND VGND VPWR VPWR _4482_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold527 _7465_/Q VGND VGND VPWR VPWR hold527/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 _4254_/X VGND VGND VPWR VPWR _6993_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6221_ _7557_/Q _6112_/X _6137_/X _7485_/Q _6220_/X VGND VGND VPWR VPWR _6221_/X
+ sky130_fd_sc_hd__a221o_1
X_3433_ hold87/A VGND VGND VPWR VPWR _3433_/Y sky130_fd_sc_hd__inv_2
Xhold549 hold549/A VGND VGND VPWR VPWR hold549/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6152_ _6158_/D _6231_/B _6392_/B _6166_/B VGND VGND VPWR VPWR _6152_/X sky130_fd_sc_hd__and4bb_4
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _5407_/B _5102_/B _4948_/A _5429_/D VGND VGND VPWR VPWR _5103_/X sky130_fd_sc_hd__a211o_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _6082_/Y _6109_/B _6065_/Y VGND VGND VPWR VPWR _6083_/X sky130_fd_sc_hd__a21o_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1205 _4239_/A1 VGND VGND VPWR VPWR hold606/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1216 _4232_/A1 VGND VGND VPWR VPWR hold696/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1227 _4236_/A1 VGND VGND VPWR VPWR hold808/A sky130_fd_sc_hd__dlygate4sd3_1
X_5034_ _5614_/A _5042_/A _5034_/C VGND VGND VPWR VPWR _5056_/B sky130_fd_sc_hd__and3_1
Xhold1238 _7309_/Q VGND VGND VPWR VPWR _5700_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1249 _5863_/X VGND VGND VPWR VPWR _7454_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6985_ _7676_/CLK _6985_/D VGND VGND VPWR VPWR _6985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5936_ hold879/X _6044_/A1 _5938_/S VGND VGND VPWR VPWR _5936_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5867_ _5903_/A _5939_/B _6038_/C VGND VGND VPWR VPWR _5875_/S sky130_fd_sc_hd__and3_4
X_7606_ _7606_/CLK _7606_/D fanout612/X VGND VGND VPWR VPWR _7606_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_139_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4818_ _5375_/A _5186_/B _5186_/C _5042_/A VGND VGND VPWR VPWR _4827_/B sky130_fd_sc_hd__nand4_1
X_5798_ hold317/X _5843_/A1 _5803_/S VGND VGND VPWR VPWR _5798_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7537_ _7584_/CLK _7537_/D fanout613/X VGND VGND VPWR VPWR _7537_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_135_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4749_ _4658_/X _4660_/Y _5027_/B _5027_/D VGND VGND VPWR VPWR _5030_/D sky130_fd_sc_hd__a2bb2oi_2
XFILLER_119_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7468_ _7606_/CLK _7468_/D fanout606/X VGND VGND VPWR VPWR _7468_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_107_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6419_ _7228_/Q _6166_/B _6427_/A3 _6428_/B1 _7080_/Q VGND VGND VPWR VPWR _6419_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_122_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7399_ _7568_/CLK _7399_/D fanout622/X VGND VGND VPWR VPWR _7399_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_103_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput103 wb_adr_i[13] VGND VGND VPWR VPWR _4585_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput114 wb_adr_i[23] VGND VGND VPWR VPWR _5096_/B sky130_fd_sc_hd__buf_2
XFILLER_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput125 wb_adr_i[4] VGND VGND VPWR VPWR _5008_/C sky130_fd_sc_hd__buf_4
XFILLER_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput136 wb_dat_i[13] VGND VGND VPWR VPWR _6845_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput147 wb_dat_i[23] VGND VGND VPWR VPWR _6852_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput158 wb_dat_i[4] VGND VGND VPWR VPWR _6843_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput169 wb_stb_i VGND VGND VPWR VPWR _4116_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_186_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_2_csclk _7236_/CLK VGND VGND VPWR VPWR _7217_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3982_ _7214_/Q _5993_/A _4529_/B _3569_/X _7594_/Q VGND VGND VPWR VPWR _3982_/X
+ sky130_fd_sc_hd__a32o_1
X_6770_ _7074_/Q _6469_/A _6562_/C _6441_/X _7124_/Q VGND VGND VPWR VPWR _6770_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_16_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5721_ hold663/X _5991_/A1 _5722_/S VGND VGND VPWR VPWR _5721_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5652_ _5869_/A1 hold193/X _5658_/S VGND VGND VPWR VPWR _5652_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4603_ _4568_/Y _4599_/Y _5015_/C _4684_/A VGND VGND VPWR VPWR _5490_/B sky130_fd_sc_hd__o22ai_4
XFILLER_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5583_ _5583_/A _5583_/B _5583_/C _5583_/D VGND VGND VPWR VPWR _5587_/A sky130_fd_sc_hd__and4_1
XFILLER_175_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4534_ hold248/X _6866_/A1 _4534_/S VGND VGND VPWR VPWR _4534_/X sky130_fd_sc_hd__mux2_1
X_7322_ _7586_/CLK _7322_/D fanout625/X VGND VGND VPWR VPWR _7322_/Q sky130_fd_sc_hd__dfstp_1
Xhold302 _5809_/X VGND VGND VPWR VPWR _7406_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold313 _7380_/Q VGND VGND VPWR VPWR hold313/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 _5807_/X VGND VGND VPWR VPWR _7404_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold335 _7467_/Q VGND VGND VPWR VPWR hold335/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4465_ _6863_/A1 hold777/X _4468_/S VGND VGND VPWR VPWR _4465_/X sky130_fd_sc_hd__mux2_1
Xhold346 _5987_/X VGND VGND VPWR VPWR _7564_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7253_ _7253_/CLK _7253_/D fanout617/X VGND VGND VPWR VPWR _7253_/Q sky130_fd_sc_hd__dfstp_1
Xhold357 _7058_/Q VGND VGND VPWR VPWR hold357/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold368 hold368/A VGND VGND VPWR VPWR hold368/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6204_ _7356_/Q _6138_/X _6196_/X _6198_/X _6203_/X VGND VGND VPWR VPWR _6204_/Y
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold379 _7070_/Q VGND VGND VPWR VPWR hold379/X sky130_fd_sc_hd__dlygate4sd3_1
X_7184_ _7231_/CLK _7184_/D fanout598/X VGND VGND VPWR VPWR _7184_/Q sky130_fd_sc_hd__dfrtp_4
X_4396_ hold411/X _5869_/A1 _4399_/S VGND VGND VPWR VPWR _4396_/X sky130_fd_sc_hd__mux2_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6135_ _7522_/Q _6131_/B _6334_/C _6180_/A2 _7442_/Q VGND VGND VPWR VPWR _6135_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_112_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1002 _4512_/X VGND VGND VPWR VPWR _7199_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1013 _7126_/Q VGND VGND VPWR VPWR _4431_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1024 hold1304/X VGND VGND VPWR VPWR _5826_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_6066_ _6109_/B _6065_/Y _7623_/Q VGND VGND VPWR VPWR _7623_/D sky130_fd_sc_hd__mux2_1
Xhold1035 _7293_/Q VGND VGND VPWR VPWR _5679_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_133_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1046 _7174_/Q VGND VGND VPWR VPWR _4482_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5017_ _5017_/A _5017_/B _5094_/D VGND VGND VPWR VPWR _5095_/C sky130_fd_sc_hd__and3_2
Xhold1057 _4488_/X VGND VGND VPWR VPWR _7179_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1068 hold1316/X VGND VGND VPWR VPWR _5979_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1079 _4560_/X VGND VGND VPWR VPWR _7239_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_54_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_208 _7450_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_219 _7071_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6968_ _7668_/CLK _6968_/D _6815_/A VGND VGND VPWR VPWR _6968_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5919_ hold752/X _5991_/A1 _5920_/S VGND VGND VPWR VPWR _5919_/X sky130_fd_sc_hd__mux2_1
X_6899_ _6899_/A _6907_/B VGND VGND VPWR VPWR _6899_/X sky130_fd_sc_hd__and2_1
XFILLER_108_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold880 _5936_/X VGND VGND VPWR VPWR _7519_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 _4496_/X VGND VGND VPWR VPWR _7186_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1580 _7636_/Q VGND VGND VPWR VPWR _6108_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1591 _7128_/Q VGND VGND VPWR VPWR hold1591/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_720 _6482_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_731 _6002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_742 _6002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4250_ _4250_/A0 _4249_/X _4258_/S VGND VGND VPWR VPWR _4250_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4181_ input84/X _4171_/D _6923_/Q VGND VGND VPWR VPWR _4181_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6822_ _3655_/Y _6822_/A1 _6823_/S VGND VGND VPWR VPWR _7670_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6753_ _7241_/Q _6694_/B _6720_/D _6474_/B _7053_/Q VGND VGND VPWR VPWR _6758_/C
+ sky130_fd_sc_hd__a32o_1
XFILLER_23_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3965_ _3922_/X _3923_/X _3965_/C _3965_/D VGND VGND VPWR VPWR _3965_/Y sky130_fd_sc_hd__nand4bb_1
XFILLER_149_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5704_ _6028_/A1 hold508/X _5704_/S VGND VGND VPWR VPWR _5704_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6684_ _6684_/A _6684_/B _6684_/C _6809_/D VGND VGND VPWR VPWR _6684_/Y sky130_fd_sc_hd__nor4_1
X_3896_ _7118_/Q _4541_/A _5680_/A _3845_/X VGND VGND VPWR VPWR _3896_/X sky130_fd_sc_hd__a31o_1
XFILLER_31_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5635_ _5635_/A0 _5697_/A0 _5636_/S VGND VGND VPWR VPWR _7259_/D sky130_fd_sc_hd__mux2_1
XFILLER_164_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5566_ _5314_/A _5566_/B _5566_/C _5566_/D VGND VGND VPWR VPWR _5567_/B sky130_fd_sc_hd__and4b_1
XFILLER_191_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold110 _5767_/X VGND VGND VPWR VPWR _7369_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7305_ _7305_/CLK _7305_/D fanout620/X VGND VGND VPWR VPWR _7305_/Q sky130_fd_sc_hd__dfrtp_1
Xhold121 _5682_/X VGND VGND VPWR VPWR _5685_/S sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_163_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold132 _6927_/Q VGND VGND VPWR VPWR hold132/X sky130_fd_sc_hd__dlygate4sd3_1
X_4517_ _5993_/A _5666_/B _5686_/D VGND VGND VPWR VPWR _4522_/S sky130_fd_sc_hd__and3_4
XFILLER_144_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5497_ _4817_/Y _4825_/Y _5189_/Y _5187_/X _4613_/X VGND VGND VPWR VPWR _5497_/X
+ sky130_fd_sc_hd__o2111a_1
Xhold143 _7491_/Q VGND VGND VPWR VPWR hold143/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 _3483_/X VGND VGND VPWR VPWR _3484_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold165 _5762_/X VGND VGND VPWR VPWR _7364_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 _7550_/Q VGND VGND VPWR VPWR hold176/X sky130_fd_sc_hd__dlygate4sd3_1
X_7236_ _7236_/CLK _7236_/D fanout603/X VGND VGND VPWR VPWR _7236_/Q sky130_fd_sc_hd__dfstp_1
X_4448_ _3902_/Y _4448_/A1 _4453_/S VGND VGND VPWR VPWR _7145_/D sky130_fd_sc_hd__mux2_1
XFILLER_104_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold187 _3505_/Y VGND VGND VPWR VPWR hold187/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout601 fanout602/X VGND VGND VPWR VPWR _6903_/A sky130_fd_sc_hd__buf_6
Xhold198 _5959_/X VGND VGND VPWR VPWR _7539_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout612 fanout633/X VGND VGND VPWR VPWR fanout612/X sky130_fd_sc_hd__buf_6
Xfanout623 fanout624/X VGND VGND VPWR VPWR fanout623/X sky130_fd_sc_hd__buf_6
XFILLER_132_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout634 fanout635/X VGND VGND VPWR VPWR _6815_/A sky130_fd_sc_hd__buf_8
XFILLER_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4379_ hold333/X _5789_/A1 _4381_/S VGND VGND VPWR VPWR _4379_/X sky130_fd_sc_hd__mux2_1
X_7167_ _7254_/CLK _7167_/D fanout619/X VGND VGND VPWR VPWR _7167_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_86_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout645 _4948_/A VGND VGND VPWR VPWR _5407_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_58_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6118_ _7338_/Q _6157_/C _6166_/C wire484/X _6117_/X VGND VGND VPWR VPWR _6118_/X
+ sky130_fd_sc_hd__a311o_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7098_ _7238_/CLK _7098_/D fanout602/X VGND VGND VPWR VPWR _7098_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_100_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__1128_ _3776_/X VGND VGND VPWR VPWR clkbuf_0__1128_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6049_ _3421_/Y _7139_/Q _7293_/Q _6048_/X _6049_/B2 VGND VGND VPWR VPWR _7618_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_86_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_82_csclk _7095_/CLK VGND VGND VPWR VPWR _7160_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_127_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_20_csclk _7202_/CLK VGND VGND VPWR VPWR _7304_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_76_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_35_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7599_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_550 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_561 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_572 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_583 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_594 _6759_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3750_ _7318_/Q _5993_/B _5682_/C _3557_/X _7574_/Q VGND VGND VPWR VPWR _3750_/X
+ sky130_fd_sc_hd__a32o_1
X_3681_ input8/X _3573_/X _3574_/X input25/X _3680_/X VGND VGND VPWR VPWR _3691_/A
+ sky130_fd_sc_hd__a221o_4
XFILLER_9_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5420_ _5093_/B _5040_/C _5313_/A _5291_/B _5291_/C VGND VGND VPWR VPWR _5425_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput204 _4148_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[36] sky130_fd_sc_hd__buf_12
X_5351_ _5476_/A _5322_/A _5233_/C _5074_/B VGND VGND VPWR VPWR _5579_/B sky130_fd_sc_hd__a31o_1
XFILLER_161_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput215 _7694_/X VGND VGND VPWR VPWR mgmt_gpio_out[11] sky130_fd_sc_hd__buf_12
XFILLER_160_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput226 _7703_/X VGND VGND VPWR VPWR mgmt_gpio_out[23] sky130_fd_sc_hd__buf_12
XFILLER_160_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput237 _4152_/X VGND VGND VPWR VPWR mgmt_gpio_out[33] sky130_fd_sc_hd__buf_12
X_4302_ hold619/X _5991_/A1 _4303_/S VGND VGND VPWR VPWR _4302_/X sky130_fd_sc_hd__mux2_1
Xoutput248 _4184_/Y VGND VGND VPWR VPWR pad_flash_clk_oeb sky130_fd_sc_hd__buf_12
Xoutput259 _7271_/Q VGND VGND VPWR VPWR pll90_sel[2] sky130_fd_sc_hd__buf_12
X_5282_ _5279_/Y _5280_/X _5281_/X _4847_/X VGND VGND VPWR VPWR _5282_/X sky130_fd_sc_hd__o31a_1
X_4233_ _3966_/X _4233_/A1 _4239_/S VGND VGND VPWR VPWR _6981_/D sky130_fd_sc_hd__mux2_1
X_7021_ _7421_/CLK _7021_/D fanout630/X VGND VGND VPWR VPWR _7021_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_114_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4164_ input1/X input2/X VGND VGND VPWR VPWR _4164_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4095_ _7257_/Q _7256_/Q _4104_/D _7258_/Q VGND VGND VPWR VPWR _4096_/S sky130_fd_sc_hd__and4b_1
XFILLER_55_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6805_ _7233_/Q _6720_/C _6536_/C _6454_/X _7193_/Q VGND VGND VPWR VPWR _6805_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_169_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4997_ _5109_/A _5025_/B _5008_/C VGND VGND VPWR VPWR _5034_/C sky130_fd_sc_hd__and3_1
XFILLER_23_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6736_ _6735_/X _7658_/Q _7140_/Q VGND VGND VPWR VPWR _6736_/X sky130_fd_sc_hd__mux2_1
X_3948_ _7299_/Q _5682_/C _5984_/B _3554_/X _7563_/Q VGND VGND VPWR VPWR _3948_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_149_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6667_ _7601_/Q _6474_/B _6464_/X _7465_/Q _6666_/X VGND VGND VPWR VPWR _6675_/B
+ sky130_fd_sc_hd__a221o_1
X_3879_ _7316_/Q _5993_/B _5682_/C hold56/A _7133_/Q VGND VGND VPWR VPWR _3879_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_109_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5618_ _5618_/A _5618_/B _5618_/C VGND VGND VPWR VPWR _5618_/Y sky130_fd_sc_hd__nand3_1
XFILLER_136_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6598_ _7590_/Q _6468_/X _6487_/X _7470_/Q _6589_/X VGND VGND VPWR VPWR _6598_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_152_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5549_ _5549_/A _5549_/B VGND VGND VPWR VPWR _5553_/A sky130_fd_sc_hd__nand2_1
XFILLER_155_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_0__f_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR _7680_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7219_ _7294_/CLK _7219_/D fanout597/X VGND VGND VPWR VPWR _7219_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout442 _5595_/D VGND VGND VPWR VPWR _5358_/B sky130_fd_sc_hd__buf_4
XFILLER_171_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout486 _6080_/Y VGND VGND VPWR VPWR _6145_/C sky130_fd_sc_hd__buf_6
XFILLER_171_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4920_ _5375_/C _4923_/B _5452_/A _4934_/C VGND VGND VPWR VPWR _4921_/B sky130_fd_sc_hd__and4_1
X_4851_ _5614_/C _4972_/C VGND VGND VPWR VPWR _4971_/C sky130_fd_sc_hd__nand2_1
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_380 _3531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_391 _4275_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3802_ _7284_/Q _5993_/B _4481_/A _3798_/X _3801_/X VGND VGND VPWR VPWR _3816_/A
+ sky130_fd_sc_hd__a311o_1
X_7570_ _7613_/CLK _7570_/D fanout625/X VGND VGND VPWR VPWR _7570_/Q sky130_fd_sc_hd__dfstp_2
X_4782_ _4785_/C _4785_/A _4786_/A _5231_/B VGND VGND VPWR VPWR _4782_/Y sky130_fd_sc_hd__nand4_2
XFILLER_20_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6521_ _7435_/Q _6099_/B _6694_/C _6458_/X _7419_/Q VGND VGND VPWR VPWR _6521_/X
+ sky130_fd_sc_hd__a32o_1
X_3733_ _7125_/Q _5903_/A _4535_/B _3574_/X input24/X VGND VGND VPWR VPWR _3733_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_146_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6452_ _6791_/B _6645_/B _6645_/C VGND VGND VPWR VPWR _6452_/X sky130_fd_sc_hd__and3_4
XFILLER_146_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3664_ _7319_/Q _5993_/B _5682_/C _3557_/X _7575_/Q VGND VGND VPWR VPWR _3664_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_134_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5403_ _5400_/X _5573_/C _5403_/C VGND VGND VPWR VPWR _5403_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_146_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3595_ _7497_/Q _5903_/A _5975_/B _3573_/X input10/X VGND VGND VPWR VPWR _3595_/X
+ sky130_fd_sc_hd__a32o_1
X_6383_ _7684_/Q _6359_/B _6309_/C _6132_/X _7118_/Q VGND VGND VPWR VPWR _6383_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_133_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5334_ _4982_/Y _5001_/Y _5212_/Y _4976_/Y _5216_/X VGND VGND VPWR VPWR _5537_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_88_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5265_ _4943_/A _4935_/C _4934_/C _5452_/C _5092_/A VGND VGND VPWR VPWR _5265_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_87_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7004_ _7307_/CLK _7004_/D _6886_/A VGND VGND VPWR VPWR _7004_/Q sky130_fd_sc_hd__dfrtp_1
X_4216_ _5669_/B _4505_/B _5680_/C VGND VGND VPWR VPWR _4230_/S sky130_fd_sc_hd__and3_2
X_5196_ _5196_/A _5614_/A VGND VGND VPWR VPWR _5196_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4147_ _4147_/A _4147_/B VGND VGND VPWR VPWR _4147_/Y sky130_fd_sc_hd__nand2_2
XFILLER_110_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4078_ _4078_/A1 _3508_/S _4043_/Y _4077_/X VGND VGND VPWR VPWR _4078_/X sky130_fd_sc_hd__a31o_1
XFILLER_43_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6719_ _7042_/Q _6451_/X _6471_/X _7047_/Q _6718_/X VGND VGND VPWR VPWR _6725_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_109_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7699_ _7699_/A VGND VGND VPWR VPWR _7699_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold709 _5775_/X VGND VGND VPWR VPWR _7376_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap439 _4901_/B VGND VGND VPWR VPWR _4866_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_170_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5050_ _5050_/A _5050_/B _5050_/C VGND VGND VPWR VPWR _5051_/A sky130_fd_sc_hd__nor3_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1409 _6982_/Q VGND VGND VPWR VPWR _4234_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_4001_ _7096_/Q _3713_/X _3716_/X _7261_/Q _4000_/X VGND VGND VPWR VPWR _4001_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_111_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5952_ _5952_/A0 _6042_/A1 _5956_/S VGND VGND VPWR VPWR _5952_/X sky130_fd_sc_hd__mux2_1
X_4903_ _5375_/C _5452_/A _5389_/B _4957_/C VGND VGND VPWR VPWR _4904_/B sky130_fd_sc_hd__nand4_1
X_5883_ hold477/X _6045_/A1 _5884_/S VGND VGND VPWR VPWR _5883_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7622_ _7680_/CLK _7622_/D _6886_/A VGND VGND VPWR VPWR _7622_/Q sky130_fd_sc_hd__dfrtp_1
X_4834_ _4704_/A _5146_/B _5000_/C VGND VGND VPWR VPWR _4865_/C sky130_fd_sc_hd__o21ai_4
XFILLER_21_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7553_ _7553_/CLK _7553_/D fanout622/X VGND VGND VPWR VPWR _7553_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_147_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4765_ _5074_/A _4948_/B VGND VGND VPWR VPWR _4810_/C sky130_fd_sc_hd__nor2_1
XFILLER_193_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6504_ _7330_/Q _6469_/X _6471_/X _7322_/Q _6490_/X VGND VGND VPWR VPWR _6504_/X
+ sky130_fd_sc_hd__a221o_1
X_3716_ _5661_/A _4340_/A _5678_/C VGND VGND VPWR VPWR _3716_/X sky130_fd_sc_hd__and3_1
X_7484_ _7497_/CLK _7484_/D fanout608/X VGND VGND VPWR VPWR _7484_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_146_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4696_ _5025_/C _5027_/B _5027_/C _5025_/B VGND VGND VPWR VPWR _5011_/B sky130_fd_sc_hd__nand4_2
X_6435_ _6428_/X _6359_/B _6426_/X _6434_/X VGND VGND VPWR VPWR _6435_/X sky130_fd_sc_hd__a211o_1
XFILLER_174_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3647_ _7576_/Q _5993_/A _5993_/B _3546_/X _7536_/Q VGND VGND VPWR VPWR _3647_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_161_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6366_ _6366_/A1 _6109_/X _6365_/X _6811_/S VGND VGND VPWR VPWR _6366_/X sky130_fd_sc_hd__o22a_1
XFILLER_136_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3578_ _5682_/A _5682_/B _6002_/B VGND VGND VPWR VPWR _4257_/S sky130_fd_sc_hd__and3_4
XFILLER_115_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5317_ _4992_/D _5512_/C _5084_/X _5316_/X _5404_/C VGND VGND VPWR VPWR _5602_/B
+ sky130_fd_sc_hd__a32o_1
X_6297_ _6686_/S _6297_/A2 _6295_/X _6296_/X VGND VGND VPWR VPWR _6297_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold14 hold14/A VGND VGND VPWR VPWR hold14/X sky130_fd_sc_hd__dlygate4sd3_1
X_5248_ _4570_/Y _4862_/Y _4871_/X _4888_/Y _5009_/Y VGND VGND VPWR VPWR _5256_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_102_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold25 hold25/A VGND VGND VPWR VPWR hold25/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A VGND VGND VPWR VPWR hold36/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold47 hold47/A VGND VGND VPWR VPWR hold47/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold58 hold58/A VGND VGND VPWR VPWR hold58/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 hold69/A VGND VGND VPWR VPWR hold69/X sky130_fd_sc_hd__clkbuf_8
XFILLER_56_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5179_ _5551_/A1 _5181_/C _5490_/B _5186_/C _4770_/A VGND VGND VPWR VPWR _5552_/A
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_56_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4550_ _4550_/A0 _6864_/A1 _4552_/S VGND VGND VPWR VPWR _4550_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3501_ hold94/X _3508_/S _3500_/X VGND VGND VPWR VPWR hold95/A sky130_fd_sc_hd__a21oi_2
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold506 _7068_/Q VGND VGND VPWR VPWR hold506/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4481_ _4481_/A hold98/A _6861_/C VGND VGND VPWR VPWR _4486_/S sky130_fd_sc_hd__and3_2
Xwire492 _5042_/C VGND VGND VPWR VPWR _5291_/B sky130_fd_sc_hd__clkbuf_2
Xhold517 _5910_/X VGND VGND VPWR VPWR _7496_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold528 _5875_/X VGND VGND VPWR VPWR _7465_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold539 _7173_/Q VGND VGND VPWR VPWR hold539/X sky130_fd_sc_hd__dlygate4sd3_1
X_6220_ _7533_/Q _6157_/C _6146_/C _6077_/X _7509_/Q VGND VGND VPWR VPWR _6220_/X
+ sky130_fd_sc_hd__a32o_1
X_3432_ _7533_/Q VGND VGND VPWR VPWR _3432_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6151_ _6158_/D _6151_/B _6392_/B _6231_/D VGND VGND VPWR VPWR _6151_/X sky130_fd_sc_hd__and4_4
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _5407_/B _5102_/B VGND VGND VPWR VPWR _5318_/C sky130_fd_sc_hd__nand2_1
XFILLER_111_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _6082_/A _6082_/B VGND VGND VPWR VPWR _6082_/Y sky130_fd_sc_hd__nand2_8
XFILLER_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1206 _4235_/A1 VGND VGND VPWR VPWR hold608/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1217 _4233_/A1 VGND VGND VPWR VPWR hold714/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1228 _6817_/A1 VGND VGND VPWR VPWR hold645/A sky130_fd_sc_hd__dlygate4sd3_1
X_5033_ _5042_/A _5311_/C _5089_/A VGND VGND VPWR VPWR _5059_/B sky130_fd_sc_hd__and3_1
Xhold1239 _7299_/Q VGND VGND VPWR VPWR _5688_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6984_ _7668_/CLK _6984_/D VGND VGND VPWR VPWR _6984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5935_ hold223/X _5935_/A1 _5938_/S VGND VGND VPWR VPWR _7518_/D sky130_fd_sc_hd__mux2_1
XFILLER_179_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5866_ hold256/X hold102/X _5866_/S VGND VGND VPWR VPWR _5866_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7605_ _7613_/CLK _7605_/D fanout626/X VGND VGND VPWR VPWR _7605_/Q sky130_fd_sc_hd__dfrtp_4
X_4817_ _5375_/A _5189_/C VGND VGND VPWR VPWR _4817_/Y sky130_fd_sc_hd__nand2_1
X_5797_ hold976/X _6040_/A1 _5803_/S VGND VGND VPWR VPWR _5797_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7536_ _7616_/CLK _7536_/D fanout611/X VGND VGND VPWR VPWR _7536_/Q sky130_fd_sc_hd__dfrtp_2
X_4748_ _5476_/A _4748_/B VGND VGND VPWR VPWR _4751_/C sky130_fd_sc_hd__nand2_1
XFILLER_107_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7467_ _7603_/CLK _7467_/D fanout611/X VGND VGND VPWR VPWR _7467_/Q sky130_fd_sc_hd__dfstp_2
X_4679_ _5015_/C _4684_/A _4668_/C VGND VGND VPWR VPWR _4740_/D sky130_fd_sc_hd__a21oi_4
X_6418_ _7238_/Q _6124_/X _6309_/C _7168_/Q _6417_/X VGND VGND VPWR VPWR _6418_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7398_ _7398_/CLK _7398_/D fanout627/X VGND VGND VPWR VPWR _7398_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_122_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6349_ _7165_/Q _6309_/C _6149_/X _7087_/Q _6348_/X VGND VGND VPWR VPWR _6349_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput104 wb_adr_i[14] VGND VGND VPWR VPWR _4585_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput115 wb_adr_i[24] VGND VGND VPWR VPWR _4113_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_88_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput126 wb_adr_i[5] VGND VGND VPWR VPWR input126/X sky130_fd_sc_hd__clkbuf_1
Xinput137 wb_dat_i[14] VGND VGND VPWR VPWR _6848_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput148 wb_dat_i[24] VGND VGND VPWR VPWR _6831_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput159 wb_dat_i[5] VGND VGND VPWR VPWR _6846_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3981_ _7131_/Q hold56/A _3574_/X input20/X _3980_/X VGND VGND VPWR VPWR _3995_/B
+ sky130_fd_sc_hd__a221o_2
X_5720_ hold958/X _6044_/A1 _5722_/S VGND VGND VPWR VPWR _5720_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5651_ _5697_/A0 _5651_/A1 _5658_/S VGND VGND VPWR VPWR _5651_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4602_ _4568_/Y _4599_/Y _5015_/C _4684_/A VGND VGND VPWR VPWR _4704_/C sky130_fd_sc_hd__o22a_2
XFILLER_191_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5582_ _4761_/A _5068_/C _4989_/X _5581_/X VGND VGND VPWR VPWR _5583_/D sky130_fd_sc_hd__a211oi_1
X_7321_ _7547_/CLK _7321_/D fanout607/X VGND VGND VPWR VPWR _7321_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_190_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4533_ hold733/X _5673_/A1 _4534_/S VGND VGND VPWR VPWR _7217_/D sky130_fd_sc_hd__mux2_1
Xhold303 _7297_/Q VGND VGND VPWR VPWR hold303/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold314 _5780_/X VGND VGND VPWR VPWR _7380_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold325 _7340_/Q VGND VGND VPWR VPWR hold325/X sky130_fd_sc_hd__dlygate4sd3_1
X_7252_ _7252_/CLK _7252_/D fanout618/X VGND VGND VPWR VPWR _7252_/Q sky130_fd_sc_hd__dfrtp_4
Xhold336 _5878_/X VGND VGND VPWR VPWR _7467_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4464_ _6862_/A1 _4464_/A1 _4468_/S VGND VGND VPWR VPWR _4464_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold347 _7572_/Q VGND VGND VPWR VPWR hold347/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold358 _4349_/X VGND VGND VPWR VPWR _7058_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6203_ _6194_/X _6309_/B _6201_/X _6200_/X _6202_/X VGND VGND VPWR VPWR _6203_/X
+ sky130_fd_sc_hd__a2111o_1
Xhold369 _7191_/Q VGND VGND VPWR VPWR hold369/X sky130_fd_sc_hd__dlygate4sd3_1
X_7183_ _7254_/CLK _7183_/D fanout618/X VGND VGND VPWR VPWR _7183_/Q sky130_fd_sc_hd__dfrtp_4
X_4395_ _4395_/A0 _6862_/A1 _4399_/S VGND VGND VPWR VPWR _4395_/X sky130_fd_sc_hd__mux2_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6134_ _7554_/Q _6131_/B _6432_/A3 _6133_/X _7474_/Q VGND VGND VPWR VPWR _6134_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1003 _7189_/Q VGND VGND VPWR VPWR _4500_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1014 _4431_/X VGND VGND VPWR VPWR _7126_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6065_ _7139_/Q _6109_/B VGND VGND VPWR VPWR _6065_/Y sky130_fd_sc_hd__nor2_2
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1025 hold1384/X VGND VGND VPWR VPWR _5781_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1036 _5679_/X VGND VGND VPWR VPWR _7293_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1047 _4482_/X VGND VGND VPWR VPWR _7174_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1058 _7056_/Q VGND VGND VPWR VPWR _4347_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5016_ _5195_/B _5476_/B _5311_/A _5249_/C VGND VGND VPWR VPWR _5047_/C sky130_fd_sc_hd__nand4_1
XFILLER_66_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1069 _7169_/Q VGND VGND VPWR VPWR _4476_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_209 _7047_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6967_ _7668_/CLK _6967_/D _6815_/A VGND VGND VPWR VPWR _6967_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_13_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5918_ hold955/X _5999_/A1 _5920_/S VGND VGND VPWR VPWR _5918_/X sky130_fd_sc_hd__mux2_1
X_6898_ _6899_/A _6907_/B VGND VGND VPWR VPWR _6898_/X sky130_fd_sc_hd__and2_1
X_5849_ _5849_/A _6029_/B VGND VGND VPWR VPWR _5857_/S sky130_fd_sc_hd__nand2_8
XFILLER_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7519_ _7599_/CLK _7519_/D fanout629/X VGND VGND VPWR VPWR _7519_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold870 _5830_/X VGND VGND VPWR VPWR _7425_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold881 _7407_/Q VGND VGND VPWR VPWR hold881/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold892 _7413_/Q VGND VGND VPWR VPWR hold892/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1570 _7663_/Q VGND VGND VPWR VPWR _6814_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1581 _6950_/Q VGND VGND VPWR VPWR _3481_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_83_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1592 _7221_/Q VGND VGND VPWR VPWR hold1592/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_710 _5007_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_721 _6506_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_732 _6002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_743 _5869_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4180_ _4092_/S _4179_/Y _3464_/X VGND VGND VPWR VPWR _6957_/D sky130_fd_sc_hd__a21o_1
XFILLER_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6821_ _3692_/Y _6821_/A1 _6823_/S VGND VGND VPWR VPWR _7669_/D sky130_fd_sc_hd__mux2_1
XFILLER_51_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6752_ _7123_/Q _6441_/X _6482_/X _7113_/Q VGND VGND VPWR VPWR _6758_/B sky130_fd_sc_hd__a22o_1
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3964_ _3937_/X _3964_/B _3964_/C _3964_/D VGND VGND VPWR VPWR _3965_/D sky130_fd_sc_hd__and4b_1
XFILLER_50_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5703_ hold50/X hold58/X _5703_/S VGND VGND VPWR VPWR hold59/A sky130_fd_sc_hd__mux2_1
XFILLER_50_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6683_ _7385_/Q _6481_/X _6680_/X _6682_/X VGND VGND VPWR VPWR _6684_/C sky130_fd_sc_hd__a211o_1
X_3895_ _7226_/Q _5628_/A hold98/A _5849_/A _7444_/Q VGND VGND VPWR VPWR _3895_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_31_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5634_ hold24/X _5669_/B _5680_/C VGND VGND VPWR VPWR _5636_/S sky130_fd_sc_hd__and3_1
XFILLER_136_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5565_ _5565_/A _5565_/B VGND VGND VPWR VPWR _5566_/C sky130_fd_sc_hd__nor2_1
XFILLER_191_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold100 _6938_/Q VGND VGND VPWR VPWR hold100/X sky130_fd_sc_hd__dlygate4sd3_1
X_7304_ _7304_/CLK _7304_/D fanout620/X VGND VGND VPWR VPWR _7304_/Q sky130_fd_sc_hd__dfrtp_1
X_4516_ hold413/X _5926_/A0 _4516_/S VGND VGND VPWR VPWR _4516_/X sky130_fd_sc_hd__mux2_1
Xhold111 _7384_/Q VGND VGND VPWR VPWR hold111/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 hold122/A VGND VGND VPWR VPWR _7295_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 _3498_/X VGND VGND VPWR VPWR hold133/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5496_ _4707_/X _4711_/X _5375_/A VGND VGND VPWR VPWR _5496_/X sky130_fd_sc_hd__o21a_1
Xhold144 _5905_/X VGND VGND VPWR VPWR _7491_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold155 _3547_/D VGND VGND VPWR VPWR _3568_/C sky130_fd_sc_hd__dlygate4sd3_1
X_7235_ _7255_/CLK _7235_/D fanout618/X VGND VGND VPWR VPWR _7235_/Q sky130_fd_sc_hd__dfrtp_1
Xhold166 _7582_/Q VGND VGND VPWR VPWR hold166/X sky130_fd_sc_hd__dlygate4sd3_1
X_4447_ _3966_/X _4447_/A1 _4453_/S VGND VGND VPWR VPWR _7144_/D sky130_fd_sc_hd__mux2_1
Xhold177 _5971_/X VGND VGND VPWR VPWR _7550_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 _3506_/X VGND VGND VPWR VPWR hold188/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 _7195_/Q VGND VGND VPWR VPWR hold199/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout602 fanout603/X VGND VGND VPWR VPWR fanout602/X sky130_fd_sc_hd__buf_8
XFILLER_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout613 fanout615/X VGND VGND VPWR VPWR fanout613/X sky130_fd_sc_hd__buf_8
Xfanout624 fanout632/X VGND VGND VPWR VPWR fanout624/X sky130_fd_sc_hd__buf_8
X_7166_ _7254_/CLK _7166_/D fanout617/X VGND VGND VPWR VPWR _7166_/Q sky130_fd_sc_hd__dfstp_1
Xfanout635 input164/X VGND VGND VPWR VPWR fanout635/X sky130_fd_sc_hd__buf_6
X_4378_ hold409/X _5869_/A1 _4381_/S VGND VGND VPWR VPWR _4378_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_1_csclk _7095_/CLK VGND VGND VPWR VPWR _7240_/CLK sky130_fd_sc_hd__clkbuf_16
Xfanout646 _4992_/A VGND VGND VPWR VPWR _4948_/A sky130_fd_sc_hd__buf_6
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6117_ _7426_/Q _6432_/A3 wire455/A _7346_/Q _6116_/X VGND VGND VPWR VPWR _6117_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7097_ _7238_/CLK _7097_/D fanout602/X VGND VGND VPWR VPWR _7097_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6048_ _4121_/Y _7142_/Q _6047_/Y VGND VGND VPWR VPWR _6048_/X sky130_fd_sc_hd__a21o_1
XFILLER_73_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_540 input81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_551 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_562 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_573 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_584 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_595 _6809_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3680_ _7375_/Q _3572_/X _4275_/S input40/X _3679_/X VGND VGND VPWR VPWR _3680_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_145_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5350_ _5350_/A _5350_/B VGND VGND VPWR VPWR _5350_/Y sky130_fd_sc_hd__nand2_1
Xoutput205 _4146_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[37] sky130_fd_sc_hd__buf_12
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput216 _7695_/X VGND VGND VPWR VPWR mgmt_gpio_out[12] sky130_fd_sc_hd__buf_12
Xoutput227 _7704_/X VGND VGND VPWR VPWR mgmt_gpio_out[24] sky130_fd_sc_hd__buf_12
XFILLER_5_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput238 _7712_/X VGND VGND VPWR VPWR mgmt_gpio_out[34] sky130_fd_sc_hd__buf_12
X_4301_ hold231/X hold85/X _4303_/S VGND VGND VPWR VPWR _4301_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput249 _4181_/X VGND VGND VPWR VPWR pad_flash_csb sky130_fd_sc_hd__buf_12
XFILLER_99_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5281_ _5407_/A _5429_/D _5189_/D _4972_/C _4972_/X VGND VGND VPWR VPWR _5281_/X
+ sky130_fd_sc_hd__a41o_1
X_7020_ _7421_/CLK _7020_/D fanout630/X VGND VGND VPWR VPWR _7020_/Q sky130_fd_sc_hd__dfrtp_1
X_4232_ _4037_/Y _4232_/A1 _4239_/S VGND VGND VPWR VPWR _6980_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4163_ _7294_/Q _4171_/C _4171_/D _6953_/Q _4162_/Y VGND VGND VPWR VPWR _4163_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_67_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4094_ _4053_/A input58/X _4094_/S VGND VGND VPWR VPWR _6921_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6804_ _7198_/Q _6457_/X _6463_/X _7228_/Q _6803_/X VGND VGND VPWR VPWR _6809_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4996_ _5614_/A _5043_/B _5614_/B _5311_/A VGND VGND VPWR VPWR _4996_/Y sky130_fd_sc_hd__nand4_1
XFILLER_168_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6735_ wire374/X _6734_/Y _7037_/Q _6759_/D VGND VGND VPWR VPWR _6735_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_189_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3947_ _7037_/Q _5682_/C _4505_/B _3530_/X _7539_/Q VGND VGND VPWR VPWR _3947_/X
+ sky130_fd_sc_hd__a32o_1
X_6666_ _7441_/Q _6099_/B _6694_/C _6480_/X _7537_/Q VGND VGND VPWR VPWR _6666_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_177_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3878_ _7572_/Q _3557_/X _5689_/A _4196_/A _3877_/X VGND VGND VPWR VPWR _3878_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_191_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5617_ _5617_/A _5617_/B _5617_/C VGND VGND VPWR VPWR _5618_/C sky130_fd_sc_hd__and3_1
XFILLER_192_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6597_ _7366_/Q _6445_/X _6463_/X _7398_/Q _6596_/X VGND VGND VPWR VPWR _6597_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_136_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5548_ _5490_/B _5485_/X _5364_/X _5171_/X _5493_/B VGND VGND VPWR VPWR _5548_/Y
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_155_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5479_ _5595_/B _5595_/D _5375_/C _4707_/X VGND VGND VPWR VPWR _5480_/A sky130_fd_sc_hd__a31o_1
X_7218_ _7312_/CLK _7218_/D _6907_/A VGND VGND VPWR VPWR _7218_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout421 _4511_/A VGND VGND VPWR VPWR _5682_/A sky130_fd_sc_hd__buf_8
XFILLER_48_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7149_ _7672_/CLK _7149_/D VGND VGND VPWR VPWR _7149_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout465 _4738_/B VGND VGND VPWR VPWR _5490_/C sky130_fd_sc_hd__buf_4
Xfanout476 _6516_/C VGND VGND VPWR VPWR _6720_/D sky130_fd_sc_hd__buf_12
Xfanout487 _6157_/C VGND VGND VPWR VPWR _6160_/D sky130_fd_sc_hd__buf_12
Xfanout498 _5611_/A2 VGND VGND VPWR VPWR _5604_/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_101_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4850_ _4959_/C _5233_/A _4972_/C VGND VGND VPWR VPWR _4850_/X sky130_fd_sc_hd__and3_1
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_370 _3514_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_381 _3531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_392 _6011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3801_ hold40/A _3519_/X _3531_/X _7485_/Q _3800_/X VGND VGND VPWR VPWR _3801_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_33_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4781_ _5008_/C _4781_/B _4781_/C _5231_/B VGND VGND VPWR VPWR _4781_/Y sky130_fd_sc_hd__nand4_2
XFILLER_20_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6520_ _7507_/Q _6484_/X _6485_/X _7547_/Q _6519_/X VGND VGND VPWR VPWR _6523_/C
+ sky130_fd_sc_hd__a221o_1
X_3732_ _7276_/Q _5650_/A _3728_/X _3729_/X _3731_/X VGND VGND VPWR VPWR _3732_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_119_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6451_ _6791_/B _6791_/C _6645_/B VGND VGND VPWR VPWR _6451_/X sky130_fd_sc_hd__and3_4
X_3663_ _7423_/Q hold24/A _5628_/A _3530_/X _7543_/Q VGND VGND VPWR VPWR _3663_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_146_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5402_ _4767_/Y _4945_/Y _5088_/Y _4854_/X _5401_/Y VGND VGND VPWR VPWR _5573_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_134_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6382_ _7108_/Q _6159_/X _6160_/X _7058_/Q _6381_/X VGND VGND VPWR VPWR _6382_/X
+ sky130_fd_sc_hd__a221o_1
X_3594_ _7465_/Q _5903_/A _5939_/B hold75/A _7513_/Q VGND VGND VPWR VPWR _3594_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_127_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5333_ _4688_/C _4977_/X _4981_/X _5089_/A _5224_/B VGND VGND VPWR VPWR _5471_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_142_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5264_ _4943_/A _4935_/C _4934_/C _5452_/C _5092_/A VGND VGND VPWR VPWR _5264_/Y
+ sky130_fd_sc_hd__a32oi_2
XFILLER_141_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7003_ _7512_/CLK _7003_/D fanout608/X VGND VGND VPWR VPWR _7003_/Q sky130_fd_sc_hd__dfrtp_1
X_4215_ _6965_/D _4215_/B _6854_/B _4215_/D VGND VGND VPWR VPWR _4215_/Y sky130_fd_sc_hd__nand4b_1
XFILLER_87_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5195_ _5196_/A _5195_/B _5476_/B VGND VGND VPWR VPWR _5195_/X sky130_fd_sc_hd__and3_2
X_4146_ _7613_/Q _4147_/A _4145_/Y VGND VGND VPWR VPWR _4146_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_leaf_81_csclk _7095_/CLK VGND VGND VPWR VPWR _7312_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_96_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4077_ _6927_/Q _6912_/Q _3500_/C _4076_/X VGND VGND VPWR VPWR _4077_/X sky130_fd_sc_hd__a31o_1
XFILLER_141_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4979_ _5196_/A _5043_/B _5030_/D _5229_/B VGND VGND VPWR VPWR _5472_/C sky130_fd_sc_hd__nand4_1
X_6718_ _7082_/Q _6645_/B _6536_/C _6463_/X _7225_/Q VGND VGND VPWR VPWR _6718_/X
+ sky130_fd_sc_hd__a32o_1
X_7698_ _7698_/A VGND VGND VPWR VPWR _7698_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6649_ _7616_/Q _6451_/X _6457_/X _7576_/Q _6648_/X VGND VGND VPWR VPWR _6649_/X
+ sky130_fd_sc_hd__a221o_2
Xclkbuf_leaf_34_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7432_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_145_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_49_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7545_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_115_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap429 _5011_/A VGND VGND VPWR VPWR _5585_/A1 sky130_fd_sc_hd__buf_4
XFILLER_143_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4000_ _7522_/Q _5993_/A _5939_/B _3710_/X _7071_/Q VGND VGND VPWR VPWR _4000_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_84_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5951_ hold935/X _6041_/A1 _5956_/S VGND VGND VPWR VPWR _5951_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4902_ _4902_/A _4902_/B _4902_/C VGND VGND VPWR VPWR _4904_/A sky130_fd_sc_hd__nor3_1
X_5882_ hold794/X _5999_/A1 _5884_/S VGND VGND VPWR VPWR _5882_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7621_ _7680_/CLK _7621_/D _6911_/A VGND VGND VPWR VPWR _7621_/Q sky130_fd_sc_hd__dfrtp_2
X_4833_ _4704_/A _5146_/B _5000_/C VGND VGND VPWR VPWR _4833_/X sky130_fd_sc_hd__o21a_1
XFILLER_61_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7552_ _7616_/CLK _7552_/D fanout611/X VGND VGND VPWR VPWR _7552_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_193_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4764_ _5233_/A _4763_/X _4762_/Y VGND VGND VPWR VPWR _4775_/A sky130_fd_sc_hd__a21oi_1
XFILLER_193_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6503_ _7578_/Q _6452_/X _6458_/X _7418_/Q _6502_/X VGND VGND VPWR VPWR _6503_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3715_ _5682_/A _5628_/A _5682_/B VGND VGND VPWR VPWR _3715_/X sky130_fd_sc_hd__and3_2
X_7483_ _7512_/CLK _7483_/D fanout608/X VGND VGND VPWR VPWR _7483_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_119_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4695_ _5000_/C _4590_/B _4660_/C _5027_/B _5027_/C VGND VGND VPWR VPWR _5197_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_174_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6434_ _7193_/Q _6138_/X _6152_/X _7203_/Q _6433_/X VGND VGND VPWR VPWR _6434_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3646_ _7560_/Q _3558_/X _4293_/S input69/X _3645_/X VGND VGND VPWR VPWR _3646_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_106_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6365_ _7037_/Q _6082_/Y _6364_/X VGND VGND VPWR VPWR _6365_/X sky130_fd_sc_hd__o21a_1
X_3577_ _5682_/A _3622_/A _3622_/B VGND VGND VPWR VPWR _5666_/B sky130_fd_sc_hd__and3_4
XFILLER_115_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5316_ _5316_/A _5318_/B _5316_/C VGND VGND VPWR VPWR _5316_/X sky130_fd_sc_hd__and3_1
XFILLER_0_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6296_ _7320_/Q _6082_/Y _7140_/Q VGND VGND VPWR VPWR _6296_/X sky130_fd_sc_hd__o21ba_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5247_ _5092_/A _5523_/A3 _4906_/B VGND VGND VPWR VPWR _5524_/A sky130_fd_sc_hd__a21oi_1
XFILLER_76_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold15 hold43/X VGND VGND VPWR VPWR hold44/A sky130_fd_sc_hd__buf_6
Xhold26 hold26/A VGND VGND VPWR VPWR hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A VGND VGND VPWR VPWR hold37/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold48 hold48/A VGND VGND VPWR VPWR hold48/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold59 hold59/A VGND VGND VPWR VPWR hold59/X sky130_fd_sc_hd__dlygate4sd3_1
X_5178_ _4681_/Y _5175_/Y _5176_/Y _5177_/X VGND VGND VPWR VPWR _5180_/A sky130_fd_sc_hd__o211a_1
XFILLER_56_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4129_ _4140_/B _6811_/S VGND VGND VPWR VPWR _4129_/X sky130_fd_sc_hd__and2b_1
XFILLER_28_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3500_ _6925_/Q _6912_/Q _3500_/C VGND VGND VPWR VPWR _3500_/X sky130_fd_sc_hd__and3_1
XFILLER_183_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4480_ hold539/X _4564_/A1 _4480_/S VGND VGND VPWR VPWR _4480_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold507 _4361_/X VGND VGND VPWR VPWR _7068_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 _7078_/Q VGND VGND VPWR VPWR hold518/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold529 hold529/A VGND VGND VPWR VPWR hold529/X sky130_fd_sc_hd__dlygate4sd3_1
X_3431_ hold46/A VGND VGND VPWR VPWR _3431_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6150_ _6231_/B _6416_/B _6231_/D _6159_/B VGND VGND VPWR VPWR _6150_/X sky130_fd_sc_hd__and4_2
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _5099_/Y _5100_/Y _5098_/X VGND VGND VPWR VPWR _5116_/D sky130_fd_sc_hd__o21ai_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6081_ _7624_/Q _7623_/Q _6151_/B _6392_/B VGND VGND VPWR VPWR _6081_/Y sky130_fd_sc_hd__nor4_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1207 _4237_/A1 VGND VGND VPWR VPWR hold628/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5032_ _5311_/C _5089_/A _5191_/C VGND VGND VPWR VPWR _5059_/A sky130_fd_sc_hd__and3_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1218 _6819_/A1 VGND VGND VPWR VPWR hold690/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1229 _6818_/A1 VGND VGND VPWR VPWR hold655/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6983_ _7676_/CLK _6983_/D VGND VGND VPWR VPWR _6983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5934_ _5934_/A0 _6042_/A1 _5938_/S VGND VGND VPWR VPWR _7517_/D sky130_fd_sc_hd__mux2_1
XFILLER_80_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5865_ hold498/X _6045_/A1 _5866_/S VGND VGND VPWR VPWR _5865_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7604_ _7606_/CLK _7604_/D fanout612/X VGND VGND VPWR VPWR _7604_/Q sky130_fd_sc_hd__dfrtp_1
X_4816_ _4992_/D _5146_/B _4822_/A VGND VGND VPWR VPWR _4816_/Y sky130_fd_sc_hd__nand3b_4
X_5796_ _5796_/A0 _6012_/A0 _5803_/S VGND VGND VPWR VPWR _5796_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7535_ _7584_/CLK _7535_/D fanout613/X VGND VGND VPWR VPWR _7535_/Q sky130_fd_sc_hd__dfrtp_1
X_4747_ _5186_/C _4747_/B _5595_/B VGND VGND VPWR VPWR _4748_/B sky130_fd_sc_hd__and3_1
X_7466_ _7613_/CLK _7466_/D fanout626/X VGND VGND VPWR VPWR _7466_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_147_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4678_ _4761_/A _4999_/B VGND VGND VPWR VPWR _5218_/C sky130_fd_sc_hd__nand2_1
XFILLER_162_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6417_ _7070_/Q _6231_/D _6427_/A3 _6428_/A2 _7213_/Q VGND VGND VPWR VPWR _6417_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_107_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3629_ _7408_/Q _5840_/A _6020_/A _3571_/X _7360_/Q VGND VGND VPWR VPWR _3629_/X
+ sky130_fd_sc_hd__a32o_1
X_7397_ _7445_/CLK _7397_/D fanout628/X VGND VGND VPWR VPWR _7397_/Q sky130_fd_sc_hd__dfrtp_4
X_6348_ _7170_/Q _6160_/D _6166_/C _6432_/A3 _7097_/Q VGND VGND VPWR VPWR _6348_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_88_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput105 wb_adr_i[15] VGND VGND VPWR VPWR _4585_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_6279_ _7392_/Q _6231_/D _6146_/C _6119_/X _7416_/Q VGND VGND VPWR VPWR _6279_/X
+ sky130_fd_sc_hd__a32o_1
Xinput116 wb_adr_i[25] VGND VGND VPWR VPWR input116/X sky130_fd_sc_hd__clkbuf_1
Xinput127 wb_adr_i[6] VGND VGND VPWR VPWR _5007_/A sky130_fd_sc_hd__buf_2
XFILLER_88_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput138 wb_dat_i[15] VGND VGND VPWR VPWR _6851_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput149 wb_dat_i[25] VGND VGND VPWR VPWR _6833_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_756 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3980_ _7688_/A _5682_/A _5661_/A _5669_/B _3979_/X VGND VGND VPWR VPWR _3980_/X
+ sky130_fd_sc_hd__a41o_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5650_ _5650_/A _5686_/D VGND VGND VPWR VPWR _5658_/S sky130_fd_sc_hd__nand2_4
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4601_ _5000_/C _4568_/Y _5025_/B VGND VGND VPWR VPWR _4668_/C sky130_fd_sc_hd__o21a_1
X_5581_ _5614_/C _4702_/X _5068_/C _5614_/A VGND VGND VPWR VPWR _5581_/X sky130_fd_sc_hd__o211a_1
XFILLER_191_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7320_ _7497_/CLK _7320_/D fanout607/X VGND VGND VPWR VPWR _7320_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_163_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4532_ _4532_/A0 _6864_/A1 _4534_/S VGND VGND VPWR VPWR _4532_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold304 _5685_/X VGND VGND VPWR VPWR _7297_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 _7420_/Q VGND VGND VPWR VPWR hold315/X sky130_fd_sc_hd__dlygate4sd3_1
X_7251_ _7253_/CLK _7251_/D fanout618/X VGND VGND VPWR VPWR _7251_/Q sky130_fd_sc_hd__dfrtp_4
X_4463_ _4463_/A _5686_/D VGND VGND VPWR VPWR _4468_/S sky130_fd_sc_hd__nand2_2
Xhold326 _5735_/X VGND VGND VPWR VPWR _7340_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 _7118_/Q VGND VGND VPWR VPWR hold337/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 _5996_/X VGND VGND VPWR VPWR _7572_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6202_ _7508_/Q _6136_/X _6144_/X _7540_/Q _6193_/X VGND VGND VPWR VPWR _6202_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold359 _7181_/Q VGND VGND VPWR VPWR hold359/X sky130_fd_sc_hd__dlygate4sd3_1
X_7182_ _7212_/CLK _7182_/D fanout619/X VGND VGND VPWR VPWR _7182_/Q sky130_fd_sc_hd__dfrtp_1
X_4394_ _5682_/A _5628_/A _5659_/C _6861_/C VGND VGND VPWR VPWR _4399_/S sky130_fd_sc_hd__and4_2
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6133_ _6151_/B _6392_/B _6416_/C _6158_/D VGND VGND VPWR VPWR _6133_/X sky130_fd_sc_hd__and4b_4
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6064_ _6064_/A _6064_/B _6064_/C VGND VGND VPWR VPWR _7622_/D sky130_fd_sc_hd__and3_1
Xhold1004 _4500_/X VGND VGND VPWR VPWR _7189_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1015 hold1246/X VGND VGND VPWR VPWR _4395_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1026 _7106_/Q VGND VGND VPWR VPWR _4407_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _4990_/A _5017_/B _5015_/C _5015_/D VGND VGND VPWR VPWR _5015_/Y sky130_fd_sc_hd__nand4bb_4
Xhold1037 hold1312/X VGND VGND VPWR VPWR _5880_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1048 hold1366/X VGND VGND VPWR VPWR _5997_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1059 _4347_/X VGND VGND VPWR VPWR _7056_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_54_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6966_ _7668_/CLK _6966_/D _6815_/A VGND VGND VPWR VPWR _6966_/Q sky130_fd_sc_hd__dfrtp_1
X_5917_ hold174/X _6043_/A1 _5920_/S VGND VGND VPWR VPWR _5917_/X sky130_fd_sc_hd__mux2_1
X_6897_ _6899_/A _6907_/B VGND VGND VPWR VPWR _6897_/X sky130_fd_sc_hd__and2_1
XFILLER_139_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5848_ hold914/X _6046_/A1 _5848_/S VGND VGND VPWR VPWR _5848_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5779_ _6040_/A1 hold975/X _5785_/S VGND VGND VPWR VPWR _5779_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7518_ _7518_/CLK _7518_/D fanout625/X VGND VGND VPWR VPWR _7518_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7449_ _7553_/CLK _7449_/D fanout624/X VGND VGND VPWR VPWR _7449_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_162_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold860 _4527_/X VGND VGND VPWR VPWR _7212_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold871 _7591_/Q VGND VGND VPWR VPWR hold871/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 _5810_/X VGND VGND VPWR VPWR _7407_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold893 _5817_/X VGND VGND VPWR VPWR _7413_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1560 _7646_/Q VGND VGND VPWR VPWR _6390_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1571 _7137_/Q VGND VGND VPWR VPWR _4443_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1582 _3481_/X VGND VGND VPWR VPWR _6950_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_700 _4116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1593 _7442_/Q VGND VGND VPWR VPWR _5850_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_711 _3516_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_722 _7438_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_733 _5452_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_744 _6454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6820_ _6820_/A0 _6820_/A1 _6823_/S VGND VGND VPWR VPWR _7668_/D sky130_fd_sc_hd__mux2_1
XFILLER_63_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6751_ _7063_/Q _6453_/X _6485_/X _7216_/Q _6750_/X VGND VGND VPWR VPWR _6758_/A
+ sky130_fd_sc_hd__a221o_1
X_3963_ _7483_/Q _3531_/X _3958_/X _3960_/X _3962_/X VGND VGND VPWR VPWR _3963_/Y
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_189_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5702_ _5999_/A1 hold653/X _5704_/S VGND VGND VPWR VPWR _5702_/X sky130_fd_sc_hd__mux2_1
X_6682_ _7617_/Q _6451_/X _6454_/X _7361_/Q _6681_/X VGND VGND VPWR VPWR _6682_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_188_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3894_ _7404_/Q _3545_/X _4382_/A _7088_/Q _3893_/X VGND VGND VPWR VPWR _3894_/X
+ sky130_fd_sc_hd__a221o_1
X_5633_ _5926_/A0 hold434/X _5633_/S VGND VGND VPWR VPWR _5633_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5564_ _5429_/A _5512_/C _5137_/A _5313_/C VGND VGND VPWR VPWR _5565_/B sky130_fd_sc_hd__o211a_1
XFILLER_176_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7303_ _7304_/CLK _7303_/D fanout620/X VGND VGND VPWR VPWR _7303_/Q sky130_fd_sc_hd__dfrtp_1
Xhold101 _4229_/X VGND VGND VPWR VPWR hold101/X sky130_fd_sc_hd__dlygate4sd3_1
X_4515_ _4515_/A0 _6865_/A1 _4516_/S VGND VGND VPWR VPWR _4515_/X sky130_fd_sc_hd__mux2_1
Xhold112 _5784_/X VGND VGND VPWR VPWR _7384_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold123 _7484_/Q VGND VGND VPWR VPWR hold123/X sky130_fd_sc_hd__dlygate4sd3_1
X_5495_ _5375_/B _4797_/C _5376_/B _5494_/Y VGND VGND VPWR VPWR _5495_/X sky130_fd_sc_hd__a211o_1
Xhold134 _3513_/D VGND VGND VPWR VPWR hold69/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 _7132_/Q VGND VGND VPWR VPWR hold145/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 _5686_/X VGND VGND VPWR VPWR _5688_/S sky130_fd_sc_hd__dlygate4sd3_1
X_4446_ _4037_/Y _4446_/A1 _4453_/S VGND VGND VPWR VPWR _7143_/D sky130_fd_sc_hd__mux2_1
X_7234_ _7252_/CLK _7234_/D fanout616/X VGND VGND VPWR VPWR _7234_/Q sky130_fd_sc_hd__dfrtp_1
Xhold167 _6007_/X VGND VGND VPWR VPWR _7582_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 _7547_/Q VGND VGND VPWR VPWR hold178/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 _3673_/C VGND VGND VPWR VPWR hold189/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout603 fanout633/X VGND VGND VPWR VPWR fanout603/X sky130_fd_sc_hd__buf_6
X_7165_ _7254_/CLK _7165_/D fanout617/X VGND VGND VPWR VPWR _7165_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout614 fanout615/X VGND VGND VPWR VPWR fanout614/X sky130_fd_sc_hd__buf_4
X_4377_ _4377_/A0 _6862_/A1 _4381_/S VGND VGND VPWR VPWR _4377_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout625 fanout632/X VGND VGND VPWR VPWR fanout625/X sky130_fd_sc_hd__buf_8
Xfanout636 _5015_/D VGND VGND VPWR VPWR _5014_/D sky130_fd_sc_hd__buf_12
Xfanout647 _4992_/A VGND VGND VPWR VPWR _5189_/A sky130_fd_sc_hd__buf_8
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6116_ _7386_/Q _6231_/D _6146_/C _6114_/X _7394_/Q VGND VGND VPWR VPWR _6116_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7096_ _7238_/CLK _7096_/D fanout602/X VGND VGND VPWR VPWR _7096_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6047_ _7142_/Q _7139_/Q VGND VGND VPWR VPWR _6047_/Y sky130_fd_sc_hd__nor2_1
XFILLER_100_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6949_ _4172_/B2 _6949_/D _6904_/X VGND VGND VPWR VPWR _6949_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_179_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold690 hold690/A VGND VGND VPWR VPWR hold690/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1390 _7046_/Q VGND VGND VPWR VPWR hold1390/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_530 input78/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_541 input81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_552 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_563 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_574 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_585 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_596 _6809_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput206 _3423_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[3] sky130_fd_sc_hd__buf_12
Xoutput217 _4168_/X VGND VGND VPWR VPWR mgmt_gpio_out[13] sky130_fd_sc_hd__buf_12
X_4300_ hold309/X _5935_/A1 _4303_/S VGND VGND VPWR VPWR _4300_/X sky130_fd_sc_hd__mux2_1
Xoutput228 _7705_/X VGND VGND VPWR VPWR mgmt_gpio_out[25] sky130_fd_sc_hd__buf_12
Xoutput239 _4153_/X VGND VGND VPWR VPWR mgmt_gpio_out[35] sky130_fd_sc_hd__buf_12
XFILLER_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5280_ _4969_/B _5512_/B _5452_/B _4972_/C _5375_/C VGND VGND VPWR VPWR _5280_/X
+ sky130_fd_sc_hd__a32o_1
X_4231_ _6815_/A _6963_/Q VGND VGND VPWR VPWR _4239_/S sky130_fd_sc_hd__nand2_4
XFILLER_141_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4162_ _7294_/Q _4171_/C _4171_/D _7325_/Q VGND VGND VPWR VPWR _4162_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_68_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4093_ _7257_/Q _7256_/Q _4104_/D _7258_/Q VGND VGND VPWR VPWR _4094_/S sky130_fd_sc_hd__and4bb_1
XFILLER_67_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6803_ _7095_/Q _6791_/D _6536_/C _6474_/B _7055_/Q VGND VGND VPWR VPWR _6803_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4995_ _4995_/A _5191_/C VGND VGND VPWR VPWR _4995_/Y sky130_fd_sc_hd__nand2_1
XFILLER_23_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6734_ _6734_/A _6734_/B _6734_/C _6809_/D VGND VGND VPWR VPWR _6734_/Y sky130_fd_sc_hd__nor4_1
XFILLER_51_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3946_ _3946_/A _3946_/B _3946_/C _3946_/D VGND VGND VPWR VPWR _3964_/B sky130_fd_sc_hd__nor4_4
XFILLER_192_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3877_ _7123_/Q _4559_/B _4535_/B _4463_/A _7161_/Q VGND VGND VPWR VPWR _3877_/X
+ sky130_fd_sc_hd__a32o_1
X_6665_ _7425_/Q _6458_/X _6483_/X _7393_/Q _6664_/X VGND VGND VPWR VPWR _6675_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5616_ _5616_/A _5616_/B _5616_/C _5616_/D VGND VGND VPWR VPWR _5617_/C sky130_fd_sc_hd__nor4_1
XFILLER_191_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6596_ _7414_/Q _6450_/X _6483_/X _7390_/Q _6595_/X VGND VGND VPWR VPWR _6596_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_164_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5547_ _5547_/A _5547_/B _5547_/C VGND VGND VPWR VPWR _5549_/A sky130_fd_sc_hd__and3_1
XFILLER_105_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5478_ _5614_/C _5233_/B _5068_/C _5475_/X _5477_/X VGND VGND VPWR VPWR _5478_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_144_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4429_ hold239/X _6866_/A1 _4429_/S VGND VGND VPWR VPWR _4429_/X sky130_fd_sc_hd__mux2_1
X_7217_ _7217_/CLK _7217_/D _6903_/A VGND VGND VPWR VPWR _7217_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_132_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout411 _3529_/X VGND VGND VPWR VPWR _5957_/B sky130_fd_sc_hd__buf_12
Xfanout433 _6908_/B VGND VGND VPWR VPWR _6911_/B sky130_fd_sc_hd__buf_4
X_7148_ _7672_/CLK _7148_/D VGND VGND VPWR VPWR _7148_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout444 _5595_/A VGND VGND VPWR VPWR _4747_/B sky130_fd_sc_hd__clkbuf_8
Xfanout477 _6516_/C VGND VGND VPWR VPWR _6563_/C sky130_fd_sc_hd__buf_8
XFILLER_86_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout488 _6161_/D VGND VGND VPWR VPWR _6416_/C sky130_fd_sc_hd__clkbuf_16
X_7079_ _7398_/CLK _7079_/D fanout619/X VGND VGND VPWR VPWR _7079_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout499 _4885_/Y VGND VGND VPWR VPWR _5611_/A2 sky130_fd_sc_hd__buf_4
XFILLER_73_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_360 _7006_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_371 _3514_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_382 _5659_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3800_ _7162_/Q _4463_/A _3703_/X _7114_/Q _3799_/X VGND VGND VPWR VPWR _3800_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_393 _6011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4780_ _5407_/A _5074_/A _4948_/B _4959_/C _5017_/B VGND VGND VPWR VPWR _4865_/B
+ sky130_fd_sc_hd__o2111ai_4
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3731_ _7454_/Q _5903_/A _6002_/A _3730_/X VGND VGND VPWR VPWR _3731_/X sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_0_csclk _7095_/CLK VGND VGND VPWR VPWR _7686_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_9_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6450_ _7631_/Q _6485_/B _6791_/D _6771_/C VGND VGND VPWR VPWR _6450_/X sky130_fd_sc_hd__and4_4
X_3662_ _7463_/Q _3549_/X _3561_/X _7527_/Q _3661_/X VGND VGND VPWR VPWR _3667_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5401_ _5401_/A _5401_/B VGND VGND VPWR VPWR _5401_/Y sky130_fd_sc_hd__nand2_1
XFILLER_146_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6381_ _7216_/Q _6151_/X _6157_/X _7103_/Q _6380_/X VGND VGND VPWR VPWR _6381_/X
+ sky130_fd_sc_hd__a221o_1
X_3593_ _7321_/Q _5993_/B _5682_/C _3546_/X _7537_/Q VGND VGND VPWR VPWR _3593_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_127_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5332_ _4759_/X _4976_/Y _4982_/Y _4987_/Y _5227_/B VGND VGND VPWR VPWR _5583_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_154_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5263_ _5263_/A _5263_/B _5263_/C VGND VGND VPWR VPWR _5263_/Y sky130_fd_sc_hd__nor3_1
XFILLER_142_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4214_ _4118_/B _4229_/S VGND VGND VPWR VPWR _4215_/D sky130_fd_sc_hd__nand2b_1
X_7002_ _7568_/CLK _7002_/D fanout622/X VGND VGND VPWR VPWR _7002_/Q sky130_fd_sc_hd__dfrtp_1
X_5194_ _4995_/Y _5018_/Y _5193_/Y _4648_/Y _5192_/X VGND VGND VPWR VPWR _5201_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_68_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4145_ _4147_/A _4145_/B VGND VGND VPWR VPWR _4145_/Y sky130_fd_sc_hd__nand2_2
XFILLER_28_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4076_ _4064_/X _4076_/B _4192_/B _4192_/C VGND VGND VPWR VPWR _4076_/X sky130_fd_sc_hd__and4b_1
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4978_ _5024_/C _5024_/D _4572_/X _5476_/D VGND VGND VPWR VPWR _5229_/B sky130_fd_sc_hd__a211oi_4
X_6717_ _7122_/Q _6441_/X _6481_/X _7210_/Q _6716_/X VGND VGND VPWR VPWR _6725_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_149_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3929_ _7379_/Q _5993_/B _5759_/B _3928_/X VGND VGND VPWR VPWR _3929_/X sky130_fd_sc_hd__a31o_1
XFILLER_177_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7697_ _7697_/A VGND VGND VPWR VPWR _7697_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_177_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6648_ _7592_/Q _6468_/X _6487_/X _7472_/Q _6637_/X VGND VGND VPWR VPWR _6648_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_137_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6579_ _7557_/Q _6453_/X _6482_/X _7485_/Q _6563_/X VGND VGND VPWR VPWR _6579_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_180_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5950_ hold970/X _6040_/A1 _5956_/S VGND VGND VPWR VPWR _7531_/D sky130_fd_sc_hd__mux2_1
XFILLER_46_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4901_ _4943_/A _4901_/B _4901_/C _4950_/C VGND VGND VPWR VPWR _4902_/A sky130_fd_sc_hd__and4_1
X_5881_ hold245/X _6043_/A1 _5884_/S VGND VGND VPWR VPWR _5881_/X sky130_fd_sc_hd__mux2_1
X_7620_ _7680_/CLK _7620_/D _6886_/A VGND VGND VPWR VPWR _7620_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4832_ _4599_/Y _4777_/Y _4830_/Y VGND VGND VPWR VPWR _4860_/B sky130_fd_sc_hd__o21ai_4
XANTENNA_190 _6837_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7551_ _7569_/CLK _7551_/D fanout614/X VGND VGND VPWR VPWR _7551_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_159_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4763_ _5186_/C _5595_/A _4801_/C VGND VGND VPWR VPWR _4763_/X sky130_fd_sc_hd__and3_1
X_6502_ _7506_/Q _6484_/X _6501_/X _7562_/Q _6489_/X VGND VGND VPWR VPWR _6502_/X
+ sky130_fd_sc_hd__a221o_2
X_3714_ _3714_/A _5686_/A _4535_/B VGND VGND VPWR VPWR _3714_/X sky130_fd_sc_hd__and3_2
X_7482_ _7512_/CLK _7482_/D fanout608/X VGND VGND VPWR VPWR _7482_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_146_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4694_ _5046_/A _5007_/D _5008_/C VGND VGND VPWR VPWR _4694_/Y sky130_fd_sc_hd__nand3_1
X_6433_ _7075_/Q _6359_/B _6334_/C _6159_/X _7110_/Q VGND VGND VPWR VPWR _6433_/X
+ sky130_fd_sc_hd__a32o_1
X_3645_ input41/X _4275_/S _3623_/X _3624_/X _3644_/X VGND VGND VPWR VPWR _3645_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3576_ _5661_/B _5659_/C _5680_/B VGND VGND VPWR VPWR _4291_/S sky130_fd_sc_hd__and3_2
X_6364_ _6351_/X _6355_/X _6363_/X VGND VGND VPWR VPWR _6364_/X sky130_fd_sc_hd__a21o_1
XFILLER_136_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5315_ _4568_/Y _5085_/Y _5314_/Y VGND VGND VPWR VPWR _5319_/C sky130_fd_sc_hd__o21ai_1
X_6295_ _6082_/B _6281_/X _6294_/X VGND VGND VPWR VPWR _6295_/X sky130_fd_sc_hd__a21o_1
XFILLER_170_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5246_ _5375_/C _4935_/C _5389_/B _5523_/A3 _5091_/B VGND VGND VPWR VPWR _5384_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_130_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold16 hold16/A VGND VGND VPWR VPWR hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 hold27/A VGND VGND VPWR VPWR hold27/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 hold38/A VGND VGND VPWR VPWR hold38/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold49 hold66/X VGND VGND VPWR VPWR hold49/X sky130_fd_sc_hd__dlygate4sd3_1
X_5177_ _4704_/D _4681_/Y _4709_/Y _4762_/B VGND VGND VPWR VPWR _5177_/X sky130_fd_sc_hd__o31a_1
XFILLER_56_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4128_ _7619_/Q _7620_/Q _7621_/Q _7622_/Q VGND VGND VPWR VPWR _4130_/B sky130_fd_sc_hd__nand4bb_2
XFILLER_28_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4059_ _4059_/A0 _4060_/A0 _4192_/B VGND VGND VPWR VPWR _6934_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_80_csclk _7095_/CLK VGND VGND VPWR VPWR _7307_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_51_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire450 wire452/X VGND VGND VPWR VPWR _6286_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_129_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold508 _7313_/Q VGND VGND VPWR VPWR hold508/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3430_ _7549_/Q VGND VGND VPWR VPWR _3430_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold519 _4373_/X VGND VGND VPWR VPWR _7078_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5100_ _5011_/C _4821_/Y _4960_/Y _5013_/Y VGND VGND VPWR VPWR _5100_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6080_ _6151_/B _6392_/B VGND VGND VPWR VPWR _6080_/Y sky130_fd_sc_hd__nor2_2
XFILLER_112_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _5109_/A _5040_/A _5313_/B VGND VGND VPWR VPWR _5107_/B sky130_fd_sc_hd__and3_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1208 _4234_/A1 VGND VGND VPWR VPWR hold630/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1219 _4461_/A1 VGND VGND VPWR VPWR hold706/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6982_ _7676_/CLK _6982_/D VGND VGND VPWR VPWR _6982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5933_ hold957/X _6041_/A1 _5938_/S VGND VGND VPWR VPWR _5933_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_33_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7549_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_15_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5864_ hold962/X _5999_/A1 _5866_/S VGND VGND VPWR VPWR _7455_/D sky130_fd_sc_hd__mux2_1
XFILLER_178_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7603_ _7603_/CLK _7603_/D fanout611/X VGND VGND VPWR VPWR _7603_/Q sky130_fd_sc_hd__dfstp_1
X_4815_ _4959_/C _5318_/A _4822_/A VGND VGND VPWR VPWR _5042_/A sky130_fd_sc_hd__and3b_4
XFILLER_166_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5795_ _5939_/B _5840_/A _6029_/B VGND VGND VPWR VPWR _5803_/S sky130_fd_sc_hd__and3_4
X_7534_ _7584_/CLK _7534_/D fanout613/X VGND VGND VPWR VPWR _7534_/Q sky130_fd_sc_hd__dfrtp_2
X_4746_ _4747_/B _5490_/C _5297_/A _5490_/B VGND VGND VPWR VPWR _4751_/B sky130_fd_sc_hd__nand4_1
Xclkbuf_leaf_48_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7602_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_147_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7465_ _7616_/CLK _7465_/D fanout612/X VGND VGND VPWR VPWR _7465_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_174_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4677_ _5007_/D _5025_/C _5025_/B _5007_/A VGND VGND VPWR VPWR _4677_/Y sky130_fd_sc_hd__nand4_1
X_6416_ _7626_/Q _6416_/B _6416_/C _7183_/Q VGND VGND VPWR VPWR _6416_/X sky130_fd_sc_hd__and4b_1
X_3628_ _7504_/Q _3562_/X _3572_/X _7376_/Q _3627_/X VGND VGND VPWR VPWR _3628_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7396_ _7562_/CLK _7396_/D fanout632/X VGND VGND VPWR VPWR _7396_/Q sky130_fd_sc_hd__dfrtp_1
X_6347_ _7077_/Q _6428_/B1 _6407_/A3 _7200_/Q VGND VGND VPWR VPWR _6347_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3559_ hold69/X _3559_/B _5659_/C VGND VGND VPWR VPWR hold70/A sky130_fd_sc_hd__and3_4
XFILLER_0_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6278_ _7344_/Q _6131_/C _6124_/X _7408_/Q _6277_/X VGND VGND VPWR VPWR _6278_/X
+ sky130_fd_sc_hd__a221o_1
Xinput106 wb_adr_i[16] VGND VGND VPWR VPWR _4584_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput117 wb_adr_i[26] VGND VGND VPWR VPWR _4110_/D sky130_fd_sc_hd__clkbuf_1
Xinput128 wb_adr_i[7] VGND VGND VPWR VPWR _5015_/D sky130_fd_sc_hd__buf_2
Xinput139 wb_dat_i[16] VGND VGND VPWR VPWR _6830_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_130_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5229_ _5229_/A _5229_/B VGND VGND VPWR VPWR _5472_/B sky130_fd_sc_hd__nand2_1
XFILLER_130_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_551 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_90 _4570_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4600_ _5189_/A _4822_/A _4992_/D _5008_/C VGND VGND VPWR VPWR _4684_/A sky130_fd_sc_hd__a31o_2
XFILLER_175_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5580_ _5580_/A _5580_/B _5580_/C _5580_/D VGND VGND VPWR VPWR _5580_/X sky130_fd_sc_hd__and4_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4531_ hold967/X _6863_/A1 _4534_/S VGND VGND VPWR VPWR _4531_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold305 _7363_/Q VGND VGND VPWR VPWR hold305/X sky130_fd_sc_hd__dlygate4sd3_1
X_7250_ _7679_/CLK _7250_/D fanout635/X VGND VGND VPWR VPWR hold60/A sky130_fd_sc_hd__dfrtp_2
Xhold316 _5825_/X VGND VGND VPWR VPWR _7420_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4462_ _3618_/Y _4462_/A1 _4462_/S VGND VGND VPWR VPWR _7158_/D sky130_fd_sc_hd__mux2_1
Xhold327 _7029_/Q VGND VGND VPWR VPWR hold327/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 _4421_/X VGND VGND VPWR VPWR _7118_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6201_ _7564_/Q _6153_/X _6159_/X _7436_/Q VGND VGND VPWR VPWR _6201_/X sky130_fd_sc_hd__a22o_1
Xhold349 _7088_/Q VGND VGND VPWR VPWR hold349/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4393_ _6866_/A1 hold775/X _4393_/S VGND VGND VPWR VPWR _4393_/X sky130_fd_sc_hd__mux2_1
X_7181_ _7254_/CLK _7181_/D fanout618/X VGND VGND VPWR VPWR _7181_/Q sky130_fd_sc_hd__dfstp_2
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6132_ _6158_/D _6231_/D _6145_/C VGND VGND VPWR VPWR _6132_/X sky130_fd_sc_hd__and3_4
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6063_ _7620_/Q _7621_/Q _7622_/Q _6063_/D VGND VGND VPWR VPWR _6064_/C sky130_fd_sc_hd__nand4_1
XFILLER_98_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1005 hold1427/X VGND VGND VPWR VPWR _4484_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_140_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1016 _7081_/Q VGND VGND VPWR VPWR _4377_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1027 _4407_/X VGND VGND VPWR VPWR _7106_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1038 _7214_/Q VGND VGND VPWR VPWR _4530_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5014_ _4990_/A _5017_/B _5015_/C _5014_/D VGND VGND VPWR VPWR _5249_/C sky130_fd_sc_hd__and4bb_4
Xhold1049 hold1325/X VGND VGND VPWR VPWR _6015_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6965_ _7668_/CLK _6965_/D _6815_/A VGND VGND VPWR VPWR _6965_/Q sky130_fd_sc_hd__dfrtp_4
X_5916_ _5916_/A0 _6042_/A1 _5920_/S VGND VGND VPWR VPWR _5916_/X sky130_fd_sc_hd__mux2_1
X_6896_ _6899_/A _6907_/B VGND VGND VPWR VPWR _6896_/X sky130_fd_sc_hd__and2_1
XFILLER_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5847_ hold718/X _5991_/A1 _5848_/S VGND VGND VPWR VPWR _5847_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5778_ _6003_/A1 hold427/X _5785_/S VGND VGND VPWR VPWR _5778_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7517_ _7613_/CLK _7517_/D fanout625/X VGND VGND VPWR VPWR _7517_/Q sky130_fd_sc_hd__dfrtp_4
X_4729_ _4738_/A _5614_/C _5358_/B _5490_/B VGND VGND VPWR VPWR _4729_/Y sky130_fd_sc_hd__nand4_1
XFILLER_135_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7448_ _7584_/CLK _7448_/D fanout613/X VGND VGND VPWR VPWR _7448_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_135_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold850 _5821_/X VGND VGND VPWR VPWR _7417_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold861 _7375_/Q VGND VGND VPWR VPWR hold861/X sky130_fd_sc_hd__dlygate4sd3_1
X_7379_ _7515_/CLK _7379_/D fanout621/X VGND VGND VPWR VPWR _7379_/Q sky130_fd_sc_hd__dfstp_2
Xhold872 _6017_/X VGND VGND VPWR VPWR _7591_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 _7599_/Q VGND VGND VPWR VPWR hold883/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold894 _7329_/Q VGND VGND VPWR VPWR hold894/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1550 _7263_/Q VGND VGND VPWR VPWR hold1550/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1561 _7546_/Q VGND VGND VPWR VPWR hold466/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1572 _7586_/Q VGND VGND VPWR VPWR hold1572/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1583 _7040_/Q VGND VGND VPWR VPWR hold228/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1594 _7136_/Q VGND VGND VPWR VPWR _4442_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_701 _4116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_712 _5666_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_723 _4196_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_734 _5666_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_745 _6454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6750_ _7221_/Q _6479_/X _6486_/X _7103_/Q VGND VGND VPWR VPWR _6750_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3962_ _7499_/Q _3562_/X _4388_/A _7092_/Q _3961_/X VGND VGND VPWR VPWR _3962_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5701_ _6043_/A1 hold147/X _5704_/S VGND VGND VPWR VPWR _5701_/X sky130_fd_sc_hd__mux2_1
X_6681_ _7513_/Q _6791_/D _6536_/C _6463_/X _7401_/Q VGND VGND VPWR VPWR _6681_/X
+ sky130_fd_sc_hd__a32o_1
X_3893_ _7348_/Q _5741_/A _5777_/A _7380_/Q _3892_/X VGND VGND VPWR VPWR _3893_/X
+ sky130_fd_sc_hd__a221o_1
X_5632_ _6865_/A1 hold985/X _5633_/S VGND VGND VPWR VPWR _5632_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5563_ _5625_/C _5626_/D VGND VGND VPWR VPWR _5567_/A sky130_fd_sc_hd__and2b_1
X_7302_ _7586_/CLK _7302_/D fanout625/X VGND VGND VPWR VPWR _7712_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_191_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4514_ hold535/X _5789_/A1 _4516_/S VGND VGND VPWR VPWR _4514_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold102 hold102/A VGND VGND VPWR VPWR hold102/X sky130_fd_sc_hd__buf_8
Xhold113 _7282_/Q VGND VGND VPWR VPWR hold113/X sky130_fd_sc_hd__dlygate4sd3_1
X_5494_ _5552_/A _5552_/B _5494_/C VGND VGND VPWR VPWR _5494_/Y sky130_fd_sc_hd__nand3_1
Xhold124 _5897_/X VGND VGND VPWR VPWR _7484_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold135 _4340_/Y VGND VGND VPWR VPWR _4345_/S sky130_fd_sc_hd__dlygate4sd3_1
X_7233_ _7233_/CLK _7233_/D fanout599/X VGND VGND VPWR VPWR _7233_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_105_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold146 _4438_/X VGND VGND VPWR VPWR _7132_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4445_ _6966_/Q _6815_/A VGND VGND VPWR VPWR _4453_/S sky130_fd_sc_hd__nand2_4
XFILLER_172_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold157 _5688_/X VGND VGND VPWR VPWR _7299_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 _7478_/Q VGND VGND VPWR VPWR hold168/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold179 _5968_/X VGND VGND VPWR VPWR _7547_/D sky130_fd_sc_hd__dlygate4sd3_1
Xfanout604 fanout606/X VGND VGND VPWR VPWR fanout604/X sky130_fd_sc_hd__buf_6
X_7164_ _7254_/CLK _7164_/D fanout617/X VGND VGND VPWR VPWR _7164_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_144_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout615 fanout633/X VGND VGND VPWR VPWR fanout615/X sky130_fd_sc_hd__buf_8
X_4376_ _6861_/A _5680_/A _6861_/C VGND VGND VPWR VPWR _4381_/S sky130_fd_sc_hd__and3_4
Xfanout626 fanout627/X VGND VGND VPWR VPWR fanout626/X sky130_fd_sc_hd__buf_6
Xfanout637 _5007_/A VGND VGND VPWR VPWR _4990_/A sky130_fd_sc_hd__buf_12
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6115_ _6151_/B _6231_/D _6126_/D VGND VGND VPWR VPWR _6115_/X sky130_fd_sc_hd__and3_4
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7095_ _7095_/CLK _7095_/D fanout599/X VGND VGND VPWR VPWR _7095_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ hold902/X _6046_/A1 _6046_/S VGND VGND VPWR VPWR _6046_/X sky130_fd_sc_hd__mux2_1
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6948_ _4172_/B2 _6948_/D _6903_/X VGND VGND VPWR VPWR _6948_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_41_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6879_ _6891_/A _6908_/B VGND VGND VPWR VPWR _6879_/X sky130_fd_sc_hd__and2_1
XFILLER_22_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold680 _7432_/Q VGND VGND VPWR VPWR hold680/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold691 hold691/A VGND VGND VPWR VPWR wb_dat_o[27] sky130_fd_sc_hd__buf_12
XFILLER_89_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1380 _5727_/X VGND VGND VPWR VPWR _7333_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1391 _7672_/Q VGND VGND VPWR VPWR hold14/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_520 _4195_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_531 input78/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_542 input81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_553 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_564 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_575 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_586 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_597 _6809_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput207 _3455_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[4] sky130_fd_sc_hd__buf_12
XFILLER_154_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput218 _7696_/X VGND VGND VPWR VPWR mgmt_gpio_out[16] sky130_fd_sc_hd__buf_12
Xoutput229 _7706_/X VGND VGND VPWR VPWR mgmt_gpio_out[26] sky130_fd_sc_hd__buf_12
XFILLER_175_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4230_ hold615/X _6028_/A1 _4230_/S VGND VGND VPWR VPWR _4230_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4161_ _7004_/Q input3/X input1/X VGND VGND VPWR VPWR _4161_/X sky130_fd_sc_hd__mux2_4
XFILLER_68_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4092_ _6922_/Q _4097_/A0 _4092_/S VGND VGND VPWR VPWR _4092_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6802_ _7120_/Q _6459_/X _6479_/X _7223_/Q _6801_/X VGND VGND VPWR VPWR _6809_/A
+ sky130_fd_sc_hd__a221o_1
X_4994_ _5189_/D _5146_/B _5311_/C VGND VGND VPWR VPWR _4994_/X sky130_fd_sc_hd__and3_2
X_6733_ _7117_/Q _6459_/X _6730_/X _6732_/X VGND VGND VPWR VPWR _6734_/C sky130_fd_sc_hd__a211o_1
X_3945_ _7419_/Q _3602_/X _3942_/X _3943_/X _3944_/X VGND VGND VPWR VPWR _3946_/D
+ sky130_fd_sc_hd__a2111o_1
X_6664_ _7585_/Q _6452_/X _6453_/X _7561_/Q _6663_/X VGND VGND VPWR VPWR _6664_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3876_ _7263_/Q _5939_/B _5678_/C _3710_/X _7073_/Q VGND VGND VPWR VPWR _3876_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_176_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5615_ _5614_/A _4702_/X _5092_/B _5614_/X VGND VGND VPWR VPWR _5616_/D sky130_fd_sc_hd__a31o_1
X_6595_ _7422_/Q _6458_/X _6469_/X _7334_/Q _6594_/X VGND VGND VPWR VPWR _6595_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_192_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5546_ _4743_/C _5358_/B _5595_/C _5545_/X _5162_/B VGND VGND VPWR VPWR _5547_/A
+ sky130_fd_sc_hd__a311oi_1
XFILLER_191_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5477_ _5068_/A _5233_/B _5476_/C _5077_/X _5233_/X VGND VGND VPWR VPWR _5477_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_160_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7216_ _7686_/CLK _7216_/D _6891_/A VGND VGND VPWR VPWR _7216_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_105_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4428_ hold717/X _5673_/A1 _4429_/S VGND VGND VPWR VPWR _7124_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_2_3__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _4172_/B2
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_120_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout434 _6908_/B VGND VGND VPWR VPWR _6907_/B sky130_fd_sc_hd__buf_4
X_7147_ _7668_/CLK _7147_/D VGND VGND VPWR VPWR _7147_/Q sky130_fd_sc_hd__dfxtp_2
Xfanout445 _5595_/A VGND VGND VPWR VPWR _4738_/A sky130_fd_sc_hd__buf_2
X_4359_ _6012_/A0 _4359_/A1 _4363_/S VGND VGND VPWR VPWR _4359_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout467 _6771_/B VGND VGND VPWR VPWR _6694_/B sky130_fd_sc_hd__buf_12
Xfanout478 _6487_/A VGND VGND VPWR VPWR _6720_/C sky130_fd_sc_hd__clkbuf_16
X_7078_ _7212_/CLK _7078_/D fanout627/X VGND VGND VPWR VPWR _7078_/Q sky130_fd_sc_hd__dfstp_1
Xfanout489 _6067_/X VGND VGND VPWR VPWR _6231_/D sky130_fd_sc_hd__buf_8
XFILLER_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6029_ _6029_/A _6029_/B VGND VGND VPWR VPWR _6037_/S sky130_fd_sc_hd__nand2_8
XFILLER_39_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_350 hold80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_361 _7269_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_372 _3514_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_383 _3543_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_394 _3637_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3730_ _7478_/Q _5903_/A _5957_/B _3560_/X _6976_/Q VGND VGND VPWR VPWR _3730_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_41_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3661_ _7479_/Q _5903_/A _5957_/B _5650_/A _7277_/Q VGND VGND VPWR VPWR _3661_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_158_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5400_ _5375_/C _4951_/A _5389_/D _4943_/B VGND VGND VPWR VPWR _5400_/X sky130_fd_sc_hd__o31a_1
X_6380_ _7128_/Q _6359_/B _6131_/C _6153_/X _7206_/Q VGND VGND VPWR VPWR _6380_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3592_ _7609_/Q _6029_/A _3589_/X _3590_/X _3591_/X VGND VGND VPWR VPWR _3592_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_161_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5331_ _5313_/C _4985_/B _5068_/C _5195_/X _5330_/X VGND VGND VPWR VPWR _5472_/A
+ sky130_fd_sc_hd__a221oi_1
XFILLER_127_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5262_ _5375_/C _5389_/B _5389_/C _5290_/A2 _5095_/C VGND VGND VPWR VPWR _5262_/X
+ sky130_fd_sc_hd__a32o_1
X_7001_ _7512_/CLK _7001_/D fanout608/X VGND VGND VPWR VPWR _7001_/Q sky130_fd_sc_hd__dfrtp_1
X_4213_ _6967_/Q _6858_/C VGND VGND VPWR VPWR _6829_/D sky130_fd_sc_hd__nand2b_2
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5193_ _5197_/B _5614_/D VGND VGND VPWR VPWR _5193_/Y sky130_fd_sc_hd__nand2_1
X_4144_ _7304_/Q input89/X _4147_/A VGND VGND VPWR VPWR _4144_/X sky130_fd_sc_hd__mux2_2
XFILLER_68_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4075_ _6927_/Q hold94/A _6925_/Q hold21/A _6928_/Q VGND VGND VPWR VPWR _4076_/B
+ sky130_fd_sc_hd__a41o_1
XFILLER_95_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_671 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_4_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_4_0_csclk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_34_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4977_ _5046_/A _5614_/A _5043_/B VGND VGND VPWR VPWR _4977_/X sky130_fd_sc_hd__and3_1
X_6716_ _7235_/Q _6807_/A2 _6483_/X _7067_/Q VGND VGND VPWR VPWR _6716_/X sky130_fd_sc_hd__a22o_1
X_3928_ _7117_/Q _3550_/B _5680_/A _3552_/X _7387_/Q VGND VGND VPWR VPWR _3928_/X
+ sky130_fd_sc_hd__a32o_1
X_7696_ _7696_/A VGND VGND VPWR VPWR _7696_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6647_ _7528_/Q _6447_/X _6474_/C _7376_/Q _6646_/X VGND VGND VPWR VPWR _6647_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_137_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3859_ _7211_/Q hold70/A _4487_/B _3585_/X _7332_/Q VGND VGND VPWR VPWR _3859_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_164_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6578_ _7445_/Q _6460_/X _6575_/X _6577_/X VGND VGND VPWR VPWR _6578_/X sky130_fd_sc_hd__a211o_1
XFILLER_192_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5529_ _5407_/C _4937_/Y _5270_/X _5274_/X _5573_/C VGND VGND VPWR VPWR _5530_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_132_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_663 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4900_ _4900_/A _4900_/B _4900_/C _4900_/D VGND VGND VPWR VPWR _4902_/B sky130_fd_sc_hd__nand4_1
XFILLER_92_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5880_ _5880_/A0 _6042_/A1 _5884_/S VGND VGND VPWR VPWR _7469_/D sky130_fd_sc_hd__mux2_1
X_4831_ _4704_/A _4599_/Y _5146_/B _4830_/Y VGND VGND VPWR VPWR _4892_/B sky130_fd_sc_hd__o31a_1
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_180 _6834_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_191 _6837_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7550_ _7614_/CLK _7550_/D fanout605/X VGND VGND VPWR VPWR _7550_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4762_ _4762_/A _4762_/B _4762_/C VGND VGND VPWR VPWR _4762_/Y sky130_fd_sc_hd__nand3_1
X_6501_ _7631_/Q _7630_/Q _6720_/C _6563_/C VGND VGND VPWR VPWR _6501_/X sky130_fd_sc_hd__and4_4
X_3713_ _3713_/A _5628_/A _5659_/C VGND VGND VPWR VPWR _3713_/X sky130_fd_sc_hd__and3_4
X_7481_ _7609_/CLK _7481_/D fanout614/X VGND VGND VPWR VPWR _7481_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_147_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4693_ _5000_/C _4836_/A _4660_/C _5014_/D VGND VGND VPWR VPWR _4693_/Y sky130_fd_sc_hd__o31ai_2
XFILLER_146_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6432_ _7065_/Q _6359_/B _6432_/A3 _6431_/X VGND VGND VPWR VPWR _6432_/X sky130_fd_sc_hd__a31o_1
X_3644_ input32/X _5669_/B _4529_/B _3643_/X VGND VGND VPWR VPWR _3644_/X sky130_fd_sc_hd__a31o_1
XFILLER_134_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6363_ _6363_/A1 _6359_/Y _6360_/X _6362_/X _6358_/X VGND VGND VPWR VPWR _6363_/X
+ sky130_fd_sc_hd__a2111o_1
X_3575_ _5661_/A _5628_/A _5661_/B VGND VGND VPWR VPWR _5849_/A sky130_fd_sc_hd__and3_4
XFILLER_114_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5314_ _5314_/A _5314_/B _5314_/C _5565_/A VGND VGND VPWR VPWR _5314_/Y sky130_fd_sc_hd__nor4_1
XFILLER_161_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6294_ _6284_/X _6309_/B _6283_/X _6285_/X _6293_/X VGND VGND VPWR VPWR _6294_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_170_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5245_ _4943_/A _4935_/C _5389_/B _5092_/A _5110_/C VGND VGND VPWR VPWR _5245_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_114_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold17 hold17/A VGND VGND VPWR VPWR hold17/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 hold28/A VGND VGND VPWR VPWR hold28/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 hold39/A VGND VGND VPWR VPWR hold39/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5176_ _5153_/C _4748_/B _5174_/X _5173_/X VGND VGND VPWR VPWR _5176_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_69_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4127_ _6791_/B _6694_/B VGND VGND VPWR VPWR _4127_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4058_ hold1/A _4059_/A0 _4192_/B VGND VGND VPWR VPWR _6935_/D sky130_fd_sc_hd__mux2_1
XFILLER_37_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7679_ _7679_/CLK _7679_/D fanout635/X VGND VGND VPWR VPWR _7679_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_138_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire440 _4791_/Y VGND VGND VPWR VPWR _4901_/B sky130_fd_sc_hd__buf_2
XFILLER_144_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold509 _5704_/X VGND VGND VPWR VPWR _7313_/D sky130_fd_sc_hd__dlygate4sd3_1
Xwire484 _6081_/Y VGND VGND VPWR VPWR wire484/X sky130_fd_sc_hd__clkbuf_2
Xwire495 _4948_/Y VGND VGND VPWR VPWR _5130_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_124_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5030_ _5061_/A _5197_/A _5311_/A _5030_/D VGND VGND VPWR VPWR _5030_/Y sky130_fd_sc_hd__nand4_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1209 _4451_/A1 VGND VGND VPWR VPWR hold642/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_65_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6981_ _7668_/CLK _6981_/D VGND VGND VPWR VPWR _6981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5932_ hold982/X _6040_/A1 _5938_/S VGND VGND VPWR VPWR _7515_/D sky130_fd_sc_hd__mux2_1
XFILLER_53_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5863_ hold251/X _6043_/A1 _5866_/S VGND VGND VPWR VPWR _5863_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7602_ _7602_/CLK _7602_/D fanout615/X VGND VGND VPWR VPWR _7602_/Q sky130_fd_sc_hd__dfstp_1
X_4814_ _4814_/A _4814_/B _4814_/C VGND VGND VPWR VPWR _4827_/A sky130_fd_sc_hd__nor3_1
X_5794_ hold867/X _6046_/A1 _5794_/S VGND VGND VPWR VPWR _5794_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7533_ _7549_/CLK _7533_/D fanout629/X VGND VGND VPWR VPWR _7533_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_21_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4745_ _4617_/X _4619_/Y _4622_/Y _4744_/Y VGND VGND VPWR VPWR _4751_/A sky130_fd_sc_hd__o31a_1
XFILLER_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7464_ _7616_/CLK _7464_/D fanout610/X VGND VGND VPWR VPWR _7464_/Q sky130_fd_sc_hd__dfrtp_1
X_4676_ _5614_/B _5025_/B _5025_/C VGND VGND VPWR VPWR _4999_/B sky130_fd_sc_hd__and3_1
XFILLER_107_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6415_ _6414_/X _6438_/A1 _6812_/S VGND VGND VPWR VPWR _6415_/X sky130_fd_sc_hd__mux2_1
X_3627_ _7336_/Q _5939_/B _5759_/B _3625_/X VGND VGND VPWR VPWR _3627_/X sky130_fd_sc_hd__a31o_1
X_7395_ _7562_/CLK _7395_/D fanout632/X VGND VGND VPWR VPWR _7395_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_134_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6346_ _7225_/Q _6334_/C _6170_/C _7047_/Q _6345_/X VGND VGND VPWR VPWR _6346_/X
+ sky130_fd_sc_hd__a221o_1
X_3558_ _5984_/A _5682_/A _5661_/A VGND VGND VPWR VPWR _3558_/X sky130_fd_sc_hd__and3_2
XFILLER_88_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6277_ _7400_/Q _6166_/B _6146_/C _6309_/C _7336_/Q VGND VGND VPWR VPWR _6277_/X
+ sky130_fd_sc_hd__a32o_1
X_3489_ hold33/X _3488_/X _4229_/S VGND VGND VPWR VPWR hold34/A sky130_fd_sc_hd__o21ba_2
Xinput107 wb_adr_i[17] VGND VGND VPWR VPWR _4584_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput118 wb_adr_i[27] VGND VGND VPWR VPWR input118/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5228_ _5614_/A _5313_/C _5042_/A _5068_/C _5195_/X VGND VGND VPWR VPWR _5230_/C
+ sky130_fd_sc_hd__a32oi_1
Xinput129 wb_adr_i[8] VGND VGND VPWR VPWR _4586_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5159_ _5186_/C _5358_/A _5181_/C _5156_/Y _5158_/X VGND VGND VPWR VPWR _5159_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_57_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_80 _3966_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_91 _5203_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4530_ _4530_/A0 _6862_/A1 _4534_/S VGND VGND VPWR VPWR _4530_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4461_ _3655_/Y _4461_/A1 _4462_/S VGND VGND VPWR VPWR _7157_/D sky130_fd_sc_hd__mux2_1
Xhold306 _5761_/X VGND VGND VPWR VPWR _7363_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold317 _7396_/Q VGND VGND VPWR VPWR hold317/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 _4315_/X VGND VGND VPWR VPWR _7029_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6200_ _7460_/Q _6145_/X _6158_/X _7492_/Q _6199_/X VGND VGND VPWR VPWR _6200_/X
+ sky130_fd_sc_hd__a221o_1
Xhold339 _7563_/Q VGND VGND VPWR VPWR hold339/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7180_ _7254_/CLK _7180_/D fanout617/X VGND VGND VPWR VPWR _7180_/Q sky130_fd_sc_hd__dfrtp_4
X_4392_ _5673_/A1 hold688/X _4393_/S VGND VGND VPWR VPWR _4392_/X sky130_fd_sc_hd__mux2_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6131_ _7466_/Q _6131_/B _6131_/C VGND VGND VPWR VPWR _6131_/X sky130_fd_sc_hd__and3_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _7620_/Q _7621_/Q _6063_/D _7622_/Q VGND VGND VPWR VPWR _6064_/B sky130_fd_sc_hd__a31o_1
XFILLER_85_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1006 _7161_/Q VGND VGND VPWR VPWR _4466_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1017 _4377_/X VGND VGND VPWR VPWR _7081_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _5017_/A _5094_/D VGND VGND VPWR VPWR _5013_/Y sky130_fd_sc_hd__nand2_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1028 hold1345/X VGND VGND VPWR VPWR _5754_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1039 _4530_/X VGND VGND VPWR VPWR _7214_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6964_ _7680_/CLK _6964_/D _6815_/A VGND VGND VPWR VPWR _6964_/Q sky130_fd_sc_hd__dfrtp_1
X_5915_ hold765/X _6041_/A1 _5920_/S VGND VGND VPWR VPWR _5915_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6895_ _6899_/A _6907_/B VGND VGND VPWR VPWR _6895_/X sky130_fd_sc_hd__and2_1
XFILLER_22_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5846_ hold837/X _6044_/A1 _5848_/S VGND VGND VPWR VPWR _5846_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5777_ _5777_/A _6029_/B VGND VGND VPWR VPWR _5785_/S sky130_fd_sc_hd__nand2_8
XFILLER_166_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4728_ _5153_/A _5358_/B VGND VGND VPWR VPWR _4728_/Y sky130_fd_sc_hd__nand2_1
X_7516_ _7558_/CLK _7516_/D fanout606/X VGND VGND VPWR VPWR _7516_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_147_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7447_ _7569_/CLK _7447_/D fanout613/X VGND VGND VPWR VPWR _7447_/Q sky130_fd_sc_hd__dfrtp_1
X_4659_ _4599_/Y _4631_/Y _4990_/A VGND VGND VPWR VPWR _4688_/B sky130_fd_sc_hd__o21bai_2
XFILLER_174_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold840 _5945_/X VGND VGND VPWR VPWR _7527_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7378_ _7518_/CLK _7378_/D fanout625/X VGND VGND VPWR VPWR _7378_/Q sky130_fd_sc_hd__dfstp_1
Xhold851 _7553_/Q VGND VGND VPWR VPWR hold851/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold862 _5774_/X VGND VGND VPWR VPWR _7375_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 _7409_/Q VGND VGND VPWR VPWR hold873/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap581 _4995_/A VGND VGND VPWR VPWR _5297_/C sky130_fd_sc_hd__clkbuf_2
X_6329_ _7116_/Q _6132_/X _6160_/X _7056_/Q _6328_/X VGND VGND VPWR VPWR _6329_/X
+ sky130_fd_sc_hd__a221o_1
Xhold884 _6026_/X VGND VGND VPWR VPWR _7599_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold895 _5722_/X VGND VGND VPWR VPWR _7329_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1540 _7241_/Q VGND VGND VPWR VPWR hold1540/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1551 _5640_/X VGND VGND VPWR VPWR _7263_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1562 _7466_/Q VGND VGND VPWR VPWR hold460/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1573 _7063_/Q VGND VGND VPWR VPWR hold1573/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1584 _7643_/Q VGND VGND VPWR VPWR _6320_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_702 _4116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1595 _7073_/Q VGND VGND VPWR VPWR hold1595/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_713 _6011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_724 _4196_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_735 _5666_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_746 _6809_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_32_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7597_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_164_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_47_csclk _7352_/CLK VGND VGND VPWR VPWR _7566_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_82_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3961_ _7185_/Q _4547_/A _5680_/A _3905_/X _7260_/Q VGND VGND VPWR VPWR _3961_/X
+ sky130_fd_sc_hd__a32o_1
X_5700_ hold9/X _5700_/A1 _5704_/S VGND VGND VPWR VPWR hold10/A sky130_fd_sc_hd__mux2_1
XFILLER_16_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6680_ _7593_/Q _6468_/X _6471_/X _7329_/Q VGND VGND VPWR VPWR _6680_/X sky130_fd_sc_hd__a22o_1
X_3892_ _7372_/Q _5984_/B _5759_/B _3567_/X _7340_/Q VGND VGND VPWR VPWR _3892_/X
+ sky130_fd_sc_hd__a32o_1
X_5631_ _5789_/A1 hold397/X _5633_/S VGND VGND VPWR VPWR _5631_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5562_ _5417_/X _4998_/Y _5288_/X _5561_/X _5414_/X VGND VGND VPWR VPWR _5626_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_129_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7301_ _7305_/CLK _7301_/D fanout620/X VGND VGND VPWR VPWR _7301_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_191_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4513_ hold446/X _5761_/A1 _4516_/S VGND VGND VPWR VPWR _4513_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold103 _4312_/X VGND VGND VPWR VPWR _7027_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5493_ _5493_/A _5493_/B _5493_/C VGND VGND VPWR VPWR _5494_/C sky130_fd_sc_hd__nor3_1
XFILLER_7_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold114 _5663_/X VGND VGND VPWR VPWR _7282_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 _7711_/A VGND VGND VPWR VPWR hold125/X sky130_fd_sc_hd__dlygate4sd3_1
X_7232_ _7233_/CLK _7232_/D fanout599/X VGND VGND VPWR VPWR _7232_/Q sky130_fd_sc_hd__dfrtp_4
Xhold136 hold136/A VGND VGND VPWR VPWR _7052_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4444_ _6028_/A1 hold514/X _4444_/S VGND VGND VPWR VPWR _4444_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold147 _7310_/Q VGND VGND VPWR VPWR hold147/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 _7483_/Q VGND VGND VPWR VPWR hold158/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold169 _5890_/X VGND VGND VPWR VPWR _7478_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7163_ _7215_/CLK _7163_/D _6903_/A VGND VGND VPWR VPWR _7163_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_125_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4375_ hold570/X _5926_/A0 _4375_/S VGND VGND VPWR VPWR _4375_/X sky130_fd_sc_hd__mux2_1
Xfanout605 fanout606/X VGND VGND VPWR VPWR fanout605/X sky130_fd_sc_hd__buf_8
Xfanout616 fanout618/X VGND VGND VPWR VPWR fanout616/X sky130_fd_sc_hd__buf_8
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6114_ _6151_/B _6166_/B _6126_/D VGND VGND VPWR VPWR _6114_/X sky130_fd_sc_hd__and3_4
Xfanout627 fanout632/X VGND VGND VPWR VPWR fanout627/X sky130_fd_sc_hd__buf_8
Xfanout638 _5017_/A VGND VGND VPWR VPWR _5015_/C sky130_fd_sc_hd__buf_12
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7094_ _7238_/CLK _7094_/D fanout602/X VGND VGND VPWR VPWR _7094_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6045_ hold479/X _6045_/A1 _6046_/S VGND VGND VPWR VPWR _6045_/X sky130_fd_sc_hd__mux2_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6947_ _4172_/B2 _6947_/D _6902_/X VGND VGND VPWR VPWR _6947_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_81_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6878_ _6911_/A _6911_/B VGND VGND VPWR VPWR _6878_/X sky130_fd_sc_hd__and2_1
XFILLER_22_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5829_ hold78/X hold50/X _5830_/S VGND VGND VPWR VPWR _5829_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold670 _4354_/X VGND VGND VPWR VPWR _7062_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold681 _5838_/X VGND VGND VPWR VPWR _7432_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 _7373_/Q VGND VGND VPWR VPWR hold692/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1370 _7517_/Q VGND VGND VPWR VPWR hold1370/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1381 hold42/A VGND VGND VPWR VPWR _4221_/S sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1392 _5859_/X VGND VGND VPWR VPWR _7450_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_510 _7714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_521 _4195_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_532 input81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_543 input81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_588 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_554 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_565 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_576 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_587 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_598 _4505_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput208 _3454_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[5] sky130_fd_sc_hd__buf_12
XFILLER_126_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput219 _7697_/X VGND VGND VPWR VPWR mgmt_gpio_out[17] sky130_fd_sc_hd__buf_12
XFILLER_5_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4160_ _4159_/X _4191_/B _6951_/Q VGND VGND VPWR VPWR _4160_/X sky130_fd_sc_hd__mux2_4
XFILLER_110_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4091_ _7258_/Q _7257_/Q _7256_/Q _4104_/D VGND VGND VPWR VPWR _4092_/S sky130_fd_sc_hd__and4_1
XFILLER_68_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6801_ _7110_/Q _6099_/B _6694_/C _6447_/X _7075_/Q VGND VGND VPWR VPWR _6801_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_91_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4993_ _5189_/D _5146_/B VGND VGND VPWR VPWR _4993_/Y sky130_fd_sc_hd__nand2_4
XFILLER_51_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6732_ _7077_/Q _6450_/X _6457_/X _7195_/Q _6731_/X VGND VGND VPWR VPWR _6732_/X
+ sky130_fd_sc_hd__a221o_1
X_3944_ _7077_/Q _5628_/A _4487_/A _4293_/S input47/X VGND VGND VPWR VPWR _3944_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_32_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6663_ _7569_/Q _6099_/B _6720_/D _6456_/X _7609_/Q VGND VGND VPWR VPWR _6663_/X
+ sky130_fd_sc_hd__a32o_1
X_3875_ _7532_/Q _5984_/A _6020_/A _3874_/X VGND VGND VPWR VPWR _3875_/X sky130_fd_sc_hd__a31o_1
XFILLER_176_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5614_ _5614_/A _5614_/B _5614_/C _5614_/D VGND VGND VPWR VPWR _5614_/X sky130_fd_sc_hd__and4_1
XFILLER_191_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6594_ _7518_/Q _6455_/C _6562_/C _6454_/X _7358_/Q VGND VGND VPWR VPWR _6594_/X
+ sky130_fd_sc_hd__a32o_1
X_5545_ _5476_/A _5375_/C _5358_/B _5358_/A VGND VGND VPWR VPWR _5545_/X sky130_fd_sc_hd__o211a_1
XFILLER_191_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_0_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR _7095_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_117_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5476_ _5476_/A _5476_/B _5476_/C _5476_/D VGND VGND VPWR VPWR _5476_/Y sky130_fd_sc_hd__nand4_1
X_4427_ _4427_/A0 _6864_/A1 _4429_/S VGND VGND VPWR VPWR _4427_/X sky130_fd_sc_hd__mux2_1
X_7215_ _7215_/CLK _7215_/D _6907_/A VGND VGND VPWR VPWR _7215_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout413 _5723_/A VGND VGND VPWR VPWR _5939_/B sky130_fd_sc_hd__buf_12
X_7146_ _7672_/CLK _7146_/D VGND VGND VPWR VPWR _7146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4358_ _4358_/A _6861_/C VGND VGND VPWR VPWR _4363_/S sky130_fd_sc_hd__nand2_2
Xfanout435 _3472_/Y VGND VGND VPWR VPWR _6908_/B sky130_fd_sc_hd__buf_2
Xfanout446 _4615_/Y VGND VGND VPWR VPWR _5595_/A sky130_fd_sc_hd__buf_4
Xfanout457 _6112_/X VGND VGND VPWR VPWR _6432_/A3 sky130_fd_sc_hd__buf_12
Xfanout468 _6446_/X VGND VGND VPWR VPWR _6536_/C sky130_fd_sc_hd__buf_8
X_7077_ _7212_/CLK _7077_/D fanout619/X VGND VGND VPWR VPWR _7077_/Q sky130_fd_sc_hd__dfrtp_4
X_4289_ hold653/X _5999_/A1 _4293_/S VGND VGND VPWR VPWR _4289_/X sky130_fd_sc_hd__mux2_1
Xfanout479 _6455_/C VGND VGND VPWR VPWR _6645_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6028_ hold602/X _6028_/A1 _6028_/S VGND VGND VPWR VPWR _6028_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_340 _6003_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_351 hold81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_362 _4347_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_373 _3550_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_384 _5813_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_395 _3667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3660_ _7455_/Q _6861_/A _6002_/A _3562_/X _7503_/Q VGND VGND VPWR VPWR _3667_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_118_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3591_ _7617_/Q hold24/A _4481_/A _3558_/X _7561_/Q VGND VGND VPWR VPWR _3591_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_186_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5330_ _5476_/A _5476_/C _5229_/B _4981_/X _5313_/C VGND VGND VPWR VPWR _5330_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_182_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5261_ _4953_/B _5429_/D _5429_/A _5261_/D VGND VGND VPWR VPWR _5261_/Y sky130_fd_sc_hd__nand4b_1
XFILLER_141_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7000_ _7553_/CLK _7000_/D fanout622/X VGND VGND VPWR VPWR _7695_/A sky130_fd_sc_hd__dfrtp_1
X_4212_ _6967_/Q _6969_/Q _6971_/Q _6970_/Q VGND VGND VPWR VPWR _6854_/B sky130_fd_sc_hd__nor4_2
X_5192_ _4570_/Y _4953_/C _4821_/Y _5011_/A VGND VGND VPWR VPWR _5192_/X sky130_fd_sc_hd__a211o_1
XFILLER_141_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4143_ _7305_/Q input91/X _4147_/A VGND VGND VPWR VPWR _4143_/X sky130_fd_sc_hd__mux2_2
XFILLER_95_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4074_ _4074_/A1 _3508_/S _4043_/Y _4073_/X VGND VGND VPWR VPWR _6929_/D sky130_fd_sc_hd__a31o_1
XFILLER_95_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4976_ _5297_/A _5061_/A VGND VGND VPWR VPWR _4976_/Y sky130_fd_sc_hd__nand2_1
X_6715_ _7200_/Q _6445_/X _6487_/X _7127_/Q _6714_/X VGND VGND VPWR VPWR _6725_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_177_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3927_ _6973_/Q _3573_/C _4505_/B _3925_/X _3926_/X VGND VGND VPWR VPWR _3927_/X
+ sky130_fd_sc_hd__a311o_1
X_7695_ _7695_/A VGND VGND VPWR VPWR _7695_/X sky130_fd_sc_hd__clkbuf_1
X_6646_ _7512_/Q _6484_/X _6645_/X _6445_/C _6639_/X VGND VGND VPWR VPWR _6646_/X
+ sky130_fd_sc_hd__a221o_1
X_3858_ _7181_/Q _4487_/A _4511_/C _3857_/X VGND VGND VPWR VPWR _3858_/X sky130_fd_sc_hd__a31o_1
XFILLER_177_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3789_ _7212_/Q _4505_/B _4511_/C _4499_/A _7192_/Q VGND VGND VPWR VPWR _3789_/X
+ sky130_fd_sc_hd__a32o_1
X_6577_ _7429_/Q _6444_/X _6459_/X _7453_/Q _6576_/X VGND VGND VPWR VPWR _6577_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_152_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5528_ _5407_/C _4854_/X _5270_/X _5570_/D _5273_/C VGND VGND VPWR VPWR _5530_/C
+ sky130_fd_sc_hd__o311a_1
XFILLER_105_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5459_ _5459_/A _5459_/B _5570_/B VGND VGND VPWR VPWR _5459_/X sky130_fd_sc_hd__and3_1
XFILLER_78_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7129_ _7207_/CLK _7129_/D fanout633/X VGND VGND VPWR VPWR _7129_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_19_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_170 _6633_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4830_ _4836_/B _5146_/B _5017_/A VGND VGND VPWR VPWR _4830_/Y sky130_fd_sc_hd__o21bai_4
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_181 _6834_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_192 _6843_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4761_ _4761_/A _5375_/B VGND VGND VPWR VPWR _4762_/C sky130_fd_sc_hd__nand2_1
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6500_ _7434_/Q _6097_/X _6771_/C _6468_/X _7586_/Q VGND VGND VPWR VPWR _6500_/X
+ sky130_fd_sc_hd__a32o_1
X_3712_ _4547_/A _5682_/A _5682_/B VGND VGND VPWR VPWR _3712_/X sky130_fd_sc_hd__and3_1
X_7480_ _7608_/CLK _7480_/D fanout610/X VGND VGND VPWR VPWR _7480_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_174_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4692_ _4743_/C _5358_/B VGND VGND VPWR VPWR _4692_/Y sky130_fd_sc_hd__nand2_1
XFILLER_174_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3643_ input18/X _5669_/B _4535_/B _3555_/X _7520_/Q VGND VGND VPWR VPWR _3643_/X
+ sky130_fd_sc_hd__a32o_1
X_6431_ _7130_/Q _6130_/X _6160_/X _7060_/Q _6430_/X VGND VGND VPWR VPWR _6431_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6362_ _7205_/Q _6153_/X _6158_/X _7240_/Q _6361_/X VGND VGND VPWR VPWR _6362_/X
+ sky130_fd_sc_hd__a221o_1
X_3574_ hold74/A _5686_/B _6020_/A VGND VGND VPWR VPWR _3574_/X sky130_fd_sc_hd__and3_4
X_5313_ _5313_/A _5313_/B _5313_/C VGND VGND VPWR VPWR _5314_/A sky130_fd_sc_hd__and3_1
X_6293_ _7472_/Q _6130_/X _6286_/X _6287_/X _6292_/X VGND VGND VPWR VPWR _6293_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_170_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5244_ _5244_/A1 _4811_/Y _4873_/Y _5004_/Y _5088_/Y VGND VGND VPWR VPWR _5259_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_142_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold18 hold18/A VGND VGND VPWR VPWR hold2/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold29 hold29/A VGND VGND VPWR VPWR hold29/X sky130_fd_sc_hd__buf_12
X_5175_ _5614_/C _5181_/C _5186_/C VGND VGND VPWR VPWR _5175_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_29_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4126_ _6469_/A _4126_/B _6485_/B VGND VGND VPWR VPWR _6771_/B sky130_fd_sc_hd__and3_4
XFILLER_29_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4057_ _4057_/A0 hold1/A _4192_/B VGND VGND VPWR VPWR _6936_/D sky130_fd_sc_hd__mux2_1
XFILLER_37_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4959_ _4948_/A _4948_/B _4959_/C _5074_/A VGND VGND VPWR VPWR _5093_/B sky130_fd_sc_hd__and4bb_1
XFILLER_177_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7678_ _7679_/CLK _7678_/D fanout635/X VGND VGND VPWR VPWR hold65/A sky130_fd_sc_hd__dfrtp_2
XFILLER_177_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6629_ _7527_/Q _6469_/A _6536_/C _6484_/X _7511_/Q VGND VGND VPWR VPWR _6629_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_165_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire441 _4787_/Y VGND VGND VPWR VPWR _4950_/C sky130_fd_sc_hd__buf_4
XFILLER_156_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire452 wire452/A VGND VGND VPWR VPWR wire452/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6980_ _7668_/CLK _6980_/D VGND VGND VPWR VPWR _6980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5931_ hold297/X _6039_/A1 _5938_/S VGND VGND VPWR VPWR _7514_/D sky130_fd_sc_hd__mux2_1
XFILLER_65_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5862_ hold644/X _5988_/A1 _5866_/S VGND VGND VPWR VPWR _7453_/D sky130_fd_sc_hd__mux2_1
XFILLER_33_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7601_ _7601_/CLK _7601_/D fanout611/X VGND VGND VPWR VPWR _7601_/Q sky130_fd_sc_hd__dfrtp_1
X_4813_ _5375_/A _4813_/B _4813_/C VGND VGND VPWR VPWR _4813_/X sky130_fd_sc_hd__and3_1
X_5793_ hold617/X _5991_/A1 _5794_/S VGND VGND VPWR VPWR _5793_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7532_ _7603_/CLK _7532_/D fanout611/X VGND VGND VPWR VPWR _7532_/Q sky130_fd_sc_hd__dfrtp_2
X_4744_ _4744_/A _4744_/B _4744_/C VGND VGND VPWR VPWR _4744_/Y sky130_fd_sc_hd__nor3_1
XFILLER_159_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4675_ _4747_/B _5490_/C _5364_/B _5614_/C VGND VGND VPWR VPWR _4742_/C sky130_fd_sc_hd__nand4_1
X_7463_ _7616_/CLK _7463_/D fanout610/X VGND VGND VPWR VPWR _7463_/Q sky130_fd_sc_hd__dfrtp_2
X_6414_ _7647_/Q _6109_/X _6413_/X _6811_/S VGND VGND VPWR VPWR _6414_/X sky130_fd_sc_hd__o22a_1
XFILLER_147_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3626_ _7416_/Q _5840_/A _5957_/B _3552_/X _7392_/Q VGND VGND VPWR VPWR _3626_/X
+ sky130_fd_sc_hd__a32o_1
X_7394_ _7586_/CLK _7394_/D fanout625/X VGND VGND VPWR VPWR _7394_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_134_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3557_ _5993_/A _5661_/A _5661_/B VGND VGND VPWR VPWR _3557_/X sky130_fd_sc_hd__and3_4
X_6345_ _7067_/Q _6231_/D _6427_/A3 _6428_/A2 _7210_/Q VGND VGND VPWR VPWR _6345_/X
+ sky130_fd_sc_hd__a32o_1
X_6276_ _7328_/Q _6067_/X _6145_/C _6112_/X _7432_/Q VGND VGND VPWR VPWR _6276_/X
+ sky130_fd_sc_hd__a32o_1
X_3488_ _4067_/A _6912_/Q _3500_/C VGND VGND VPWR VPWR _3488_/X sky130_fd_sc_hd__and3_1
XFILLER_130_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput108 wb_adr_i[18] VGND VGND VPWR VPWR _4584_/D sky130_fd_sc_hd__clkbuf_2
X_5227_ _5227_/A _5227_/B _5227_/C VGND VGND VPWR VPWR _5230_/B sky130_fd_sc_hd__and3_1
Xinput119 wb_adr_i[28] VGND VGND VPWR VPWR input119/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5158_ _4747_/B _5595_/B _5358_/B _5153_/C _5157_/X VGND VGND VPWR VPWR _5158_/X
+ sky130_fd_sc_hd__a41o_1
X_4109_ _5143_/A _4109_/B VGND VGND VPWR VPWR _4573_/A sky130_fd_sc_hd__nand2_2
XFILLER_57_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5089_ _5089_/A _5091_/B VGND VGND VPWR VPWR _5127_/C sky130_fd_sc_hd__nand2_1
XFILLER_72_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_70 _3676_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_81 _4009_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_92 _5249_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4460_ _3692_/Y _4460_/A1 _4462_/S VGND VGND VPWR VPWR _7156_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold307 _7523_/Q VGND VGND VPWR VPWR hold307/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold318 _5798_/X VGND VGND VPWR VPWR _7396_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold329 _7332_/Q VGND VGND VPWR VPWR hold329/X sky130_fd_sc_hd__dlygate4sd3_1
X_4391_ _6864_/A1 _4391_/A1 _4393_/S VGND VGND VPWR VPWR _4391_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6130_ _6158_/D _6160_/D _6145_/C VGND VGND VPWR VPWR _6130_/X sky130_fd_sc_hd__and3_4
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _6064_/A _6061_/B _6061_/C VGND VGND VPWR VPWR _7621_/D sky130_fd_sc_hd__and3_1
XFILLER_98_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1007 _4466_/X VGND VGND VPWR VPWR _7161_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5012_ _4990_/A _5014_/D _5017_/A VGND VGND VPWR VPWR _5012_/X sky130_fd_sc_hd__and3b_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1018 _7159_/Q VGND VGND VPWR VPWR _4464_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1029 _7693_/A VGND VGND VPWR VPWR _4294_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6963_ _7668_/CLK _6963_/D _6815_/A VGND VGND VPWR VPWR _6963_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5914_ _5914_/A0 _6031_/A0 _5920_/S VGND VGND VPWR VPWR _5914_/X sky130_fd_sc_hd__mux2_1
X_6894_ _6899_/A _6907_/B VGND VGND VPWR VPWR _6894_/X sky130_fd_sc_hd__and2_1
X_5845_ hold552/X _5926_/A0 _5848_/S VGND VGND VPWR VPWR _5845_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5776_ _6046_/A1 hold863/X _5776_/S VGND VGND VPWR VPWR _5776_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7515_ _7515_/CLK _7515_/D fanout623/X VGND VGND VPWR VPWR _7515_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_159_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4727_ _4727_/A _4727_/B _4727_/C VGND VGND VPWR VPWR _4727_/Y sky130_fd_sc_hd__nor3_1
XFILLER_147_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7446_ _7602_/CLK hold20/X fanout615/X VGND VGND VPWR VPWR _7446_/Q sky130_fd_sc_hd__dfrtp_2
X_4658_ _4599_/Y _4660_/C _4990_/A VGND VGND VPWR VPWR _4658_/X sky130_fd_sc_hd__o21ba_1
XFILLER_190_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput90 spimemio_flash_io2_oeb VGND VGND VPWR VPWR _4147_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_123_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold830 _6014_/X VGND VGND VPWR VPWR _7588_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3609_ _7545_/Q _3530_/X _3554_/X _7569_/Q _3608_/X VGND VGND VPWR VPWR _3617_/C
+ sky130_fd_sc_hd__a221o_1
Xhold841 _7048_/Q VGND VGND VPWR VPWR hold841/X sky130_fd_sc_hd__dlygate4sd3_1
X_7377_ _7553_/CLK _7377_/D fanout624/X VGND VGND VPWR VPWR _7377_/Q sky130_fd_sc_hd__dfrtp_1
X_4589_ _4990_/A _5014_/D _5015_/C VGND VGND VPWR VPWR _4590_/B sky130_fd_sc_hd__nand3_1
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold852 _5974_/X VGND VGND VPWR VPWR _7553_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap571 wire572/X VGND VGND VPWR VPWR _5512_/D sky130_fd_sc_hd__clkbuf_2
Xhold863 _7377_/Q VGND VGND VPWR VPWR hold863/X sky130_fd_sc_hd__dlygate4sd3_1
X_6328_ _7061_/Q _6359_/B _6432_/A3 _6153_/X _7204_/Q VGND VGND VPWR VPWR _6328_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_107_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold874 _5812_/X VGND VGND VPWR VPWR _7409_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap582 _4884_/Y VGND VGND VPWR VPWR _4995_/A sky130_fd_sc_hd__clkbuf_2
Xhold885 _7521_/Q VGND VGND VPWR VPWR hold885/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 _7401_/Q VGND VGND VPWR VPWR hold896/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6259_ _7383_/Q _6077_/X _6254_/X _6256_/X _6258_/X VGND VGND VPWR VPWR _6259_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_88_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1530 _6415_/X VGND VGND VPWR VPWR _7648_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1541 _4562_/X VGND VGND VPWR VPWR _7241_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1552 _7635_/Q VGND VGND VPWR VPWR _6106_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1563 _7258_/Q VGND VGND VPWR VPWR _3467_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1574 _4355_/X VGND VGND VPWR VPWR _7063_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1585 _7271_/Q VGND VGND VPWR VPWR _5649_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_703 _4116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1596 hold60/A VGND VGND VPWR VPWR _5627_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_714 _4969_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_725 _4196_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_736 _5666_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_747 _6451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3960_ _7292_/Q _3623_/X _3695_/X _7047_/Q _3959_/X VGND VGND VPWR VPWR _3960_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_51_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3891_ _7612_/Q _3580_/X _3887_/X _3889_/X _3890_/X VGND VGND VPWR VPWR _3901_/C
+ sky130_fd_sc_hd__a2111o_1
XFILLER_43_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5630_ _5761_/A1 hold458/X _5633_/S VGND VGND VPWR VPWR _5630_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5561_ _5604_/B1 _5415_/X _4991_/Y _5287_/X _5413_/X VGND VGND VPWR VPWR _5561_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_129_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7300_ _7305_/CLK _7300_/D fanout620/X VGND VGND VPWR VPWR _7300_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_157_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4512_ _4512_/A0 _6012_/A0 _4516_/S VGND VGND VPWR VPWR _4512_/X sky130_fd_sc_hd__mux2_1
X_5492_ _5490_/B _5490_/C _5490_/A _5491_/Y VGND VGND VPWR VPWR _5493_/C sky130_fd_sc_hd__a31o_1
Xhold104 _7245_/Q VGND VGND VPWR VPWR hold104/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_156_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold115 _7690_/A VGND VGND VPWR VPWR hold115/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold126 _4303_/X VGND VGND VPWR VPWR _7019_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7231_ _7231_/CLK _7231_/D fanout599/X VGND VGND VPWR VPWR _7231_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_105_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4443_ hold50/X _4443_/A1 _4444_/S VGND VGND VPWR VPWR hold57/A sky130_fd_sc_hd__mux2_1
XFILLER_132_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold137 _7047_/Q VGND VGND VPWR VPWR hold137/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold148 _5701_/X VGND VGND VPWR VPWR _7310_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 _5896_/X VGND VGND VPWR VPWR _7483_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7162_ _7215_/CLK _7162_/D _6903_/A VGND VGND VPWR VPWR _7162_/Q sky130_fd_sc_hd__dfstp_2
X_4374_ _4374_/A0 _6865_/A1 _4375_/S VGND VGND VPWR VPWR _4374_/X sky130_fd_sc_hd__mux2_1
Xfanout606 fanout612/X VGND VGND VPWR VPWR fanout606/X sky130_fd_sc_hd__clkbuf_16
Xfanout617 fanout618/X VGND VGND VPWR VPWR fanout617/X sky130_fd_sc_hd__buf_8
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6113_ _7624_/Q _7623_/Q _6151_/B _6126_/D VGND VGND VPWR VPWR _6113_/Y sky130_fd_sc_hd__nor4_2
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7093_ _7240_/CLK _7093_/D fanout599/X VGND VGND VPWR VPWR _7093_/Q sky130_fd_sc_hd__dfstp_1
Xfanout628 fanout631/X VGND VGND VPWR VPWR fanout628/X sky130_fd_sc_hd__buf_8
Xfanout639 input126/X VGND VGND VPWR VPWR _5017_/A sky130_fd_sc_hd__buf_8
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6044_ hold951/X _6044_/A1 _6046_/S VGND VGND VPWR VPWR _6044_/X sky130_fd_sc_hd__mux2_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6946_ _4172_/B2 _6946_/D _6901_/X VGND VGND VPWR VPWR _6946_/Q sky130_fd_sc_hd__dfrtn_1
X_6877_ _6911_/A _6911_/B VGND VGND VPWR VPWR _6877_/X sky130_fd_sc_hd__and2_1
X_5828_ hold933/X _6044_/A1 _5830_/S VGND VGND VPWR VPWR _5828_/X sky130_fd_sc_hd__mux2_1
X_5759_ _5975_/B _5759_/B _6029_/B VGND VGND VPWR VPWR _5767_/S sky130_fd_sc_hd__and3_4
XFILLER_162_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7429_ _7432_/CLK _7429_/D fanout631/X VGND VGND VPWR VPWR _7429_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_163_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold660 _5873_/X VGND VGND VPWR VPWR _7463_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 _7298_/Q VGND VGND VPWR VPWR hold671/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold682 _7209_/Q VGND VGND VPWR VPWR hold682/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 _5772_/X VGND VGND VPWR VPWR _7373_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1360 _7228_/Q VGND VGND VPWR VPWR hold593/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_523 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1371 _7331_/Q VGND VGND VPWR VPWR hold980/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1382 _5654_/X VGND VGND VPWR VPWR _7275_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1393 _7280_/Q VGND VGND VPWR VPWR hold887/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_500 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_511 _7714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_522 _4195_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_533 input81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_544 input81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_555 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_566 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_577 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_588 _4185_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_599 _6002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput209 _3453_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[6] sky130_fd_sc_hd__buf_12
XFILLER_153_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4090_ _4090_/A0 _4096_/A0 _4097_/S VGND VGND VPWR VPWR _6923_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6800_ _6800_/A _6800_/B _6800_/C _6800_/D VGND VGND VPWR VPWR _6800_/Y sky130_fd_sc_hd__nor4_1
XFILLER_91_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4992_ _4992_/A _4992_/B _4992_/C _4992_/D VGND VGND VPWR VPWR _5002_/B sky130_fd_sc_hd__nor4_2
XFILLER_63_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6731_ _7107_/Q _6099_/B _6694_/C _6469_/X _7165_/Q VGND VGND VPWR VPWR _6731_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_189_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3943_ _7252_/Q _5840_/A hold70/A _3545_/X _7403_/Q VGND VGND VPWR VPWR _3943_/X
+ sky130_fd_sc_hd__a32o_1
X_6662_ _6661_/X _6686_/A1 _6812_/S VGND VGND VPWR VPWR _7656_/D sky130_fd_sc_hd__mux2_1
X_3874_ _7216_/Q _4547_/A _4529_/B _3714_/X _7221_/Q VGND VGND VPWR VPWR _3874_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_176_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5613_ _5613_/A1 wire535/X _5612_/Y _5599_/X VGND VGND VPWR VPWR _7249_/D sky130_fd_sc_hd__a211o_1
X_6593_ _7526_/Q _6447_/X _6474_/C _7374_/Q _6590_/X VGND VGND VPWR VPWR _6593_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_191_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5544_ _5079_/B _5233_/X _5544_/C _5544_/D VGND VGND VPWR VPWR _5580_/C sky130_fd_sc_hd__and4bb_1
XFILLER_129_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5475_ _5476_/A _5233_/B _5233_/C _5074_/B _5474_/X VGND VGND VPWR VPWR _5475_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_117_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7214_ _7217_/CLK _7214_/D _6903_/A VGND VGND VPWR VPWR _7214_/Q sky130_fd_sc_hd__dfrtp_4
X_4426_ hold757/X _6863_/A1 _4429_/S VGND VGND VPWR VPWR _4426_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout403 _5682_/C VGND VGND VPWR VPWR _5678_/C sky130_fd_sc_hd__clkbuf_8
Xfanout414 _4295_/A VGND VGND VPWR VPWR _5975_/B sky130_fd_sc_hd__buf_12
X_7145_ _7676_/CLK _7145_/D VGND VGND VPWR VPWR _7145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4357_ hold568/X _4564_/A1 _4357_/S VGND VGND VPWR VPWR _4357_/X sky130_fd_sc_hd__mux2_1
Xfanout425 _5261_/D VGND VGND VPWR VPWR _5452_/A sky130_fd_sc_hd__buf_4
XFILLER_86_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout458 _6097_/X VGND VGND VPWR VPWR _6099_/B sky130_fd_sc_hd__buf_12
X_4288_ _4287_/X hold492/X _4294_/S VGND VGND VPWR VPWR _4288_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7076_ _7398_/CLK _7076_/D fanout619/X VGND VGND VPWR VPWR _7076_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout469 _6446_/X VGND VGND VPWR VPWR _6562_/C sky130_fd_sc_hd__buf_6
X_6027_ hold763/X _6045_/A1 _6028_/S VGND VGND VPWR VPWR _6027_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6929_ _4183_/A1 _6929_/D _6884_/X VGND VGND VPWR VPWR _6929_/Q sky130_fd_sc_hd__dfrtp_2
Xclkbuf_leaf_31_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7613_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_120_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_46_csclk _7352_/CLK VGND VGND VPWR VPWR _7611_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_89_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold490 _7087_/Q VGND VGND VPWR VPWR hold490/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1190 hold1465/X VGND VGND VPWR VPWR _4403_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_330 _5988_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_341 _6159_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_352 hold81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_363 _5753_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_374 _3550_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_385 _3553_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_396 _3702_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3590_ _7481_/Q _6861_/A _5957_/B _3557_/X _7577_/Q VGND VGND VPWR VPWR _3590_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_173_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5260_ _5526_/A _5260_/B _5527_/A _5260_/D VGND VGND VPWR VPWR _5263_/C sky130_fd_sc_hd__nand4_1
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4211_ _6969_/Q _6971_/Q _6970_/Q VGND VGND VPWR VPWR _6858_/C sky130_fd_sc_hd__nor3_4
XFILLER_142_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5191_ _5195_/B _5476_/B _5191_/C _5249_/C VGND VGND VPWR VPWR _5203_/B sky130_fd_sc_hd__nand4_1
XFILLER_141_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4142_ _6917_/Q _4192_/B _3464_/X VGND VGND VPWR VPWR _6953_/D sky130_fd_sc_hd__a21oi_1
XFILLER_96_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4073_ _4078_/A1 _6912_/Q _3500_/C _4072_/X VGND VGND VPWR VPWR _4073_/X sky130_fd_sc_hd__a31o_1
XFILLER_68_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4975_ _5027_/D _4800_/Y _6970_/Q VGND VGND VPWR VPWR _4975_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_149_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6714_ _7190_/Q _6454_/X _6468_/X _7175_/Q _6713_/X VGND VGND VPWR VPWR _6714_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_149_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3926_ _7451_/Q _6861_/A wire401/X _3580_/X _7611_/Q VGND VGND VPWR VPWR _3926_/X
+ sky130_fd_sc_hd__a32o_1
X_7694_ _7694_/A VGND VGND VPWR VPWR _7694_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_177_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6645_ _7328_/Q _6645_/B _6645_/C VGND VGND VPWR VPWR _6645_/X sky130_fd_sc_hd__and3_1
X_3857_ _7078_/Q _5840_/A _4487_/A _3581_/X _7364_/Q VGND VGND VPWR VPWR _3857_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_20_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6576_ _7533_/Q _6487_/A _6562_/C _6481_/X _7381_/Q VGND VGND VPWR VPWR _6576_/X
+ sky130_fd_sc_hd__a32o_1
X_3788_ _7288_/Q _3623_/X _3674_/X _7269_/Q _3787_/X VGND VGND VPWR VPWR _3788_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_192_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5527_ _5527_/A _5527_/B _5527_/C _5527_/D VGND VGND VPWR VPWR _5530_/B sky130_fd_sc_hd__and4_1
XFILLER_117_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5458_ _5021_/B _5404_/B _5571_/B1 _5074_/A _4963_/X VGND VGND VPWR VPWR _5459_/B
+ sky130_fd_sc_hd__a221oi_1
XFILLER_160_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4409_ _4409_/A0 _4556_/A1 _4411_/S VGND VGND VPWR VPWR _4409_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5389_ _5452_/A _5389_/B _5389_/C _5389_/D VGND VGND VPWR VPWR _5389_/X sky130_fd_sc_hd__and4_1
XFILLER_120_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7128_ _7686_/CLK _7128_/D _6891_/A VGND VGND VPWR VPWR _7128_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_59_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7059_ _7192_/CLK _7059_/D fanout617/X VGND VGND VPWR VPWR _7059_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_101_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_160 _6487_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_171 _6633_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_182 _6834_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_193 _6843_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4760_ _4801_/C _4760_/B _4760_/C _4760_/D VGND VGND VPWR VPWR _5375_/B sky130_fd_sc_hd__and4_1
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3711_ _4547_/A _5661_/B _5682_/B VGND VGND VPWR VPWR _3711_/X sky130_fd_sc_hd__and3_1
X_4691_ _4760_/C _4760_/B _4760_/D VGND VGND VPWR VPWR _4691_/X sky130_fd_sc_hd__a21bo_1
X_6430_ _7085_/Q _6359_/B _6115_/X _6157_/X _7105_/Q VGND VGND VPWR VPWR _6430_/X
+ sky130_fd_sc_hd__a32o_1
X_3642_ _7424_/Q _3602_/X _3640_/X _3641_/X VGND VGND VPWR VPWR _3654_/C sky130_fd_sc_hd__a211o_1
X_6361_ _7117_/Q _6359_/B _6170_/C _6159_/X _7107_/Q VGND VGND VPWR VPWR _6361_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_127_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3573_ _5661_/A _3717_/B _3573_/C VGND VGND VPWR VPWR _3573_/X sky130_fd_sc_hd__and3_2
X_5312_ _5313_/B _5130_/B _5452_/C _5311_/X VGND VGND VPWR VPWR _5314_/B sky130_fd_sc_hd__a31o_1
XFILLER_161_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6292_ _7440_/Q _6159_/X _6290_/X _6291_/X _6289_/X VGND VGND VPWR VPWR _6292_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_170_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5243_ _4570_/Y _4873_/Y _4910_/Y _5001_/Y _4888_/Y VGND VGND VPWR VPWR _5259_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_142_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold19 hold2/X VGND VGND VPWR VPWR hold19/X sky130_fd_sc_hd__buf_6
X_5174_ _5153_/A _5490_/C _5297_/A _4946_/A _4748_/B VGND VGND VPWR VPWR _5174_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_69_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4125_ _7628_/Q _7629_/Q VGND VGND VPWR VPWR _6469_/A sky130_fd_sc_hd__and2b_4
XFILLER_68_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4056_ _4056_/A0 _4057_/A0 _4192_/B VGND VGND VPWR VPWR _6937_/D sky130_fd_sc_hd__mux2_1
XFILLER_43_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4958_ _4966_/A _5021_/B _4946_/B _5401_/A _5404_/B VGND VGND VPWR VPWR _5570_/A
+ sky130_fd_sc_hd__a32oi_1
XFILLER_51_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3909_ _7042_/Q _4529_/B _6038_/B _7467_/Q _3528_/X VGND VGND VPWR VPWR _3909_/X
+ sky130_fd_sc_hd__a32o_1
X_7677_ _7679_/CLK _7677_/D fanout635/X VGND VGND VPWR VPWR hold89/A sky130_fd_sc_hd__dfrtp_2
X_4889_ _5375_/C _5389_/B VGND VGND VPWR VPWR _4889_/Y sky130_fd_sc_hd__nand2_1
XFILLER_137_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6628_ _7559_/Q _6453_/X _6457_/X _7575_/Q VGND VGND VPWR VPWR _6628_/X sky130_fd_sc_hd__a22o_1
XFILLER_124_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6559_ _6686_/S _6559_/A2 _6557_/X _6558_/X VGND VGND VPWR VPWR _6559_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5930_ _5984_/A _6002_/A _6029_/B VGND VGND VPWR VPWR _5938_/S sky130_fd_sc_hd__and3_4
XFILLER_65_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5861_ _5861_/A0 hold81/X _5866_/S VGND VGND VPWR VPWR hold82/A sky130_fd_sc_hd__mux2_1
X_7600_ _7603_/CLK _7600_/D fanout611/X VGND VGND VPWR VPWR _7600_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_61_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4812_ _4943_/A _5375_/C _4813_/B _5375_/A VGND VGND VPWR VPWR _4814_/B sky130_fd_sc_hd__o211a_1
X_5792_ hold926/X _6044_/A1 _5794_/S VGND VGND VPWR VPWR _5792_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7531_ _7553_/CLK _7531_/D fanout624/X VGND VGND VPWR VPWR _7531_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_187_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4743_ _5490_/C _5297_/A _4743_/C VGND VGND VPWR VPWR _4744_/B sky130_fd_sc_hd__and3_1
XFILLER_159_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7462_ _7462_/CLK _7462_/D fanout604/X VGND VGND VPWR VPWR _7462_/Q sky130_fd_sc_hd__dfrtp_4
X_4674_ _4992_/D _5233_/A VGND VGND VPWR VPWR _4674_/Y sky130_fd_sc_hd__nand2_2
XFILLER_119_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6413_ _7039_/Q _6082_/Y _6399_/X _6412_/X VGND VGND VPWR VPWR _6413_/X sky130_fd_sc_hd__o22a_2
X_3625_ _7384_/Q _5993_/B _5759_/B _3567_/X _7344_/Q VGND VGND VPWR VPWR _3625_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_135_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7393_ _7568_/CLK _7393_/D fanout622/X VGND VGND VPWR VPWR _7393_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_134_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6344_ _6343_/X _6366_/A1 _6812_/S VGND VGND VPWR VPWR _6344_/X sky130_fd_sc_hd__mux2_1
X_3556_ _3713_/A _5661_/A _5628_/A VGND VGND VPWR VPWR _3556_/X sky130_fd_sc_hd__and3_4
XFILLER_143_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6275_ _6274_/X _6297_/A2 _6611_/S VGND VGND VPWR VPWR _6275_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3487_ _3508_/S hold32/X VGND VGND VPWR VPWR hold33/A sky130_fd_sc_hd__and2_1
XFILLER_102_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput109 wb_adr_i[19] VGND VGND VPWR VPWR _4584_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_102_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5226_ _4761_/A _5068_/C _4989_/X VGND VGND VPWR VPWR _5227_/C sky130_fd_sc_hd__a21oi_1
XFILLER_69_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5157_ _5153_/C _4946_/A _4740_/D _4747_/B _5358_/B VGND VGND VPWR VPWR _5157_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_111_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4108_ _5096_/B _5096_/C VGND VGND VPWR VPWR _5143_/A sky130_fd_sc_hd__nor2_4
X_5088_ _5313_/B _5088_/B VGND VGND VPWR VPWR _5088_/Y sky130_fd_sc_hd__nand2_8
XFILLER_72_727 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4039_ _3967_/S _4037_/Y _4038_/X _3904_/S VGND VGND VPWR VPWR _6942_/D sky130_fd_sc_hd__o211a_1
XFILLER_37_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_60 _3562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_71 _3700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_82 _4036_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_93 _5625_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_532 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold308 _5941_/X VGND VGND VPWR VPWR _7523_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold319 _7348_/Q VGND VGND VPWR VPWR hold319/X sky130_fd_sc_hd__dlygate4sd3_1
X_4390_ _6863_/A1 hold729/X _4393_/S VGND VGND VPWR VPWR _4390_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _7620_/Q _6063_/D _7621_/Q VGND VGND VPWR VPWR _6061_/C sky130_fd_sc_hd__a21o_1
XFILLER_140_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1008 _7171_/Q VGND VGND VPWR VPWR _4478_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5011_ _5011_/A _5011_/B _5011_/C VGND VGND VPWR VPWR _5048_/B sky130_fd_sc_hd__nor3_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1019 _4464_/X VGND VGND VPWR VPWR _7159_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6962_ _7668_/CLK _6962_/D _6815_/A VGND VGND VPWR VPWR _6962_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_53_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5913_ hold534/X _6039_/A1 _5920_/S VGND VGND VPWR VPWR _5913_/X sky130_fd_sc_hd__mux2_1
X_6893_ _6903_/A _6907_/B VGND VGND VPWR VPWR _6893_/X sky130_fd_sc_hd__and2_1
X_5844_ _5844_/A0 _6042_/A1 _5848_/S VGND VGND VPWR VPWR _5844_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5775_ _5991_/A1 hold708/X _5776_/S VGND VGND VPWR VPWR _5775_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7514_ _7614_/CLK _7514_/D fanout606/X VGND VGND VPWR VPWR _7514_/Q sky130_fd_sc_hd__dfstp_2
X_4726_ _5297_/A _4743_/C _5358_/B VGND VGND VPWR VPWR _4727_/B sky130_fd_sc_hd__and3_1
XFILLER_21_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7445_ _7445_/CLK _7445_/D fanout628/X VGND VGND VPWR VPWR _7445_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_147_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4657_ _4660_/C _4653_/Y _4655_/Y _4651_/Y VGND VGND VPWR VPWR _4657_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_175_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput80 spi_sck VGND VGND VPWR VPWR input80/X sky130_fd_sc_hd__buf_4
X_3608_ _7505_/Q _3516_/X _5984_/B _3607_/X VGND VGND VPWR VPWR _3608_/X sky130_fd_sc_hd__a31o_1
Xhold820 _4371_/X VGND VGND VPWR VPWR _7076_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput91 spimemio_flash_io3_do VGND VGND VPWR VPWR input91/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7376_ _7568_/CLK _7376_/D fanout622/X VGND VGND VPWR VPWR _7376_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_174_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4588_ _4990_/A _5015_/C VGND VGND VPWR VPWR _4836_/A sky130_fd_sc_hd__nand2_8
Xhold831 _7449_/Q VGND VGND VPWR VPWR hold831/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold842 _4337_/X VGND VGND VPWR VPWR _7048_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold853 _7537_/Q VGND VGND VPWR VPWR hold853/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6327_ _7066_/Q _6115_/X _6322_/X _6324_/X _6326_/X VGND VGND VPWR VPWR _6327_/X
+ sky130_fd_sc_hd__a2111o_1
Xhold864 _5776_/X VGND VGND VPWR VPWR _7377_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3539_ _3714_/A hold74/X _5993_/B VGND VGND VPWR VPWR hold75/A sky130_fd_sc_hd__and3_4
XFILLER_116_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmgmt_gpio_15_buff_inst _4166_/X VGND VGND VPWR VPWR mgmt_gpio_out[15] sky130_fd_sc_hd__clkbuf_8
Xhold875 _7367_/Q VGND VGND VPWR VPWR hold875/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold886 _5938_/X VGND VGND VPWR VPWR _7521_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold897 _5803_/X VGND VGND VPWR VPWR _7401_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6258_ _7399_/Q _6114_/X _6149_/X _7423_/Q _6257_/X VGND VGND VPWR VPWR _6258_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5209_ _5209_/A _5209_/B _5209_/C VGND VGND VPWR VPWR _5215_/A sky130_fd_sc_hd__nor3_1
X_6189_ _7340_/Q _6131_/C _6149_/X _7420_/Q _6188_/X VGND VGND VPWR VPWR _6189_/X
+ sky130_fd_sc_hd__a221o_1
Xhold1520 _4055_/X VGND VGND VPWR VPWR _6938_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1531 _7133_/Q VGND VGND VPWR VPWR hold1531/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1542 _7640_/Q VGND VGND VPWR VPWR _6252_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1553 _7650_/Q VGND VGND VPWR VPWR _6510_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1564 _7362_/Q VGND VGND VPWR VPWR _5760_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1575 _7322_/Q VGND VGND VPWR VPWR hold812/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1586 _7162_/Q VGND VGND VPWR VPWR hold725/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_704 _4116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1597 _7647_/Q VGND VGND VPWR VPWR _6391_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_83_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_715 _4969_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_726 _4196_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_737 _5666_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_748 _6451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3890_ _7053_/Q _5680_/B _5678_/B _6011_/A _7588_/Q VGND VGND VPWR VPWR _3890_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_188_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5560_ _5560_/A _5560_/B _5560_/C _5560_/D VGND VGND VPWR VPWR _5625_/C sky130_fd_sc_hd__nand4_1
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4511_ _4511_/A _5659_/C _4511_/C _6861_/C VGND VGND VPWR VPWR _4516_/S sky130_fd_sc_hd__and4_4
XFILLER_184_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5491_ _4772_/Y _5484_/Y _5174_/X VGND VGND VPWR VPWR _5491_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_172_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7230_ _7233_/CLK _7230_/D fanout599/X VGND VGND VPWR VPWR _7230_/Q sky130_fd_sc_hd__dfrtp_2
Xhold105 hold189/X VGND VGND VPWR VPWR _3622_/A sky130_fd_sc_hd__buf_6
X_4442_ hold85/X _4442_/A1 _4444_/S VGND VGND VPWR VPWR hold91/A sky130_fd_sc_hd__mux2_1
Xhold116 _4286_/X VGND VGND VPWR VPWR _7007_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 _7244_/Q VGND VGND VPWR VPWR hold127/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 _4336_/X VGND VGND VPWR VPWR _7047_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 _7507_/Q VGND VGND VPWR VPWR hold149/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7161_ _7215_/CLK _7161_/D _6891_/A VGND VGND VPWR VPWR _7161_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_113_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4373_ hold518/X _5789_/A1 _4375_/S VGND VGND VPWR VPWR _4373_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout607 fanout609/X VGND VGND VPWR VPWR fanout607/X sky130_fd_sc_hd__buf_8
X_6112_ _6151_/B _6392_/B _6166_/B VGND VGND VPWR VPWR _6112_/X sky130_fd_sc_hd__and3_4
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout618 fanout633/X VGND VGND VPWR VPWR fanout618/X sky130_fd_sc_hd__buf_8
X_7092_ _7233_/CLK _7092_/D fanout599/X VGND VGND VPWR VPWR _7092_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout629 fanout630/X VGND VGND VPWR VPWR fanout629/X sky130_fd_sc_hd__buf_8
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ hold162/X _6043_/A1 _6046_/S VGND VGND VPWR VPWR _6043_/X sky130_fd_sc_hd__mux2_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6945_ _4172_/B2 _6945_/D _6900_/X VGND VGND VPWR VPWR _6945_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_54_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6876_ _6911_/A _6911_/B VGND VGND VPWR VPWR _6876_/X sky130_fd_sc_hd__and2_1
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5827_ hold226/X _5926_/A0 _5830_/S VGND VGND VPWR VPWR _5827_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5758_ hold857/X _6046_/A1 _5758_/S VGND VGND VPWR VPWR _5758_/X sky130_fd_sc_hd__mux2_1
X_4709_ _5407_/A _5404_/A _5429_/D VGND VGND VPWR VPWR _4709_/Y sky130_fd_sc_hd__nand3_4
X_5689_ _5689_/A hold29/X VGND VGND VPWR VPWR _5695_/S sky130_fd_sc_hd__nand2_4
XFILLER_175_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7428_ _7557_/CLK _7428_/D fanout627/X VGND VGND VPWR VPWR _7428_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_162_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold650 _4366_/X VGND VGND VPWR VPWR _7072_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7359_ _7445_/CLK _7359_/D fanout628/X VGND VGND VPWR VPWR _7359_/Q sky130_fd_sc_hd__dfrtp_4
Xhold661 hold661/A VGND VGND VPWR VPWR hold661/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold672 _5687_/X VGND VGND VPWR VPWR _7298_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold683 _4524_/X VGND VGND VPWR VPWR _7209_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold694 _7408_/Q VGND VGND VPWR VPWR hold694/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_134_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1350 _3657_/X VGND VGND VPWR VPWR _6948_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1361 _7501_/Q VGND VGND VPWR VPWR hold1361/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1372 _5725_/X VGND VGND VPWR VPWR _7331_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1383 _7044_/Q VGND VGND VPWR VPWR hold966/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_501 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1394 _7423_/Q VGND VGND VPWR VPWR hold933/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_512 _7714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_523 _4195_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_534 input81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_545 input81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_556 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_567 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_578 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_589 _4116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4991_ _5109_/A _5040_/A VGND VGND VPWR VPWR _4991_/Y sky130_fd_sc_hd__nand2_2
XFILLER_51_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6730_ _7097_/Q _6444_/X _6460_/X _7252_/Q VGND VGND VPWR VPWR _6730_/X sky130_fd_sc_hd__a22o_1
X_3942_ _7427_/Q _3556_/X _5849_/A _7443_/Q _3906_/X VGND VGND VPWR VPWR _3942_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_177_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6661_ _6660_/X _6661_/A1 _6686_/S VGND VGND VPWR VPWR _6661_/X sky130_fd_sc_hd__mux2_1
X_3873_ _7460_/Q _3549_/X _3715_/X _7108_/Q _3872_/X VGND VGND VPWR VPWR _3883_/C
+ sky130_fd_sc_hd__a221o_1
X_5612_ _5626_/D _5626_/C _5611_/X _5603_/Y VGND VGND VPWR VPWR _5612_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_177_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6592_ _7326_/Q _6471_/X _6501_/X _7566_/Q _6591_/X VGND VGND VPWR VPWR _6592_/X
+ sky130_fd_sc_hd__a221o_1
X_5543_ _4709_/Y _4800_/Y _4821_/Y _5476_/Y _5235_/X VGND VGND VPWR VPWR _5544_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_157_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5474_ _5233_/B _5068_/C _5250_/X _5473_/Y VGND VGND VPWR VPWR _5474_/X sky130_fd_sc_hd__a31o_1
XFILLER_172_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7213_ _7255_/CLK _7213_/D fanout618/X VGND VGND VPWR VPWR _7213_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_172_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4425_ _4425_/A0 _6862_/A1 _4429_/S VGND VGND VPWR VPWR _4425_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout404 hold36/X VGND VGND VPWR VPWR _5682_/C sky130_fd_sc_hd__buf_8
X_7144_ _7676_/CLK _7144_/D VGND VGND VPWR VPWR _7144_/Q sky130_fd_sc_hd__dfxtp_1
X_4356_ _4356_/A0 _6865_/A1 _4357_/S VGND VGND VPWR VPWR _4356_/X sky130_fd_sc_hd__mux2_1
Xfanout415 _3581_/B VGND VGND VPWR VPWR _5661_/A sky130_fd_sc_hd__buf_8
XFILLER_99_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout426 _5233_/B VGND VGND VPWR VPWR _5322_/A sky130_fd_sc_hd__buf_6
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7075_ _7686_/CLK _7075_/D _6891_/A VGND VGND VPWR VPWR _7075_/Q sky130_fd_sc_hd__dfrtp_2
X_4287_ hold147/X _6043_/A1 _4293_/S VGND VGND VPWR VPWR _4287_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6026_ hold883/X _6044_/A1 _6028_/S VGND VGND VPWR VPWR _6026_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6928_ _6950_/CLK _6928_/D _6883_/X VGND VGND VPWR VPWR _6928_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6859_ _7681_/Q _6967_/Q _6858_/X VGND VGND VPWR VPWR _6859_/X sky130_fd_sc_hd__o21a_1
XFILLER_50_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold480 _6045_/X VGND VGND VPWR VPWR _7616_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 _4384_/X VGND VGND VPWR VPWR _7087_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1180 hold1550/X VGND VGND VPWR VPWR _5640_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1191 _7182_/Q VGND VGND VPWR VPWR _4491_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_320 _6427_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_331 _5988_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_342 fanout612/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_353 hold85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_364 _5807_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_375 _3525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_386 _3571_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_397 _3702_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4210_ _4210_/A _4210_/B _4210_/C _4209_/Y VGND VGND VPWR VPWR _4215_/B sky130_fd_sc_hd__nor4b_1
X_5190_ _5188_/X _5189_/Y _4613_/X VGND VGND VPWR VPWR _5190_/X sky130_fd_sc_hd__a21bo_1
XFILLER_141_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4141_ _4130_/B _6811_/S _6109_/B _4139_/X VGND VGND VPWR VPWR _7140_/D sky130_fd_sc_hd__a211o_1
XFILLER_68_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4072_ _6929_/Q _4064_/X _4065_/Y _4085_/B VGND VGND VPWR VPWR _4072_/X sky130_fd_sc_hd__o211a_1
XFILLER_83_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4974_ _4658_/X _4660_/Y _4688_/C _5229_/A _5043_/B VGND VGND VPWR VPWR _5476_/C
+ sky130_fd_sc_hd__o221a_4
XFILLER_189_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6713_ _7087_/Q _6458_/X _6474_/B _7052_/Q VGND VGND VPWR VPWR _6713_/X sky130_fd_sc_hd__a22o_1
X_3925_ _7339_/Q _3567_/X _3585_/X _7331_/Q _3924_/X VGND VGND VPWR VPWR _3925_/X
+ sky130_fd_sc_hd__a221o_1
X_7693_ _7693_/A VGND VGND VPWR VPWR _7693_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6644_ _7568_/Q _6097_/X _6516_/C _6466_/X _7408_/Q VGND VGND VPWR VPWR _6644_/X
+ sky130_fd_sc_hd__a32o_1
X_3856_ _7388_/Q _3552_/X _3556_/X _7428_/Q _3842_/X VGND VGND VPWR VPWR _3856_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_149_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6575_ hold40/A _6694_/B _6563_/C _6464_/X _7461_/Q VGND VGND VPWR VPWR _6575_/X
+ sky130_fd_sc_hd__a32o_1
X_3787_ _6975_/Q _3560_/X _4275_/S input38/X _3786_/X VGND VGND VPWR VPWR _3787_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5526_ _5526_/A _5526_/B _5526_/C VGND VGND VPWR VPWR _5527_/D sky130_fd_sc_hd__and3_1
XFILLER_117_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5457_ _5404_/X _5457_/B _5570_/D VGND VGND VPWR VPWR _5459_/A sky130_fd_sc_hd__and3b_1
XFILLER_160_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4408_ hold418/X _5869_/A1 _4411_/S VGND VGND VPWR VPWR _4408_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5388_ _4953_/B _4859_/Y _4949_/Y _5387_/X _4880_/Y VGND VGND VPWR VPWR _5392_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7127_ _7312_/CLK _7127_/D _6891_/A VGND VGND VPWR VPWR _7127_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_87_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4339_ hold213/X _6866_/A1 _4339_/S VGND VGND VPWR VPWR _7050_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7058_ _7207_/CLK _7058_/D fanout616/X VGND VGND VPWR VPWR _7058_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_86_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6009_ hold788/X _6045_/A1 _6010_/S VGND VGND VPWR VPWR _6009_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_150 _6474_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_161 _6487_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_172 _6651_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_183 _6834_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_194 _6843_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3710_ _3714_/A _5686_/A hold98/A VGND VGND VPWR VPWR _3710_/X sky130_fd_sc_hd__and3_2
XFILLER_14_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4690_ _4760_/C _4760_/B _4760_/D VGND VGND VPWR VPWR _5595_/D sky130_fd_sc_hd__a21boi_4
XFILLER_186_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_587 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3641_ _7584_/Q _6002_/A _6038_/B _3554_/X _7568_/Q VGND VGND VPWR VPWR _3641_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6360_ _7072_/Q _6359_/B _6334_/C _6160_/X _7057_/Q VGND VGND VPWR VPWR _6360_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_127_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3572_ _3905_/B _5661_/B _4511_/C VGND VGND VPWR VPWR _3572_/X sky130_fd_sc_hd__and3_4
XFILLER_155_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5311_ _5311_/A _5313_/C _5311_/C VGND VGND VPWR VPWR _5311_/X sky130_fd_sc_hd__and3_1
X_6291_ _7360_/Q _6159_/B _6137_/X _6157_/X _7504_/Q VGND VGND VPWR VPWR _6291_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_142_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5242_ _5244_/A1 _4811_/Y _4871_/X _5001_/Y _5088_/Y VGND VGND VPWR VPWR _5527_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_88_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__1128_ clkbuf_0__1128_/X VGND VGND VPWR VPWR _4459_/A0 sky130_fd_sc_hd__clkbuf_16
XFILLER_69_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_30_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7518_/CLK sky130_fd_sc_hd__clkbuf_16
X_5173_ _5358_/A _5490_/C _5153_/C _5172_/Y VGND VGND VPWR VPWR _5173_/X sky130_fd_sc_hd__a31o_1
XFILLER_96_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4124_ _4126_/B _6485_/B VGND VGND VPWR VPWR _6791_/C sky130_fd_sc_hd__and2_4
XFILLER_56_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput1 debug_mode VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__clkbuf_2
X_4055_ _4055_/A0 hold48/A _4192_/B VGND VGND VPWR VPWR _4055_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_45_csclk _7352_/CLK VGND VGND VPWR VPWR _7435_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_71_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4957_ _4966_/A _4957_/B _4957_/C VGND VGND VPWR VPWR _5404_/B sky130_fd_sc_hd__and3_2
XFILLER_51_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3908_ input21/X _3574_/X _3706_/X _7102_/Q _3907_/X VGND VGND VPWR VPWR _3908_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_177_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7676_ _7676_/CLK _7676_/D fanout635/X VGND VGND VPWR VPWR hold17/A sky130_fd_sc_hd__dfrtp_1
X_4888_ _5401_/A _5313_/B VGND VGND VPWR VPWR _4888_/Y sky130_fd_sc_hd__nand2_2
XFILLER_192_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3839_ _3838_/Y _6945_/Q _3967_/S VGND VGND VPWR VPWR _3839_/X sky130_fd_sc_hd__mux2_1
X_6627_ _7455_/Q _6459_/X _6468_/X _7591_/Q _6626_/X VGND VGND VPWR VPWR _6632_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_137_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6558_ _7316_/Q _6759_/D _6686_/S VGND VGND VPWR VPWR _6558_/X sky130_fd_sc_hd__o21ba_1
XFILLER_152_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5509_ _5285_/X _5412_/X _4949_/Y _5015_/Y _5604_/B1 VGND VGND VPWR VPWR _5560_/A
+ sky130_fd_sc_hd__a311o_1
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6489_ _7450_/Q _6459_/X _6486_/X _7498_/Q VGND VGND VPWR VPWR _6489_/X sky130_fd_sc_hd__a22o_1
XFILLER_106_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire410 hold54/X VGND VGND VPWR VPWR hold55/A sky130_fd_sc_hd__clkbuf_1
XFILLER_11_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_616 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5860_ hold996/X _6040_/A1 _5866_/S VGND VGND VPWR VPWR _7451_/D sky130_fd_sc_hd__mux2_1
XFILLER_34_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4811_ _4992_/D _4813_/C VGND VGND VPWR VPWR _4811_/Y sky130_fd_sc_hd__nand2_8
XFILLER_92_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5791_ hold218/X _5935_/A1 _5794_/S VGND VGND VPWR VPWR _5791_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4742_ _4742_/A _5218_/C _4742_/C _4742_/D VGND VGND VPWR VPWR _4744_/C sky130_fd_sc_hd__nand4_1
X_7530_ _7603_/CLK _7530_/D fanout611/X VGND VGND VPWR VPWR _7530_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_193_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7461_ _7616_/CLK hold13/X fanout610/X VGND VGND VPWR VPWR _7461_/Q sky130_fd_sc_hd__dfrtp_4
X_4673_ _5189_/A _4992_/B _5146_/A VGND VGND VPWR VPWR _4673_/X sky130_fd_sc_hd__and3_1
XFILLER_174_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6412_ _7104_/Q _6158_/D _6127_/X _6405_/X _6411_/X VGND VGND VPWR VPWR _6412_/X
+ sky130_fd_sc_hd__a311o_1
X_3624_ _7662_/Q _7291_/Q _7292_/Q VGND VGND VPWR VPWR _3624_/X sky130_fd_sc_hd__mux2_4
X_7392_ _7445_/CLK _7392_/D fanout628/X VGND VGND VPWR VPWR _7392_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_174_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6343_ _6811_/S _7644_/Q _6341_/X _6342_/X VGND VGND VPWR VPWR _6343_/X sky130_fd_sc_hd__a22o_1
X_3555_ _3714_/A _5686_/A _6002_/A VGND VGND VPWR VPWR _3555_/X sky130_fd_sc_hd__and3_4
XFILLER_127_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6274_ _6686_/S _7641_/Q _6272_/X _6273_/X VGND VGND VPWR VPWR _6274_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3486_ hold42/X hold72/X _3484_/X VGND VGND VPWR VPWR _3547_/D sky130_fd_sc_hd__a21oi_4
XFILLER_143_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5225_ _4625_/Y _5585_/A1 _4759_/X _4984_/Y _4987_/Y VGND VGND VPWR VPWR _5227_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_130_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5156_ _5156_/A _5156_/B _5597_/D VGND VGND VPWR VPWR _5156_/Y sky130_fd_sc_hd__nand3_1
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4107_ _4884_/A _5096_/A VGND VGND VPWR VPWR _4109_/B sky130_fd_sc_hd__nand2_1
XFILLER_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5087_ _5189_/D _5112_/B _5313_/B VGND VGND VPWR VPWR _5091_/B sky130_fd_sc_hd__and3_2
XFILLER_110_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4038_ _6917_/Q _6913_/Q _4193_/B _4038_/B1 VGND VGND VPWR VPWR _4038_/X sky130_fd_sc_hd__a31o_1
XFILLER_72_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5989_ hold407/X _6043_/A1 hold63/X VGND VGND VPWR VPWR _5989_/X sky130_fd_sc_hd__mux2_1
XFILLER_169_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_671 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_50 hold70/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7659_ _7662_/CLK _7659_/D fanout598/X VGND VGND VPWR VPWR _7659_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_61 _3562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 _3701_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_83 _4036_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_94 _5893_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput190 _3436_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[23] sky130_fd_sc_hd__buf_12
XFILLER_121_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold309 _7708_/A VGND VGND VPWR VPWR hold309/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _5042_/A _5311_/C _5111_/D VGND VGND VPWR VPWR _5048_/A sky130_fd_sc_hd__and3_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1009 _4478_/X VGND VGND VPWR VPWR _7171_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6961_ _7668_/CLK _6961_/D _6815_/A VGND VGND VPWR VPWR _6961_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_81_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5912_ _6861_/A _5984_/B _6038_/C VGND VGND VPWR VPWR _5920_/S sky130_fd_sc_hd__and3_4
X_6892_ _6903_/A _6907_/B VGND VGND VPWR VPWR _6892_/X sky130_fd_sc_hd__and2_1
XFILLER_34_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5843_ hold371/X _5843_/A1 _5848_/S VGND VGND VPWR VPWR _5843_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5774_ _6044_/A1 hold861/X _5776_/S VGND VGND VPWR VPWR _5774_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7513_ _7616_/CLK _7513_/D fanout610/X VGND VGND VPWR VPWR _7513_/Q sky130_fd_sc_hd__dfrtp_4
X_4725_ _5196_/A _4743_/C _5358_/B VGND VGND VPWR VPWR _4727_/A sky130_fd_sc_hd__and3_1
XFILLER_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7444_ _7602_/CLK _7444_/D fanout613/X VGND VGND VPWR VPWR _7444_/Q sky130_fd_sc_hd__dfrtp_2
X_4656_ _4704_/A _5316_/C _4653_/Y _4655_/Y _4651_/Y VGND VGND VPWR VPWR _5043_/B
+ sky130_fd_sc_hd__o311a_2
XFILLER_190_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput70 mgmt_gpio_in[7] VGND VGND VPWR VPWR _4198_/B sky130_fd_sc_hd__buf_2
X_3607_ input19/X _3573_/C _4535_/B _3555_/X _7521_/Q VGND VGND VPWR VPWR _3607_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_135_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput81 spi_sdo VGND VGND VPWR VPWR input81/X sky130_fd_sc_hd__buf_4
Xhold810 _7511_/Q VGND VGND VPWR VPWR hold810/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_174_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4587_ _4587_/A _4587_/B VGND VGND VPWR VPWR _4785_/A sky130_fd_sc_hd__nor2_8
X_7375_ _7553_/CLK _7375_/D fanout624/X VGND VGND VPWR VPWR _7375_/Q sky130_fd_sc_hd__dfrtp_2
Xhold821 _7359_/Q VGND VGND VPWR VPWR hold821/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold832 _5857_/X VGND VGND VPWR VPWR _7449_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput92 spimemio_flash_io3_oeb VGND VGND VPWR VPWR _4145_/B sky130_fd_sc_hd__clkbuf_1
Xhold843 hold843/A VGND VGND VPWR VPWR hold843/X sky130_fd_sc_hd__dlygate4sd3_1
X_3538_ _5661_/A _3573_/C _5661_/B VGND VGND VPWR VPWR hold56/A sky130_fd_sc_hd__and3_4
Xhold854 _5956_/X VGND VGND VPWR VPWR _7537_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6326_ _7179_/Q wire452/A _6149_/X _7086_/Q _6325_/X VGND VGND VPWR VPWR _6326_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_116_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold865 _7337_/Q VGND VGND VPWR VPWR hold865/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap573 _5137_/C VGND VGND VPWR VPWR _5517_/A2 sky130_fd_sc_hd__clkbuf_2
Xhold876 _5765_/X VGND VGND VPWR VPWR _7367_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 hold887/A VGND VGND VPWR VPWR hold887/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold898 _7371_/Q VGND VGND VPWR VPWR hold898/X sky130_fd_sc_hd__dlygate4sd3_1
X_6257_ _7327_/Q _6067_/X _6145_/C _6119_/X _7415_/Q VGND VGND VPWR VPWR _6257_/X
+ sky130_fd_sc_hd__a32o_1
X_3469_ _3469_/A _3469_/B VGND VGND VPWR VPWR _7257_/D sky130_fd_sc_hd__nor2_1
XFILLER_131_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5208_ _5614_/A _5002_/B _5007_/Y _4761_/A _5005_/C VGND VGND VPWR VPWR _5209_/C
+ sky130_fd_sc_hd__a32o_1
XFILLER_190_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6188_ _7348_/Q _6302_/B1 _6141_/X _7364_/Q VGND VGND VPWR VPWR _6188_/X sky130_fd_sc_hd__a22o_1
Xhold1510 _7236_/Q VGND VGND VPWR VPWR hold1510/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1521 _7338_/Q VGND VGND VPWR VPWR hold487/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1532 _4439_/X VGND VGND VPWR VPWR _7133_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5139_ _5074_/A _4704_/A _5085_/Y _5138_/Y VGND VGND VPWR VPWR _5139_/Y sky130_fd_sc_hd__o31ai_1
Xhold1543 _7652_/Q VGND VGND VPWR VPWR _6560_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1554 hold4/A VGND VGND VPWR VPWR _4061_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1565 hold48/A VGND VGND VPWR VPWR _4056_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1576 _7506_/Q VGND VGND VPWR VPWR _5922_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_83_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1587 _7418_/Q VGND VGND VPWR VPWR hold1587/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_705 _5669_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1598 _6963_/Q VGND VGND VPWR VPWR _4210_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_716 _6082_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_727 _4196_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_738 _5282_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4510_ hold278/X _6866_/A1 _4510_/S VGND VGND VPWR VPWR _4510_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5490_ _5490_/A _5490_/B _5490_/C VGND VGND VPWR VPWR _5490_/X sky130_fd_sc_hd__and3_1
XFILLER_8_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold106 _3905_/B VGND VGND VPWR VPWR _3586_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4441_ _6866_/A1 hold191/X _4444_/S VGND VGND VPWR VPWR _4441_/X sky130_fd_sc_hd__mux2_1
Xhold117 hold117/A VGND VGND VPWR VPWR hold117/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 _3509_/Y VGND VGND VPWR VPWR hold128/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold139 _7022_/Q VGND VGND VPWR VPWR hold139/X sky130_fd_sc_hd__dlygate4sd3_1
X_7160_ _7160_/CLK _7160_/D _6891_/A VGND VGND VPWR VPWR _7160_/Q sky130_fd_sc_hd__dfrtp_2
X_4372_ hold564/X _5761_/A1 _4375_/S VGND VGND VPWR VPWR _4372_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6111_ _7624_/Q _7623_/Q _6166_/C VGND VGND VPWR VPWR _6131_/C sky130_fd_sc_hd__and3_4
Xfanout608 fanout609/X VGND VGND VPWR VPWR fanout608/X sky130_fd_sc_hd__buf_8
XFILLER_98_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7091_ _7238_/CLK _7091_/D fanout602/X VGND VGND VPWR VPWR _7091_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_140_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout619 fanout633/X VGND VGND VPWR VPWR fanout619/X sky130_fd_sc_hd__buf_8
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6042_ _6042_/A0 _6042_/A1 _6046_/S VGND VGND VPWR VPWR _7613_/D sky130_fd_sc_hd__mux2_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6944_ _4172_/B2 _6944_/D _6899_/X VGND VGND VPWR VPWR _6944_/Q sky130_fd_sc_hd__dfrtn_1
X_6875_ _6911_/A _6911_/B VGND VGND VPWR VPWR _6875_/X sky130_fd_sc_hd__and2_1
XFILLER_169_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5826_ _5826_/A0 _6042_/A1 _5830_/S VGND VGND VPWR VPWR _5826_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5757_ hold773/X _5991_/A1 _5758_/S VGND VGND VPWR VPWR _5757_/X sky130_fd_sc_hd__mux2_1
X_4708_ _4992_/B _4992_/D _4822_/A _5189_/A VGND VGND VPWR VPWR _4708_/X sky130_fd_sc_hd__and4bb_2
X_5688_ _5688_/A0 _5869_/A1 _5688_/S VGND VGND VPWR VPWR _5688_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7427_ _7515_/CLK _7427_/D fanout632/X VGND VGND VPWR VPWR _7427_/Q sky130_fd_sc_hd__dfstp_1
X_4639_ _4785_/A _5046_/A _4786_/A _4794_/D VGND VGND VPWR VPWR _4639_/Y sky130_fd_sc_hd__nand4_4
XFILLER_162_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold640 _7129_/Q VGND VGND VPWR VPWR hold640/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold651 hold651/A VGND VGND VPWR VPWR hold651/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7358_ _7613_/CLK _7358_/D fanout626/X VGND VGND VPWR VPWR _7358_/Q sky130_fd_sc_hd__dfrtp_4
Xhold662 hold662/A VGND VGND VPWR VPWR wb_dat_o[0] sky130_fd_sc_hd__buf_12
XFILLER_89_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold673 hold673/A VGND VGND VPWR VPWR hold673/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold684 hold684/A VGND VGND VPWR VPWR hold684/X sky130_fd_sc_hd__dlygate4sd3_1
X_6309_ _7465_/Q _6309_/B _6309_/C VGND VGND VPWR VPWR _6309_/X sky130_fd_sc_hd__and3_1
XFILLER_143_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold695 _5811_/X VGND VGND VPWR VPWR _7408_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7289_ _7289_/CLK _7289_/D fanout597/X VGND VGND VPWR VPWR _7289_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_89_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1340 _7101_/Q VGND VGND VPWR VPWR hold1340/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1351 _7355_/Q VGND VGND VPWR VPWR hold988/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1362 _5916_/X VGND VGND VPWR VPWR _7501_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1373 _7512_/Q VGND VGND VPWR VPWR hold556/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1384 _7381_/Q VGND VGND VPWR VPWR hold1384/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1395 _5828_/X VGND VGND VPWR VPWR _7423_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_502 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_513 _7714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_524 _4195_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_535 input81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_546 input81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_557 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_568 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_579 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4990_ _4990_/A _5040_/A _5007_/D VGND VGND VPWR VPWR _5089_/A sky130_fd_sc_hd__and3_4
XFILLER_90_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3941_ _7515_/Q _3555_/X _3571_/X _7355_/Q _3940_/X VGND VGND VPWR VPWR _3946_/C
+ sky130_fd_sc_hd__a221o_2
XFILLER_31_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6660_ _6651_/Y wire367/X _7320_/Q _6759_/D VGND VGND VPWR VPWR _6660_/X sky130_fd_sc_hd__o2bb2a_1
X_3872_ _7684_/Q _4559_/B hold98/A _3561_/X _7524_/Q VGND VGND VPWR VPWR _3872_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_176_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5611_ _4816_/Y _5611_/A2 _5015_/Y _5610_/Y VGND VGND VPWR VPWR _5611_/X sky130_fd_sc_hd__o31a_1
XFILLER_149_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6591_ _7510_/Q _6791_/D _6536_/C _6807_/A2 _7406_/Q VGND VGND VPWR VPWR _6591_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_192_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5542_ _5551_/A1 _5322_/A _5071_/C _5541_/Y VGND VGND VPWR VPWR _5542_/X sky130_fd_sc_hd__a31o_1
X_5473_ _5473_/A _5583_/B _5580_/A VGND VGND VPWR VPWR _5473_/Y sky130_fd_sc_hd__nand3_1
XFILLER_172_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4424_ _4559_/B _4535_/B _5680_/C VGND VGND VPWR VPWR _4429_/S sky130_fd_sc_hd__and3_2
XFILLER_144_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7212_ _7212_/CLK _7212_/D fanout619/X VGND VGND VPWR VPWR _7212_/Q sky130_fd_sc_hd__dfrtp_1
X_4355_ _4355_/A0 _6864_/A1 _4357_/S VGND VGND VPWR VPWR _4355_/X sky130_fd_sc_hd__mux2_1
X_7143_ _7668_/CLK _7143_/D VGND VGND VPWR VPWR _7143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout416 _5993_/A VGND VGND VPWR VPWR _4547_/A sky130_fd_sc_hd__buf_6
XFILLER_59_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7074_ _7312_/CLK _7074_/D _6891_/A VGND VGND VPWR VPWR _7074_/Q sky130_fd_sc_hd__dfrtp_4
X_4286_ _4285_/X hold115/X _4294_/S VGND VGND VPWR VPWR _4286_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6025_ hold429/X _6043_/A1 _6028_/S VGND VGND VPWR VPWR _6025_/X sky130_fd_sc_hd__mux2_1
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6927_ _6950_/CLK _6927_/D _6882_/X VGND VGND VPWR VPWR _6927_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6858_ _6965_/Q _6968_/Q _6858_/C _6858_/D VGND VGND VPWR VPWR _6858_/X sky130_fd_sc_hd__and4bb_1
XFILLER_167_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5809_ hold301/X _5935_/A1 _5812_/S VGND VGND VPWR VPWR _5809_/X sky130_fd_sc_hd__mux2_1
X_6789_ _7065_/Q _6453_/X _6465_/X _7183_/Q _6788_/X VGND VGND VPWR VPWR _6789_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold470 _5955_/X VGND VGND VPWR VPWR _7536_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 _7028_/Q VGND VGND VPWR VPWR hold481/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold492 _7691_/A VGND VGND VPWR VPWR hold492/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1170 hold1425/X VGND VGND VPWR VPWR _4550_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1181 hold1620/X VGND VGND VPWR VPWR _5681_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1192 _4491_/X VGND VGND VPWR VPWR _7182_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_310 _6759_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_321 _6694_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_332 _5988_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_343 _7662_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_354 _4511_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_365 _5025_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_376 _3525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_387 _3583_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_398 _3788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4140_ _6811_/S _4140_/B VGND VGND VPWR VPWR _4140_/Y sky130_fd_sc_hd__nand2_1
XFILLER_110_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4071_ _4074_/A1 _3490_/X _4085_/B _4064_/X _4070_/Y VGND VGND VPWR VPWR _6930_/D
+ sky130_fd_sc_hd__a41oi_1
XFILLER_49_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4973_ _4972_/X _4971_/Y _4848_/Y VGND VGND VPWR VPWR _4973_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_51_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6712_ _6711_/X _6712_/A1 _6812_/S VGND VGND VPWR VPWR _6712_/X sky130_fd_sc_hd__mux2_1
X_3924_ _7087_/Q _4541_/A _4529_/B _4358_/A _7067_/Q VGND VGND VPWR VPWR _3924_/X
+ sky130_fd_sc_hd__a32o_1
X_7692_ _7692_/A VGND VGND VPWR VPWR _7692_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_189_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6643_ _7416_/Q _6450_/X _6483_/X _7392_/Q _6642_/X VGND VGND VPWR VPWR _6651_/B
+ sky130_fd_sc_hd__a221o_1
X_3855_ _7176_/Q _4481_/A hold98/A _3854_/X VGND VGND VPWR VPWR _3855_/X sky130_fd_sc_hd__a31o_1
XFILLER_149_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3786_ _7039_/Q _5678_/C _4505_/B _3785_/X VGND VGND VPWR VPWR _3786_/X sky130_fd_sc_hd__a31o_1
X_6574_ _7349_/Q _6465_/X _6566_/X _6571_/X _6573_/X VGND VGND VPWR VPWR _6574_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_117_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5525_ _5261_/D _5452_/B _5089_/A _4933_/A _5263_/B VGND VGND VPWR VPWR _5526_/C
+ sky130_fd_sc_hd__a311oi_2
XFILLER_145_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5456_ _4709_/Y _4882_/Y _4854_/X _5407_/C VGND VGND VPWR VPWR _5570_/D sky130_fd_sc_hd__a211o_1
XFILLER_172_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4407_ _4407_/A0 _6862_/A1 _4411_/S VGND VGND VPWR VPWR _4407_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5387_ _4709_/Y _4882_/Y _4859_/Y _4953_/B VGND VGND VPWR VPWR _5387_/X sky130_fd_sc_hd__a211o_1
XFILLER_99_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7126_ _7130_/CLK _7126_/D fanout602/X VGND VGND VPWR VPWR _7126_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_115_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4338_ hold452/X _5673_/A1 _4339_/S VGND VGND VPWR VPWR _7049_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7057_ _7207_/CLK _7057_/D fanout616/X VGND VGND VPWR VPWR _7057_/Q sky130_fd_sc_hd__dfrtp_4
X_4269_ hold363/X _5935_/A1 _4275_/S VGND VGND VPWR VPWR _4269_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6008_ hold224/X hold85/X _6010_/S VGND VGND VPWR VPWR _6008_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_140 _6453_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_151 _6474_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_162 _6487_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_173 _6742_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_184 _6834_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_195 _6843_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3640_ _7488_/Q _3531_/X _6011_/A _7592_/Q _3639_/X VGND VGND VPWR VPWR _3640_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_159_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3571_ _5768_/C _5768_/B hold24/A VGND VGND VPWR VPWR _3571_/X sky130_fd_sc_hd__and3_4
X_5310_ _5310_/A _5310_/B _5310_/C VGND VGND VPWR VPWR _5314_/C sky130_fd_sc_hd__nand3_1
XFILLER_142_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6290_ _7448_/Q _6082_/B _6416_/C _6166_/C VGND VGND VPWR VPWR _6290_/X sky130_fd_sc_hd__o211a_1
XFILLER_154_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5241_ _4570_/Y _4871_/X _4910_/Y _4998_/Y _4888_/Y VGND VGND VPWR VPWR _5260_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_142_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5172_ _4669_/Y _5165_/X _5169_/X _5170_/X VGND VGND VPWR VPWR _5172_/Y sky130_fd_sc_hd__o211ai_1
X_4123_ _7632_/Q _7633_/Q VGND VGND VPWR VPWR _6791_/B sky130_fd_sc_hd__and2b_4
XFILLER_84_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4054_ _4053_/Y _4051_/Y _4048_/Y _4054_/B2 VGND VGND VPWR VPWR _6939_/D sky130_fd_sc_hd__a2bb2o_1
Xinput2 debug_oeb VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4956_ _4961_/A _5401_/A VGND VGND VPWR VPWR _4964_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3907_ _7160_/Q _4535_/B _6038_/B _3583_/X input53/X VGND VGND VPWR VPWR _3907_/X
+ sky130_fd_sc_hd__a32o_1
X_7675_ _7676_/CLK _7675_/D fanout635/X VGND VGND VPWR VPWR hold11/A sky130_fd_sc_hd__dfrtp_1
X_4887_ _5404_/A _5112_/B _5313_/B VGND VGND VPWR VPWR _5092_/A sky130_fd_sc_hd__and3_2
XFILLER_20_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6626_ _7415_/Q _6450_/X _6474_/B _7599_/Q VGND VGND VPWR VPWR _6626_/X sky130_fd_sc_hd__a22o_1
X_3838_ _3796_/X _3838_/B _3838_/C VGND VGND VPWR VPWR _3838_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_118_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6557_ _7404_/Q _6807_/A2 _6541_/X _6548_/X _6556_/X VGND VGND VPWR VPWR _6557_/X
+ sky130_fd_sc_hd__a2111o_2
X_3769_ _7422_/Q _3602_/X _3697_/X _7168_/Q _3768_/X VGND VGND VPWR VPWR _3769_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5508_ _5011_/C _4816_/Y _4953_/C _5064_/Y VGND VGND VPWR VPWR _5560_/D sky130_fd_sc_hd__a31o_1
XFILLER_193_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6488_ _7426_/Q _6444_/X _6482_/X _7482_/Q VGND VGND VPWR VPWR _6488_/X sky130_fd_sc_hd__a22o_1
XFILLER_10_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5439_ _5439_/A1 _6829_/D _5354_/X _5437_/X VGND VGND VPWR VPWR _7246_/D sky130_fd_sc_hd__o22a_1
XFILLER_121_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7109_ _7207_/CLK _7109_/D fanout633/X VGND VGND VPWR VPWR _7109_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_113_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire400 wire401/X VGND VGND VPWR VPWR _5786_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_128_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire455 wire455/A VGND VGND VPWR VPWR wire455/X sky130_fd_sc_hd__clkbuf_2
XFILLER_171_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4810_ _5407_/A _4959_/C _4810_/C VGND VGND VPWR VPWR _5375_/C sky130_fd_sc_hd__and3_4
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5790_ _5790_/A0 _6006_/A1 _5794_/S VGND VGND VPWR VPWR _5790_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4741_ _4741_/A _4741_/B VGND VGND VPWR VPWR _4742_/A sky130_fd_sc_hd__nor2_1
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7460_ _7614_/CLK _7460_/D fanout605/X VGND VGND VPWR VPWR _7460_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_147_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4672_ _4948_/B _4959_/C VGND VGND VPWR VPWR _5102_/B sky130_fd_sc_hd__nand2b_4
XFILLER_147_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6411_ _6158_/D _6400_/X _6406_/X _6410_/X VGND VGND VPWR VPWR _6411_/X sky130_fd_sc_hd__a211o_1
X_3623_ _4340_/A _4493_/C _5678_/C VGND VGND VPWR VPWR _3623_/X sky130_fd_sc_hd__and3_2
X_7391_ _7408_/CLK _7391_/D fanout628/X VGND VGND VPWR VPWR _7391_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_162_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6342_ _7036_/Q _6082_/Y _7140_/Q VGND VGND VPWR VPWR _6342_/X sky130_fd_sc_hd__o21ba_1
XFILLER_127_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3554_ _5984_/A _3905_/B _5661_/B VGND VGND VPWR VPWR _3554_/X sky130_fd_sc_hd__and3_4
XFILLER_127_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6273_ _7319_/Q _6082_/Y _6686_/S VGND VGND VPWR VPWR _6273_/X sky130_fd_sc_hd__o21ba_1
X_3485_ hold42/X hold72/X _3484_/X VGND VGND VPWR VPWR hold73/A sky130_fd_sc_hd__a21o_4
XFILLER_143_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5224_ _5224_/A _5224_/B _5224_/C VGND VGND VPWR VPWR _5227_/A sky130_fd_sc_hd__nor3_1
XFILLER_130_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5155_ wire428/X _5020_/X _5595_/A VGND VGND VPWR VPWR _5597_/D sky130_fd_sc_hd__o21ai_1
XFILLER_84_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4106_ _7635_/Q _7287_/Q _7292_/Q VGND VGND VPWR VPWR _4140_/B sky130_fd_sc_hd__mux2_8
X_5086_ _4795_/Y _4823_/Y _4987_/Y _5085_/Y _4568_/Y VGND VGND VPWR VPWR _5566_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_2_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4037_ _4037_/A _4037_/B _4037_/C VGND VGND VPWR VPWR _4037_/Y sky130_fd_sc_hd__nand3_4
XFILLER_56_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5988_ hold673/X _5988_/A1 hold63/X VGND VGND VPWR VPWR _7565_/D sky130_fd_sc_hd__mux2_1
X_4939_ _4943_/B VGND VGND VPWR VPWR _4939_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_40 _3546_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7658_ _7662_/CLK _7658_/D fanout598/X VGND VGND VPWR VPWR _7658_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_51 hold70/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_62 _3569_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 _3702_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6609_ _6592_/X _6600_/X _6608_/X _6759_/D _7318_/Q VGND VGND VPWR VPWR _6609_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA_84 _6791_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7589_ _7613_/CLK _7589_/D fanout626/X VGND VGND VPWR VPWR _7589_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_95 _5920_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput180 _3445_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[14] sky130_fd_sc_hd__buf_12
Xoutput191 _3435_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[24] sky130_fd_sc_hd__buf_12
XFILLER_153_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_44_csclk _7352_/CLK VGND VGND VPWR VPWR _7607_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_109_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_59_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7601_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6960_ _7680_/CLK _6960_/D _6815_/A VGND VGND VPWR VPWR hold42/A sky130_fd_sc_hd__dfrtp_4
XFILLER_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5911_ hold566/X _6028_/A1 _5911_/S VGND VGND VPWR VPWR _5911_/X sky130_fd_sc_hd__mux2_1
X_6891_ _6891_/A _6907_/B VGND VGND VPWR VPWR _6891_/X sky130_fd_sc_hd__and2_1
XFILLER_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5842_ hold995/X _6040_/A1 _5848_/S VGND VGND VPWR VPWR _5842_/X sky130_fd_sc_hd__mux2_1
XFILLER_167_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5773_ _5935_/A1 hold209/X _5776_/S VGND VGND VPWR VPWR _5773_/X sky130_fd_sc_hd__mux2_1
X_7512_ _7512_/CLK _7512_/D fanout609/X VGND VGND VPWR VPWR _7512_/Q sky130_fd_sc_hd__dfrtp_4
X_4724_ _4724_/A _4724_/B _5203_/C VGND VGND VPWR VPWR _4727_/C sky130_fd_sc_hd__nand3_1
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7443_ _7611_/CLK _7443_/D fanout621/X VGND VGND VPWR VPWR _7443_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_174_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4655_ _5000_/C _4660_/C _5015_/C VGND VGND VPWR VPWR _4655_/Y sky130_fd_sc_hd__o21ai_2
Xinput60 mgmt_gpio_in[31] VGND VGND VPWR VPWR input60/X sky130_fd_sc_hd__clkbuf_1
Xhold800 _7508_/Q VGND VGND VPWR VPWR hold800/X sky130_fd_sc_hd__dlygate4sd3_1
X_3606_ _7425_/Q _3602_/X _3603_/X _3605_/X _3601_/X VGND VGND VPWR VPWR _3617_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_190_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold811 _5927_/X VGND VGND VPWR VPWR _7511_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput71 mgmt_gpio_in[8] VGND VGND VPWR VPWR input71/X sky130_fd_sc_hd__buf_2
X_7374_ _7518_/CLK _7374_/D fanout626/X VGND VGND VPWR VPWR _7374_/Q sky130_fd_sc_hd__dfrtp_4
X_4586_ _4586_/A _4586_/B _4586_/C _4586_/D VGND VGND VPWR VPWR _4587_/B sky130_fd_sc_hd__nand4_4
Xinput82 spi_sdoenb VGND VGND VPWR VPWR _4149_/A sky130_fd_sc_hd__buf_2
Xinput93 trap VGND VGND VPWR VPWR input93/X sky130_fd_sc_hd__clkbuf_4
Xhold822 _5756_/X VGND VGND VPWR VPWR _7359_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold833 hold833/A VGND VGND VPWR VPWR hold833/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 hold844/A VGND VGND VPWR VPWR wb_dat_o[16] sky130_fd_sc_hd__buf_12
X_6325_ _7169_/Q _6157_/C _6166_/C _6428_/B1 _7076_/Q VGND VGND VPWR VPWR _6325_/X
+ sky130_fd_sc_hd__a32o_1
X_3537_ _3622_/A _5661_/B hold23/X VGND VGND VPWR VPWR _5993_/B sky130_fd_sc_hd__and3_4
Xhold855 _7385_/Q VGND VGND VPWR VPWR hold855/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 _5731_/X VGND VGND VPWR VPWR _7337_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap574 _5137_/C VGND VGND VPWR VPWR _5040_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_143_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold877 _7335_/Q VGND VGND VPWR VPWR hold877/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 _7481_/Q VGND VGND VPWR VPWR hold888/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold899 _5770_/X VGND VGND VPWR VPWR _7371_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6256_ _7343_/Q _6131_/C _6309_/C _7335_/Q _6255_/X VGND VGND VPWR VPWR _6256_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_170_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3468_ _3470_/B _3470_/A _3468_/B1 VGND VGND VPWR VPWR _3469_/B sky130_fd_sc_hd__a21oi_1
XFILLER_130_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5207_ _5196_/A _5614_/A _5027_/X _5007_/Y _4985_/B VGND VGND VPWR VPWR _5209_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_69_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6187_ _7404_/Q _6124_/X _6309_/C _7332_/Q _6186_/X VGND VGND VPWR VPWR _6187_/X
+ sky130_fd_sc_hd__a221o_1
Xhold1500 _7651_/Q VGND VGND VPWR VPWR _6559_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1511 _4556_/X VGND VGND VPWR VPWR _7236_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1522 _5733_/X VGND VGND VPWR VPWR _7338_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1533 _7645_/Q VGND VGND VPWR VPWR _6366_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5138_ _5138_/A _5138_/B _5138_/C VGND VGND VPWR VPWR _5138_/Y sky130_fd_sc_hd__nor3_1
Xhold1544 _7649_/Q VGND VGND VPWR VPWR _6439_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_184_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1555 hold7/A VGND VGND VPWR VPWR _4059_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1566 _6976_/Q VGND VGND VPWR VPWR hold222/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1577 _7217_/Q VGND VGND VPWR VPWR hold733/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1588 _7461_/Q VGND VGND VPWR VPWR _5871_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5069_ _5297_/A _5071_/B _5071_/C VGND VGND VPWR VPWR _5069_/X sky130_fd_sc_hd__and3_1
Xhold1599 _6929_/Q VGND VGND VPWR VPWR _4074_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_706 _6694_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_717 _6082_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_728 _4196_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_739 _6464_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4440_ _5673_/A1 hold400/X _4444_/S VGND VGND VPWR VPWR _7134_/D sky130_fd_sc_hd__mux2_1
XFILLER_156_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold107 _3553_/X VGND VGND VPWR VPWR hold107/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold118 _7246_/Q VGND VGND VPWR VPWR _3502_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold129 _5682_/B VGND VGND VPWR VPWR _4493_/C sky130_fd_sc_hd__buf_6
XFILLER_144_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4371_ hold819/X _6003_/A1 _4375_/S VGND VGND VPWR VPWR _4371_/X sky130_fd_sc_hd__mux2_1
X_6110_ _6811_/S _4140_/B _6109_/X VGND VGND VPWR VPWR _6611_/S sky130_fd_sc_hd__a21oi_4
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout609 fanout612/X VGND VGND VPWR VPWR fanout609/X sky130_fd_sc_hd__buf_4
XFILLER_98_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7090_ _7253_/CLK _7090_/D fanout617/X VGND VGND VPWR VPWR _7090_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_152_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6041_ hold847/X _6041_/A1 _6046_/S VGND VGND VPWR VPWR _6041_/X sky130_fd_sc_hd__mux2_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6943_ _6950_/CLK _6943_/D _6898_/X VGND VGND VPWR VPWR _6943_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_35_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6874_ _6911_/A _6911_/B VGND VGND VPWR VPWR _6874_/X sky130_fd_sc_hd__and2_1
XFILLER_62_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5825_ hold315/X _5843_/A1 _5830_/S VGND VGND VPWR VPWR _5825_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5756_ hold821/X _6044_/A1 _5758_/S VGND VGND VPWR VPWR _5756_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4707_ _4943_/A _5186_/C _5364_/B VGND VGND VPWR VPWR _4707_/X sky130_fd_sc_hd__and3_1
XFILLER_148_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5687_ hold671/X _6862_/A1 _5688_/S VGND VGND VPWR VPWR _5687_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7426_ _7518_/CLK _7426_/D fanout627/X VGND VGND VPWR VPWR _7426_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_147_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4638_ _5143_/B _4595_/B _5229_/A _4785_/A _4785_/C VGND VGND VPWR VPWR _5024_/D
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_190_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold630 hold630/A VGND VGND VPWR VPWR hold630/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7357_ _7421_/CLK _7357_/D fanout630/X VGND VGND VPWR VPWR _7357_/Q sky130_fd_sc_hd__dfrtp_4
Xhold641 _4434_/X VGND VGND VPWR VPWR _7129_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4569_ _4948_/A _5316_/A _5429_/D VGND VGND VPWR VPWR _4569_/X sky130_fd_sc_hd__and3_2
XFILLER_162_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold652 hold652/A VGND VGND VPWR VPWR wb_dat_o[1] sky130_fd_sc_hd__buf_12
XFILLER_89_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap371 _4291_/S VGND VGND VPWR VPWR _4293_/S sky130_fd_sc_hd__buf_12
Xhold663 _7328_/Q VGND VGND VPWR VPWR hold663/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 hold674/A VGND VGND VPWR VPWR hold674/X sky130_fd_sc_hd__dlygate4sd3_1
X_6308_ _7457_/Q _6131_/B _6170_/C _6159_/X _7441_/Q VGND VGND VPWR VPWR _6308_/X
+ sky130_fd_sc_hd__a32o_1
Xhold685 hold685/A VGND VGND VPWR VPWR wb_dat_o[3] sky130_fd_sc_hd__buf_12
X_7288_ _7291_/CLK _7288_/D fanout596/X VGND VGND VPWR VPWR _7288_/Q sky130_fd_sc_hd__dfrtp_1
Xhold696 hold696/A VGND VGND VPWR VPWR hold696/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6239_ _7446_/Q _6082_/B _6416_/C _6166_/C VGND VGND VPWR VPWR _6239_/X sky130_fd_sc_hd__o211a_1
XFILLER_77_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1330 _7219_/Q VGND VGND VPWR VPWR hold1330/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1341 _7427_/Q VGND VGND VPWR VPWR hold981/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1352 _5752_/X VGND VGND VPWR VPWR _7355_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1363 _7269_/Q VGND VGND VPWR VPWR hold529/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1374 _7613_/Q VGND VGND VPWR VPWR hold1374/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1385 _5781_/X VGND VGND VPWR VPWR _7381_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_503 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1396 _7594_/Q VGND VGND VPWR VPWR hold504/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_514 _7714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_525 _4195_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_536 input81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_547 input81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_558 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_569 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3940_ _7435_/Q _5840_/A _5984_/B _3581_/X _7363_/Q VGND VGND VPWR VPWR _3940_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_189_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3871_ _7236_/Q _5628_/A _5678_/B _3870_/X VGND VGND VPWR VPWR _3883_/B sky130_fd_sc_hd__a31o_1
XFILLER_176_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5610_ _5610_/A _5610_/B _5610_/C _5610_/D VGND VGND VPWR VPWR _5610_/Y sky130_fd_sc_hd__nor4_1
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6590_ _7438_/Q _6097_/X _6445_/C _6474_/A _7342_/Q VGND VGND VPWR VPWR _6590_/X
+ sky130_fd_sc_hd__a32o_1
X_5541_ _5580_/A _5618_/A _5583_/C _5580_/B VGND VGND VPWR VPWR _5541_/Y sky130_fd_sc_hd__nand4_1
XFILLER_157_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5472_ _5472_/A _5472_/B _5472_/C VGND VGND VPWR VPWR _5580_/A sky130_fd_sc_hd__and3_1
X_7211_ _7254_/CLK _7211_/D fanout618/X VGND VGND VPWR VPWR _7211_/Q sky130_fd_sc_hd__dfstp_1
X_4423_ _5926_/A0 hold401/X _4423_/S VGND VGND VPWR VPWR _4423_/X sky130_fd_sc_hd__mux2_1
X_7142_ _7680_/CLK _7142_/D _6907_/A VGND VGND VPWR VPWR _7142_/Q sky130_fd_sc_hd__dfrtp_4
X_4354_ hold669/X _6863_/A1 _4357_/S VGND VGND VPWR VPWR _4354_/X sky130_fd_sc_hd__mux2_1
Xfanout406 _3543_/X VGND VGND VPWR VPWR _4529_/B sky130_fd_sc_hd__buf_12
Xfanout417 _5984_/A VGND VGND VPWR VPWR _5993_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7073_ _7686_/CLK _7073_/D fanout599/X VGND VGND VPWR VPWR _7073_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_59_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4285_ _5700_/A1 hold9/X _4293_/S VGND VGND VPWR VPWR _4285_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6024_ _6024_/A0 _6042_/A1 _6028_/S VGND VGND VPWR VPWR _6024_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6926_ _7258_/CLK _6926_/D _6881_/X VGND VGND VPWR VPWR hold94/A sky130_fd_sc_hd__dfrtp_2
XFILLER_81_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6857_ _6970_/Q _6857_/A2 _6856_/X VGND VGND VPWR VPWR _6857_/X sky130_fd_sc_hd__a21o_1
XFILLER_80_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5808_ _5808_/A0 _6006_/A1 _5812_/S VGND VGND VPWR VPWR _5808_/X sky130_fd_sc_hd__mux2_1
X_6788_ _7085_/Q _6645_/B _6536_/C _6468_/X _7178_/Q VGND VGND VPWR VPWR _6788_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_183_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5739_ hold589/X _5991_/A1 _5740_/S VGND VGND VPWR VPWR _5739_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7409_ _7553_/CLK _7409_/D fanout622/X VGND VGND VPWR VPWR _7409_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_163_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold460 hold460/A VGND VGND VPWR VPWR hold460/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold471 hold471/A VGND VGND VPWR VPWR hold471/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold482 _4314_/X VGND VGND VPWR VPWR _7028_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold493 _4288_/X VGND VGND VPWR VPWR _7008_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1160 hold1591/X VGND VGND VPWR VPWR _4433_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1171 _7306_/Q VGND VGND VPWR VPWR _5697_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1182 hold1646/X VGND VGND VPWR VPWR _4437_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_300 input96/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1193 _7079_/Q VGND VGND VPWR VPWR _4374_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_311 _6809_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_322 _6694_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_333 _4556_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_344 _4167_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_355 hold455/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_366 hold73/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_377 _3525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_388 _3583_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_399 _3838_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_2__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _6950_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4070_ _4070_/A1 _4085_/B _4064_/X _3491_/X VGND VGND VPWR VPWR _4070_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_96_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4972_ _5189_/D _5112_/B _4972_/C VGND VGND VPWR VPWR _4972_/X sky130_fd_sc_hd__and3_1
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6711_ _6710_/X _7657_/Q _7140_/Q VGND VGND VPWR VPWR _6711_/X sky130_fd_sc_hd__mux2_1
X_3923_ _7082_/Q _4559_/B _5680_/A _5689_/A input62/X VGND VGND VPWR VPWR _3923_/X
+ sky130_fd_sc_hd__a32o_1
X_7691_ _7691_/A VGND VGND VPWR VPWR _7691_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_177_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6642_ _7368_/Q _6694_/B _6445_/C _6463_/X _7400_/Q VGND VGND VPWR VPWR _6642_/X
+ sky130_fd_sc_hd__a32o_1
X_3854_ input37/X _5984_/B _6038_/B input13/X _3542_/X VGND VGND VPWR VPWR _3854_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_20_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6573_ _7613_/Q _6451_/X _6457_/X _7573_/Q _6572_/X VGND VGND VPWR VPWR _6573_/X
+ sky130_fd_sc_hd__a221o_1
X_3785_ input95/X _5975_/B _5682_/C _3695_/X _7049_/Q VGND VGND VPWR VPWR _3785_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_158_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5524_ _5524_/A _5524_/B _5524_/C _5524_/D VGND VGND VPWR VPWR _5621_/B sky130_fd_sc_hd__and4_1
XFILLER_118_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5455_ _5455_/A _5573_/B _5573_/C VGND VGND VPWR VPWR _5457_/B sky130_fd_sc_hd__and3_1
XFILLER_117_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4406_ _5628_/A _5666_/B _6861_/C VGND VGND VPWR VPWR _4411_/S sky130_fd_sc_hd__and3_2
X_5386_ _4867_/X _4889_/Y _5009_/Y _5088_/Y _5385_/X VGND VGND VPWR VPWR _5524_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_120_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7125_ _7312_/CLK _7125_/D _6891_/A VGND VGND VPWR VPWR _7125_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_99_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4337_ hold841/X _4556_/A1 _4339_/S VGND VGND VPWR VPWR _4337_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7056_ _7242_/CLK _7056_/D fanout616/X VGND VGND VPWR VPWR _7056_/Q sky130_fd_sc_hd__dfrtp_2
X_4268_ _4267_/X hold949/X _4274_/S VGND VGND VPWR VPWR _4268_/X sky130_fd_sc_hd__mux2_1
X_6007_ hold166/X _6043_/A1 _6010_/S VGND VGND VPWR VPWR _6007_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4199_ _7299_/Q _4199_/B VGND VGND VPWR VPWR _4199_/X sky130_fd_sc_hd__and2_2
XFILLER_27_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6909_ _6911_/A _6911_/B VGND VGND VPWR VPWR _6909_/X sky130_fd_sc_hd__and2_1
XFILLER_24_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold290 _4297_/X VGND VGND VPWR VPWR _7013_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_130 _6370_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_141 _6454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_152 _6471_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_163 _6487_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_174 _6785_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_185 _6834_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_196 _6843_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3570_ _3581_/B _5661_/B _5759_/B VGND VGND VPWR VPWR _5777_/A sky130_fd_sc_hd__and3_4
XFILLER_6_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5240_ _5244_/A1 _4811_/Y _4867_/X _4998_/Y _5088_/Y VGND VGND VPWR VPWR _5526_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_115_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5171_ _5358_/A _4946_/A _4934_/C _4744_/B VGND VGND VPWR VPWR _5171_/X sky130_fd_sc_hd__a31o_1
X_4122_ _3421_/Y _4121_/Y _3422_/Y _7139_/Q VGND VGND VPWR VPWR _7139_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_68_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4053_ _4053_/A _6956_/Q _6957_/Q _6955_/Q VGND VGND VPWR VPWR _4053_/Y sky130_fd_sc_hd__nor4b_1
Xinput3 debug_out VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4955_ _4955_/A _5572_/A _4955_/C _4955_/D VGND VGND VPWR VPWR _4964_/A sky130_fd_sc_hd__nor4_1
X_3906_ _7180_/Q _4535_/B _4511_/C _3696_/X _7200_/Q VGND VGND VPWR VPWR _3906_/X
+ sky130_fd_sc_hd__a32o_1
X_7674_ _7676_/CLK _7674_/D _6815_/A VGND VGND VPWR VPWR _7674_/Q sky130_fd_sc_hd__dfrtp_1
X_4886_ _5143_/A _5112_/B _4983_/C VGND VGND VPWR VPWR _5090_/B sky130_fd_sc_hd__and3_1
X_6625_ _7607_/Q _6456_/X _6471_/X _7327_/Q _6624_/X VGND VGND VPWR VPWR _6632_/A
+ sky130_fd_sc_hd__a221o_1
X_3837_ _3837_/A _3837_/B _3837_/C _3837_/D VGND VGND VPWR VPWR _3838_/C sky130_fd_sc_hd__nor4_2
XFILLER_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6556_ _7380_/Q _6481_/X _6552_/X _6555_/X _6809_/D VGND VGND VPWR VPWR _6556_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_146_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3768_ _7090_/Q _4541_/A _4529_/B _3767_/X VGND VGND VPWR VPWR _3768_/X sky130_fd_sc_hd__a31o_1
XFILLER_146_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5507_ _5429_/A _5512_/B _5311_/C _5295_/X _5506_/X VGND VGND VPWR VPWR _5610_/C
+ sky130_fd_sc_hd__a311o_1
X_6487_ _6487_/A _6563_/C _6645_/C VGND VGND VPWR VPWR _6487_/X sky130_fd_sc_hd__and3_4
XFILLER_3_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3699_ _3717_/B _5659_/C _5680_/B VGND VGND VPWR VPWR _4463_/A sky130_fd_sc_hd__and3_2
XFILLER_105_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5438_ _5285_/X _4993_/Y _4960_/Y _5604_/B1 _4991_/Y VGND VGND VPWR VPWR _5438_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_10_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput340 hold686/X VGND VGND VPWR VPWR hold687/A sky130_fd_sc_hd__buf_12
XFILLER_121_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5369_ _5595_/A _5196_/A _5375_/B _4770_/A _4711_/X VGND VGND VPWR VPWR _5369_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_120_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7108_ _7217_/CLK _7108_/D _6903_/A VGND VGND VPWR VPWR _7108_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7039_ _7294_/CLK _7039_/D fanout597/X VGND VGND VPWR VPWR _7039_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_19_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire401 wire401/A VGND VGND VPWR VPWR wire401/X sky130_fd_sc_hd__clkbuf_2
XFILLER_129_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire423 _5601_/Y VGND VGND VPWR VPWR _5603_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_128_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4740_ _4747_/B _5490_/C _5297_/A _4740_/D VGND VGND VPWR VPWR _4741_/A sky130_fd_sc_hd__and4_1
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4671_ _4822_/A _4959_/C VGND VGND VPWR VPWR _5146_/A sky130_fd_sc_hd__and2b_4
XFILLER_159_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6410_ _7217_/Q _6151_/X _6160_/X _7059_/Q _6409_/X VGND VGND VPWR VPWR _6410_/X
+ sky130_fd_sc_hd__a221o_1
X_3622_ _3622_/A _3622_/B _4340_/A VGND VGND VPWR VPWR _3622_/X sky130_fd_sc_hd__and3_1
X_7390_ _7518_/CLK _7390_/D fanout627/X VGND VGND VPWR VPWR _7390_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_162_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6341_ _6159_/B _6327_/X _6340_/X VGND VGND VPWR VPWR _6341_/X sky130_fd_sc_hd__a21o_2
X_3553_ hold69/X _3559_/B _3586_/A VGND VGND VPWR VPWR _3553_/X sky130_fd_sc_hd__and3_4
XFILLER_128_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6272_ _6082_/B _6259_/X _6271_/X VGND VGND VPWR VPWR _6272_/X sky130_fd_sc_hd__a21o_1
X_3484_ hold42/X _3484_/B VGND VGND VPWR VPWR _3484_/X sky130_fd_sc_hd__and2b_1
XFILLER_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5223_ _5476_/A _5614_/A _4758_/X _5059_/A VGND VGND VPWR VPWR _5224_/C sky130_fd_sc_hd__a31o_1
XFILLER_142_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5154_ _5153_/A _5358_/B _4946_/A _4727_/B VGND VGND VPWR VPWR _5162_/B sky130_fd_sc_hd__a31o_1
XFILLER_111_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4105_ _4105_/A0 input58/X _4105_/S VGND VGND VPWR VPWR _6915_/D sky130_fd_sc_hd__mux2_1
XFILLER_111_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5085_ _5313_/C _5146_/C VGND VGND VPWR VPWR _5085_/Y sky130_fd_sc_hd__nand2_1
XFILLER_110_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4036_ _4036_/A _4036_/B _4036_/C _4036_/D VGND VGND VPWR VPWR _4037_/C sky130_fd_sc_hd__nor4_2
XFILLER_112_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5987_ hold345/X hold81/X hold63/X VGND VGND VPWR VPWR _5987_/X sky130_fd_sc_hd__mux2_1
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4938_ _4957_/B _5452_/A _5389_/C VGND VGND VPWR VPWR _4943_/B sky130_fd_sc_hd__and3_1
XANTENNA_30 _5682_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_41 _3553_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7657_ _7657_/CLK _7657_/D fanout607/X VGND VGND VPWR VPWR _7657_/Q sky130_fd_sc_hd__dfrtp_1
X_4869_ _5181_/C _5452_/A _5389_/B _4957_/C VGND VGND VPWR VPWR _4904_/C sky130_fd_sc_hd__nand4_1
XANTENNA_52 hold70/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_63 _3569_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_74 _3704_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6608_ _7382_/Q _6481_/X _6603_/X _6607_/X _6809_/D VGND VGND VPWR VPWR _6608_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA_85 _6791_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7588_ _7612_/CLK _7588_/D fanout606/X VGND VGND VPWR VPWR _7588_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_96 hold76/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6539_ _7612_/Q _6451_/X _6487_/X _7468_/Q VGND VGND VPWR VPWR _6539_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput181 _3444_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[15] sky130_fd_sc_hd__buf_12
Xoutput192 _3434_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[25] sky130_fd_sc_hd__buf_12
XFILLER_47_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5910_ hold516/X _6045_/A1 _5911_/S VGND VGND VPWR VPWR _5910_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6890_ _6891_/A _6908_/B VGND VGND VPWR VPWR _6890_/X sky130_fd_sc_hd__and2_1
XFILLER_34_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5841_ _5841_/A0 _6012_/A0 _5848_/S VGND VGND VPWR VPWR _5841_/X sky130_fd_sc_hd__mux2_1
X_5772_ _6042_/A1 hold692/X _5776_/S VGND VGND VPWR VPWR _5772_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4723_ _4747_/B _5364_/B _5614_/C _5595_/D VGND VGND VPWR VPWR _4724_/B sky130_fd_sc_hd__nand4_1
X_7511_ _7601_/CLK _7511_/D fanout609/X VGND VGND VPWR VPWR _7511_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_147_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7442_ _7568_/CLK hold45/X fanout623/X VGND VGND VPWR VPWR _7442_/Q sky130_fd_sc_hd__dfstp_2
X_4654_ _5297_/A _5108_/B VGND VGND VPWR VPWR _4654_/Y sky130_fd_sc_hd__nand2_1
XFILLER_175_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput50 mgmt_gpio_in[22] VGND VGND VPWR VPWR input50/X sky130_fd_sc_hd__buf_2
XFILLER_116_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3605_ _7489_/Q _3531_/X _3545_/X _7409_/Q _3604_/X VGND VGND VPWR VPWR _3605_/X
+ sky130_fd_sc_hd__a221o_1
Xinput61 mgmt_gpio_in[32] VGND VGND VPWR VPWR input61/X sky130_fd_sc_hd__buf_2
X_7373_ _7445_/CLK _7373_/D fanout628/X VGND VGND VPWR VPWR _7373_/Q sky130_fd_sc_hd__dfrtp_4
X_4585_ _4585_/A _4585_/B _4585_/C _4585_/D VGND VGND VPWR VPWR _4587_/A sky130_fd_sc_hd__nand4_4
Xhold801 _5924_/X VGND VGND VPWR VPWR _7508_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput72 mgmt_gpio_in[9] VGND VGND VPWR VPWR input72/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold812 hold812/A VGND VGND VPWR VPWR hold812/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_174_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold823 _6996_/Q VGND VGND VPWR VPWR hold823/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput83 spimemio_flash_clk VGND VGND VPWR VPWR input83/X sky130_fd_sc_hd__clkbuf_4
Xinput94 uart_enabled VGND VGND VPWR VPWR _4195_/B sky130_fd_sc_hd__clkbuf_1
X_6324_ _7209_/Q _6428_/A2 _6124_/X _7234_/Q _6323_/X VGND VGND VPWR VPWR _6324_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_116_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold834 hold834/A VGND VGND VPWR VPWR wb_dat_o[28] sky130_fd_sc_hd__buf_12
X_3536_ _5669_/B _5661_/B _4493_/C VGND VGND VPWR VPWR _5650_/A sky130_fd_sc_hd__and3_4
XFILLER_143_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold845 _7025_/Q VGND VGND VPWR VPWR hold845/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 _5785_/X VGND VGND VPWR VPWR _7385_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 _7393_/Q VGND VGND VPWR VPWR hold867/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap586 _4631_/Y VGND VGND VPWR VPWR _4660_/C sky130_fd_sc_hd__buf_8
Xhold878 _5729_/X VGND VGND VPWR VPWR _7335_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold889 _5893_/X VGND VGND VPWR VPWR _7481_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6255_ _7391_/Q _6067_/X _6146_/C _6124_/X _7407_/Q VGND VGND VPWR VPWR _6255_/X
+ sky130_fd_sc_hd__a32o_1
X_3467_ _3467_/A _3469_/A VGND VGND VPWR VPWR _7258_/D sky130_fd_sc_hd__xor2_1
X_5206_ _5206_/A _5206_/B _5206_/C VGND VGND VPWR VPWR _5209_/A sky130_fd_sc_hd__nand3_1
X_6186_ _7388_/Q _6231_/D _6146_/C _6432_/A3 _7428_/Q VGND VGND VPWR VPWR _6186_/X
+ sky130_fd_sc_hd__a32o_1
Xhold1501 _6535_/X VGND VGND VPWR VPWR _7651_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1512 _7570_/Q VGND VGND VPWR VPWR hold448/A sky130_fd_sc_hd__dlygate4sd3_1
X_5137_ _5137_/A _5452_/C _5137_/C VGND VGND VPWR VPWR _5138_/B sky130_fd_sc_hd__and3_1
Xhold1523 hold17/A VGND VGND VPWR VPWR _6844_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1534 _6344_/X VGND VGND VPWR VPWR _7645_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1545 _7152_/Q VGND VGND VPWR VPWR _4456_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1556 _7216_/Q VGND VGND VPWR VPWR hold1556/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1567 _6968_/Q VGND VGND VPWR VPWR _6965_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5068_ _5068_/A _5322_/A _5068_/C VGND VGND VPWR VPWR _5073_/A sky130_fd_sc_hd__and3_1
Xhold1578 _6966_/Q VGND VGND VPWR VPWR _4210_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1589 _7163_/Q VGND VGND VPWR VPWR hold563/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_177_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_707 _6407_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4019_ _7354_/Q _3571_/X _5689_/A input61/X _4018_/X VGND VGND VPWR VPWR _4019_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_718 _6645_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_729 _6759_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7709_ _7709_/A VGND VGND VPWR VPWR _7709_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold108 _5914_/X VGND VGND VPWR VPWR _7499_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_156_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold119 _3502_/Y VGND VGND VPWR VPWR hold119/X sky130_fd_sc_hd__dlygate4sd3_1
X_4370_ _4541_/A _4487_/A _6861_/C VGND VGND VPWR VPWR _4375_/S sky130_fd_sc_hd__and3_2
XFILLER_98_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ hold987/X _6040_/A1 _6046_/S VGND VGND VPWR VPWR _7611_/D sky130_fd_sc_hd__mux2_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_663 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6942_ _6950_/CLK _6942_/D _6897_/X VGND VGND VPWR VPWR _6942_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6873_ _6899_/A _6911_/B VGND VGND VPWR VPWR _6873_/X sky130_fd_sc_hd__and2_1
XFILLER_35_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5824_ hold965/X _6040_/A1 _5830_/S VGND VGND VPWR VPWR _5824_/X sky130_fd_sc_hd__mux2_1
XFILLER_167_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5755_ hold276/X _5935_/A1 _5758_/S VGND VGND VPWR VPWR _5755_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4706_ _4760_/D _4706_/B _4760_/C _4706_/D VGND VGND VPWR VPWR _4706_/Y sky130_fd_sc_hd__nand4_1
X_5686_ _5686_/A _5686_/B _5984_/B _5686_/D VGND VGND VPWR VPWR _5686_/X sky130_fd_sc_hd__and4_1
XFILLER_148_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7425_ _7553_/CLK _7425_/D fanout622/X VGND VGND VPWR VPWR _7425_/Q sky130_fd_sc_hd__dfrtp_1
X_4637_ _4637_/A _4884_/A VGND VGND VPWR VPWR _5024_/C sky130_fd_sc_hd__nand2_2
XFILLER_190_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold620 _4302_/X VGND VGND VPWR VPWR _7018_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4568_ _5189_/A _4822_/A _4992_/D VGND VGND VPWR VPWR _4568_/Y sky130_fd_sc_hd__nand3_4
Xhold631 hold631/A VGND VGND VPWR VPWR wb_dat_o[10] sky130_fd_sc_hd__buf_12
X_7356_ _7562_/CLK _7356_/D fanout621/X VGND VGND VPWR VPWR _7356_/Q sky130_fd_sc_hd__dfrtp_4
Xhold642 hold642/A VGND VGND VPWR VPWR hold642/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold653 _7311_/Q VGND VGND VPWR VPWR hold653/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3519_ _3714_/A hold74/A _5975_/B VGND VGND VPWR VPWR _3519_/X sky130_fd_sc_hd__and3_2
X_6307_ _7537_/Q _6160_/D _6427_/A3 _6137_/X _7489_/Q VGND VGND VPWR VPWR _6307_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_116_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold664 _5721_/X VGND VGND VPWR VPWR _7328_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7287_ _7293_/CLK _7287_/D fanout596/X VGND VGND VPWR VPWR _7287_/Q sky130_fd_sc_hd__dfrtp_2
Xhold675 hold675/A VGND VGND VPWR VPWR wb_dat_o[2] sky130_fd_sc_hd__buf_12
XFILLER_143_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold686 hold686/A VGND VGND VPWR VPWR hold686/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4499_ _4499_/A hold29/X VGND VGND VPWR VPWR _4504_/S sky130_fd_sc_hd__nand2_4
Xhold697 hold697/A VGND VGND VPWR VPWR wb_dat_o[8] sky130_fd_sc_hd__buf_12
XFILLER_104_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6238_ _7534_/Q _6160_/D _6427_/A3 _6427_/B1 _7486_/Q VGND VGND VPWR VPWR _6238_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_89_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ _6212_/C1 _6166_/X _6168_/X _6165_/X _6159_/B VGND VGND VPWR VPWR _6169_/X
+ sky130_fd_sc_hd__o41a_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1320 _7365_/Q VGND VGND VPWR VPWR hold1320/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1331 _6944_/Q VGND VGND VPWR VPWR _3903_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1342 _5833_/X VGND VGND VPWR VPWR _7427_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1353 _7341_/Q VGND VGND VPWR VPWR hold1353/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1364 _5647_/X VGND VGND VPWR VPWR _7269_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1375 _7403_/Q VGND VGND VPWR VPWR hold977/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1386 _7518_/Q VGND VGND VPWR VPWR hold223/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1397 _7196_/Q VGND VGND VPWR VPWR hold1397/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_504 _6968_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_515 _7714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_526 input78/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_43_csclk _7352_/CLK VGND VGND VPWR VPWR _7617_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_537 input81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_548 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_559 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_58_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7547_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_185_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3870_ _7171_/Q _4475_/A _5678_/B _3713_/X _7098_/Q VGND VGND VPWR VPWR _3870_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_149_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5540_ _4660_/C _4633_/Y _5011_/A _5350_/A _5539_/Y VGND VGND VPWR VPWR _5580_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_192_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5471_ _5471_/A _5471_/B VGND VGND VPWR VPWR _5583_/B sky130_fd_sc_hd__nor2_1
XFILLER_172_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7210_ _7210_/CLK _7210_/D fanout618/X VGND VGND VPWR VPWR _7210_/Q sky130_fd_sc_hd__dfrtp_2
X_4422_ _6865_/A1 _4422_/A1 _4423_/S VGND VGND VPWR VPWR _4422_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7141_ _7680_/CLK _7141_/D _6886_/A VGND VGND VPWR VPWR _7141_/Q sky130_fd_sc_hd__dfrtp_4
X_4353_ _4353_/A0 _6012_/A0 _4357_/S VGND VGND VPWR VPWR _4353_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout407 _4487_/A VGND VGND VPWR VPWR _4535_/B sky130_fd_sc_hd__buf_12
Xfanout418 hold62/X VGND VGND VPWR VPWR _5984_/A sky130_fd_sc_hd__buf_12
XFILLER_113_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7072_ _7686_/CLK _7072_/D fanout599/X VGND VGND VPWR VPWR _7072_/Q sky130_fd_sc_hd__dfrtp_2
X_4284_ _4283_/X hold953/X _4294_/S VGND VGND VPWR VPWR _4284_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6023_ hold771/X _6041_/A1 _6028_/S VGND VGND VPWR VPWR _6023_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6925_ _4183_/A1 _6925_/D _6880_/X VGND VGND VPWR VPWR _6925_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_82_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6856_ _6969_/Q _6825_/A _6827_/B _6971_/Q VGND VGND VPWR VPWR _6856_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5807_ hold323/X _5843_/A1 _5812_/S VGND VGND VPWR VPWR _5807_/X sky130_fd_sc_hd__mux2_1
X_3999_ _7562_/Q _4547_/A _5984_/B _3998_/X VGND VGND VPWR VPWR _3999_/X sky130_fd_sc_hd__a31o_1
X_6787_ _6786_/X _6787_/A1 _6812_/S VGND VGND VPWR VPWR _7661_/D sky130_fd_sc_hd__mux2_1
XFILLER_183_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5738_ hold929/X _6044_/A1 _5740_/S VGND VGND VPWR VPWR _5738_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5669_ _5975_/B _5669_/B VGND VGND VPWR VPWR _5669_/Y sky130_fd_sc_hd__nand2_1
XFILLER_129_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7408_ _7408_/CLK _7408_/D fanout628/X VGND VGND VPWR VPWR _7408_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_191_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold450 hold450/A VGND VGND VPWR VPWR hold450/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 _7558_/Q VGND VGND VPWR VPWR hold461/X sky130_fd_sc_hd__dlygate4sd3_1
X_7339_ _7515_/CLK _7339_/D fanout621/X VGND VGND VPWR VPWR _7339_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_150_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold472 hold472/A VGND VGND VPWR VPWR hold472/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold483 _7712_/A VGND VGND VPWR VPWR hold483/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 _7090_/Q VGND VGND VPWR VPWR hold494/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1150 _7268_/Q VGND VGND VPWR VPWR _5646_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1161 _7289_/Q VGND VGND VPWR VPWR _5674_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1172 _5697_/X VGND VGND VPWR VPWR _7306_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1183 hold1640/X VGND VGND VPWR VPWR _4220_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_301 input97/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1194 _4374_/X VGND VGND VPWR VPWR _7079_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_312 _6809_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_323 _6694_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_334 _5789_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_345 _4172_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_356 hold571/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_367 _3713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_378 _3529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_389 _3584_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4971_ _4971_/A _4971_/B _4971_/C _4971_/D VGND VGND VPWR VPWR _4971_/Y sky130_fd_sc_hd__nand4_1
XFILLER_64_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6710_ _6700_/Y _6709_/Y _7036_/Q _6759_/D VGND VGND VPWR VPWR _6710_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_32_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3922_ _7175_/Q _6038_/B hold98/A _3712_/X _7205_/Q VGND VGND VPWR VPWR _3922_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_189_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7690_ _7690_/A VGND VGND VPWR VPWR _7690_/X sky130_fd_sc_hd__clkbuf_2
X_3853_ _7516_/Q _3555_/X _3704_/X _7196_/Q _3852_/X VGND VGND VPWR VPWR _3853_/X
+ sky130_fd_sc_hd__a221o_1
X_6641_ _7360_/Q _6454_/X _6469_/X _7336_/Q _6640_/X VGND VGND VPWR VPWR _6651_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_149_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6572_ _7589_/Q _6468_/X _6487_/X _7469_/Q _6561_/X VGND VGND VPWR VPWR _6572_/X
+ sky130_fd_sc_hd__a221o_1
X_3784_ _7064_/Q _3702_/X _3782_/X _3783_/X VGND VGND VPWR VPWR _3784_/X sky130_fd_sc_hd__a211o_1
XFILLER_118_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5523_ _5452_/A _5452_/B _5523_/A3 _4906_/A VGND VGND VPWR VPWR _5524_/D sky130_fd_sc_hd__a31oi_1
XFILLER_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5454_ _5454_/A _5454_/B VGND VGND VPWR VPWR _5455_/A sky130_fd_sc_hd__nor2_1
XFILLER_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4405_ hold549/X _4564_/A1 _4405_/S VGND VGND VPWR VPWR _4405_/X sky130_fd_sc_hd__mux2_1
X_5385_ _4769_/Y _4953_/C _4862_/Y _4867_/X VGND VGND VPWR VPWR _5385_/X sky130_fd_sc_hd__a211o_1
X_4336_ hold137/X _5869_/A1 _4339_/S VGND VGND VPWR VPWR _4336_/X sky130_fd_sc_hd__mux2_1
X_7124_ _7215_/CLK _7124_/D _6903_/A VGND VGND VPWR VPWR _7124_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_99_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7055_ _7231_/CLK _7055_/D fanout598/X VGND VGND VPWR VPWR _7055_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_86_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4267_ hold665/X _5988_/A1 _4275_/S VGND VGND VPWR VPWR _4267_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6006_ _6006_/A0 _6006_/A1 _6010_/S VGND VGND VPWR VPWR _6006_/X sky130_fd_sc_hd__mux2_1
X_4198_ _7298_/Q _4198_/B VGND VGND VPWR VPWR _4198_/X sky130_fd_sc_hd__and2_2
XFILLER_67_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6908_ _6911_/A _6908_/B VGND VGND VPWR VPWR _6908_/X sky130_fd_sc_hd__and2_1
XFILLER_35_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6839_ _6971_/Q _6839_/A2 _6839_/B1 _6970_/Q VGND VGND VPWR VPWR _6839_/X sky130_fd_sc_hd__a22o_1
XFILLER_11_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold280 hold280/A VGND VGND VPWR VPWR hold280/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold291 _7577_/Q VGND VGND VPWR VPWR hold291/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_120 _6151_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_131 _6371_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_142 _6454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_153 _6478_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_164 _6487_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_175 _6785_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_186 _6834_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_197 _6843_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5170_ _4619_/Y _4660_/C _4669_/Y _4912_/Y _4617_/X VGND VGND VPWR VPWR _5170_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4121_ _7619_/Q _7620_/Q _6107_/C VGND VGND VPWR VPWR _4121_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_68_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4052_ _4050_/X _4048_/Y _4052_/B1 _4051_/Y VGND VGND VPWR VPWR _6940_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput4 mask_rev_in[0] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4954_ _4966_/A _4957_/B _5021_/B _5389_/C VGND VGND VPWR VPWR _4955_/C sky130_fd_sc_hd__and4_1
X_3905_ _5682_/A _3905_/B _5669_/B VGND VGND VPWR VPWR _3905_/X sky130_fd_sc_hd__and3_1
X_7673_ _7676_/CLK _7673_/D _6815_/A VGND VGND VPWR VPWR _7673_/Q sky130_fd_sc_hd__dfrtp_1
X_4885_ _5143_/A _4983_/C VGND VGND VPWR VPWR _4885_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6624_ _7463_/Q _6464_/X _6479_/X _7543_/Q VGND VGND VPWR VPWR _6624_/X sky130_fd_sc_hd__a22o_1
XFILLER_165_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3836_ _7437_/Q _5840_/A _5984_/B _3832_/X _3835_/X VGND VGND VPWR VPWR _3837_/D
+ sky130_fd_sc_hd__a311o_1
XFILLER_192_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6555_ _7476_/Q _6441_/X _6482_/X _7484_/Q _6554_/X VGND VGND VPWR VPWR _6555_/X
+ sky130_fd_sc_hd__a221o_1
X_3767_ _7120_/Q _4541_/A _5680_/A _3579_/X _7438_/Q VGND VGND VPWR VPWR _3767_/X
+ sky130_fd_sc_hd__a32o_1
X_5506_ _5099_/Y _5297_/C _4985_/B _5095_/C _5297_/X VGND VGND VPWR VPWR _5506_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3698_ _3717_/B _4493_/C _4511_/C VGND VGND VPWR VPWR _4499_/A sky130_fd_sc_hd__and3_4
X_6486_ _6791_/C _6720_/C _6563_/C VGND VGND VPWR VPWR _6486_/X sky130_fd_sc_hd__and3_4
XFILLER_118_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput330 hold790/X VGND VGND VPWR VPWR hold791/A sky130_fd_sc_hd__buf_12
X_5437_ _4613_/X _5378_/Y _5408_/X _4847_/X _5436_/X VGND VGND VPWR VPWR _5437_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_160_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput341 hold712/X VGND VGND VPWR VPWR hold713/A sky130_fd_sc_hd__buf_12
XFILLER_10_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5368_ _4570_/Y _4622_/Y _4769_/Y _4685_/Y _4704_/D VGND VGND VPWR VPWR _5371_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7107_ _7130_/CLK _7107_/D fanout602/X VGND VGND VPWR VPWR _7107_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4319_ hold798/X _5999_/A1 _4321_/S VGND VGND VPWR VPWR _4319_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5299_ _5015_/Y _5018_/Y _5604_/B1 _5285_/X VGND VGND VPWR VPWR _5299_/X sky130_fd_sc_hd__a211o_1
XFILLER_19_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7038_ _7294_/CLK _7038_/D fanout597/X VGND VGND VPWR VPWR _7038_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire424 _4953_/Y VGND VGND VPWR VPWR _5572_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_183_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout590 input99/X VGND VGND VPWR VPWR _4992_/B sky130_fd_sc_hd__buf_4
XFILLER_80_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4670_ _4747_/B _5490_/C _5196_/A _5364_/B VGND VGND VPWR VPWR _4742_/D sky130_fd_sc_hd__nand4_1
XFILLER_186_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3621_ _3621_/A0 _3620_/X _3904_/S VGND VGND VPWR VPWR _3621_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6340_ _6330_/X _6158_/D _6329_/X _6331_/X _6339_/X VGND VGND VPWR VPWR _6340_/X
+ sky130_fd_sc_hd__a2111o_1
X_3552_ hold73/A _5768_/C _6002_/A VGND VGND VPWR VPWR _3552_/X sky130_fd_sc_hd__and3_4
XFILLER_174_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6271_ _6265_/X _6131_/B _6261_/X _6270_/X _6263_/X VGND VGND VPWR VPWR _6271_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_170_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3483_ hold132/X hold153/X _3508_/S VGND VGND VPWR VPWR _3483_/X sky130_fd_sc_hd__mux2_1
X_5222_ _5043_/B _5614_/B _5195_/X _5089_/A _4985_/B VGND VGND VPWR VPWR _5224_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_142_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5153_ _5153_/A _5358_/B _5153_/C VGND VGND VPWR VPWR _5162_/A sky130_fd_sc_hd__and3_1
X_4104_ _7258_/Q _7257_/Q _7256_/Q _4104_/D VGND VGND VPWR VPWR _4105_/S sky130_fd_sc_hd__and4b_1
X_5084_ _5131_/A _5131_/B _5137_/A VGND VGND VPWR VPWR _5084_/X sky130_fd_sc_hd__and3_1
XFILLER_56_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4035_ _7314_/Q hold37/A _4029_/X _4032_/X _4034_/X VGND VGND VPWR VPWR _4036_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_25_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5986_ hold339/X _6031_/A0 hold63/X VGND VGND VPWR VPWR _5986_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4937_ _4957_/B _5389_/C VGND VGND VPWR VPWR _4937_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_20 _4295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7656_ _7657_/CLK _7656_/D fanout608/X VGND VGND VPWR VPWR _7656_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_31 _3535_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4868_ _4943_/A _5389_/B _4926_/B VGND VGND VPWR VPWR _4906_/B sky130_fd_sc_hd__and3_1
XANTENNA_42 _3554_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_53 hold70/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6607_ _7486_/Q _6482_/X _6604_/X _6605_/X _6606_/X VGND VGND VPWR VPWR _6607_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA_64 _3569_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3819_ input14/X _3542_/X _3544_/X input29/X _3818_/X VGND VGND VPWR VPWR _3819_/X
+ sky130_fd_sc_hd__a221o_2
XANTENNA_75 _3704_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7587_ _7602_/CLK hold6/X fanout614/X VGND VGND VPWR VPWR _7587_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA_86 _6791_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4799_ _4799_/A _5476_/D _5024_/D VGND VGND VPWR VPWR _5233_/B sky130_fd_sc_hd__and3_2
XANTENNA_97 _6010_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6538_ _7436_/Q _6099_/B _6694_/C _6474_/A _7340_/Q VGND VGND VPWR VPWR _6538_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_119_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6469_ _6469_/A _6771_/C _6645_/C VGND VGND VPWR VPWR _6469_/X sky130_fd_sc_hd__and3_4
XFILLER_106_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput171 _4197_/X VGND VGND VPWR VPWR debug_in sky130_fd_sc_hd__buf_12
XFILLER_133_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput182 _3443_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[16] sky130_fd_sc_hd__buf_12
Xoutput193 _3433_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[26] sky130_fd_sc_hd__buf_12
XFILLER_121_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5840_ _5840_/A _5984_/B _6029_/B VGND VGND VPWR VPWR _5848_/S sky130_fd_sc_hd__and3_4
XFILLER_179_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5771_ _5843_/A1 hold355/X _5776_/S VGND VGND VPWR VPWR _5771_/X sky130_fd_sc_hd__mux2_1
X_7510_ _7566_/CLK _7510_/D fanout621/X VGND VGND VPWR VPWR _7510_/Q sky130_fd_sc_hd__dfrtp_2
X_4722_ _4722_/A _4722_/B _4722_/C VGND VGND VPWR VPWR _4724_/A sky130_fd_sc_hd__nor3_1
XFILLER_175_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7441_ _7617_/CLK _7441_/D fanout624/X VGND VGND VPWR VPWR _7441_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_30_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4653_ _5025_/B _5008_/C VGND VGND VPWR VPWR _4653_/Y sky130_fd_sc_hd__nand2_1
XFILLER_175_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput40 mgmt_gpio_in[13] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__clkbuf_1
X_3604_ _7417_/Q _5840_/A _3529_/X _3514_/X _7553_/Q VGND VGND VPWR VPWR _3604_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_162_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput51 mgmt_gpio_in[23] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__clkbuf_1
X_7372_ _7611_/CLK _7372_/D fanout621/X VGND VGND VPWR VPWR _7372_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_162_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput62 mgmt_gpio_in[33] VGND VGND VPWR VPWR input62/X sky130_fd_sc_hd__clkbuf_4
X_4584_ _4584_/A _4584_/B _4584_/C _4584_/D VGND VGND VPWR VPWR _4584_/Y sky130_fd_sc_hd__nand4_4
Xhold802 _7262_/Q VGND VGND VPWR VPWR hold802/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput73 pad_flash_io0_di VGND VGND VPWR VPWR _4190_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_128_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput84 spimemio_flash_csb VGND VGND VPWR VPWR input84/X sky130_fd_sc_hd__clkbuf_4
Xhold813 _7383_/Q VGND VGND VPWR VPWR hold813/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput95 usr1_vcc_pwrgood VGND VGND VPWR VPWR input95/X sky130_fd_sc_hd__clkbuf_4
Xhold824 _4262_/X VGND VGND VPWR VPWR _6996_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6323_ _7046_/Q _6231_/D _6166_/C _6309_/C _7164_/Q VGND VGND VPWR VPWR _6323_/X
+ sky130_fd_sc_hd__a32o_1
X_3535_ hold69/X _3559_/B _5682_/B VGND VGND VPWR VPWR _3535_/X sky130_fd_sc_hd__and3_4
Xhold835 _7561_/Q VGND VGND VPWR VPWR hold835/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 _4310_/X VGND VGND VPWR VPWR _7025_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap554 _3968_/S VGND VGND VPWR VPWR _3904_/S sky130_fd_sc_hd__buf_2
Xhold857 _7361_/Q VGND VGND VPWR VPWR hold857/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold868 _5794_/X VGND VGND VPWR VPWR _7393_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold879 _7519_/Q VGND VGND VPWR VPWR hold879/X sky130_fd_sc_hd__dlygate4sd3_1
X_3466_ _3470_/B _7256_/Q _7257_/Q VGND VGND VPWR VPWR _3469_/A sky130_fd_sc_hd__and3_1
X_6254_ _7431_/Q _6112_/X _6141_/X _7367_/Q VGND VGND VPWR VPWR _6254_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5205_ _4994_/X _5111_/D _5027_/X _4761_/A VGND VGND VPWR VPWR _5206_/C sky130_fd_sc_hd__a22oi_1
X_6185_ _6184_/X _6206_/A1 _6812_/S VGND VGND VPWR VPWR _6185_/X sky130_fd_sc_hd__mux2_1
Xhold1502 _7538_/Q VGND VGND VPWR VPWR hold555/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1513 _7653_/Q VGND VGND VPWR VPWR _6610_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5136_ _5512_/B _5291_/C _5137_/C VGND VGND VPWR VPWR _5138_/A sky130_fd_sc_hd__and3_1
Xhold1524 _7658_/Q VGND VGND VPWR VPWR _6712_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1535 _7134_/Q VGND VGND VPWR VPWR hold400/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1546 _7113_/Q VGND VGND VPWR VPWR hold1546/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1557 _4532_/X VGND VGND VPWR VPWR _7216_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5067_ _4756_/Y _4800_/Y _4953_/C _5066_/Y VGND VGND VPWR VPWR _5073_/C sky130_fd_sc_hd__o31ai_1
Xhold1568 _7270_/Q VGND VGND VPWR VPWR hold236/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1579 _7674_/Q VGND VGND VPWR VPWR _6838_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4018_ _7189_/Q _4499_/A _3780_/X input98/X _3975_/X VGND VGND VPWR VPWR _4018_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_708 _5926_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_719 _6464_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5969_ hold753/X _6041_/A1 _5974_/S VGND VGND VPWR VPWR _5969_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7708_ _7708_/A VGND VGND VPWR VPWR _7708_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7639_ _7657_/CLK _7639_/D fanout607/X VGND VGND VPWR VPWR _7639_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_180_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold109 _7369_/Q VGND VGND VPWR VPWR hold109/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_137_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6941_ _4183_/A1 _6941_/D _6896_/X VGND VGND VPWR VPWR _6941_/Q sky130_fd_sc_hd__dfrtp_1
X_6872_ _6899_/A _6907_/B VGND VGND VPWR VPWR _6872_/X sky130_fd_sc_hd__and2_1
XFILLER_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5823_ _5823_/A0 _6012_/A0 _5830_/S VGND VGND VPWR VPWR _7418_/D sky130_fd_sc_hd__mux2_1
XFILLER_167_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5754_ _5754_/A0 _6042_/A1 _5758_/S VGND VGND VPWR VPWR _5754_/X sky130_fd_sc_hd__mux2_1
X_4705_ _4760_/D _4706_/B _4760_/C _4706_/D VGND VGND VPWR VPWR _4813_/B sky130_fd_sc_hd__and4_1
X_5685_ hold303/X _6039_/A1 _5685_/S VGND VGND VPWR VPWR _5685_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7424_ _7445_/CLK _7424_/D fanout628/X VGND VGND VPWR VPWR _7424_/Q sky130_fd_sc_hd__dfrtp_4
X_4636_ _4785_/C _4785_/A _5046_/A _4786_/A VGND VGND VPWR VPWR _4637_/A sky130_fd_sc_hd__nand4_4
XFILLER_148_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold610 _7301_/Q VGND VGND VPWR VPWR hold610/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7355_ _7435_/CLK _7355_/D fanout623/X VGND VGND VPWR VPWR _7355_/Q sky130_fd_sc_hd__dfstp_1
Xhold621 _7368_/Q VGND VGND VPWR VPWR hold621/X sky130_fd_sc_hd__dlygate4sd3_1
X_4567_ _4948_/B _4959_/C VGND VGND VPWR VPWR _4704_/A sky130_fd_sc_hd__nand2_8
Xhold632 hold632/A VGND VGND VPWR VPWR hold632/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold643 hold643/A VGND VGND VPWR VPWR wb_dat_o[21] sky130_fd_sc_hd__buf_12
Xhold654 _5702_/X VGND VGND VPWR VPWR _7311_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6306_ _7473_/Q _6130_/X _6136_/X _7513_/Q _6305_/X VGND VGND VPWR VPWR _6306_/X
+ sky130_fd_sc_hd__a221o_1
Xmax_cap362 _4311_/S VGND VGND VPWR VPWR _4312_/S sky130_fd_sc_hd__clkbuf_2
X_3518_ _5682_/A _3622_/A hold23/X VGND VGND VPWR VPWR _4295_/A sky130_fd_sc_hd__and3_4
XFILLER_104_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold665 _7031_/Q VGND VGND VPWR VPWR hold665/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold676 _7283_/Q VGND VGND VPWR VPWR hold676/X sky130_fd_sc_hd__dlygate4sd3_1
X_7286_ _7286_/CLK _7286_/D fanout598/X VGND VGND VPWR VPWR _7688_/A sky130_fd_sc_hd__dfrtp_4
X_4498_ _4564_/A1 hold993/X _4498_/S VGND VGND VPWR VPWR _4498_/X sky130_fd_sc_hd__mux2_1
Xhold687 hold687/A VGND VGND VPWR VPWR wb_dat_o[4] sky130_fd_sc_hd__buf_12
XFILLER_143_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold698 hold698/A VGND VGND VPWR VPWR hold698/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6237_ _6231_/X _6233_/X _6236_/X _6159_/B VGND VGND VPWR VPWR _6237_/X sky130_fd_sc_hd__o31a_2
X_3449_ _7397_/Q VGND VGND VPWR VPWR _3449_/Y sky130_fd_sc_hd__inv_2
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ _7427_/Q _6112_/X _6115_/X _7387_/Q _6167_/X VGND VGND VPWR VPWR _6168_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1310 _7437_/Q VGND VGND VPWR VPWR hold1310/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1321 _5763_/X VGND VGND VPWR VPWR _7365_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1332 _3840_/X VGND VGND VPWR VPWR _6945_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1343 _7104_/Q VGND VGND VPWR VPWR hold716/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5119_ _5401_/A _5038_/B _5110_/X _5118_/Y VGND VGND VPWR VPWR _5119_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1354 _5736_/X VGND VGND VPWR VPWR _7341_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6099_ _7632_/Q _6099_/B VGND VGND VPWR VPWR _6099_/Y sky130_fd_sc_hd__nand2_1
XFILLER_27_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1365 _7565_/Q VGND VGND VPWR VPWR hold673/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1376 _5806_/X VGND VGND VPWR VPWR _7403_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1387 _7451_/Q VGND VGND VPWR VPWR hold996/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1398 _4508_/X VGND VGND VPWR VPWR _7196_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_505 input13/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_516 _7714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_527 input78/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_538 input81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_549 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5470_ _4761_/A _4758_/X _5089_/A _4994_/X _5469_/X VGND VGND VPWR VPWR _5471_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4421_ _5789_/A1 hold337/X _4423_/S VGND VGND VPWR VPWR _4421_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7140_ _7680_/CLK _7140_/D _6886_/A VGND VGND VPWR VPWR _7140_/Q sky130_fd_sc_hd__dfrtp_4
X_4352_ _4547_/A _5682_/A _5659_/C _5680_/C VGND VGND VPWR VPWR _4357_/S sky130_fd_sc_hd__and4_4
XFILLER_125_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout408 _3573_/C VGND VGND VPWR VPWR _5669_/B sky130_fd_sc_hd__buf_6
X_7071_ _7312_/CLK _7071_/D _6891_/A VGND VGND VPWR VPWR _7071_/Q sky130_fd_sc_hd__dfrtp_4
X_4283_ hold727/X _6041_/A1 _4293_/S VGND VGND VPWR VPWR _4283_/X sky130_fd_sc_hd__mux2_1
Xfanout419 _6611_/S VGND VGND VPWR VPWR _6812_/S sky130_fd_sc_hd__buf_8
XFILLER_59_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6022_ hold353/X _6031_/A0 _6028_/S VGND VGND VPWR VPWR _6022_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6924_ _7258_/CLK _6924_/D _6879_/X VGND VGND VPWR VPWR hold21/A sky130_fd_sc_hd__dfrtp_2
XFILLER_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6855_ _4118_/B _6965_/D _6854_/Y _6855_/B1 VGND VGND VPWR VPWR _7680_/D sky130_fd_sc_hd__o31ai_2
X_5806_ hold977/X _6040_/A1 _5812_/S VGND VGND VPWR VPWR _5806_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6786_ _6785_/X _6786_/A1 _6811_/S VGND VGND VPWR VPWR _6786_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3998_ input71/X _4275_/S _3623_/X _7618_/Q _3997_/X VGND VGND VPWR VPWR _3998_/X
+ sky130_fd_sc_hd__a221o_1
X_5737_ hold234/X _5935_/A1 _5740_/S VGND VGND VPWR VPWR _5737_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5668_ _5682_/A _5661_/A _5669_/B hold904/X VGND VGND VPWR VPWR _5668_/X sky130_fd_sc_hd__a31o_1
XFILLER_135_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7407_ _7599_/CLK _7407_/D fanout629/X VGND VGND VPWR VPWR _7407_/Q sky130_fd_sc_hd__dfrtp_1
X_4619_ _4706_/D _4836_/A _4604_/Y _5007_/D VGND VGND VPWR VPWR _4619_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_151_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5599_ _5580_/X _5587_/Y _5598_/Y _5578_/X VGND VGND VPWR VPWR _5599_/X sky130_fd_sc_hd__a211o_1
XFILLER_2_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold440 _7205_/Q VGND VGND VPWR VPWR hold440/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7338_ _7430_/CLK _7338_/D fanout627/X VGND VGND VPWR VPWR _7338_/Q sky130_fd_sc_hd__dfstp_1
Xhold451 hold451/A VGND VGND VPWR VPWR hold451/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 _5980_/X VGND VGND VPWR VPWR _7558_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold473 _7210_/Q VGND VGND VPWR VPWR hold473/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 _5692_/X VGND VGND VPWR VPWR _7302_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold495 _4387_/X VGND VGND VPWR VPWR _7090_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7269_ _7291_/CLK _7269_/D fanout596/X VGND VGND VPWR VPWR _7269_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_38_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1140 hold1572/X VGND VGND VPWR VPWR _6012_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1151 _5646_/X VGND VGND VPWR VPWR _7268_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1162 _5674_/X VGND VGND VPWR VPWR _7289_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1173 _7111_/Q VGND VGND VPWR VPWR _4413_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1184 _7285_/Q VGND VGND VPWR VPWR _5667_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_302 input164/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1195 _7227_/Q VGND VGND VPWR VPWR _4545_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_313 _6809_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_324 _6694_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_335 _5869_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_346 hold9/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_357 hold615/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_368 _3905_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_379 _3531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4970_ _4625_/Y _4800_/Y _5407_/D _4969_/Y VGND VGND VPWR VPWR _4971_/B sky130_fd_sc_hd__o31a_1
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3921_ _7315_/Q _5993_/B _5682_/C _3915_/X _3920_/X VGND VGND VPWR VPWR _3921_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_189_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6640_ _7520_/Q _6645_/B _6536_/C _6458_/X _7424_/Q VGND VGND VPWR VPWR _6640_/X
+ sky130_fd_sc_hd__a32o_1
X_3852_ _7268_/Q _3674_/X _3711_/X _7186_/Q _3851_/X VGND VGND VPWR VPWR _3852_/X
+ sky130_fd_sc_hd__a221o_1
X_6571_ _7517_/Q _6455_/C _6562_/C _6570_/X VGND VGND VPWR VPWR _6571_/X sky130_fd_sc_hd__a31o_1
X_3783_ _7129_/Q _6861_/A _4553_/B _3562_/X _7501_/Q VGND VGND VPWR VPWR _3783_/X
+ sky130_fd_sc_hd__a32o_1
X_5522_ _5614_/C _4972_/C _5280_/X _5407_/Y _5521_/X VGND VGND VPWR VPWR _5522_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_117_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5453_ _4946_/A _4943_/B _5265_/X _5452_/X _5382_/X VGND VGND VPWR VPWR _5454_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_133_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4404_ hold716/X _5673_/A1 _4405_/S VGND VGND VPWR VPWR _7104_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_42_csclk _7352_/CLK VGND VGND VPWR VPWR _7553_/CLK sky130_fd_sc_hd__clkbuf_16
X_5384_ _5384_/A _5384_/B VGND VGND VPWR VPWR _5442_/B sky130_fd_sc_hd__nor2_1
XFILLER_99_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7123_ _7160_/CLK _7123_/D _6891_/A VGND VGND VPWR VPWR _7123_/Q sky130_fd_sc_hd__dfstp_2
X_4335_ _4335_/A0 _5697_/A0 _4339_/S VGND VGND VPWR VPWR _7046_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7054_ _7289_/CLK _7054_/D fanout598/X VGND VGND VPWR VPWR _7054_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_140_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4266_ _4265_/X hold638/X _4274_/S VGND VGND VPWR VPWR _4266_/X sky130_fd_sc_hd__mux2_1
X_6005_ hold761/X _6041_/A1 _6010_/S VGND VGND VPWR VPWR _6005_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_57_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7497_/CLK sky130_fd_sc_hd__clkbuf_16
X_4197_ _4197_/A input1/X VGND VGND VPWR VPWR _4197_/X sky130_fd_sc_hd__and2_1
XFILLER_67_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6907_ _6907_/A _6907_/B VGND VGND VPWR VPWR _6907_/X sky130_fd_sc_hd__and2_1
XFILLER_23_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6838_ _6838_/A0 _6837_/X _6853_/S VGND VGND VPWR VPWR _7674_/D sky130_fd_sc_hd__mux2_1
XFILLER_11_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6769_ _7227_/Q _6463_/X _6807_/A2 _7237_/Q _6768_/X VGND VGND VPWR VPWR _6775_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_108_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold270 _5834_/X VGND VGND VPWR VPWR _7428_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold281 hold281/A VGND VGND VPWR VPWR hold281/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 _6001_/X VGND VGND VPWR VPWR _7577_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_110 _6133_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_121 _6152_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_132 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_143 _6454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_154 _6479_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_165 _6533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_176 _6785_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_187 _6837_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_198 _6843_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4120_ _7621_/Q _7622_/Q VGND VGND VPWR VPWR _6107_/C sky130_fd_sc_hd__nor2_1
XFILLER_96_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4051_ _4048_/B _3419_/Y _4049_/B VGND VGND VPWR VPWR _4051_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_83_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput5 mask_rev_in[10] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4953_ _4953_/A _4953_/B _4953_/C _4953_/D VGND VGND VPWR VPWR _4953_/Y sky130_fd_sc_hd__nor4_1
XFILLER_189_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3904_ _3904_/A0 _3903_/X _3904_/S VGND VGND VPWR VPWR _6944_/D sky130_fd_sc_hd__mux2_1
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7672_ _7672_/CLK _7672_/D fanout635/X VGND VGND VPWR VPWR _7672_/Q sky130_fd_sc_hd__dfrtp_1
X_4884_ _4884_/A _5096_/A _5096_/B _5096_/C VGND VGND VPWR VPWR _4884_/Y sky130_fd_sc_hd__nor4_2
XFILLER_60_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6623_ _6623_/A _6623_/B _6623_/C _6623_/D VGND VGND VPWR VPWR _6633_/C sky130_fd_sc_hd__nor4_1
X_3835_ _7119_/Q _4541_/A _5680_/A _3833_/X _3834_/X VGND VGND VPWR VPWR _3835_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_165_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6554_ _7556_/Q _6453_/X _6474_/B _7596_/Q _6553_/X VGND VGND VPWR VPWR _6554_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_192_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3766_ _7228_/Q _4541_/A _4541_/B _3556_/X _7430_/Q VGND VGND VPWR VPWR _3774_/C
+ sky130_fd_sc_hd__a32o_1
X_5505_ _5313_/B _5110_/C _5416_/X _5425_/B _5290_/X VGND VGND VPWR VPWR _5625_/B
+ sky130_fd_sc_hd__a311o_1
X_6485_ _7631_/Q _6485_/B _6645_/B _6563_/C VGND VGND VPWR VPWR _6485_/X sky130_fd_sc_hd__and4_4
XFILLER_173_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3697_ _5768_/C hold98/A _5768_/B VGND VGND VPWR VPWR _3697_/X sky130_fd_sc_hd__and3_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5436_ _6829_/D _5602_/C _5434_/X _5501_/B VGND VGND VPWR VPWR _5436_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_145_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput320 hold606/X VGND VGND VPWR VPWR hold607/A sky130_fd_sc_hd__buf_12
Xoutput331 hold645/X VGND VGND VPWR VPWR hold646/A sky130_fd_sc_hd__buf_12
XFILLER_160_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput342 hold706/X VGND VGND VPWR VPWR hold707/A sky130_fd_sc_hd__buf_12
XFILLER_161_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5367_ _5358_/A _5490_/C _5153_/C _5366_/X _5365_/X VGND VGND VPWR VPWR _5367_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_87_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7106_ _7130_/CLK _7106_/D fanout602/X VGND VGND VPWR VPWR _7106_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4318_ hold363/X _5935_/A1 _4321_/S VGND VGND VPWR VPWR _4318_/X sky130_fd_sc_hd__mux2_1
X_5298_ _5291_/C _5130_/B _5249_/C _5297_/X VGND VGND VPWR VPWR _5298_/X sky130_fd_sc_hd__a31o_1
XFILLER_87_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7037_ _7231_/CLK _7037_/D fanout597/X VGND VGND VPWR VPWR _7037_/Q sky130_fd_sc_hd__dfrtp_1
X_4249_ _4308_/A1 _6006_/A1 _4257_/S VGND VGND VPWR VPWR _4249_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout580 _4884_/Y VGND VGND VPWR VPWR _5311_/C sky130_fd_sc_hd__buf_6
Xfanout591 _6911_/A VGND VGND VPWR VPWR _6886_/A sky130_fd_sc_hd__buf_6
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3620_ _3618_/Y _6949_/Q _3967_/S VGND VGND VPWR VPWR _3620_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3551_ hold69/X _3559_/B _3622_/A _3622_/B VGND VGND VPWR VPWR _3551_/Y sky130_fd_sc_hd__nor4_2
XFILLER_155_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6270_ _7551_/Q _6151_/X _6269_/X _6268_/X _6267_/X VGND VGND VPWR VPWR _6270_/X
+ sky130_fd_sc_hd__a2111o_1
X_3482_ _7258_/Q _7257_/Q _7256_/Q VGND VGND VPWR VPWR _3968_/S sky130_fd_sc_hd__nor3_2
XFILLER_142_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5221_ _5221_/A _5221_/B _5536_/A VGND VGND VPWR VPWR _5224_/A sky130_fd_sc_hd__nand3_1
XFILLER_142_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5152_ _5189_/A _4992_/B _5146_/A _5181_/C VGND VGND VPWR VPWR _5153_/C sky130_fd_sc_hd__a31o_2
XFILLER_69_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4103_ input58/X _3968_/S _4104_/D _4102_/Y VGND VGND VPWR VPWR _6916_/D sky130_fd_sc_hd__a31o_1
XFILLER_29_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5083_ _5079_/Y _5081_/X _5082_/Y _4975_/Y VGND VGND VPWR VPWR _5083_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_111_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4034_ _7458_/Q _3549_/X _3715_/X _7106_/Q _4033_/X VGND VGND VPWR VPWR _4034_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5985_ _5985_/A0 hold44/X hold63/X VGND VGND VPWR VPWR hold64/A sky130_fd_sc_hd__mux2_1
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4936_ _4936_/A _4936_/B _4936_/C VGND VGND VPWR VPWR _4941_/B sky130_fd_sc_hd__nand3_1
XFILLER_178_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_10 hold24/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7655_ _7657_/CLK _7655_/D fanout608/X VGND VGND VPWR VPWR _7655_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_21 _5723_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4867_ _5000_/C _4777_/Y _4830_/Y _4859_/Y VGND VGND VPWR VPWR _4867_/X sky130_fd_sc_hd__a211o_2
XANTENNA_32 hold75/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_43 _3555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6606_ _7494_/Q _6694_/B _6720_/D _6474_/B _7598_/Q VGND VGND VPWR VPWR _6606_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_54 hold70/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3818_ _7232_/Q _5993_/A _5678_/B _3530_/X hold46/A VGND VGND VPWR VPWR _3818_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_193_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_65 _3569_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7586_ _7586_/CLK _7586_/D fanout625/X VGND VGND VPWR VPWR _7586_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA_76 _3780_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4798_ _5182_/A _4797_/X _4992_/B VGND VGND VPWR VPWR _4798_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_87 _6771_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_98 _6010_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6537_ _7500_/Q _6791_/C _6720_/C _6720_/D VGND VGND VPWR VPWR _6537_/X sky130_fd_sc_hd__and4_1
XFILLER_192_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3749_ _7590_/Q _6011_/A _3712_/X _7208_/Q _3748_/X VGND VGND VPWR VPWR _3749_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6468_ _6791_/B _6469_/A _6645_/C VGND VGND VPWR VPWR _6468_/X sky130_fd_sc_hd__and3_4
XFILLER_97_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5419_ _5452_/B _5040_/C _5313_/A _5110_/C _5291_/C VGND VGND VPWR VPWR _5425_/A
+ sky130_fd_sc_hd__o311a_1
X_6399_ _6392_/X _6394_/X _6398_/X _6159_/B VGND VGND VPWR VPWR _6399_/X sky130_fd_sc_hd__o31a_1
Xoutput172 _7688_/X VGND VGND VPWR VPWR irq[0] sky130_fd_sc_hd__buf_12
XFILLER_161_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput183 _3442_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[17] sky130_fd_sc_hd__buf_12
Xoutput194 _3432_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[27] sky130_fd_sc_hd__buf_12
XFILLER_102_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5770_ _6040_/A1 hold898/X _5776_/S VGND VGND VPWR VPWR _5770_/X sky130_fd_sc_hd__mux2_1
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4721_ _4721_/A _4721_/B _5156_/A _5156_/B VGND VGND VPWR VPWR _4722_/C sky130_fd_sc_hd__nand4_1
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7440_ _7568_/CLK _7440_/D fanout623/X VGND VGND VPWR VPWR _7440_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_147_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4652_ _5015_/C _5017_/B VGND VGND VPWR VPWR _5108_/B sky130_fd_sc_hd__and2b_4
XFILLER_147_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput30 mask_rev_in[4] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__clkbuf_1
X_3603_ _7279_/Q _3573_/C _5680_/A _3567_/X _7345_/Q VGND VGND VPWR VPWR _3603_/X
+ sky130_fd_sc_hd__a32o_1
X_7371_ _7611_/CLK _7371_/D fanout621/X VGND VGND VPWR VPWR _7371_/Q sky130_fd_sc_hd__dfstp_1
Xinput41 mgmt_gpio_in[14] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__clkbuf_4
X_4583_ _4584_/A _4584_/B _4584_/C _4584_/D VGND VGND VPWR VPWR _4785_/C sky130_fd_sc_hd__and4_4
Xinput52 mgmt_gpio_in[24] VGND VGND VPWR VPWR input52/X sky130_fd_sc_hd__buf_2
XFILLER_116_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput63 mgmt_gpio_in[34] VGND VGND VPWR VPWR _4196_/A sky130_fd_sc_hd__buf_4
Xmax_cap500 _5146_/C VGND VGND VPWR VPWR _5137_/A sky130_fd_sc_hd__clkbuf_2
Xhold803 _5639_/X VGND VGND VPWR VPWR _7262_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput74 pad_flash_io1_di VGND VGND VPWR VPWR _4191_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6322_ _7224_/Q _6166_/B _6427_/A3 _6432_/A3 _7096_/Q VGND VGND VPWR VPWR _6322_/X
+ sky130_fd_sc_hd__a32o_1
Xhold814 _5783_/X VGND VGND VPWR VPWR _7383_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3534_ _4229_/S hold22/X hold128/X _3622_/A VGND VGND VPWR VPWR _5682_/B sky130_fd_sc_hd__o211a_4
Xhold825 _7569_/Q VGND VGND VPWR VPWR hold825/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput85 spimemio_flash_io0_do VGND VGND VPWR VPWR input85/X sky130_fd_sc_hd__clkbuf_4
Xinput96 usr1_vdd_pwrgood VGND VGND VPWR VPWR input96/X sky130_fd_sc_hd__clkbuf_4
Xhold836 _5983_/X VGND VGND VPWR VPWR _7561_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 _7612_/Q VGND VGND VPWR VPWR hold847/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold858 _5758_/X VGND VGND VPWR VPWR _7361_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6253_ _6252_/X _6253_/A1 _6812_/S VGND VGND VPWR VPWR _7641_/D sky130_fd_sc_hd__mux2_1
Xhold869 _7425_/Q VGND VGND VPWR VPWR hold869/X sky130_fd_sc_hd__dlygate4sd3_1
X_3465_ _6913_/Q _6914_/Q VGND VGND VPWR VPWR _3470_/B sky130_fd_sc_hd__nand2b_1
XFILLER_88_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5204_ _4625_/Y _5585_/A1 _5011_/B _4984_/Y _5009_/Y VGND VGND VPWR VPWR _5206_/B
+ sky130_fd_sc_hd__o32a_1
X_6184_ _7637_/Q _6109_/X _6183_/X _6686_/S VGND VGND VPWR VPWR _6184_/X sky130_fd_sc_hd__o22a_1
Xhold1503 _7232_/Q VGND VGND VPWR VPWR hold471/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5135_ _4756_/Y _4888_/Y _5132_/Y _5514_/C VGND VGND VPWR VPWR _5138_/C sky130_fd_sc_hd__o211ai_1
XFILLER_29_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1514 _6586_/X VGND VGND VPWR VPWR _7653_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1525 _6712_/X VGND VGND VPWR VPWR _7658_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1536 _7402_/Q VGND VGND VPWR VPWR hold451/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1547 _4415_/X VGND VGND VPWR VPWR _7113_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1558 hold79/A VGND VGND VPWR VPWR _4060_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5066_ _5066_/A _5066_/B _5066_/C VGND VGND VPWR VPWR _5066_/Y sky130_fd_sc_hd__nor3_1
Xhold1569 hold65/A VGND VGND VPWR VPWR _6850_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_4017_ _7036_/Q _5682_/C _4505_/B _3584_/X _7578_/Q VGND VGND VPWR VPWR _4017_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_84_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_709 _6039_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5968_ hold178/X _6031_/A0 _5974_/S VGND VGND VPWR VPWR _5968_/X sky130_fd_sc_hd__mux2_1
X_7707_ _7707_/A VGND VGND VPWR VPWR _7707_/X sky130_fd_sc_hd__clkbuf_1
X_4919_ _4923_/B _5452_/A _4925_/C VGND VGND VPWR VPWR _4921_/A sky130_fd_sc_hd__and3_1
XFILLER_178_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5899_ hold233/X _6043_/A1 hold25/X VGND VGND VPWR VPWR _5899_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7638_ _7657_/CLK _7638_/D fanout606/X VGND VGND VPWR VPWR _7638_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_166_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7569_ _7569_/CLK _7569_/D fanout614/X VGND VGND VPWR VPWR _7569_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6940_ _6950_/CLK _6940_/D _6895_/X VGND VGND VPWR VPWR _6940_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_66_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6871_ _6899_/A _6907_/B VGND VGND VPWR VPWR _6871_/X sky130_fd_sc_hd__and2_1
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5822_ hold24/X _5840_/A _6029_/B VGND VGND VPWR VPWR _5830_/S sky130_fd_sc_hd__and3_4
XFILLER_179_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5753_ hold321/X _5843_/A1 _5758_/S VGND VGND VPWR VPWR _5753_/X sky130_fd_sc_hd__mux2_1
X_4704_ _4704_/A _5404_/C _4704_/C _4704_/D VGND VGND VPWR VPWR _4704_/Y sky130_fd_sc_hd__nor4_1
XFILLER_148_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5684_ hold151/X _6031_/A0 _5685_/S VGND VGND VPWR VPWR _5684_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7423_ _7568_/CLK _7423_/D fanout623/X VGND VGND VPWR VPWR _7423_/Q sky130_fd_sc_hd__dfrtp_4
X_4635_ _5046_/A _4786_/A VGND VGND VPWR VPWR _5027_/D sky130_fd_sc_hd__nand2_2
XFILLER_135_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold600 _6997_/Q VGND VGND VPWR VPWR hold600/X sky130_fd_sc_hd__dlygate4sd3_1
X_7354_ _7613_/CLK _7354_/D fanout626/X VGND VGND VPWR VPWR _7354_/Q sky130_fd_sc_hd__dfstp_2
Xhold611 _5691_/X VGND VGND VPWR VPWR _7301_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4566_ _4948_/B _4959_/C VGND VGND VPWR VPWR _5316_/A sky130_fd_sc_hd__and2_4
Xhold622 _5766_/X VGND VGND VPWR VPWR _7368_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 hold633/A VGND VGND VPWR VPWR wb_dat_o[30] sky130_fd_sc_hd__buf_12
X_6305_ _7529_/Q _6309_/B _6334_/C _6144_/X _7545_/Q VGND VGND VPWR VPWR _6305_/X
+ sky130_fd_sc_hd__a32o_1
Xhold644 hold644/A VGND VGND VPWR VPWR hold644/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3517_ _3622_/A hold23/X VGND VGND VPWR VPWR _3581_/B sky130_fd_sc_hd__and2_4
XFILLER_104_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7285_ _7307_/CLK _7285_/D _6886_/A VGND VGND VPWR VPWR _7285_/Q sky130_fd_sc_hd__dfrtp_1
Xhold655 hold655/A VGND VGND VPWR VPWR hold655/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4497_ _6865_/A1 _4497_/A1 _4498_/S VGND VGND VPWR VPWR _4497_/X sky130_fd_sc_hd__mux2_1
Xhold666 _4317_/X VGND VGND VPWR VPWR _7031_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 _5664_/X VGND VGND VPWR VPWR _7283_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold688 _7094_/Q VGND VGND VPWR VPWR hold688/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold699 hold699/A VGND VGND VPWR VPWR wb_dat_o[18] sky130_fd_sc_hd__buf_12
X_6236_ _7350_/Q wire455/X _6234_/X _6235_/X VGND VGND VPWR VPWR _6236_/X sky130_fd_sc_hd__a211o_1
XFILLER_103_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3448_ _7405_/Q VGND VGND VPWR VPWR _3448_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6167_ _7323_/Q _6231_/D _6145_/C _6077_/X _7379_/Q VGND VGND VPWR VPWR _6167_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1300 _7405_/Q VGND VGND VPWR VPWR hold1300/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1311 _5844_/X VGND VGND VPWR VPWR _7437_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1322 _7443_/Q VGND VGND VPWR VPWR hold983/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _4949_/Y _5039_/Y _5090_/Y _5004_/Y _5117_/Y VGND VGND VPWR VPWR _5118_/Y
+ sky130_fd_sc_hd__o221ai_1
Xhold1333 _7261_/Q VGND VGND VPWR VPWR hold1333/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1344 _7515_/Q VGND VGND VPWR VPWR hold982/A sky130_fd_sc_hd__dlygate4sd3_1
X_6098_ _7141_/Q _6099_/B _6093_/X _7632_/Q VGND VGND VPWR VPWR _6098_/Y sky130_fd_sc_hd__a211oi_1
Xhold1355 _6948_/Q VGND VGND VPWR VPWR _3621_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1366 _7573_/Q VGND VGND VPWR VPWR hold1366/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1377 _7435_/Q VGND VGND VPWR VPWR hold995/A sky130_fd_sc_hd__dlygate4sd3_1
X_5049_ _5011_/A _4823_/Y _5009_/Y _5043_/Y _5048_/Y VGND VGND VPWR VPWR _5050_/C
+ sky130_fd_sc_hd__o311ai_1
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1388 _7124_/Q VGND VGND VPWR VPWR hold717/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1399 _7530_/Q VGND VGND VPWR VPWR hold520/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_506 input46/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_517 _7714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_528 input78/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_539 input81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4420_ _5761_/A1 hold403/X _4423_/S VGND VGND VPWR VPWR _4420_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_702 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4351_ _5926_/A0 hold431/X _4351_/S VGND VGND VPWR VPWR _4351_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout409 hold55/X VGND VGND VPWR VPWR _3573_/C sky130_fd_sc_hd__buf_8
XFILLER_113_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7070_ _7254_/CLK _7070_/D fanout617/X VGND VGND VPWR VPWR _7070_/Q sky130_fd_sc_hd__dfrtp_2
X_4282_ _4281_/X hold991/X _4292_/S VGND VGND VPWR VPWR _4282_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6021_ hold504/X _6039_/A1 _6028_/S VGND VGND VPWR VPWR _7594_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6923_ _7258_/CLK _6923_/D _6878_/X VGND VGND VPWR VPWR _6923_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6854_ _6854_/A _6854_/B VGND VGND VPWR VPWR _6854_/Y sky130_fd_sc_hd__nand2_2
XFILLER_22_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5805_ hold451/X _6003_/A1 _5812_/S VGND VGND VPWR VPWR _5805_/X sky130_fd_sc_hd__mux2_1
X_6785_ wire373/X _6784_/Y _7039_/Q _6478_/Y VGND VGND VPWR VPWR _6785_/X sky130_fd_sc_hd__o2bb2a_2
X_3997_ _7051_/Q _5680_/B _5678_/B _6972_/Q _3560_/X VGND VGND VPWR VPWR _3997_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5736_ _5736_/A0 _6006_/A1 _5740_/S VGND VGND VPWR VPWR _5736_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5667_ _5667_/A0 _5697_/A0 _5667_/S VGND VGND VPWR VPWR _5667_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7406_ _7557_/CLK _7406_/D fanout627/X VGND VGND VPWR VPWR _7406_/Q sky130_fd_sc_hd__dfrtp_2
X_4618_ _5000_/C _4568_/Y _4836_/A _4604_/Y _5007_/D VGND VGND VPWR VPWR _4738_/B
+ sky130_fd_sc_hd__o311a_2
XFILLER_135_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5598_ _5591_/X _5597_/X _5589_/Y VGND VGND VPWR VPWR _5598_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_190_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold430 _6025_/X VGND VGND VPWR VPWR _7598_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7337_ _7553_/CLK _7337_/D fanout622/X VGND VGND VPWR VPWR _7337_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_151_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4549_ hold742/X _6863_/A1 _4552_/S VGND VGND VPWR VPWR _4549_/X sky130_fd_sc_hd__mux2_1
Xhold441 _4519_/X VGND VGND VPWR VPWR _7205_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 hold452/A VGND VGND VPWR VPWR hold452/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold463 _7175_/Q VGND VGND VPWR VPWR hold463/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold474 _4525_/X VGND VGND VPWR VPWR _7210_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 _7488_/Q VGND VGND VPWR VPWR hold485/X sky130_fd_sc_hd__dlygate4sd3_1
X_7268_ _7291_/CLK _7268_/D fanout596/X VGND VGND VPWR VPWR _7268_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_104_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold496 _7560_/Q VGND VGND VPWR VPWR hold496/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6219_ _7357_/Q _6138_/X _6153_/X _7565_/Q _6218_/X VGND VGND VPWR VPWR _6219_/X
+ sky130_fd_sc_hd__a221o_1
X_7199_ _7685_/CLK _7199_/D fanout617/X VGND VGND VPWR VPWR _7199_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1130 _4557_/X VGND VGND VPWR VPWR _7237_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1141 hold1526/X VGND VGND VPWR VPWR _5841_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1152 _7685_/Q VGND VGND VPWR VPWR _6865_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_161_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1163 _7197_/Q VGND VGND VPWR VPWR _4509_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_161_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1174 _4413_/X VGND VGND VPWR VPWR _7111_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1185 _5667_/X VGND VGND VPWR VPWR _7285_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1196 _4545_/X VGND VGND VPWR VPWR _7227_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_303 _4116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_314 _4505_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_325 _6694_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_336 _6031_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_347 hold44/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_358 hold676/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_369 _3514_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3920_ _7282_/Q _5993_/B _6002_/B _3918_/X _3919_/X VGND VGND VPWR VPWR _3920_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_17_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3851_ _7038_/Q _5678_/C _4505_/B _3850_/X VGND VGND VPWR VPWR _3851_/X sky130_fd_sc_hd__a31o_1
XFILLER_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6570_ _7421_/Q _6458_/X _6567_/X _6569_/X VGND VGND VPWR VPWR _6570_/X sky130_fd_sc_hd__a211o_1
X_3782_ _7054_/Q _4481_/A _4553_/B _3781_/X VGND VGND VPWR VPWR _3782_/X sky130_fd_sc_hd__a31o_1
X_5521_ _5021_/B _5404_/B _5452_/B _4961_/A _4963_/X VGND VGND VPWR VPWR _5521_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_157_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5452_ _5452_/A _5452_/B _5452_/C VGND VGND VPWR VPWR _5452_/X sky130_fd_sc_hd__and3_1
XFILLER_117_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4403_ _4403_/A0 _6864_/A1 _4405_/S VGND VGND VPWR VPWR _4403_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5383_ _5181_/C _5021_/B _4935_/C _5389_/B VGND VGND VPWR VPWR _5384_/B sky130_fd_sc_hd__o211a_1
X_7122_ _7312_/CLK _7122_/D _6891_/A VGND VGND VPWR VPWR _7122_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_132_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4334_ _5680_/A _5678_/C _5680_/C VGND VGND VPWR VPWR _4339_/S sky130_fd_sc_hd__and3_2
XFILLER_99_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7053_ _7459_/CLK _7053_/D fanout600/X VGND VGND VPWR VPWR _7053_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_86_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4265_ hold366/X _5843_/A1 _4275_/S VGND VGND VPWR VPWR _4265_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6004_ hold160/X _6031_/A0 _6010_/S VGND VGND VPWR VPWR _6004_/X sky130_fd_sc_hd__mux2_1
X_4196_ _4196_/A _4196_/B VGND VGND VPWR VPWR _4196_/X sky130_fd_sc_hd__and2_1
XFILLER_55_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6906_ _6911_/A _6911_/B VGND VGND VPWR VPWR _6906_/X sky130_fd_sc_hd__and2_1
XFILLER_23_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6837_ _6969_/Q _6837_/A2 _6837_/B1 wire537/X _6836_/X VGND VGND VPWR VPWR _6837_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_168_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6768_ _7167_/Q _6469_/X _6479_/X _7222_/Q VGND VGND VPWR VPWR _6768_/X sky130_fd_sc_hd__a22o_1
XFILLER_136_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5719_ hold286/X _5935_/A1 _5722_/S VGND VGND VPWR VPWR _5719_/X sky130_fd_sc_hd__mux2_1
X_6699_ _7086_/Q _6458_/X _6459_/X _7116_/Q _6698_/X VGND VGND VPWR VPWR _6700_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_149_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold260 _7287_/Q VGND VGND VPWR VPWR hold260/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold271 _7318_/Q VGND VGND VPWR VPWR hold271/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 _7609_/Q VGND VGND VPWR VPWR hold282/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 hold293/A VGND VGND VPWR VPWR hold293/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_100 _6516_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_111 _6136_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_122 _6157_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_133 _6444_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_144 _6454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_155 _6482_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_166 _6533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_177 _6831_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_188 _6837_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_199 _6843_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4050_ _6940_/Q _6939_/Q _4049_/B _4049_/Y VGND VGND VPWR VPWR _4050_/X sky130_fd_sc_hd__o31a_1
Xinput6 mask_rev_in[11] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4952_ _4767_/Y _4945_/Y _4951_/Y _4947_/Y VGND VGND VPWR VPWR _4955_/D sky130_fd_sc_hd__o211ai_1
XFILLER_51_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3903_ _3902_/Y _3903_/A1 _3967_/S VGND VGND VPWR VPWR _3903_/X sky130_fd_sc_hd__mux2_1
X_7671_ _7676_/CLK _7671_/D VGND VGND VPWR VPWR _7671_/Q sky130_fd_sc_hd__dfxtp_2
X_4883_ _4884_/A _5096_/A VGND VGND VPWR VPWR _4983_/C sky130_fd_sc_hd__nor2_1
XFILLER_177_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6622_ _7535_/Q _6480_/X _6487_/X _7471_/Q _6621_/X VGND VGND VPWR VPWR _6623_/D
+ sky130_fd_sc_hd__a221o_1
X_3834_ _7254_/Q _4541_/A _4505_/B _3581_/X _7365_/Q VGND VGND VPWR VPWR _3834_/X
+ sky130_fd_sc_hd__a32o_1
X_6553_ _7540_/Q _6479_/X _6485_/X _7548_/Q _6537_/X VGND VGND VPWR VPWR _6553_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3765_ _7080_/Q _4541_/A _4535_/B _5813_/A _7414_/Q VGND VGND VPWR VPWR _3774_/B
+ sky130_fd_sc_hd__a32o_1
X_5504_ _5313_/B _5092_/B _5416_/X _5425_/A _5289_/X VGND VGND VPWR VPWR _5625_/A
+ sky130_fd_sc_hd__a311o_1
XFILLER_173_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6484_ _6485_/B _6563_/C _6791_/D _7631_/Q VGND VGND VPWR VPWR _6484_/X sky130_fd_sc_hd__and4b_4
X_3696_ _3713_/A _5659_/C _4511_/C VGND VGND VPWR VPWR _3696_/X sky130_fd_sc_hd__and3_2
Xpad_flashh_clk_buff_inst _4183_/X VGND VGND VPWR VPWR pad_flash_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_133_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5435_ _5404_/A _5137_/A _5512_/B wire535/X VGND VGND VPWR VPWR _5501_/B sky130_fd_sc_hd__a31o_1
XFILLER_173_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput310 _4191_/X VGND VGND VPWR VPWR spimemio_flash_io1_di sky130_fd_sc_hd__buf_12
Xoutput321 hold843/X VGND VGND VPWR VPWR hold844/A sky130_fd_sc_hd__buf_12
XFILLER_10_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput332 hold655/X VGND VGND VPWR VPWR hold656/A sky130_fd_sc_hd__buf_12
XFILLER_145_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput343 hold710/X VGND VGND VPWR VPWR hold711/A sky130_fd_sc_hd__buf_12
XFILLER_133_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5366_ _5551_/A1 _5196_/A _5490_/C _5358_/A VGND VGND VPWR VPWR _5366_/X sky130_fd_sc_hd__o211a_1
XFILLER_113_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7105_ _7215_/CLK _7105_/D _6903_/A VGND VGND VPWR VPWR _7105_/Q sky130_fd_sc_hd__dfrtp_4
X_4317_ hold665/X _5988_/A1 _4321_/S VGND VGND VPWR VPWR _4317_/X sky130_fd_sc_hd__mux2_1
X_5297_ _5297_/A _5512_/B _5297_/C VGND VGND VPWR VPWR _5297_/X sky130_fd_sc_hd__and3_1
XFILLER_141_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7036_ _7289_/CLK _7036_/D fanout597/X VGND VGND VPWR VPWR _7036_/Q sky130_fd_sc_hd__dfrtp_2
X_4248_ hold475/X _4247_/X _4258_/S VGND VGND VPWR VPWR _4248_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4179_ _4179_/A _4179_/B VGND VGND VPWR VPWR _4179_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout570 hold42/X VGND VGND VPWR VPWR _4229_/S sky130_fd_sc_hd__buf_12
Xfanout592 _6907_/A VGND VGND VPWR VPWR _6911_/A sky130_fd_sc_hd__buf_6
XFILLER_59_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_csclk _7352_/CLK VGND VGND VPWR VPWR _7568_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_56_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7512_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_186_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3550_ _5661_/A _3550_/B _3717_/B VGND VGND VPWR VPWR _5813_/A sky130_fd_sc_hd__and3_4
XFILLER_128_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3481_ _3481_/A1 _4192_/B _3478_/X _3480_/Y VGND VGND VPWR VPWR _3481_/X sky130_fd_sc_hd__o31a_1
X_5220_ _4994_/X _5034_/C _4744_/A VGND VGND VPWR VPWR _5536_/A sky130_fd_sc_hd__a21oi_1
XFILLER_170_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5151_ _4829_/Y _4973_/Y _5150_/Y _4565_/Y VGND VGND VPWR VPWR _7244_/D sky130_fd_sc_hd__a31oi_1
XFILLER_123_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4102_ _3968_/S _4104_/D hold1633/X VGND VGND VPWR VPWR _4102_/Y sky130_fd_sc_hd__a21boi_1
X_5082_ _5196_/A _5476_/B _5476_/C _5476_/D VGND VGND VPWR VPWR _5082_/Y sky130_fd_sc_hd__nand4_1
XFILLER_96_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4033_ _7234_/Q _5628_/A _4553_/B _3700_/X _7169_/Q VGND VGND VPWR VPWR _4033_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_49_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5984_ _5984_/A _5984_/B _6029_/B VGND VGND VPWR VPWR hold63/A sky130_fd_sc_hd__and3_4
XFILLER_80_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4935_ _4943_/A _4935_/B _4935_/C _5007_/D VGND VGND VPWR VPWR _4936_/C sky130_fd_sc_hd__nand4_1
Xclkbuf_3_7_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_7_0_csclk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_33_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7654_ _7657_/CLK _7654_/D fanout607/X VGND VGND VPWR VPWR _7654_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_11 hold24/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4866_ _4866_/A _4957_/C _4950_/C VGND VGND VPWR VPWR _4926_/B sky130_fd_sc_hd__and3_1
XANTENNA_22 _5723_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_33 hold75/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6605_ _7558_/Q _6453_/X _6485_/X _7550_/Q VGND VGND VPWR VPWR _6605_/X sky130_fd_sc_hd__a22o_1
XANTENNA_44 _3555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_55 hold70/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3817_ _7207_/Q _5984_/A _5666_/B _3514_/X _7549_/Q VGND VGND VPWR VPWR _3817_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_177_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7585_ _7617_/CLK _7585_/D fanout624/X VGND VGND VPWR VPWR _7585_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_66 _5666_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4797_ _5186_/C _4801_/C _4797_/C VGND VGND VPWR VPWR _4797_/X sky130_fd_sc_hd__and3_1
XFILLER_165_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_77 _3815_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_88 hold5/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3748_ _3673_/C _4340_/A _5669_/B _3544_/X input30/X VGND VGND VPWR VPWR _3748_/X
+ sky130_fd_sc_hd__a32o_1
X_6536_ _7508_/Q _6791_/D _6536_/C VGND VGND VPWR VPWR _6536_/X sky130_fd_sc_hd__and3_1
XANTENNA_99 _6487_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3679_ _7607_/Q _3529_/X _6002_/B _3580_/X _7615_/Q VGND VGND VPWR VPWR _3679_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_133_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6467_ _7631_/Q _7632_/Q _6562_/B _6485_/B VGND VGND VPWR VPWR _6467_/X sky130_fd_sc_hd__and4bb_1
XFILLER_118_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5418_ _5313_/B _5092_/B _5416_/X _5289_/X VGND VGND VPWR VPWR _5418_/X sky130_fd_sc_hd__a31o_1
X_6398_ _7089_/Q _6149_/X _6396_/X _6397_/X VGND VGND VPWR VPWR _6398_/X sky130_fd_sc_hd__a211o_1
XFILLER_133_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput173 _4198_/X VGND VGND VPWR VPWR irq[1] sky130_fd_sc_hd__buf_12
XFILLER_133_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5349_ _4761_/A _4999_/B _5002_/X _5348_/X VGND VGND VPWR VPWR _5537_/B sky130_fd_sc_hd__a211oi_1
Xoutput184 _3441_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[18] sky130_fd_sc_hd__buf_12
Xoutput195 _3431_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[28] sky130_fd_sc_hd__buf_12
XFILLER_102_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7019_ _7583_/CLK _7019_/D fanout629/X VGND VGND VPWR VPWR _7711_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4720_ _4943_/A _4813_/B _4770_/A VGND VGND VPWR VPWR _5156_/B sky130_fd_sc_hd__nand3_1
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4651_ _5429_/D _4706_/D _4649_/X VGND VGND VPWR VPWR _4651_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_147_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput20 mask_rev_in[24] VGND VGND VPWR VPWR input20/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3602_ _5682_/A _3905_/B _5628_/A VGND VGND VPWR VPWR _3602_/X sky130_fd_sc_hd__and3_4
Xinput31 mask_rev_in[5] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__clkbuf_1
X_4582_ _5189_/A _4822_/A _4992_/D _5017_/B VGND VGND VPWR VPWR _4706_/D sky130_fd_sc_hd__nand4_4
X_7370_ _7518_/CLK _7370_/D fanout626/X VGND VGND VPWR VPWR _7370_/Q sky130_fd_sc_hd__dfstp_2
Xinput42 mgmt_gpio_in[15] VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput53 mgmt_gpio_in[25] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__clkbuf_4
Xmax_cap501 _5071_/B VGND VGND VPWR VPWR _5146_/C sky130_fd_sc_hd__clkbuf_2
Xinput64 mgmt_gpio_in[35] VGND VGND VPWR VPWR input64/X sky130_fd_sc_hd__clkbuf_2
X_3533_ hold69/X _3559_/B VGND VGND VPWR VPWR _5661_/B sky130_fd_sc_hd__and2_4
Xhold804 _7479_/Q VGND VGND VPWR VPWR hold804/X sky130_fd_sc_hd__dlygate4sd3_1
X_6321_ _6320_/X _6321_/A1 _6812_/S VGND VGND VPWR VPWR _7644_/D sky130_fd_sc_hd__mux2_1
Xinput75 porb VGND VGND VPWR VPWR input75/X sky130_fd_sc_hd__clkbuf_1
Xhold815 _7084_/Q VGND VGND VPWR VPWR hold815/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput86 spimemio_flash_io0_oeb VGND VGND VPWR VPWR _4185_/B sky130_fd_sc_hd__clkbuf_4
Xhold826 _5992_/X VGND VGND VPWR VPWR _7569_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput97 usr2_vcc_pwrgood VGND VGND VPWR VPWR input97/X sky130_fd_sc_hd__clkbuf_4
XFILLER_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold837 _7439_/Q VGND VGND VPWR VPWR hold837/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold848 _6041_/X VGND VGND VPWR VPWR _7612_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6252_ _6252_/A1 _6109_/X _6251_/X _6686_/S VGND VGND VPWR VPWR _6252_/X sky130_fd_sc_hd__o22a_1
X_3464_ _6913_/Q _6914_/Q VGND VGND VPWR VPWR _3464_/X sky130_fd_sc_hd__and2b_1
Xhold859 _7212_/Q VGND VGND VPWR VPWR hold859/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5203_ _5203_/A _5203_/B _5203_/C VGND VGND VPWR VPWR _5206_/A sky130_fd_sc_hd__and3_1
X_6183_ _7315_/Q _6082_/Y _6169_/X _6182_/X VGND VGND VPWR VPWR _6183_/X sky130_fd_sc_hd__o22a_2
XFILLER_130_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5134_ _5512_/B _5322_/C _5512_/D _5131_/X _5452_/B VGND VGND VPWR VPWR _5602_/A
+ sky130_fd_sc_hd__a32o_1
Xhold1504 _7656_/Q VGND VGND VPWR VPWR _6686_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1515 _7149_/Q VGND VGND VPWR VPWR _4452_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1526 _7434_/Q VGND VGND VPWR VPWR hold1526/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5065_ _5297_/A _5313_/C _5322_/A VGND VGND VPWR VPWR _5066_/B sky130_fd_sc_hd__and3_1
Xhold1537 _5805_/X VGND VGND VPWR VPWR _7402_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1548 _7641_/Q VGND VGND VPWR VPWR _6253_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1559 _6959_/Q VGND VGND VPWR VPWR _4208_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_4016_ _7229_/Q _4547_/A _5678_/B _3695_/X _7046_/Q VGND VGND VPWR VPWR _4016_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5967_ hold466/X _6003_/A1 _5974_/S VGND VGND VPWR VPWR _7546_/D sky130_fd_sc_hd__mux2_1
X_7706_ _7706_/A VGND VGND VPWR VPWR _7706_/X sky130_fd_sc_hd__clkbuf_1
X_4918_ _4918_/A _4918_/B _4918_/C VGND VGND VPWR VPWR _4921_/C sky130_fd_sc_hd__nand3_1
X_5898_ _5898_/A0 hold9/X hold25/X VGND VGND VPWR VPWR hold26/A sky130_fd_sc_hd__mux2_1
XFILLER_166_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7637_ _7662_/CLK _7637_/D fanout606/X VGND VGND VPWR VPWR _7637_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4849_ _4966_/A _4860_/B _4877_/C _4957_/B VGND VGND VPWR VPWR _4972_/C sky130_fd_sc_hd__and4_2
XFILLER_148_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7568_ _7568_/CLK _7568_/D fanout622/X VGND VGND VPWR VPWR _7568_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_4_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6519_ _7459_/Q _6464_/X _6469_/X _7331_/Q VGND VGND VPWR VPWR _6519_/X sky130_fd_sc_hd__a22o_1
XFILLER_107_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7499_ _7614_/CLK _7499_/D fanout605/X VGND VGND VPWR VPWR _7499_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_180_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_616 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6870_ _6899_/A _6911_/B VGND VGND VPWR VPWR _6870_/X sky130_fd_sc_hd__and2_1
XFILLER_19_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5821_ _6046_/A1 hold849/X _5821_/S VGND VGND VPWR VPWR _5821_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5752_ hold988/X _6040_/A1 _5758_/S VGND VGND VPWR VPWR _5752_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4703_ _5316_/A _5146_/B VGND VGND VPWR VPWR _5011_/C sky130_fd_sc_hd__nand2_8
XFILLER_187_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5683_ _5683_/A0 hold81/X _5685_/S VGND VGND VPWR VPWR _5683_/X sky130_fd_sc_hd__mux2_1
X_7422_ _7518_/CLK _7422_/D fanout625/X VGND VGND VPWR VPWR _7422_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4634_ _4990_/A _5014_/D _5094_/A _5046_/A VGND VGND VPWR VPWR _5229_/A sky130_fd_sc_hd__and4_2
XFILLER_163_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold601 _4264_/X VGND VGND VPWR VPWR _6997_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7353_ _7607_/CLK _7353_/D fanout624/X VGND VGND VPWR VPWR _7353_/Q sky130_fd_sc_hd__dfrtp_1
X_4565_ _7244_/Q _6829_/D VGND VGND VPWR VPWR _4565_/Y sky130_fd_sc_hd__nor2_1
XFILLER_156_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold612 hold612/A VGND VGND VPWR VPWR hold612/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold623 _7400_/Q VGND VGND VPWR VPWR hold623/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold634 hold634/A VGND VGND VPWR VPWR hold634/X sky130_fd_sc_hd__dlygate4sd3_1
X_6304_ _7409_/Q _6124_/X _6299_/X _6301_/X _6303_/X VGND VGND VPWR VPWR _6304_/X
+ sky130_fd_sc_hd__a2111o_1
X_3516_ hold34/X hold61/X hold74/A VGND VGND VPWR VPWR _3516_/X sky130_fd_sc_hd__and3b_4
XFILLER_89_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold645 hold645/A VGND VGND VPWR VPWR hold645/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap364 _4294_/S VGND VGND VPWR VPWR _4292_/S sky130_fd_sc_hd__buf_4
X_4496_ _4556_/A1 hold890/X _4498_/S VGND VGND VPWR VPWR _4496_/X sky130_fd_sc_hd__mux2_1
X_7284_ _7497_/CLK hold31/X fanout608/X VGND VGND VPWR VPWR _7284_/Q sky130_fd_sc_hd__dfrtp_4
Xhold656 hold656/A VGND VGND VPWR VPWR wb_dat_o[26] sky130_fd_sc_hd__buf_12
Xhold667 hold667/A VGND VGND VPWR VPWR hold667/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold678 _7683_/Q VGND VGND VPWR VPWR hold678/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold689 _4392_/X VGND VGND VPWR VPWR _7094_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3447_ _7413_/Q VGND VGND VPWR VPWR _3447_/Y sky130_fd_sc_hd__inv_2
X_6235_ _7406_/Q _6160_/D _6427_/A3 _6170_/C _7326_/Q VGND VGND VPWR VPWR _6235_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_131_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6166_ _7331_/Q _6166_/B _6166_/C VGND VGND VPWR VPWR _6166_/X sky130_fd_sc_hd__and3_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1301 _5808_/X VGND VGND VPWR VPWR _7405_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1312 _7469_/Q VGND VGND VPWR VPWR hold1312/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5117_ _5092_/A _5093_/C _5093_/X _5116_/Y VGND VGND VPWR VPWR _5117_/Y sky130_fd_sc_hd__a211oi_1
Xhold1323 _7504_/Q VGND VGND VPWR VPWR hold752/A sky130_fd_sc_hd__dlygate4sd3_1
X_6097_ _7631_/Q _6485_/B _6720_/C VGND VGND VPWR VPWR _6097_/X sky130_fd_sc_hd__and3_4
Xhold1334 _7071_/Q VGND VGND VPWR VPWR hold1334/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1345 _7357_/Q VGND VGND VPWR VPWR hold1345/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1356 _3621_/X VGND VGND VPWR VPWR _6949_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1367 _7455_/Q VGND VGND VPWR VPWR hold962/A sky130_fd_sc_hd__dlygate4sd3_1
X_5048_ _5048_/A _5048_/B _5048_/C VGND VGND VPWR VPWR _5048_/Y sky130_fd_sc_hd__nor3_1
XFILLER_38_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1378 _5842_/X VGND VGND VPWR VPWR _7435_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1389 _7259_/Q VGND VGND VPWR VPWR hold1389/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_507 input48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_518 _7714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_529 input78/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6999_ _7553_/CLK _6999_/D fanout624/X VGND VGND VPWR VPWR _7694_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_671 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4350_ _6865_/A1 _4350_/A1 _4351_/S VGND VGND VPWR VPWR _4350_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4281_ hold736/X _6863_/A1 _4291_/S VGND VGND VPWR VPWR _4281_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6020_ _6020_/A _6038_/B _6038_/C VGND VGND VPWR VPWR _6028_/S sky130_fd_sc_hd__and3_4
XFILLER_140_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6922_ _4183_/A1 _6922_/D _6877_/X VGND VGND VPWR VPWR _6922_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6853_ _6853_/A0 _6852_/X _6853_/S VGND VGND VPWR VPWR _7679_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5804_ _5840_/A _6020_/A _6029_/B VGND VGND VPWR VPWR _5812_/S sky130_fd_sc_hd__and3_4
X_6784_ _6784_/A _6784_/B _6784_/C _6809_/D VGND VGND VPWR VPWR _6784_/Y sky130_fd_sc_hd__nor4_1
XFILLER_167_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3996_ _7610_/Q hold24/A _5680_/B _5650_/A _7272_/Q VGND VGND VPWR VPWR _3996_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_22_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5735_ hold325/X _5843_/A1 _5740_/S VGND VGND VPWR VPWR _5735_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5666_ _5669_/B _5666_/B _5680_/C VGND VGND VPWR VPWR _5667_/S sky130_fd_sc_hd__and3_1
XFILLER_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7405_ _7421_/CLK _7405_/D fanout630/X VGND VGND VPWR VPWR _7405_/Q sky130_fd_sc_hd__dfrtp_4
X_4617_ _4597_/B _4597_/C _4704_/C _4614_/X VGND VGND VPWR VPWR _4617_/X sky130_fd_sc_hd__a211o_1
XFILLER_163_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5597_ _5597_/A _5597_/B _5597_/C _5597_/D VGND VGND VPWR VPWR _5597_/X sky130_fd_sc_hd__and4_1
XFILLER_135_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold420 hold420/A VGND VGND VPWR VPWR hold420/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 hold431/A VGND VGND VPWR VPWR hold431/X sky130_fd_sc_hd__dlygate4sd3_1
X_7336_ _7568_/CLK _7336_/D fanout628/X VGND VGND VPWR VPWR _7336_/Q sky130_fd_sc_hd__dfrtp_1
X_4548_ _4548_/A0 _5697_/A0 _4552_/S VGND VGND VPWR VPWR _7229_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold442 _7213_/Q VGND VGND VPWR VPWR hold442/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold453 _7704_/A VGND VGND VPWR VPWR hold453/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold464 _4483_/X VGND VGND VPWR VPWR _7175_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold475 _7698_/A VGND VGND VPWR VPWR hold475/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 _5901_/X VGND VGND VPWR VPWR _7488_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7267_ _7293_/CLK _7267_/D _6886_/A VGND VGND VPWR VPWR _7267_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_143_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4479_ _4479_/A0 _6865_/A1 _4480_/S VGND VGND VPWR VPWR _4479_/X sky130_fd_sc_hd__mux2_1
Xhold497 _5982_/X VGND VGND VPWR VPWR _7560_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6218_ hold87/A _6213_/B _6114_/X _6161_/X _7349_/Q VGND VGND VPWR VPWR _6218_/X
+ sky130_fd_sc_hd__a32o_1
X_7198_ _7459_/CLK _7198_/D fanout600/X VGND VGND VPWR VPWR _7198_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1120 _7699_/A VGND VGND VPWR VPWR _4250_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6149_ _6231_/B _6392_/B _6231_/D VGND VGND VPWR VPWR _6149_/X sky130_fd_sc_hd__and3_4
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1131 _7242_/Q VGND VGND VPWR VPWR _4563_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1142 hold1493/X VGND VGND VPWR VPWR _5796_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1153 _6865_/X VGND VGND VPWR VPWR _7685_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1164 _4509_/X VGND VGND VPWR VPWR _7197_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1175 hold1397/X VGND VGND VPWR VPWR _4508_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1186 hold1330/X VGND VGND VPWR VPWR _4536_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_304 _4116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1197 hold1510/X VGND VGND VPWR VPWR _4556_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_315 _4529_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_326 _5311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_337 _5761_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_348 hold31/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_359 _7003_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3850_ input97/X _5975_/B _5678_/C _3544_/X input26/X VGND VGND VPWR VPWR _3850_/X
+ sky130_fd_sc_hd__a32o_1
X_3781_ _7084_/Q _6861_/A _5680_/A _5689_/A input64/X VGND VGND VPWR VPWR _3781_/X
+ sky130_fd_sc_hd__a32o_1
X_5520_ _5520_/A1 wire535/A _5519_/X _5500_/Y VGND VGND VPWR VPWR _7247_/D sky130_fd_sc_hd__a211o_1
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5451_ _5451_/A _5451_/B VGND VGND VPWR VPWR _5454_/A sky130_fd_sc_hd__nand2_1
XFILLER_173_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4402_ hold796/X _6863_/A1 _4405_/S VGND VGND VPWR VPWR _4402_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5382_ _4935_/C _4934_/C _5389_/D _5263_/A VGND VGND VPWR VPWR _5382_/X sky130_fd_sc_hd__a31o_1
XFILLER_132_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7121_ _7215_/CLK _7121_/D _6903_/A VGND VGND VPWR VPWR _7121_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_113_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4333_ hold614/X _5926_/A0 _4333_/S VGND VGND VPWR VPWR _7045_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7052_ _7286_/CLK _7052_/D fanout604/X VGND VGND VPWR VPWR _7052_/Q sky130_fd_sc_hd__dfrtp_4
X_4264_ _4263_/X hold600/X _4274_/S VGND VGND VPWR VPWR _4264_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6003_ hold818/X _6003_/A1 _6010_/S VGND VGND VPWR VPWR _7578_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4195_ _4195_/A _4195_/B VGND VGND VPWR VPWR _4195_/X sky130_fd_sc_hd__and2_1
XFILLER_39_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6905_ _6907_/A _6908_/B VGND VGND VPWR VPWR _6905_/X sky130_fd_sc_hd__and2_1
XFILLER_54_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6836_ _6971_/Q _6836_/A2 _6836_/B1 _6970_/Q VGND VGND VPWR VPWR _6836_/X sky130_fd_sc_hd__a22o_1
XFILLER_168_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6767_ _7079_/Q _6450_/X _6452_/X _7187_/Q _6766_/X VGND VGND VPWR VPWR _6775_/B
+ sky130_fd_sc_hd__a221o_1
X_3979_ input93/X _3573_/C _5984_/B _3546_/X _7530_/Q VGND VGND VPWR VPWR _3979_/X
+ sky130_fd_sc_hd__a32o_1
X_5718_ _5718_/A0 _6006_/A1 _5722_/S VGND VGND VPWR VPWR _5718_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6698_ _7169_/Q _6474_/A _6464_/X _7682_/Q VGND VGND VPWR VPWR _6698_/X sky130_fd_sc_hd__a22o_1
X_5649_ _5649_/A0 hold85/X _5649_/S VGND VGND VPWR VPWR hold99/A sky130_fd_sc_hd__mux2_1
XFILLER_163_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold250 _6034_/X VGND VGND VPWR VPWR _7606_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 _5672_/X VGND VGND VPWR VPWR _7287_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7319_ _7497_/CLK _7319_/D fanout607/X VGND VGND VPWR VPWR _7319_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold272 _5710_/X VGND VGND VPWR VPWR _7318_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 _6037_/X VGND VGND VPWR VPWR _7609_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 _7590_/Q VGND VGND VPWR VPWR hold294/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_101 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_112 _6136_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_123 _6158_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_134 _6447_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_145 _6459_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_156 _6484_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_167 _6557_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_178 _6831_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_189 _6837_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput7 mask_rev_in[12] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4951_ _4951_/A _5401_/B VGND VGND VPWR VPWR _4951_/Y sky130_fd_sc_hd__nand2_1
XFILLER_189_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3902_ _3863_/X _3902_/B _3902_/C VGND VGND VPWR VPWR _3902_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_189_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7670_ _7672_/CLK _7670_/D VGND VGND VPWR VPWR _7670_/Q sky130_fd_sc_hd__dfxtp_2
X_4882_ _5404_/A _5112_/B VGND VGND VPWR VPWR _4882_/Y sky130_fd_sc_hd__nand2_4
XANTENNA_690 input80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6621_ _7495_/Q _6694_/B _6516_/C _6458_/X _7423_/Q VGND VGND VPWR VPWR _6621_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_32_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3833_ _7059_/Q _4487_/B _5666_/B _3585_/X _7333_/Q VGND VGND VPWR VPWR _3833_/X
+ sky130_fd_sc_hd__a32o_1
X_6552_ _7452_/Q _6459_/X _6549_/X _6551_/X VGND VGND VPWR VPWR _6552_/X sky130_fd_sc_hd__a211o_1
X_3764_ _7406_/Q _3545_/X _3565_/X _7326_/Q _3763_/X VGND VGND VPWR VPWR _3774_/A
+ sky130_fd_sc_hd__a221o_1
X_5503_ _5604_/B1 _4998_/Y _5415_/X _5288_/X VGND VGND VPWR VPWR _5503_/X sky130_fd_sc_hd__o31a_1
XFILLER_185_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6483_ _6485_/B _6645_/B _6771_/C _7631_/Q VGND VGND VPWR VPWR _6483_/X sky130_fd_sc_hd__and4b_4
X_3695_ _5661_/B _5682_/B _5678_/C VGND VGND VPWR VPWR _3695_/X sky130_fd_sc_hd__and3_1
XFILLER_145_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput300 _7284_/Q VGND VGND VPWR VPWR pwr_ctrl_out[3] sky130_fd_sc_hd__buf_12
X_5434_ _5313_/C _5137_/A _5042_/A _5433_/Y VGND VGND VPWR VPWR _5434_/X sky130_fd_sc_hd__a31o_1
XFILLER_133_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput311 _7714_/X VGND VGND VPWR VPWR spimemio_flash_io2_di sky130_fd_sc_hd__buf_12
Xoutput322 hold704/X VGND VGND VPWR VPWR hold705/A sky130_fd_sc_hd__buf_12
XFILLER_133_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput333 hold690/X VGND VGND VPWR VPWR hold691/A sky130_fd_sc_hd__buf_12
Xoutput344 hold696/X VGND VGND VPWR VPWR hold697/A sky130_fd_sc_hd__buf_12
X_5365_ _5490_/C _4801_/C _5490_/A _5364_/X _5363_/X VGND VGND VPWR VPWR _5365_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_99_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_3_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_3_0_csclk/X sky130_fd_sc_hd__clkbuf_8
X_7104_ _7130_/CLK _7104_/D fanout602/X VGND VGND VPWR VPWR _7104_/Q sky130_fd_sc_hd__dfrtp_4
X_4316_ hold366/X _5843_/A1 _4321_/S VGND VGND VPWR VPWR _4316_/X sky130_fd_sc_hd__mux2_1
X_5296_ _5311_/A _5311_/C _5291_/B _5111_/D _4981_/X VGND VGND VPWR VPWR _5296_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_87_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7035_ _7512_/CLK _7035_/D fanout608/X VGND VGND VPWR VPWR _7035_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4247_ hold139/X _5789_/A1 _4257_/S VGND VGND VPWR VPWR _4247_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4178_ _6919_/Q _6920_/Q VGND VGND VPWR VPWR _4179_/B sky130_fd_sc_hd__nand2b_1
XFILLER_67_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6819_ _3838_/Y _6819_/A1 _6823_/S VGND VGND VPWR VPWR _7667_/D sky130_fd_sc_hd__mux2_1
Xwire405 hold35/X VGND VGND VPWR VPWR hold36/A sky130_fd_sc_hd__clkbuf_1
XFILLER_183_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire427 _4969_/B VGND VGND VPWR VPWR _4966_/A sky130_fd_sc_hd__buf_2
XFILLER_137_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout560 _7627_/Q VGND VGND VPWR VPWR _6359_/B sky130_fd_sc_hd__buf_6
Xfanout593 _6907_/A VGND VGND VPWR VPWR _6899_/A sky130_fd_sc_hd__buf_4
XFILLER_120_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3480_ _4192_/B _3478_/X _6917_/Q VGND VGND VPWR VPWR _3480_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_170_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5150_ _5147_/Y _5148_/X wire535/X _5083_/Y VGND VGND VPWR VPWR _5150_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4101_ _4101_/A0 input58/X _4101_/S VGND VGND VPWR VPWR _6917_/D sky130_fd_sc_hd__mux2_1
XFILLER_69_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5081_ _4800_/Y _4821_/Y _4960_/Y _5080_/Y VGND VGND VPWR VPWR _5081_/X sky130_fd_sc_hd__o31a_1
X_4032_ _7490_/Q _3519_/X _3706_/X _7101_/Q _4031_/X VGND VGND VPWR VPWR _4032_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_96_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5983_ hold835/X _6028_/A1 _5983_/S VGND VGND VPWR VPWR _5983_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4934_ _5595_/A _5181_/C _4934_/C _5186_/B VGND VGND VPWR VPWR _4936_/B sky130_fd_sc_hd__nand4_4
X_7653_ _7657_/CLK _7653_/D fanout607/X VGND VGND VPWR VPWR _7653_/Q sky130_fd_sc_hd__dfrtp_1
X_4865_ _5025_/B _4865_/B _4865_/C VGND VGND VPWR VPWR _4957_/C sky130_fd_sc_hd__and3_2
XANTENNA_12 hold24/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 _5723_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6604_ _7542_/Q _6479_/X _6486_/X _7502_/Q _6587_/X VGND VGND VPWR VPWR _6604_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_34 hold75/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3816_ _3816_/A _3816_/B _3816_/C wire357/X VGND VGND VPWR VPWR _3816_/Y sky130_fd_sc_hd__nor4b_1
X_7584_ _7584_/CLK _7584_/D fanout613/X VGND VGND VPWR VPWR _7584_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_45 _3555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_56 hold70/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4796_ _5189_/A _5404_/A _5231_/C VGND VGND VPWR VPWR _4797_/C sky130_fd_sc_hd__and3_1
XANTENNA_67 _4275_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_78 _3901_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6535_ _6534_/X _6559_/A2 _6611_/S VGND VGND VPWR VPWR _6535_/X sky130_fd_sc_hd__mux2_1
XANTENNA_89 _4357_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3747_ _7218_/Q _5993_/A _4529_/B _3745_/X _3746_/X VGND VGND VPWR VPWR _3753_/C
+ sky130_fd_sc_hd__a311o_1
X_6466_ _6485_/B _6720_/C _6771_/C _7631_/Q VGND VGND VPWR VPWR _6466_/X sky130_fd_sc_hd__and4b_4
XFILLER_118_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3678_ _3678_/A _3678_/B _3678_/C _3678_/D VGND VGND VPWR VPWR _3692_/B sky130_fd_sc_hd__nor4_2
XFILLER_173_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5417_ _4816_/Y _4953_/C _5604_/B1 VGND VGND VPWR VPWR _5417_/X sky130_fd_sc_hd__a21o_1
X_6397_ _7237_/Q _6160_/D _6146_/C _6170_/C _7049_/Q VGND VGND VPWR VPWR _6397_/X
+ sky130_fd_sc_hd__a32o_1
Xoutput174 _4199_/X VGND VGND VPWR VPWR irq[2] sky130_fd_sc_hd__buf_12
XFILLER_0_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5348_ _5614_/C _5311_/A _4999_/B _5614_/A VGND VGND VPWR VPWR _5348_/X sky130_fd_sc_hd__o211a_1
Xoutput185 _3440_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[19] sky130_fd_sc_hd__buf_12
Xoutput196 _3430_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[29] sky130_fd_sc_hd__buf_12
X_5279_ _5279_/A _5279_/B _5279_/C VGND VGND VPWR VPWR _5279_/Y sky130_fd_sc_hd__nand3_1
XFILLER_101_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7018_ _7583_/CLK _7018_/D fanout629/X VGND VGND VPWR VPWR _7710_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_102_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout390 _6861_/A VGND VGND VPWR VPWR _5903_/A sky130_fd_sc_hd__buf_6
XFILLER_120_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4650_ _5429_/D _5000_/C _4568_/Y _4649_/X VGND VGND VPWR VPWR _5025_/C sky130_fd_sc_hd__o31a_2
XFILLER_187_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3457__1 _4183_/A1 VGND VGND VPWR VPWR _6953_/CLK sky130_fd_sc_hd__inv_2
Xinput10 mask_rev_in[15] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__clkbuf_1
X_3601_ _7393_/Q _3552_/X _5777_/A _7385_/Q _3600_/X VGND VGND VPWR VPWR _3601_/X
+ sky130_fd_sc_hd__a221o_1
Xinput21 mask_rev_in[25] VGND VGND VPWR VPWR input21/X sky130_fd_sc_hd__clkbuf_2
XFILLER_175_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4581_ _5189_/A _4822_/A _4992_/D _5017_/B VGND VGND VPWR VPWR _4581_/X sky130_fd_sc_hd__and4_1
Xinput32 mask_rev_in[6] VGND VGND VPWR VPWR input32/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput43 mgmt_gpio_in[16] VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__buf_2
XFILLER_174_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput54 mgmt_gpio_in[26] VGND VGND VPWR VPWR input54/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6320_ _6686_/S _6320_/A2 _6318_/X _6319_/X VGND VGND VPWR VPWR _6320_/X sky130_fd_sc_hd__a22o_1
XFILLER_116_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap502 _5231_/C VGND VGND VPWR VPWR _5071_/B sky130_fd_sc_hd__clkbuf_2
Xinput65 mgmt_gpio_in[36] VGND VGND VPWR VPWR _7714_/A sky130_fd_sc_hd__buf_4
X_3532_ hold73/A hold34/X hold61/A hold53/X VGND VGND VPWR VPWR hold54/A sky130_fd_sc_hd__nor4_1
Xhold805 _5891_/X VGND VGND VPWR VPWR _7479_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput76 qspi_enabled VGND VGND VPWR VPWR _4147_/A sky130_fd_sc_hd__buf_6
Xhold816 _4380_/X VGND VGND VPWR VPWR _7084_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput87 spimemio_flash_io1_do VGND VGND VPWR VPWR _7713_/A sky130_fd_sc_hd__clkbuf_4
Xinput98 usr2_vdd_pwrgood VGND VGND VPWR VPWR input98/X sky130_fd_sc_hd__clkbuf_2
Xhold827 _7575_/Q VGND VGND VPWR VPWR hold827/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold838 _5846_/X VGND VGND VPWR VPWR _7439_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6251_ _7318_/Q _6082_/Y _6237_/X _6250_/X VGND VGND VPWR VPWR _6251_/X sky130_fd_sc_hd__o22a_1
Xhold849 _7417_/Q VGND VGND VPWR VPWR hold849/X sky130_fd_sc_hd__dlygate4sd3_1
X_3463_ _5017_/B VGND VGND VPWR VPWR _5000_/C sky130_fd_sc_hd__inv_8
XFILLER_103_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5202_ _5196_/A _5614_/A _5476_/C _5045_/X VGND VGND VPWR VPWR _5202_/Y sky130_fd_sc_hd__a31oi_1
X_6182_ _7435_/Q _6159_/X _6170_/X _6172_/X _6181_/X VGND VGND VPWR VPWR _6182_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_130_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5133_ _5512_/B _5322_/C _5512_/D _5131_/X _5452_/B VGND VGND VPWR VPWR _5514_/C
+ sky130_fd_sc_hd__a32oi_2
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1505 _7661_/Q VGND VGND VPWR VPWR _6787_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1516 _7654_/Q VGND VGND VPWR VPWR _6611_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1527 _5841_/X VGND VGND VPWR VPWR _7434_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1538 _6930_/Q VGND VGND VPWR VPWR _4067_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5064_ _5313_/B _5111_/D VGND VGND VPWR VPWR _5064_/Y sky130_fd_sc_hd__nand2_1
XFILLER_123_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1549 _7277_/Q VGND VGND VPWR VPWR _5656_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_4015_ _7418_/Q _3602_/X _4007_/X _4008_/X _4014_/X VGND VGND VPWR VPWR _4036_/A
+ sky130_fd_sc_hd__a2111o_2
XFILLER_65_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5966_ _5984_/A hold24/X _6038_/C VGND VGND VPWR VPWR _5974_/S sky130_fd_sc_hd__and3_4
XFILLER_52_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7705_ _7705_/A VGND VGND VPWR VPWR _7705_/X sky130_fd_sc_hd__clkbuf_1
X_4917_ _4943_/A _5452_/A _5389_/C _4934_/C VGND VGND VPWR VPWR _4918_/C sky130_fd_sc_hd__nand4_1
X_5897_ hold123/X hold81/X hold25/X VGND VGND VPWR VPWR _5897_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7636_ _7680_/CLK _7636_/D _6886_/A VGND VGND VPWR VPWR _7636_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_166_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4848_ _5407_/C _5407_/D _4953_/C _6971_/Q VGND VGND VPWR VPWR _4848_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_165_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7567_ _7569_/CLK _7567_/D fanout614/X VGND VGND VPWR VPWR _7567_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_165_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4779_ _4948_/A _5074_/A _4822_/A _4959_/C _5017_/B VGND VGND VPWR VPWR _4779_/X
+ sky130_fd_sc_hd__o2111a_2
XFILLER_193_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6518_ _7587_/Q _6468_/X _6516_/X _6517_/X _6515_/X VGND VGND VPWR VPWR _6523_/B
+ sky130_fd_sc_hd__a2111o_1
X_7498_ _7498_/CLK _7498_/D fanout615/X VGND VGND VPWR VPWR _7498_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_134_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6449_ _6720_/C _6771_/C _6645_/C VGND VGND VPWR VPWR _6474_/A sky130_fd_sc_hd__and3_4
XFILLER_106_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_55_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7616_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_44_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5820_ _5991_/A1 hold591/X _5821_/S VGND VGND VPWR VPWR _5820_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_726 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5751_ hold449/X _6003_/A1 _5758_/S VGND VGND VPWR VPWR _5751_/X sky130_fd_sc_hd__mux2_1
X_4702_ _4822_/A _4959_/C _5146_/B VGND VGND VPWR VPWR _4702_/X sky130_fd_sc_hd__and3_2
XFILLER_147_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5682_ _5682_/A _5682_/B _5682_/C hold29/X VGND VGND VPWR VPWR _5682_/X sky130_fd_sc_hd__and4_1
XFILLER_147_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7421_ _7421_/CLK _7421_/D fanout630/X VGND VGND VPWR VPWR _7421_/Q sky130_fd_sc_hd__dfrtp_4
X_4633_ _4990_/A _5014_/D _5017_/A _5017_/B VGND VGND VPWR VPWR _4633_/Y sky130_fd_sc_hd__nand4_4
XFILLER_147_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7352_ _7352_/CLK _7352_/D fanout631/X VGND VGND VPWR VPWR _7352_/Q sky130_fd_sc_hd__dfrtp_1
X_4564_ hold598/X _4564_/A1 _4564_/S VGND VGND VPWR VPWR _4564_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold602 _7601_/Q VGND VGND VPWR VPWR hold602/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_118_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold613 hold613/A VGND VGND VPWR VPWR wb_dat_o[19] sky130_fd_sc_hd__buf_12
XFILLER_116_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6303_ _7433_/Q _6112_/X _6119_/X _7417_/Q _6302_/X VGND VGND VPWR VPWR _6303_/X
+ sky130_fd_sc_hd__a221o_1
Xhold624 _5802_/X VGND VGND VPWR VPWR _7400_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3515_ hold73/X hold53/X VGND VGND VPWR VPWR hold74/A sky130_fd_sc_hd__nor2_8
Xhold635 hold635/A VGND VGND VPWR VPWR wb_dat_o[29] sky130_fd_sc_hd__buf_12
X_7283_ _7497_/CLK _7283_/D fanout608/X VGND VGND VPWR VPWR _7283_/Q sky130_fd_sc_hd__dfrtp_4
X_4495_ _5869_/A1 _4495_/A1 _4498_/S VGND VGND VPWR VPWR _4495_/X sky130_fd_sc_hd__mux2_1
Xhold646 hold646/A VGND VGND VPWR VPWR wb_dat_o[25] sky130_fd_sc_hd__buf_12
Xhold657 hold657/A VGND VGND VPWR VPWR hold657/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold668 hold668/A VGND VGND VPWR VPWR wb_dat_o[31] sky130_fd_sc_hd__buf_12
Xmax_cap376 _6477_/X VGND VGND VPWR VPWR _6809_/D sky130_fd_sc_hd__buf_12
Xhold679 _6863_/X VGND VGND VPWR VPWR _7683_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6234_ _7342_/Q _6160_/D _6145_/C _6230_/X VGND VGND VPWR VPWR _6234_/X sky130_fd_sc_hd__a31o_1
X_3446_ _7421_/Q VGND VGND VPWR VPWR _3446_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ _7339_/Q _6131_/C _6119_/X _7411_/Q _6164_/X VGND VGND VPWR VPWR _6165_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1302 _7114_/Q VGND VGND VPWR VPWR hold426/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5116_ _5116_/A _5116_/B _5116_/C _5116_/D VGND VGND VPWR VPWR _5116_/Y sky130_fd_sc_hd__nand4_1
Xhold1313 _7445_/Q VGND VGND VPWR VPWR hold1313/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1324 _5919_/X VGND VGND VPWR VPWR _7504_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6096_ _6109_/B _6791_/C _6720_/C _6094_/Y _7631_/Q VGND VGND VPWR VPWR _7631_/D
+ sky130_fd_sc_hd__a32o_1
Xhold1335 _7060_/Q VGND VGND VPWR VPWR hold431/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1346 _5754_/X VGND VGND VPWR VPWR _7357_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1357 _6942_/Q VGND VGND VPWR VPWR _4038_/B1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1368 _6946_/Q VGND VGND VPWR VPWR _3777_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5047_ _5047_/A _5047_/B _5047_/C _5047_/D VGND VGND VPWR VPWR _5048_/C sky130_fd_sc_hd__nand4_1
XFILLER_72_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1379 _7333_/Q VGND VGND VPWR VPWR hold1379/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_508 _7714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_519 _7714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6998_ _7617_/CLK _6998_/D fanout624/X VGND VGND VPWR VPWR _6998_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_41_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5949_ hold520/X _6039_/A1 _5956_/S VGND VGND VPWR VPWR _7530_/D sky130_fd_sc_hd__mux2_1
XFILLER_166_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7619_ _7680_/CLK _7619_/D _6911_/A VGND VGND VPWR VPWR _7619_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_166_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4280_ _4279_/X _4280_/A1 _4292_/S VGND VGND VPWR VPWR _4280_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6921_ _7258_/CLK _6921_/D _6876_/X VGND VGND VPWR VPWR _6921_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6852_ _6969_/Q _6852_/A2 _6852_/B1 wire537/X _6851_/X VGND VGND VPWR VPWR _6852_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5803_ hold896/X _6046_/A1 _5803_/S VGND VGND VPWR VPWR _5803_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6783_ _7254_/Q _6460_/X _6780_/X _6782_/X VGND VGND VPWR VPWR _6784_/C sky130_fd_sc_hd__a211o_1
X_3995_ _3995_/A _3995_/B _3995_/C _3995_/D VGND VGND VPWR VPWR _3995_/Y sky130_fd_sc_hd__nor4_1
X_5734_ hold971/X _6040_/A1 _5740_/S VGND VGND VPWR VPWR _5734_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5665_ hold9/X _5665_/A1 hold30/X VGND VGND VPWR VPWR hold31/A sky130_fd_sc_hd__mux2_1
XFILLER_30_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7404_ _7562_/CLK _7404_/D fanout632/X VGND VGND VPWR VPWR _7404_/Q sky130_fd_sc_hd__dfrtp_4
X_4616_ _4597_/B _4597_/C _4704_/C _4614_/X VGND VGND VPWR VPWR _5358_/A sky130_fd_sc_hd__a211oi_4
XFILLER_135_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5596_ _4660_/C _4685_/Y _4691_/X _5592_/X _5595_/Y VGND VGND VPWR VPWR _5597_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_191_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold410 _4378_/X VGND VGND VPWR VPWR _7082_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7335_ _7599_/CLK _7335_/D fanout629/X VGND VGND VPWR VPWR _7335_/Q sky130_fd_sc_hd__dfrtp_1
X_4547_ _4547_/A _5678_/B _5680_/C VGND VGND VPWR VPWR _4552_/S sky130_fd_sc_hd__and3_2
Xhold421 hold421/A VGND VGND VPWR VPWR hold421/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 _7559_/Q VGND VGND VPWR VPWR hold432/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 _4528_/X VGND VGND VPWR VPWR _7213_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 _4296_/X VGND VGND VPWR VPWR _7012_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold465 hold465/A VGND VGND VPWR VPWR hold465/X sky130_fd_sc_hd__dlygate4sd3_1
X_7266_ _7293_/CLK _7266_/D fanout596/X VGND VGND VPWR VPWR _7266_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_89_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold476 _4248_/X VGND VGND VPWR VPWR _6990_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4478_ _4478_/A0 _4556_/A1 _4480_/S VGND VGND VPWR VPWR _4478_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold487 hold487/A VGND VGND VPWR VPWR hold487/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold498 _7456_/Q VGND VGND VPWR VPWR hold498/X sky130_fd_sc_hd__dlygate4sd3_1
X_6217_ _7445_/Q wire484/X _6146_/X _7517_/Q _6216_/X VGND VGND VPWR VPWR _6217_/X
+ sky130_fd_sc_hd__a221o_1
X_3429_ _7557_/Q VGND VGND VPWR VPWR _3429_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7197_ _7197_/CLK _7197_/D fanout618/X VGND VGND VPWR VPWR _7197_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6148_ _7538_/Q _6131_/B _6428_/B1 _6147_/X VGND VGND VPWR VPWR _6148_/X sky130_fd_sc_hd__a31o_1
Xhold1110 _7692_/A VGND VGND VPWR VPWR _4290_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1121 _4250_/X VGND VGND VPWR VPWR _6991_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1132 _4563_/X VGND VGND VPWR VPWR _7242_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1143 _7187_/Q VGND VGND VPWR VPWR _4497_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1154 _7119_/Q VGND VGND VPWR VPWR _4422_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_6079_ _6078_/Y _6109_/B _6075_/X _6151_/B _6065_/Y VGND VGND VPWR VPWR _7626_/D
+ sky130_fd_sc_hd__a32o_1
Xhold1165 hold1531/X VGND VGND VPWR VPWR _4439_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1176 hold1546/X VGND VGND VPWR VPWR _4415_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1187 hold1327/X VGND VGND VPWR VPWR _4548_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_305 _4116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1198 _7202_/Q VGND VGND VPWR VPWR _4515_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_316 _4535_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_327 _6043_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_338 _6039_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_349 hold50/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3780_ _5682_/A _5661_/A _5682_/C VGND VGND VPWR VPWR _3780_/X sky130_fd_sc_hd__and3_2
XFILLER_185_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5450_ _4871_/X _5381_/X _5449_/X _5260_/B _5527_/A VGND VGND VPWR VPWR _5451_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4401_ _4401_/A0 _6862_/A1 _4405_/S VGND VGND VPWR VPWR _7101_/D sky130_fd_sc_hd__mux2_1
X_5381_ _4769_/Y _4953_/C _5014_/D _4907_/A VGND VGND VPWR VPWR _5381_/X sky130_fd_sc_hd__a211o_1
X_7120_ _7242_/CLK _7120_/D fanout616/X VGND VGND VPWR VPWR _7120_/Q sky130_fd_sc_hd__dfrtp_4
X_4332_ hold966/X _5988_/A1 _4333_/S VGND VGND VPWR VPWR _7044_/D sky130_fd_sc_hd__mux2_1
XFILLER_5_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7051_ _7286_/CLK _7051_/D fanout598/X VGND VGND VPWR VPWR _7051_/Q sky130_fd_sc_hd__dfrtp_2
X_4263_ hold327/X _6031_/A0 _4275_/S VGND VGND VPWR VPWR _4263_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6002_ _6002_/A _6002_/B _6038_/C VGND VGND VPWR VPWR _6010_/S sky130_fd_sc_hd__and3_4
XFILLER_141_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4194_ _4202_/A _6971_/Q VGND VGND VPWR VPWR _6962_/D sky130_fd_sc_hd__and2_1
XFILLER_39_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6904_ _6907_/A _6907_/B VGND VGND VPWR VPWR _6904_/X sky130_fd_sc_hd__and2_1
XFILLER_82_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6835_ _6835_/A0 _6834_/X _6853_/S VGND VGND VPWR VPWR _7673_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6766_ _7084_/Q _6455_/C _6562_/C _6481_/X _7212_/Q VGND VGND VPWR VPWR _6766_/X
+ sky130_fd_sc_hd__a32o_1
X_3978_ input11/X _3542_/X _4257_/S input43/X _3977_/X VGND VGND VPWR VPWR _3995_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_10_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5717_ hold207/X _5789_/A1 _5722_/S VGND VGND VPWR VPWR _5717_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6697_ _7076_/Q _6450_/X _6452_/X _7184_/Q _6696_/X VGND VGND VPWR VPWR _6700_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_109_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_1__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _4183_/A1
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_164_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5648_ hold236/X _6866_/A1 _5649_/S VGND VGND VPWR VPWR _7270_/D sky130_fd_sc_hd__mux2_1
XFILLER_164_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5579_ _5579_/A _5579_/B VGND VGND VPWR VPWR _5580_/D sky130_fd_sc_hd__nor2_1
XFILLER_163_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold240 _4429_/X VGND VGND VPWR VPWR _7125_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7318_ _7541_/CLK _7318_/D fanout605/X VGND VGND VPWR VPWR _7318_/Q sky130_fd_sc_hd__dfrtp_2
Xhold251 hold251/A VGND VGND VPWR VPWR hold251/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold262 _7415_/Q VGND VGND VPWR VPWR hold262/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 _7276_/Q VGND VGND VPWR VPWR hold273/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold284 _7430_/Q VGND VGND VPWR VPWR hold284/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 _6016_/X VGND VGND VPWR VPWR _7590_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7249_ _7679_/CLK _7249_/D fanout635/X VGND VGND VPWR VPWR hold52/A sky130_fd_sc_hd__dfrtp_4
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_102 _6115_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_113 _6136_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_124 _6158_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_135 _6447_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_146 _6459_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_157 _6484_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_168 _6633_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_179 _6834_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput8 mask_rev_in[13] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4950_ _5407_/D _4953_/A _4950_/C _4950_/D VGND VGND VPWR VPWR _5401_/B sky130_fd_sc_hd__and4b_1
XFILLER_64_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3901_ _3901_/A _3901_/B _3901_/C _3901_/D VGND VGND VPWR VPWR _3901_/Y sky130_fd_sc_hd__nor4_1
X_4881_ _4992_/A _4992_/D _4992_/C _4992_/B VGND VGND VPWR VPWR _5401_/A sky130_fd_sc_hd__and4bb_4
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_680 input64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_691 input80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6620_ _7367_/Q _6445_/X _6452_/X _7583_/Q _6619_/X VGND VGND VPWR VPWR _6623_/C
+ sky130_fd_sc_hd__a221o_1
X_3832_ _7227_/Q _5840_/A _4541_/B _5849_/A _7445_/Q VGND VGND VPWR VPWR _3832_/X
+ sky130_fd_sc_hd__a32o_1
X_6551_ _7428_/Q _6444_/X _6464_/X _7460_/Q _6550_/X VGND VGND VPWR VPWR _6551_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_192_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3763_ _7366_/Q _5975_/B _5759_/B _3572_/X _7374_/Q VGND VGND VPWR VPWR _3763_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_146_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5502_ _4987_/Y _5417_/X _5438_/X _5310_/A VGND VGND VPWR VPWR _5605_/C sky130_fd_sc_hd__o211a_1
XFILLER_145_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6482_ _6791_/C _6645_/B _6563_/C VGND VGND VPWR VPWR _6482_/X sky130_fd_sc_hd__and3_4
X_3694_ _3777_/A1 _3693_/X _3904_/S VGND VGND VPWR VPWR _6947_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5433_ _5316_/X _5433_/B _5566_/D VGND VGND VPWR VPWR _5433_/Y sky130_fd_sc_hd__nand3b_1
Xoutput301 _3970_/Y VGND VGND VPWR VPWR reset sky130_fd_sc_hd__buf_12
XFILLER_10_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput312 _7715_/X VGND VGND VPWR VPWR spimemio_flash_io3_di sky130_fd_sc_hd__buf_12
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput323 hold698/X VGND VGND VPWR VPWR hold699/A sky130_fd_sc_hd__buf_12
Xoutput334 hold833/X VGND VGND VPWR VPWR hold834/A sky130_fd_sc_hd__buf_12
X_5364_ _5490_/C _5364_/B _5490_/A VGND VGND VPWR VPWR _5364_/X sky130_fd_sc_hd__and3_1
Xoutput345 hold714/X VGND VGND VPWR VPWR hold715/A sky130_fd_sc_hd__buf_12
XFILLER_126_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7103_ _7160_/CLK _7103_/D _6891_/A VGND VGND VPWR VPWR _7103_/Q sky130_fd_sc_hd__dfstp_2
X_4315_ hold327/X _6031_/A0 _4321_/S VGND VGND VPWR VPWR _4315_/X sky130_fd_sc_hd__mux2_1
X_5295_ _5071_/C _5137_/C wire572/X _5512_/B _4981_/X VGND VGND VPWR VPWR _5295_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_99_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7034_ _7568_/CLK _7034_/D fanout622/X VGND VGND VPWR VPWR _7034_/Q sky130_fd_sc_hd__dfrtp_1
X_4246_ _4246_/A0 _4245_/X _4258_/S VGND VGND VPWR VPWR _4246_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4177_ _6912_/Q _3500_/C _4192_/C _4176_/Y _6913_/Q VGND VGND VPWR VPWR _6956_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_83_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6818_ _3902_/Y _6818_/A1 _6823_/S VGND VGND VPWR VPWR _7666_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6749_ _7181_/Q _6465_/X _6740_/X _6744_/X _6748_/X VGND VGND VPWR VPWR _6749_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_149_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire428 _4704_/Y VGND VGND VPWR VPWR wire428/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout550 hold29/X VGND VGND VPWR VPWR _6038_/C sky130_fd_sc_hd__buf_8
XFILLER_59_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout561 _6213_/B VGND VGND VPWR VPWR _6158_/D sky130_fd_sc_hd__buf_6
XFILLER_65_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout583 _5021_/A VGND VGND VPWR VPWR _5512_/B sky130_fd_sc_hd__buf_6
XFILLER_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout594 _6907_/A VGND VGND VPWR VPWR _6891_/A sky130_fd_sc_hd__buf_6
XFILLER_59_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_586 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4100_ _7258_/Q _7257_/Q _7256_/Q _4104_/D VGND VGND VPWR VPWR _4101_/S sky130_fd_sc_hd__and4bb_1
X_5080_ _5476_/B _5614_/C _5476_/C _5476_/D VGND VGND VPWR VPWR _5080_/Y sky130_fd_sc_hd__nand4_2
XFILLER_96_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4031_ _7121_/Q _4559_/B _4487_/A _4030_/X VGND VGND VPWR VPWR _4031_/X sky130_fd_sc_hd__a31o_1
XFILLER_84_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5982_ hold496/X _6045_/A1 _5983_/S VGND VGND VPWR VPWR _5982_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4933_ _4933_/A _4933_/B _4933_/C VGND VGND VPWR VPWR _4936_/A sky130_fd_sc_hd__nor3_1
XFILLER_33_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7652_ _7657_/CLK _7652_/D fanout607/X VGND VGND VPWR VPWR _7652_/Q sky130_fd_sc_hd__dfrtp_1
X_4864_ _4946_/A _4935_/C _5389_/B VGND VGND VPWR VPWR _4906_/A sky130_fd_sc_hd__and3_1
XFILLER_178_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_13 hold24/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6603_ _7582_/Q _6452_/X _6464_/X _7462_/Q _6602_/X VGND VGND VPWR VPWR _6603_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_24 _3717_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3815_ _3815_/A _3815_/B _3815_/C _3815_/D VGND VGND VPWR VPWR _3815_/Y sky130_fd_sc_hd__nor4_1
XANTENNA_35 _4487_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7583_ _7583_/CLK _7583_/D fanout630/X VGND VGND VPWR VPWR _7583_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_46 _3555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4795_ _5143_/A _5143_/B VGND VGND VPWR VPWR _4795_/Y sky130_fd_sc_hd__nand2_1
XFILLER_165_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_57 hold70/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6534_ _6533_/X _7650_/Q _6686_/S VGND VGND VPWR VPWR _6534_/X sky130_fd_sc_hd__mux2_1
XANTENNA_68 _3588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_79 _3917_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3746_ _7105_/Q _6861_/A _5666_/B hold75/A _7510_/Q VGND VGND VPWR VPWR _3746_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_173_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6465_ _6791_/C _6791_/D _6771_/C VGND VGND VPWR VPWR _6465_/X sky130_fd_sc_hd__and3_4
X_3677_ _7415_/Q _5813_/A _5849_/A _7447_/Q _3676_/X VGND VGND VPWR VPWR _3678_/D
+ sky130_fd_sc_hd__a221o_1
X_5416_ _4948_/B _4959_/C _5112_/B _5042_/A VGND VGND VPWR VPWR _5416_/X sky130_fd_sc_hd__a31o_1
XFILLER_133_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6396_ _7212_/Q _6416_/C _6146_/C _6395_/X VGND VGND VPWR VPWR _6396_/X sky130_fd_sc_hd__a31o_1
XFILLER_99_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5347_ _5472_/A _5583_/A _5347_/C VGND VGND VPWR VPWR _5350_/B sky130_fd_sc_hd__and3_1
Xoutput175 _4165_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[0] sky130_fd_sc_hd__buf_12
Xoutput186 _4163_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[1] sky130_fd_sc_hd__buf_12
Xoutput197 _3456_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[2] sky130_fd_sc_hd__buf_12
XFILLER_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5278_ _4966_/A _4946_/B _4948_/Y _5276_/X VGND VGND VPWR VPWR _5278_/X sky130_fd_sc_hd__a31o_1
XFILLER_102_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7017_ _7583_/CLK _7017_/D fanout629/X VGND VGND VPWR VPWR _7709_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_101_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4229_ hold100/X _6853_/A0 _4229_/S VGND VGND VPWR VPWR _4229_/X sky130_fd_sc_hd__mux2_2
XFILLER_28_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout380 _6002_/B VGND VGND VPWR VPWR _4481_/A sky130_fd_sc_hd__buf_12
Xfanout391 _6861_/A VGND VGND VPWR VPWR _4559_/B sky130_fd_sc_hd__buf_8
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3600_ _7449_/Q _5840_/A _5993_/B _3572_/X _7377_/Q VGND VGND VPWR VPWR _3600_/X
+ sky130_fd_sc_hd__a32o_1
Xinput11 mask_rev_in[16] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput22 mask_rev_in[26] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__clkbuf_2
X_4580_ _4781_/B _4781_/C VGND VGND VPWR VPWR _4580_/Y sky130_fd_sc_hd__nand2_1
Xinput33 mask_rev_in[7] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__buf_2
XFILLER_128_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput44 mgmt_gpio_in[17] VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__clkbuf_4
Xinput55 mgmt_gpio_in[27] VGND VGND VPWR VPWR input55/X sky130_fd_sc_hd__clkbuf_1
X_3531_ _3714_/A hold24/A hold74/A VGND VGND VPWR VPWR _3531_/X sky130_fd_sc_hd__and3_4
Xinput66 mgmt_gpio_in[37] VGND VGND VPWR VPWR _7715_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput77 ser_tx VGND VGND VPWR VPWR input77/X sky130_fd_sc_hd__clkbuf_1
Xhold806 _7492_/Q VGND VGND VPWR VPWR hold806/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold817 hold817/A VGND VGND VPWR VPWR hold817/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold828 _5999_/X VGND VGND VPWR VPWR _7575_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap536 _6854_/B VGND VGND VPWR VPWR wire535/A sky130_fd_sc_hd__clkbuf_2
Xinput88 spimemio_flash_io1_oeb VGND VGND VPWR VPWR _4187_/B sky130_fd_sc_hd__clkbuf_4
Xinput99 wb_adr_i[0] VGND VGND VPWR VPWR input99/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold839 _7527_/Q VGND VGND VPWR VPWR hold839/X sky130_fd_sc_hd__dlygate4sd3_1
X_6250_ _7454_/Q _6132_/X _6240_/X _6243_/X _6249_/X VGND VGND VPWR VPWR _6250_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3462_ _5015_/C VGND VGND VPWR VPWR _5025_/B sky130_fd_sc_hd__inv_6
X_5201_ _5201_/A _5586_/A _5463_/A _5201_/D VGND VGND VPWR VPWR _5203_/A sky130_fd_sc_hd__and4_1
XFILLER_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6181_ _6178_/X _6131_/B _6174_/X _6180_/X _6176_/X VGND VGND VPWR VPWR _6181_/X
+ sky130_fd_sc_hd__a2111o_1
X_5132_ _5021_/B _5131_/X _5130_/X _5129_/Y VGND VGND VPWR VPWR _5132_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_97_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1506 _7522_/Q VGND VGND VPWR VPWR hold399/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1517 _7143_/Q VGND VGND VPWR VPWR _4446_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5063_ _4756_/Y _4982_/Y _4985_/Y _5062_/Y VGND VGND VPWR VPWR _5066_/C sky130_fd_sc_hd__o211ai_1
Xhold1528 _7639_/Q VGND VGND VPWR VPWR _6228_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1539 _6864_/X VGND VGND VPWR VPWR _7684_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4014_ _7394_/Q _3525_/X _4010_/X _4011_/X _4013_/X VGND VGND VPWR VPWR _4014_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_38_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5965_ hold908/X _6028_/A1 _5965_/S VGND VGND VPWR VPWR _5965_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7704_ _7704_/A VGND VGND VPWR VPWR _7704_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4916_ _5181_/C _5452_/A _5389_/C _4934_/C VGND VGND VPWR VPWR _4918_/B sky130_fd_sc_hd__nand4_1
X_5896_ hold158/X _6031_/A0 hold25/X VGND VGND VPWR VPWR _5896_/X sky130_fd_sc_hd__mux2_1
X_7635_ _7680_/CLK _7635_/D _6886_/A VGND VGND VPWR VPWR _7635_/Q sky130_fd_sc_hd__dfrtp_1
X_4847_ _5407_/C _5407_/D _4953_/C _6971_/Q VGND VGND VPWR VPWR _4847_/X sky130_fd_sc_hd__o31a_1
XFILLER_165_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7566_ _7566_/CLK _7566_/D fanout615/X VGND VGND VPWR VPWR _7566_/Q sky130_fd_sc_hd__dfrtp_2
X_4778_ _4948_/B _4959_/C _5017_/B VGND VGND VPWR VPWR _4836_/B sky130_fd_sc_hd__nand3_4
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3729_ _7614_/Q hold24/A _5680_/B _3674_/X _7270_/Q VGND VGND VPWR VPWR _3729_/X
+ sky130_fd_sc_hd__a32o_1
X_6517_ _7491_/Q _6694_/B _6720_/D _6479_/X _7539_/Q VGND VGND VPWR VPWR _6517_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_134_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7497_ _7497_/CLK _7497_/D fanout608/X VGND VGND VPWR VPWR _7497_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_180_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6448_ _7631_/Q _7630_/Q VGND VGND VPWR VPWR _6645_/C sky130_fd_sc_hd__nor2_8
XFILLER_134_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6379_ _6375_/X _6376_/X _6378_/X _6374_/X _6370_/X VGND VGND VPWR VPWR _6379_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_88_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5750_ hold24/X _5759_/B _6029_/B VGND VGND VPWR VPWR _5758_/S sky130_fd_sc_hd__and3_4
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4701_ _5407_/A _5429_/D VGND VGND VPWR VPWR _5404_/C sky130_fd_sc_hd__nand2b_4
X_5681_ _5681_/A0 _5697_/A0 _5681_/S VGND VGND VPWR VPWR _7294_/D sky130_fd_sc_hd__mux2_1
XFILLER_148_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4632_ _4990_/A _5014_/D _5015_/C _5008_/C VGND VGND VPWR VPWR _4786_/A sky130_fd_sc_hd__and4_4
X_7420_ _7562_/CLK _7420_/D fanout632/X VGND VGND VPWR VPWR _7420_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_175_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4563_ _4563_/A0 _6865_/A1 _4564_/S VGND VGND VPWR VPWR _4563_/X sky130_fd_sc_hd__mux2_1
X_7351_ _7432_/CLK _7351_/D fanout631/X VGND VGND VPWR VPWR _7351_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_190_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold603 _6028_/X VGND VGND VPWR VPWR _7601_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3514_ _3714_/A _5686_/A hold24/A VGND VGND VPWR VPWR _3514_/X sky130_fd_sc_hd__and3_4
X_6302_ _7401_/Q _6166_/B _6427_/A3 _6302_/B1 _7353_/Q VGND VGND VPWR VPWR _6302_/X
+ sky130_fd_sc_hd__a32o_1
Xhold614 hold614/A VGND VGND VPWR VPWR hold614/X sky130_fd_sc_hd__dlygate4sd3_1
X_7282_ _7497_/CLK _7282_/D fanout608/X VGND VGND VPWR VPWR _7282_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_116_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold625 hold625/A VGND VGND VPWR VPWR hold625/X sky130_fd_sc_hd__dlygate4sd3_1
X_4494_ _6862_/A1 hold922/X _4498_/S VGND VGND VPWR VPWR _4494_/X sky130_fd_sc_hd__mux2_1
Xhold636 _7695_/A VGND VGND VPWR VPWR hold636/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 _7460_/Q VGND VGND VPWR VPWR hold647/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 hold658/A VGND VGND VPWR VPWR wb_dat_o[22] sky130_fd_sc_hd__buf_12
XFILLER_171_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6233_ _7430_/Q _6432_/A3 _6309_/C _7334_/Q _6232_/X VGND VGND VPWR VPWR _6233_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_171_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold669 _7062_/Q VGND VGND VPWR VPWR hold669/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3445_ _7429_/Q VGND VGND VPWR VPWR _3445_/Y sky130_fd_sc_hd__inv_2
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6164_ _7395_/Q _6166_/B _6146_/C _6124_/X _7403_/Q VGND VGND VPWR VPWR _6164_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5115_ _5611_/A2 _4949_/Y _5015_/Y _5013_/Y _4888_/Y VGND VGND VPWR VPWR _5116_/C
+ sky130_fd_sc_hd__o32a_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1303 _4416_/X VGND VGND VPWR VPWR _7114_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1314 _7387_/Q VGND VGND VPWR VPWR hold979/A sky130_fd_sc_hd__dlygate4sd3_1
X_6095_ _6485_/B _6092_/X _6094_/Y VGND VGND VPWR VPWR _7630_/D sky130_fd_sc_hd__o21a_1
Xhold1325 _7589_/Q VGND VGND VPWR VPWR hold1325/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1336 _4351_/X VGND VGND VPWR VPWR _7060_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1347 _7531_/Q VGND VGND VPWR VPWR hold970/A sky130_fd_sc_hd__dlygate4sd3_1
X_5046_ _5046_/A _5046_/B _5233_/C VGND VGND VPWR VPWR _5047_/B sky130_fd_sc_hd__nand3_1
Xhold1358 _3968_/X VGND VGND VPWR VPWR _6943_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1369 _7317_/Q VGND VGND VPWR VPWR _5709_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_509 _7714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6997_ _7569_/CLK _6997_/D fanout613/X VGND VGND VPWR VPWR _6997_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5948_ _5984_/A _6020_/A hold29/X VGND VGND VPWR VPWR _5956_/S sky130_fd_sc_hd__and3_4
XFILLER_179_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5879_ hold755/X _6041_/A1 _5884_/S VGND VGND VPWR VPWR _5879_/X sky130_fd_sc_hd__mux2_1
X_7618_ _7680_/CLK _7618_/D _6911_/A VGND VGND VPWR VPWR _7618_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_193_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7549_ _7549_/CLK _7549_/D fanout629/X VGND VGND VPWR VPWR _7549_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_181_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6920_ _4183_/A1 _6920_/D _6875_/X VGND VGND VPWR VPWR _6920_/Q sky130_fd_sc_hd__dfrtp_1
X_6851_ _6971_/Q _6851_/A2 _6851_/B1 _6970_/Q VGND VGND VPWR VPWR _6851_/X sky130_fd_sc_hd__a22o_1
XFILLER_23_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5802_ hold623/X _5991_/A1 _5803_/S VGND VGND VPWR VPWR _5802_/X sky130_fd_sc_hd__mux2_1
X_3994_ _7586_/Q _6011_/A _3989_/X _3992_/X _3993_/X VGND VGND VPWR VPWR _3995_/D
+ sky130_fd_sc_hd__a2111o_1
X_6782_ _7054_/Q _6474_/B _6482_/X _7114_/Q _6781_/X VGND VGND VPWR VPWR _6782_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5733_ hold487/X _6003_/A1 _5740_/S VGND VGND VPWR VPWR _5733_/X sky130_fd_sc_hd__mux2_1
X_5664_ _6041_/A1 hold676/X hold30/X VGND VGND VPWR VPWR _5664_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7403_ _7515_/CLK _7403_/D fanout632/X VGND VGND VPWR VPWR _7403_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_148_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_54_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7608_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_129_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4615_ _4597_/B _4597_/C _4614_/X VGND VGND VPWR VPWR _4615_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_135_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5595_ _5595_/A _5595_/B _5595_/C _5595_/D VGND VGND VPWR VPWR _5595_/Y sky130_fd_sc_hd__nand4_1
XFILLER_190_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold400 hold400/A VGND VGND VPWR VPWR hold400/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold411 _7097_/Q VGND VGND VPWR VPWR hold411/X sky130_fd_sc_hd__dlygate4sd3_1
X_4546_ hold593/X _5926_/A0 _4546_/S VGND VGND VPWR VPWR _7228_/D sky130_fd_sc_hd__mux2_1
X_7334_ _7518_/CLK _7334_/D fanout625/X VGND VGND VPWR VPWR _7334_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_191_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold422 _7370_/Q VGND VGND VPWR VPWR hold422/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold433 _5981_/X VGND VGND VPWR VPWR _7559_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 _7288_/Q VGND VGND VPWR VPWR hold444/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold455 hold455/A VGND VGND VPWR VPWR hold455/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 hold466/A VGND VGND VPWR VPWR hold466/X sky130_fd_sc_hd__dlygate4sd3_1
X_7265_ _7293_/CLK _7265_/D _6886_/A VGND VGND VPWR VPWR _7265_/Q sky130_fd_sc_hd__dfrtp_2
X_4477_ hold424/X _5869_/A1 _4480_/S VGND VGND VPWR VPWR _4477_/X sky130_fd_sc_hd__mux2_1
Xhold477 _7472_/Q VGND VGND VPWR VPWR hold477/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold488 _7552_/Q VGND VGND VPWR VPWR hold488/X sky130_fd_sc_hd__dlygate4sd3_1
X_3428_ _7565_/Q VGND VGND VPWR VPWR _3428_/Y sky130_fd_sc_hd__inv_2
Xhold499 _5865_/X VGND VGND VPWR VPWR _7456_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_69_csclk _7236_/CLK VGND VGND VPWR VPWR _7194_/CLK sky130_fd_sc_hd__clkbuf_16
X_6216_ _7373_/Q _6159_/B _6127_/X _6144_/X hold46/A VGND VGND VPWR VPWR _6216_/X
+ sky130_fd_sc_hd__a32o_1
X_7196_ _7459_/CLK _7196_/D fanout600/X VGND VGND VPWR VPWR _7196_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_58_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6147_ _7514_/Q _6309_/B _6115_/X _6145_/X _7458_/Q VGND VGND VPWR VPWR _6147_/X
+ sky130_fd_sc_hd__a32o_1
Xhold1100 _5693_/X VGND VGND VPWR VPWR _7303_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1111 _4290_/X VGND VGND VPWR VPWR _7009_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1122 hold1334/X VGND VGND VPWR VPWR _4365_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1133 _7109_/Q VGND VGND VPWR VPWR _4410_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1144 _4497_/X VGND VGND VPWR VPWR _7187_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6078_ _6416_/C _6146_/C VGND VGND VPWR VPWR _6078_/Y sky130_fd_sc_hd__nand2_1
XFILLER_57_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1155 _4422_/X VGND VGND VPWR VPWR _7119_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1166 _7036_/Q VGND VGND VPWR VPWR _4323_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1177 hold1634/X VGND VGND VPWR VPWR _4217_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5029_ _4658_/X _4660_/Y _4688_/C _5229_/A _5614_/D VGND VGND VPWR VPWR _5068_/C
+ sky130_fd_sc_hd__o221a_4
Xhold1188 hold1437/X VGND VGND VPWR VPWR _4427_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_306 _4157_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1199 _4515_/X VGND VGND VPWR VPWR _7202_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_317 _5669_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_328 _5926_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_339 _6003_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_671 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4400_ _4559_/B _5666_/B _5686_/D VGND VGND VPWR VPWR _4405_/S sky130_fd_sc_hd__and3_2
X_5380_ _5407_/A _5429_/D _5189_/D _5021_/B VGND VGND VPWR VPWR _5389_/D sky130_fd_sc_hd__a31o_1
XFILLER_173_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4331_ hold377/X hold81/X _4333_/S VGND VGND VPWR VPWR _4331_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7050_ _7291_/CLK _7050_/D fanout596/X VGND VGND VPWR VPWR _7050_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_140_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4262_ _4261_/X hold823/X _4274_/S VGND VGND VPWR VPWR _4262_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6001_ hold291/X hold102/X _6001_/S VGND VGND VPWR VPWR _6001_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4193_ _4192_/C _4193_/B _6913_/Q VGND VGND VPWR VPWR _4193_/X sky130_fd_sc_hd__and3b_1
XFILLER_79_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6903_ _6903_/A _6907_/B VGND VGND VPWR VPWR _6903_/X sky130_fd_sc_hd__and2_1
XFILLER_23_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6834_ _6969_/Q _6834_/A2 _6834_/B1 wire537/X _6833_/X VGND VGND VPWR VPWR _6834_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_50_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6765_ _7172_/Q _6474_/A _6453_/X _7064_/Q _6764_/X VGND VGND VPWR VPWR _6775_/A
+ sky130_fd_sc_hd__a221o_1
X_3977_ _7602_/Q _5957_/B _4481_/A _3583_/X input52/X VGND VGND VPWR VPWR _3977_/X
+ sky130_fd_sc_hd__a32o_1
X_5716_ hold978/X _6040_/A1 _5722_/S VGND VGND VPWR VPWR _5716_/X sky130_fd_sc_hd__mux2_1
X_6696_ _7081_/Q _6645_/B _6536_/C _6479_/X _7219_/Q VGND VGND VPWR VPWR _6696_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_148_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5647_ hold529/X _5673_/A1 _5649_/S VGND VGND VPWR VPWR _5647_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5578_ _5557_/Y _5575_/Y _5577_/X _5573_/X VGND VGND VPWR VPWR _5578_/X sky130_fd_sc_hd__o31a_2
XFILLER_123_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold230 _5728_/X VGND VGND VPWR VPWR _7334_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 _7024_/Q VGND VGND VPWR VPWR hold241/X sky130_fd_sc_hd__dlygate4sd3_1
X_7317_ _7580_/CLK hold39/X fanout605/X VGND VGND VPWR VPWR _7317_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_144_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4529_ _4547_/A _4529_/B _5680_/C VGND VGND VPWR VPWR _4534_/S sky130_fd_sc_hd__and3_2
XFILLER_116_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold252 _7412_/Q VGND VGND VPWR VPWR hold252/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold263 _5819_/X VGND VGND VPWR VPWR _7415_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 _7223_/Q VGND VGND VPWR VPWR hold274/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold285 _5836_/X VGND VGND VPWR VPWR _7430_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 hold296/A VGND VGND VPWR VPWR hold296/X sky130_fd_sc_hd__dlygate4sd3_1
X_7248_ _7679_/CLK _7248_/D fanout635/X VGND VGND VPWR VPWR hold72/A sky130_fd_sc_hd__dfrtp_4
XFILLER_131_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7179_ _7254_/CLK _7179_/D fanout617/X VGND VGND VPWR VPWR _7179_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_103 _6115_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_114 _6138_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_125 _6159_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_136 _6645_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_147 _6459_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_158 _6484_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_169 _6633_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput9 mask_rev_in[14] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3900_ _7166_/Q _4511_/C _4469_/B _3894_/X _3899_/X VGND VGND VPWR VPWR _3901_/D
+ sky130_fd_sc_hd__a311o_2
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_670 _7222_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4880_ _4953_/D _4953_/A _5021_/B _4899_/C VGND VGND VPWR VPWR _4880_/Y sky130_fd_sc_hd__nand4b_2
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_681 _7714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_692 input80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3831_ _7341_/Q _3567_/X _3697_/X _7167_/Q _3830_/X VGND VGND VPWR VPWR _3837_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6550_ _7492_/Q _6694_/B _6720_/D _6452_/X _7580_/Q VGND VGND VPWR VPWR _6550_/X
+ sky130_fd_sc_hd__a32o_1
X_3762_ _7085_/Q _4559_/B _5680_/A _3707_/X _3761_/X VGND VGND VPWR VPWR _3775_/B
+ sky130_fd_sc_hd__a311oi_2
XFILLER_13_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5501_ _5602_/C _5501_/B VGND VGND VPWR VPWR _5501_/Y sky130_fd_sc_hd__nor2_1
XFILLER_158_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3693_ _3692_/Y _3693_/A1 _3967_/S VGND VGND VPWR VPWR _3693_/X sky130_fd_sc_hd__mux2_1
X_6481_ _6485_/B _6791_/D _6771_/C _7631_/Q VGND VGND VPWR VPWR _6481_/X sky130_fd_sc_hd__and4b_4
XFILLER_146_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5432_ _5452_/B _5040_/C _5095_/C _5291_/C VGND VGND VPWR VPWR _5432_/X sky130_fd_sc_hd__o211a_1
Xoutput302 _4195_/X VGND VGND VPWR VPWR ser_rx sky130_fd_sc_hd__buf_12
Xoutput313 hold941/X VGND VGND VPWR VPWR hold942/A sky130_fd_sc_hd__buf_12
Xoutput324 hold612/X VGND VGND VPWR VPWR hold613/A sky130_fd_sc_hd__buf_12
X_5363_ _5595_/B _5357_/X _5358_/X _5362_/X VGND VGND VPWR VPWR _5363_/X sky130_fd_sc_hd__a211o_1
Xoutput335 hold634/X VGND VGND VPWR VPWR hold635/A sky130_fd_sc_hd__buf_12
XFILLER_114_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7102_ _7160_/CLK _7102_/D _6891_/A VGND VGND VPWR VPWR _7102_/Q sky130_fd_sc_hd__dfrtp_4
X_4314_ hold481/X _6039_/A1 _4321_/S VGND VGND VPWR VPWR _4314_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5294_ _5404_/A _5112_/B _5111_/D _5512_/B _5551_/A1 VGND VGND VPWR VPWR _5294_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_59_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7033_ _7512_/CLK _7033_/D fanout608/X VGND VGND VPWR VPWR _7033_/Q sky130_fd_sc_hd__dfrtp_1
X_4245_ hold214/X _6040_/A1 _4257_/S VGND VGND VPWR VPWR _4245_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4176_ _6941_/Q _6940_/Q _6939_/Q _4193_/B VGND VGND VPWR VPWR _4176_/Y sky130_fd_sc_hd__nand4bb_1
XFILLER_142_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6817_ _3966_/X _6817_/A1 _6823_/S VGND VGND VPWR VPWR _7665_/D sky130_fd_sc_hd__mux2_1
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6748_ _7236_/Q _6807_/A2 _6501_/X _7206_/Q _6747_/X VGND VGND VPWR VPWR _6748_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_167_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6679_ _7449_/Q _6460_/X _6486_/X _7505_/Q _6678_/X VGND VGND VPWR VPWR _6684_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_164_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout540 hold5/X VGND VGND VPWR VPWR _6031_/A0 sky130_fd_sc_hd__buf_8
XFILLER_104_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout551 hold29/X VGND VGND VPWR VPWR _6861_/C sky130_fd_sc_hd__buf_12
XFILLER_116_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout562 _7627_/Q VGND VGND VPWR VPWR _6213_/B sky130_fd_sc_hd__buf_6
Xmgmt_gpio_14_buff_inst _4167_/X VGND VGND VPWR VPWR mgmt_gpio_out[14] sky130_fd_sc_hd__clkbuf_8
Xfanout584 _4708_/X VGND VGND VPWR VPWR _4946_/A sky130_fd_sc_hd__buf_8
Xfanout595 fanout603/X VGND VGND VPWR VPWR _6907_/A sky130_fd_sc_hd__buf_4
XFILLER_59_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4030_ _7466_/Q _3516_/X _6020_/A _3557_/X _7570_/Q VGND VGND VPWR VPWR _4030_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5981_ hold432/X hold85/X _5983_/S VGND VGND VPWR VPWR _5981_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4932_ _5375_/C _4935_/C _4934_/C VGND VGND VPWR VPWR _4933_/B sky130_fd_sc_hd__and3_1
XFILLER_33_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7651_ _7657_/CLK _7651_/D fanout605/X VGND VGND VPWR VPWR _7651_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_178_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4863_ _5595_/A _5595_/D _5181_/C _5186_/B VGND VGND VPWR VPWR _4908_/C sky130_fd_sc_hd__nand4_4
XANTENNA_14 _3514_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6602_ _7430_/Q _6444_/X _6588_/X _6601_/X VGND VGND VPWR VPWR _6602_/X sky130_fd_sc_hd__a211o_1
X_3814_ _7317_/Q hold37/A _3573_/X input6/X _3813_/X VGND VGND VPWR VPWR _3815_/D
+ sky130_fd_sc_hd__a221o_4
XANTENNA_25 _3528_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7582_ _7614_/CLK _7582_/D fanout604/X VGND VGND VPWR VPWR _7582_/Q sky130_fd_sc_hd__dfrtp_2
X_4794_ _4884_/A _5096_/B _5096_/C _4794_/D VGND VGND VPWR VPWR _5231_/C sky130_fd_sc_hd__nor4_2
XANTENNA_36 _4487_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_47 _3555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 hold70/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_69 _3623_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6533_ _6523_/Y wire368/X _7315_/Q _6759_/D VGND VGND VPWR VPWR _6533_/X sky130_fd_sc_hd__o2bb2a_2
X_3745_ _7163_/Q _4463_/A _3743_/X _3744_/X VGND VGND VPWR VPWR _3745_/X sky130_fd_sc_hd__a211o_1
XFILLER_192_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6464_ _6469_/A _6563_/C _6645_/C VGND VGND VPWR VPWR _6464_/X sky130_fd_sc_hd__and3_4
X_3676_ input17/X _5669_/B _4535_/B _3544_/X input31/X VGND VGND VPWR VPWR _3676_/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_146_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5415_ _5407_/A _5429_/D _4704_/A _4816_/Y VGND VGND VPWR VPWR _5415_/X sky130_fd_sc_hd__o31a_1
XFILLER_133_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6395_ _7172_/Q _6160_/D _6166_/C _6119_/X _7079_/Q VGND VGND VPWR VPWR _6395_/X
+ sky130_fd_sc_hd__a32o_1
X_5346_ _5471_/A _5537_/A _5346_/C _5536_/B VGND VGND VPWR VPWR _5347_/C sky130_fd_sc_hd__and4b_1
XFILLER_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput176 _3449_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[10] sky130_fd_sc_hd__buf_12
Xoutput187 _3439_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[20] sky130_fd_sc_hd__buf_12
Xoutput198 _3429_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[30] sky130_fd_sc_hd__buf_12
XFILLER_141_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5277_ _4966_/A _4946_/B _4951_/A _5276_/X VGND VGND VPWR VPWR _5279_/C sky130_fd_sc_hd__a31oi_1
XFILLER_102_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7016_ _7549_/CLK _7016_/D fanout629/X VGND VGND VPWR VPWR _7708_/A sky130_fd_sc_hd__dfrtp_1
X_4228_ _4228_/A0 hold50/X _4230_/S VGND VGND VPWR VPWR hold71/A sky130_fd_sc_hd__mux2_1
XFILLER_102_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4159_ _4158_/X input38/X _6954_/Q VGND VGND VPWR VPWR _4159_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout381 _5759_/B VGND VGND VPWR VPWR _4511_/C sky130_fd_sc_hd__buf_6
Xfanout392 _3516_/X VGND VGND VPWR VPWR _6861_/A sky130_fd_sc_hd__buf_12
XFILLER_46_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput12 mask_rev_in[17] VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__clkbuf_1
Xinput23 mask_rev_in[27] VGND VGND VPWR VPWR input23/X sky130_fd_sc_hd__clkbuf_1
Xinput34 mask_rev_in[8] VGND VGND VPWR VPWR input34/X sky130_fd_sc_hd__clkbuf_2
Xinput45 mgmt_gpio_in[18] VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3530_ _5984_/A _5661_/A _3717_/B VGND VGND VPWR VPWR _3530_/X sky130_fd_sc_hd__and3_4
XFILLER_128_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput56 mgmt_gpio_in[28] VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__clkbuf_4
Xhold807 _5906_/X VGND VGND VPWR VPWR _7492_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput67 mgmt_gpio_in[3] VGND VGND VPWR VPWR _4171_/D sky130_fd_sc_hd__buf_12
Xinput78 spi_csb VGND VGND VPWR VPWR input78/X sky130_fd_sc_hd__buf_4
XFILLER_6_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold818 hold818/A VGND VGND VPWR VPWR hold818/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput89 spimemio_flash_io2_do VGND VGND VPWR VPWR input89/X sky130_fd_sc_hd__clkbuf_2
X_3461_ _5014_/D VGND VGND VPWR VPWR _5007_/D sky130_fd_sc_hd__clkinv_8
Xhold829 _7588_/Q VGND VGND VPWR VPWR hold829/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5200_ _5046_/A _5229_/B _5233_/C _5195_/X _5476_/C VGND VGND VPWR VPWR _5201_/D
+ sky130_fd_sc_hd__a32oi_2
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6180_ _7443_/Q _6180_/A2 _6133_/X _7475_/Q _6179_/X VGND VGND VPWR VPWR _6180_/X
+ sky130_fd_sc_hd__a221o_1
X_5131_ _5131_/A _5131_/B _5291_/C VGND VGND VPWR VPWR _5131_/X sky130_fd_sc_hd__and3_1
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1507 _7485_/Q VGND VGND VPWR VPWR _5898_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5062_ _5061_/A _4989_/D _5061_/X _5060_/Y VGND VGND VPWR VPWR _5062_/Y sky130_fd_sc_hd__a211oi_1
Xhold1518 _6915_/Q VGND VGND VPWR VPWR _4105_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1529 _7648_/Q VGND VGND VPWR VPWR _6438_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_4013_ _7370_/Q _3572_/X _4382_/A _7086_/Q _4012_/X VGND VGND VPWR VPWR _4013_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_37_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5964_ hold583/X _6045_/A1 _5965_/S VGND VGND VPWR VPWR _5964_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7703_ _7703_/A VGND VGND VPWR VPWR _7703_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4915_ _4915_/A _4915_/B _4915_/C VGND VGND VPWR VPWR _4918_/A sky130_fd_sc_hd__nor3_1
XFILLER_178_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5895_ hold365/X _6039_/A1 hold25/X VGND VGND VPWR VPWR _7482_/D sky130_fd_sc_hd__mux2_1
X_7634_ _7662_/CLK _7634_/D fanout604/X VGND VGND VPWR VPWR _7634_/Q sky130_fd_sc_hd__dfrtp_1
X_4846_ _5316_/A _5112_/B VGND VGND VPWR VPWR _4953_/C sky130_fd_sc_hd__nand2_8
XFILLER_178_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7565_ _7611_/CLK _7565_/D fanout621/X VGND VGND VPWR VPWR _7565_/Q sky130_fd_sc_hd__dfrtp_4
X_4777_ _5407_/A _5074_/A _4948_/B _4959_/C VGND VGND VPWR VPWR _4777_/Y sky130_fd_sc_hd__o211ai_4
X_6516_ _7467_/Q _6720_/C _6516_/C _6645_/C VGND VGND VPWR VPWR _6516_/X sky130_fd_sc_hd__and4_1
XFILLER_107_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3728_ input16/X _3542_/X _3723_/X _3724_/X _3727_/X VGND VGND VPWR VPWR _3728_/X
+ sky130_fd_sc_hd__a2111o_1
X_7496_ _7497_/CLK _7496_/D fanout608/X VGND VGND VPWR VPWR _7496_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6447_ _6485_/B _6469_/A _6563_/C _7631_/Q VGND VGND VPWR VPWR _6447_/X sky130_fd_sc_hd__and4b_4
XFILLER_173_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3659_ _5678_/C _5678_/B _3658_/X _3560_/X _6977_/Q VGND VGND VPWR VPWR _3667_/A
+ sky130_fd_sc_hd__a32o_2
XFILLER_122_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6378_ _7093_/Q _6428_/A2 _6334_/C _7073_/Q _6377_/X VGND VGND VPWR VPWR _6378_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5329_ _5316_/C _5313_/C _5231_/B _5322_/A _5328_/X VGND VGND VPWR VPWR _5350_/A
+ sky130_fd_sc_hd__a41oi_2
XFILLER_87_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4700_ _4948_/A _5074_/A VGND VGND VPWR VPWR _5318_/A sky130_fd_sc_hd__nor2_2
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5680_ _5680_/A _5680_/B _5680_/C VGND VGND VPWR VPWR _5681_/S sky130_fd_sc_hd__and3_1
XFILLER_175_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4631_ _5189_/A _4992_/B _4822_/A _4992_/D VGND VGND VPWR VPWR _4631_/Y sky130_fd_sc_hd__nand4_4
XFILLER_30_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7350_ _7518_/CLK _7350_/D fanout627/X VGND VGND VPWR VPWR _7350_/Q sky130_fd_sc_hd__dfrtp_2
X_4562_ _4562_/A0 _6864_/A1 _4564_/S VGND VGND VPWR VPWR _4562_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold604 _7026_/Q VGND VGND VPWR VPWR hold604/X sky130_fd_sc_hd__dlygate4sd3_1
X_6301_ _7345_/Q _6131_/C _6115_/X _7393_/Q _6300_/X VGND VGND VPWR VPWR _6301_/X
+ sky130_fd_sc_hd__a221o_1
X_3513_ _3559_/B _3673_/C hold23/X _3513_/D VGND VGND VPWR VPWR hold24/A sky130_fd_sc_hd__and4bb_4
Xhold615 _6979_/Q VGND VGND VPWR VPWR hold615/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 _7305_/Q VGND VGND VPWR VPWR hold626/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7281_ _7497_/CLK _7281_/D fanout608/X VGND VGND VPWR VPWR _7281_/Q sky130_fd_sc_hd__dfrtp_4
X_4493_ _4547_/A _5661_/B _4493_/C _5680_/C VGND VGND VPWR VPWR _4493_/Y sky130_fd_sc_hd__nand4_4
XFILLER_171_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold637 _4270_/X VGND VGND VPWR VPWR _7000_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 _5870_/X VGND VGND VPWR VPWR _7460_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold659 _7463_/Q VGND VGND VPWR VPWR hold659/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6232_ _7390_/Q _6231_/D _6146_/C _6114_/X _7398_/Q VGND VGND VPWR VPWR _6232_/X
+ sky130_fd_sc_hd__a32o_1
X_3444_ _7437_/Q VGND VGND VPWR VPWR _3444_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6163_ _6163_/A1 _6812_/S _6162_/X VGND VGND VPWR VPWR _7637_/D sky130_fd_sc_hd__a21o_1
XFILLER_170_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5114_ _5611_/A2 _5094_/Y _5111_/Y _5112_/Y VGND VGND VPWR VPWR _5116_/B sky130_fd_sc_hd__o211a_1
XFILLER_97_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1304 _7421_/Q VGND VGND VPWR VPWR hold1304/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ _6485_/B _6092_/X _6093_/X VGND VGND VPWR VPWR _6094_/Y sky130_fd_sc_hd__a21oi_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1315 _5788_/X VGND VGND VPWR VPWR _7387_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1326 _7568_/Q VGND VGND VPWR VPWR hold726/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1337 _6935_/Q VGND VGND VPWR VPWR hold1/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1348 _7347_/Q VGND VGND VPWR VPWR hold984/A sky130_fd_sc_hd__dlygate4sd3_1
X_5045_ _5297_/A _5229_/B _5233_/C VGND VGND VPWR VPWR _5045_/X sky130_fd_sc_hd__and3_1
XFILLER_85_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1359 _7611_/Q VGND VGND VPWR VPWR hold987/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6996_ _7569_/CLK _6996_/D fanout613/X VGND VGND VPWR VPWR _6996_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_43_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5947_ hold299/X hold102/X _5947_/S VGND VGND VPWR VPWR _5947_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5878_ hold335/X _6031_/A0 _5884_/S VGND VGND VPWR VPWR _5878_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7617_ _7617_/CLK _7617_/D fanout624/X VGND VGND VPWR VPWR _7617_/Q sky130_fd_sc_hd__dfrtp_1
X_4829_ _4828_/X _4827_/Y _4613_/X VGND VGND VPWR VPWR _4829_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_193_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7548_ _7606_/CLK _7548_/D fanout606/X VGND VGND VPWR VPWR _7548_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_4_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7479_ _7547_/CLK _7479_/D fanout607/X VGND VGND VPWR VPWR _7479_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_134_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_752 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1 hold1/A VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6850_ _6850_/A0 _6849_/X _6853_/S VGND VGND VPWR VPWR _7678_/D sky130_fd_sc_hd__mux2_1
XFILLER_62_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5801_ hold934/X _6044_/A1 _5803_/S VGND VGND VPWR VPWR _5801_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6781_ _7109_/Q _6099_/B _6771_/C _6474_/C _7059_/Q VGND VGND VPWR VPWR _6781_/X
+ sky130_fd_sc_hd__a32o_1
X_3993_ _7266_/Q _5682_/C hold98/A _3701_/X _7239_/Q VGND VGND VPWR VPWR _3993_/X
+ sky130_fd_sc_hd__a32o_1
X_5732_ _6020_/A _5759_/B _6029_/B VGND VGND VPWR VPWR _5740_/S sky130_fd_sc_hd__and3_4
XFILLER_176_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5663_ _6031_/A0 hold113/X hold30/X VGND VGND VPWR VPWR _5663_/X sky130_fd_sc_hd__mux2_1
X_7402_ _7613_/CLK _7402_/D fanout625/X VGND VGND VPWR VPWR _7402_/Q sky130_fd_sc_hd__dfstp_1
X_4614_ _4573_/A _4573_/B _5143_/B _4595_/B VGND VGND VPWR VPWR _4614_/X sky130_fd_sc_hd__a211o_2
XFILLER_191_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5594_ _5595_/B _5357_/X _5486_/X _5593_/Y VGND VGND VPWR VPWR _5594_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_191_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold401 _7120_/Q VGND VGND VPWR VPWR hold401/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_163_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7333_ _7421_/CLK _7333_/D fanout630/X VGND VGND VPWR VPWR _7333_/Q sky130_fd_sc_hd__dfrtp_4
X_4545_ _4545_/A0 _6865_/A1 _4546_/S VGND VGND VPWR VPWR _4545_/X sky130_fd_sc_hd__mux2_1
Xhold412 _4396_/X VGND VGND VPWR VPWR _7097_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold423 _5769_/X VGND VGND VPWR VPWR _7370_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 _7255_/Q VGND VGND VPWR VPWR hold434/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold445 _5673_/X VGND VGND VPWR VPWR _7288_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7264_ _7293_/CLK _7264_/D _6886_/A VGND VGND VPWR VPWR _7264_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_89_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold456 _7051_/Q VGND VGND VPWR VPWR hold456/X sky130_fd_sc_hd__dlygate4sd3_1
X_4476_ _4476_/A0 _6012_/A0 _4480_/S VGND VGND VPWR VPWR _4476_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold467 _7464_/Q VGND VGND VPWR VPWR hold467/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 _5883_/X VGND VGND VPWR VPWR _7472_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold489 _5973_/X VGND VGND VPWR VPWR _7552_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6215_ _7469_/Q _6130_/X _6158_/X hold40/A _6214_/X VGND VGND VPWR VPWR _6215_/X
+ sky130_fd_sc_hd__a221o_1
X_3427_ _7573_/Q VGND VGND VPWR VPWR _3427_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7195_ _7459_/CLK _7195_/D fanout600/X VGND VGND VPWR VPWR _7195_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6146_ _6213_/B _6231_/D _6146_/C VGND VGND VPWR VPWR _6146_/X sky130_fd_sc_hd__and3_4
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1101 _7093_/Q VGND VGND VPWR VPWR _4391_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1112 _7172_/Q VGND VGND VPWR VPWR _4479_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1123 _7089_/Q VGND VGND VPWR VPWR _4386_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1134 _4410_/X VGND VGND VPWR VPWR _7109_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6077_ _6151_/B _6416_/C _6126_/D VGND VGND VPWR VPWR _6077_/X sky130_fd_sc_hd__and3_4
XFILLER_73_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1145 _7059_/Q VGND VGND VPWR VPWR _4350_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1156 hold1434/X VGND VGND VPWR VPWR _5644_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1167 _4323_/X VGND VGND VPWR VPWR _7036_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1178 _7038_/Q VGND VGND VPWR VPWR _4325_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5028_ _4654_/Y _4655_/Y _5025_/C VGND VGND VPWR VPWR _5614_/D sky130_fd_sc_hd__a21oi_4
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1189 hold1333/X VGND VGND VPWR VPWR _5638_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_307 _7262_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_318 _5682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_329 _5988_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6979_ _7289_/CLK _6979_/D fanout598/X VGND VGND VPWR VPWR _6979_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold990 _4274_/X VGND VGND VPWR VPWR _7002_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_95_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4330_ hold375/X _5869_/A1 _4333_/S VGND VGND VPWR VPWR _4330_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4261_ hold481/X _6039_/A1 _4275_/S VGND VGND VPWR VPWR _4261_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6000_ hold559/X _6045_/A1 _6001_/S VGND VGND VPWR VPWR _6000_/X sky130_fd_sc_hd__mux2_1
X_4192_ _6916_/Q _4192_/B _4192_/C VGND VGND VPWR VPWR _6952_/D sky130_fd_sc_hd__and3_1
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6902_ _6903_/A _6907_/B VGND VGND VPWR VPWR _6902_/X sky130_fd_sc_hd__and2_1
XFILLER_63_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6833_ _6971_/Q _6833_/A2 _6833_/B1 _6970_/Q VGND VGND VPWR VPWR _6833_/X sky130_fd_sc_hd__a22o_1
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6764_ _7192_/Q _6454_/X _6464_/X _7685_/Q _6763_/X VGND VGND VPWR VPWR _6764_/X
+ sky130_fd_sc_hd__a221o_1
X_3976_ _7682_/Q _4559_/B hold98/A VGND VGND VPWR VPWR _3976_/X sky130_fd_sc_hd__and3_1
XFILLER_149_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5715_ hold812/X _6003_/A1 _5722_/S VGND VGND VPWR VPWR _7322_/D sky130_fd_sc_hd__mux2_1
XFILLER_148_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6695_ _7179_/Q _6465_/X _6694_/X _6693_/X _6692_/X VGND VGND VPWR VPWR _6700_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_109_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5646_ _5646_/A0 _6864_/A1 _5649_/S VGND VGND VPWR VPWR _5646_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5577_ _5261_/D _5262_/X _5389_/X _5249_/X _5576_/Y VGND VGND VPWR VPWR _5577_/X
+ sky130_fd_sc_hd__a2111o_1
Xhold220 _7388_/Q VGND VGND VPWR VPWR hold220/X sky130_fd_sc_hd__dlygate4sd3_1
X_7316_ _7580_/CLK _7316_/D fanout605/X VGND VGND VPWR VPWR _7316_/Q sky130_fd_sc_hd__dfrtp_1
Xhold231 _7709_/A VGND VGND VPWR VPWR hold231/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4528_ _5926_/A0 hold442/X _4528_/S VGND VGND VPWR VPWR _4528_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold242 _4309_/X VGND VGND VPWR VPWR _7024_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 _5816_/X VGND VGND VPWR VPWR _7412_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 _7574_/Q VGND VGND VPWR VPWR hold264/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 _4540_/X VGND VGND VPWR VPWR _7223_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7247_ _7672_/CLK _7247_/D fanout635/X VGND VGND VPWR VPWR hold68/A sky130_fd_sc_hd__dfrtp_4
X_4459_ _4459_/A0 _4459_/A1 _4462_/S VGND VGND VPWR VPWR _7155_/D sky130_fd_sc_hd__mux2_1
Xhold286 _7326_/Q VGND VGND VPWR VPWR hold286/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 hold297/A VGND VGND VPWR VPWR hold297/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7178_ _7194_/CLK _7178_/D fanout602/X VGND VGND VPWR VPWR _7178_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_105_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6129_ _6118_/X _6123_/X _6128_/X _6159_/B VGND VGND VPWR VPWR _6129_/X sky130_fd_sc_hd__o31a_4
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_104 _6115_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_115 _6138_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 _6192_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_137 _6450_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_148 _6464_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_159 _6485_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_53_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7559_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_45_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_660 _6465_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_671 _7222_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_682 input80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_693 input80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3830_ _7182_/Q _4535_/B _4487_/B _5777_/A _7381_/Q VGND VGND VPWR VPWR _3830_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_189_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_68_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7498_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_177_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3761_ _7714_/A _5689_/A _3754_/X _3757_/X _3760_/X VGND VGND VPWR VPWR _3761_/X
+ sky130_fd_sc_hd__a2111o_2
X_5500_ _5459_/X _5460_/X _5499_/Y VGND VGND VPWR VPWR _5500_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_158_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6480_ _7629_/Q _7628_/Q _6562_/C VGND VGND VPWR VPWR _6480_/X sky130_fd_sc_hd__and3_4
X_3692_ _3692_/A _3692_/B _3692_/C VGND VGND VPWR VPWR _3692_/Y sky130_fd_sc_hd__nand3_4
XFILLER_187_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5431_ _4756_/Y _5285_/X _5611_/A2 _5566_/B _5428_/X VGND VGND VPWR VPWR _5433_/B
+ sky130_fd_sc_hd__o311a_1
Xoutput303 _4140_/B VGND VGND VPWR VPWR serial_clock sky130_fd_sc_hd__buf_12
Xoutput314 hold661/X VGND VGND VPWR VPWR hold662/A sky130_fd_sc_hd__buf_12
XFILLER_126_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5362_ _4743_/C _5595_/D _5595_/C _5361_/X VGND VGND VPWR VPWR _5362_/X sky130_fd_sc_hd__a31o_1
Xoutput325 hold651/X VGND VGND VPWR VPWR hold652/A sky130_fd_sc_hd__buf_12
XFILLER_99_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput336 hold674/X VGND VGND VPWR VPWR hold675/A sky130_fd_sc_hd__buf_12
X_7101_ _7215_/CLK _7101_/D _6903_/A VGND VGND VPWR VPWR _7101_/Q sky130_fd_sc_hd__dfrtp_4
X_4313_ _7294_/Q _4171_/C _4171_/D _4275_/S _6038_/C VGND VGND VPWR VPWR _4321_/S
+ sky130_fd_sc_hd__o311a_4
X_5293_ _5017_/B _5291_/C _5130_/B _5292_/X VGND VGND VPWR VPWR _5293_/X sky130_fd_sc_hd__a31o_1
XFILLER_87_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7032_ _7553_/CLK _7032_/D fanout622/X VGND VGND VPWR VPWR _7032_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4244_ hold748/X _4243_/X _4258_/S VGND VGND VPWR VPWR _4244_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4175_ _4192_/C _4104_/D _4179_/A _4174_/Y VGND VGND VPWR VPWR _6955_/D sky130_fd_sc_hd__a31o_1
XFILLER_95_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6816_ _4037_/Y _6816_/A1 _6823_/S VGND VGND VPWR VPWR _7664_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6747_ _7048_/Q _6471_/X _6484_/X _7093_/Q _6746_/X VGND VGND VPWR VPWR _6747_/X
+ sky130_fd_sc_hd__a221o_1
X_3959_ _7555_/Q _4547_/A _5975_/B _3704_/X _7195_/Q VGND VGND VPWR VPWR _3959_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_109_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6678_ _7369_/Q _6771_/B _6694_/C _6450_/X _7417_/Q VGND VGND VPWR VPWR _6678_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_164_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5629_ _6012_/A0 _5629_/A1 _5633_/S VGND VGND VPWR VPWR _5629_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout530 hold81/X VGND VGND VPWR VPWR _4556_/A1 sky130_fd_sc_hd__buf_4
Xfanout541 _5761_/A1 VGND VGND VPWR VPWR _6040_/A1 sky130_fd_sc_hd__buf_6
Xfanout552 hold29/X VGND VGND VPWR VPWR _6029_/B sky130_fd_sc_hd__buf_12
XFILLER_116_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout563 _6231_/B VGND VGND VPWR VPWR _6151_/B sky130_fd_sc_hd__buf_4
XFILLER_59_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout585 _5318_/A VGND VGND VPWR VPWR _5146_/B sky130_fd_sc_hd__buf_12
Xfanout596 fanout597/X VGND VGND VPWR VPWR fanout596/X sky130_fd_sc_hd__buf_6
XFILLER_19_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5980_ hold461/X _6043_/A1 _5983_/S VGND VGND VPWR VPWR _5980_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4931_ _4946_/A _4935_/C _4934_/C VGND VGND VPWR VPWR _4933_/A sky130_fd_sc_hd__and3_1
XFILLER_33_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7650_ _7657_/CLK _7650_/D fanout606/X VGND VGND VPWR VPWR _7650_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4862_ _4907_/A _4907_/C VGND VGND VPWR VPWR _4862_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_490 _7358_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6601_ _7534_/Q _6720_/C _6536_/C _6460_/X _7446_/Q VGND VGND VPWR VPWR _6601_/X
+ sky130_fd_sc_hd__a32o_1
X_3813_ input23/X _3546_/C _5669_/B hold56/A _7134_/Q VGND VGND VPWR VPWR _3813_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_177_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7581_ _7583_/CLK _7581_/D fanout629/X VGND VGND VPWR VPWR _7581_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_32_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_15 _3516_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 _3529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4793_ _4783_/X _4786_/Y _4884_/A _4572_/X VGND VGND VPWR VPWR _5407_/C sky130_fd_sc_hd__a211o_4
XFILLER_193_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_37 _4487_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 _3555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6532_ _6532_/A _6532_/B _6532_/C _6809_/D VGND VGND VPWR VPWR _6532_/Y sky130_fd_sc_hd__nor4_1
X_3744_ _7526_/Q _5984_/A _5939_/B _3546_/X _7534_/Q VGND VGND VPWR VPWR _3744_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_59 hold70/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6463_ _6485_/B _6469_/A _6771_/C _7631_/Q VGND VGND VPWR VPWR _6463_/X sky130_fd_sc_hd__and4b_4
X_3675_ _7511_/Q hold75/A _3674_/X _7271_/Q _3672_/X VGND VGND VPWR VPWR _3678_/C
+ sky130_fd_sc_hd__a221o_2
XFILLER_106_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5414_ _5285_/X _4993_/Y _4960_/Y _5604_/B1 _5001_/Y VGND VGND VPWR VPWR _5414_/X
+ sky130_fd_sc_hd__a311o_1
X_6394_ _7099_/Q _6112_/X _6309_/C _7167_/Q _6393_/X VGND VGND VPWR VPWR _6394_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_133_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5345_ _4677_/Y _4976_/Y _4982_/Y _4998_/Y _5221_/B VGND VGND VPWR VPWR _5536_/B
+ sky130_fd_sc_hd__o221a_1
Xoutput177 _3448_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[11] sky130_fd_sc_hd__buf_12
Xoutput188 _3438_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[21] sky130_fd_sc_hd__buf_12
XFILLER_87_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput199 _3428_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[31] sky130_fd_sc_hd__buf_12
X_5276_ _5407_/A _5404_/A _5404_/B _4963_/X VGND VGND VPWR VPWR _5276_/X sky130_fd_sc_hd__a31o_1
XFILLER_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7015_ _7597_/CLK _7015_/D fanout629/X VGND VGND VPWR VPWR _7707_/A sky130_fd_sc_hd__dfrtp_1
X_4227_ hold48/X hold65/X _4229_/S VGND VGND VPWR VPWR hold66/A sky130_fd_sc_hd__mux2_1
XFILLER_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4158_ _7005_/Q _6949_/Q _6911_/B VGND VGND VPWR VPWR _4158_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4089_ _7256_/Q _4104_/D _7258_/Q _7257_/Q VGND VGND VPWR VPWR _4097_/S sky130_fd_sc_hd__and4b_1
XFILLER_43_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout382 _5759_/B VGND VGND VPWR VPWR _4487_/B sky130_fd_sc_hd__clkbuf_4
Xfanout393 hold97/X VGND VGND VPWR VPWR hold98/A sky130_fd_sc_hd__buf_12
XFILLER_46_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput13 mask_rev_in[18] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput24 mask_rev_in[28] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput35 mask_rev_in[9] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__clkbuf_1
Xinput46 mgmt_gpio_in[19] VGND VGND VPWR VPWR input46/X sky130_fd_sc_hd__buf_2
Xinput57 mgmt_gpio_in[29] VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__clkbuf_1
Xinput68 mgmt_gpio_in[5] VGND VGND VPWR VPWR _4195_/A sky130_fd_sc_hd__buf_4
XFILLER_128_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold808 hold808/A VGND VGND VPWR VPWR hold808/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput79 spi_enabled VGND VGND VPWR VPWR _4196_/B sky130_fd_sc_hd__buf_6
Xhold819 _7076_/Q VGND VGND VPWR VPWR hold819/X sky130_fd_sc_hd__dlygate4sd3_1
X_3460_ _5074_/A VGND VGND VPWR VPWR _3460_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_182_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5130_ _5311_/C _5130_/B _5452_/C VGND VGND VPWR VPWR _5130_/X sky130_fd_sc_hd__and3_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1508 _7156_/Q VGND VGND VPWR VPWR _4460_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5061_ _5061_/A _5311_/A _5068_/C VGND VGND VPWR VPWR _5061_/X sky130_fd_sc_hd__and3_1
XFILLER_96_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1519 _6938_/Q VGND VGND VPWR VPWR _4055_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4012_ _7126_/Q _6861_/A _4553_/B _3581_/X _7362_/Q VGND VGND VPWR VPWR _4012_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_65_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5963_ hold997/X _5999_/A1 _5965_/S VGND VGND VPWR VPWR _5963_/X sky130_fd_sc_hd__mux2_1
X_7702_ _7702_/A VGND VGND VPWR VPWR _7702_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_40_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4914_ _5375_/C _5452_/A _5389_/C _4934_/C VGND VGND VPWR VPWR _4915_/B sky130_fd_sc_hd__and4_1
X_5894_ hold24/X _6861_/A _6038_/C VGND VGND VPWR VPWR hold25/A sky130_fd_sc_hd__and3_4
XFILLER_80_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4845_ _5407_/A _5074_/A _4948_/B _4959_/C VGND VGND VPWR VPWR _5021_/B sky130_fd_sc_hd__and4b_4
X_7633_ _4167_/A1 _7633_/D fanout620/X VGND VGND VPWR VPWR _7633_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7564_ _7569_/CLK _7564_/D fanout614/X VGND VGND VPWR VPWR _7564_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_178_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4776_ _5189_/A _4992_/B _4822_/A _4992_/D VGND VGND VPWR VPWR _5231_/B sky130_fd_sc_hd__o211a_4
XFILLER_148_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6515_ _7603_/Q _6456_/X _6481_/X _7379_/Q _6514_/X VGND VGND VPWR VPWR _6515_/X
+ sky130_fd_sc_hd__a221o_1
X_3727_ _7486_/Q _3531_/X _3702_/X _7065_/Q _3726_/X VGND VGND VPWR VPWR _3727_/X
+ sky130_fd_sc_hd__a221o_1
X_7495_ _7497_/CLK _7495_/D fanout608/X VGND VGND VPWR VPWR _7495_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_146_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6446_ _6485_/B _7633_/Q _7632_/Q _7631_/Q VGND VGND VPWR VPWR _6446_/X sky130_fd_sc_hd__and4bb_4
X_3658_ _7649_/Q hold92/A _7292_/Q VGND VGND VPWR VPWR _3658_/X sky130_fd_sc_hd__mux2_4
XFILLER_173_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6377_ _7231_/Q _6160_/D _6427_/A3 _6082_/B VGND VGND VPWR VPWR _6377_/X sky130_fd_sc_hd__a31o_1
X_3589_ input51/X _4257_/S _3583_/X input60/X _3588_/X VGND VGND VPWR VPWR _3589_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5328_ _5196_/A _5297_/A _4758_/X _5322_/A VGND VGND VPWR VPWR _5328_/X sky130_fd_sc_hd__o211a_1
XFILLER_88_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5259_ _5259_/A _5259_/B _5259_/C VGND VGND VPWR VPWR _5260_/D sky130_fd_sc_hd__and3_1
XFILLER_87_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4630_ _5189_/A _5074_/A _4822_/A _4992_/D VGND VGND VPWR VPWR _5046_/A sky130_fd_sc_hd__and4_4
XFILLER_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4561_ hold243/X _5869_/A1 _4564_/S VGND VGND VPWR VPWR _4561_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6300_ _7329_/Q _6067_/X _6145_/C _6077_/X _7385_/Q VGND VGND VPWR VPWR _6300_/X
+ sky130_fd_sc_hd__a32o_1
X_3512_ _3622_/A _3622_/B VGND VGND VPWR VPWR _3905_/B sky130_fd_sc_hd__nor2_8
XFILLER_155_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold605 _4311_/X VGND VGND VPWR VPWR _7026_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7280_ _7286_/CLK _7280_/D fanout604/X VGND VGND VPWR VPWR _7280_/Q sky130_fd_sc_hd__dfstp_1
Xhold616 _4230_/X VGND VGND VPWR VPWR _6979_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4492_ hold389/X _5926_/A0 _4492_/S VGND VGND VPWR VPWR _4492_/X sky130_fd_sc_hd__mux2_1
Xhold627 _5695_/X VGND VGND VPWR VPWR _7305_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 _6998_/Q VGND VGND VPWR VPWR hold638/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold649 _7072_/Q VGND VGND VPWR VPWR hold649/X sky130_fd_sc_hd__dlygate4sd3_1
X_6231_ _7422_/Q _6231_/B _6416_/B _6231_/D VGND VGND VPWR VPWR _6231_/X sky130_fd_sc_hd__and4_1
XFILLER_89_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3443_ _7445_/Q VGND VGND VPWR VPWR _3443_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _7314_/Q _6082_/Y _6129_/X _6156_/X _6109_/X VGND VGND VPWR VPWR _6162_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_124_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _5316_/A _5090_/B _5249_/C _5095_/X VGND VGND VPWR VPWR _5610_/A sky130_fd_sc_hd__a31o_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6093_ _6109_/B _7139_/Q VGND VGND VPWR VPWR _6093_/X sky130_fd_sc_hd__and2b_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1305 _5826_/X VGND VGND VPWR VPWR _7421_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1316 _7557_/Q VGND VGND VPWR VPWR hold1316/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1327 _7229_/Q VGND VGND VPWR VPWR hold1327/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _5042_/A _5191_/C _5095_/C _5614_/A VGND VGND VPWR VPWR _5047_/A sky130_fd_sc_hd__o211ai_1
XFILLER_38_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1338 _4223_/X VGND VGND VPWR VPWR hold18/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1349 _6947_/Q VGND VGND VPWR VPWR _3693_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6995_ _7583_/CLK _6995_/D fanout629/X VGND VGND VPWR VPWR _7703_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_80_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5946_ hold575/X _6045_/A1 _5947_/S VGND VGND VPWR VPWR _5946_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5877_ hold460/X _6003_/A1 _5884_/S VGND VGND VPWR VPWR _7466_/D sky130_fd_sc_hd__mux2_1
XFILLER_21_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7616_ _7616_/CLK _7616_/D fanout610/X VGND VGND VPWR VPWR _7616_/Q sky130_fd_sc_hd__dfrtp_1
X_4828_ _5375_/A _5189_/C _5181_/C VGND VGND VPWR VPWR _4828_/X sky130_fd_sc_hd__and3_1
XFILLER_193_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7547_ _7547_/CLK _7547_/D fanout607/X VGND VGND VPWR VPWR _7547_/Q sky130_fd_sc_hd__dfstp_2
X_4759_ _4654_/Y _4655_/Y _4750_/Y _4651_/Y VGND VGND VPWR VPWR _4759_/X sky130_fd_sc_hd__a211o_1
XFILLER_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7478_ _7614_/CLK _7478_/D fanout605/X VGND VGND VPWR VPWR _7478_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_108_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6429_ _7125_/Q _6359_/B _6429_/A3 _6153_/X _7208_/Q VGND VGND VPWR VPWR _6429_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_122_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2 hold2/A VGND VGND VPWR VPWR hold2/X sky130_fd_sc_hd__buf_6
XFILLER_66_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_607 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5800_ hold625/X _5926_/A0 _5803_/S VGND VGND VPWR VPWR _7398_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6780_ _7242_/Q _6694_/B _6563_/C _6459_/X _7119_/Q VGND VGND VPWR VPWR _6780_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_62_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3992_ _7554_/Q _5984_/A _5975_/B _3991_/X VGND VGND VPWR VPWR _3992_/X sky130_fd_sc_hd__a31o_1
X_5731_ hold865/X _6046_/A1 _5731_/S VGND VGND VPWR VPWR _5731_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5662_ _6039_/A1 hold298/X hold30/X VGND VGND VPWR VPWR _5662_/X sky130_fd_sc_hd__mux2_1
X_7401_ _7435_/CLK _7401_/D fanout623/X VGND VGND VPWR VPWR _7401_/Q sky130_fd_sc_hd__dfrtp_1
X_4613_ _4570_/Y _4704_/C _4704_/D _4597_/Y _6969_/Q VGND VGND VPWR VPWR _4613_/X
+ sky130_fd_sc_hd__o41a_2
XFILLER_191_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5593_ _4619_/Y _4680_/X _5484_/Y _5166_/X VGND VGND VPWR VPWR _5593_/Y sky130_fd_sc_hd__o31ai_1
X_7332_ _7562_/CLK _7332_/D fanout621/X VGND VGND VPWR VPWR _7332_/Q sky130_fd_sc_hd__dfrtp_1
X_4544_ hold530/X _5789_/A1 _4546_/S VGND VGND VPWR VPWR _4544_/X sky130_fd_sc_hd__mux2_1
Xhold402 _4423_/X VGND VGND VPWR VPWR _7120_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 _7203_/Q VGND VGND VPWR VPWR hold413/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold424 _7170_/Q VGND VGND VPWR VPWR hold424/X sky130_fd_sc_hd__dlygate4sd3_1
X_7263_ _7293_/CLK _7263_/D _6886_/A VGND VGND VPWR VPWR _7263_/Q sky130_fd_sc_hd__dfstp_2
Xhold435 _5633_/X VGND VGND VPWR VPWR _7255_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4475_ _4475_/A _4553_/B _6861_/C VGND VGND VPWR VPWR _4480_/S sky130_fd_sc_hd__and3_2
Xhold446 _7200_/Q VGND VGND VPWR VPWR hold446/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 _4341_/X VGND VGND VPWR VPWR _7051_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 _5874_/X VGND VGND VPWR VPWR _7464_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6214_ _7501_/Q _6213_/B _6127_/X _6133_/X _7477_/Q VGND VGND VPWR VPWR _6214_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_171_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3426_ _7581_/Q VGND VGND VPWR VPWR _3426_/Y sky130_fd_sc_hd__inv_2
Xhold479 _7616_/Q VGND VGND VPWR VPWR hold479/X sky130_fd_sc_hd__dlygate4sd3_1
X_7194_ _7194_/CLK _7194_/D fanout603/X VGND VGND VPWR VPWR _7194_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6145_ _6213_/B _6166_/B _6145_/C VGND VGND VPWR VPWR _6145_/X sky130_fd_sc_hd__and3_4
XFILLER_38_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1102 _4391_/X VGND VGND VPWR VPWR _7093_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1113 _4479_/X VGND VGND VPWR VPWR _7172_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1124 _4386_/X VGND VGND VPWR VPWR _7089_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_161_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6076_ _6126_/D _6151_/B VGND VGND VPWR VPWR _6076_/X sky130_fd_sc_hd__and2_1
Xhold1135 _7099_/Q VGND VGND VPWR VPWR _4398_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 _4350_/X VGND VGND VPWR VPWR _7059_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1157 hold1400/X VGND VGND VPWR VPWR _4206_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5027_ _5043_/B _5027_/B _5027_/C _5027_/D VGND VGND VPWR VPWR _5027_/X sky130_fd_sc_hd__and4_1
Xhold1168 hold1390/X VGND VGND VPWR VPWR _4335_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1179 _4325_/X VGND VGND VPWR VPWR _7038_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_308 _6978_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_319 _6099_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6978_ _7289_/CLK hold71/X fanout598/X VGND VGND VPWR VPWR _6978_/Q sky130_fd_sc_hd__dfstp_4
X_5929_ _6028_/A1 hold521/X hold76/X VGND VGND VPWR VPWR _5929_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold980 hold980/A VGND VGND VPWR VPWR hold980/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold991 _7005_/Q VGND VGND VPWR VPWR hold991/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_559 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4260_ _4275_/S _4240_/X _4259_/Y _6038_/C VGND VGND VPWR VPWR _4276_/S sky130_fd_sc_hd__o211ai_4
XFILLER_180_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4191_ _6951_/Q _4191_/B VGND VGND VPWR VPWR _4191_/X sky130_fd_sc_hd__and2b_4
XFILLER_67_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6901_ _6903_/A _6907_/B VGND VGND VPWR VPWR _6901_/X sky130_fd_sc_hd__and2_1
XFILLER_82_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6832_ hold14/A _6831_/X _6853_/S VGND VGND VPWR VPWR _7672_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3975_ _7280_/Q _5682_/A _5669_/B _5659_/C VGND VGND VPWR VPWR _3975_/X sky130_fd_sc_hd__and4_2
XFILLER_50_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6763_ _7094_/Q _6791_/D _6562_/C _6458_/X _7089_/Q VGND VGND VPWR VPWR _6763_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_149_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5714_ _5786_/B _5759_/B _6029_/B VGND VGND VPWR VPWR _5722_/S sky130_fd_sc_hd__and3_4
XFILLER_50_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6694_ _7199_/Q _6694_/B _6694_/C VGND VGND VPWR VPWR _6694_/X sky130_fd_sc_hd__and3_1
XFILLER_176_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5645_ hold781/X _6863_/A1 _5649_/S VGND VGND VPWR VPWR _5645_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5576_ _4859_/Y _4960_/Y _5015_/Y _5446_/X _4875_/X VGND VGND VPWR VPWR _5576_/Y
+ sky130_fd_sc_hd__o311ai_1
XFILLER_156_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold210 _5773_/X VGND VGND VPWR VPWR _7374_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7315_ _7547_/CLK _7315_/D fanout607/X VGND VGND VPWR VPWR _7315_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold221 _5789_/X VGND VGND VPWR VPWR _7388_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4527_ _5988_/A1 hold859/X _4528_/S VGND VGND VPWR VPWR _4527_/X sky130_fd_sc_hd__mux2_1
Xhold232 _4301_/X VGND VGND VPWR VPWR _7017_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold243 _7240_/Q VGND VGND VPWR VPWR hold243/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold254 _7055_/Q VGND VGND VPWR VPWR hold254/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 _5998_/X VGND VGND VPWR VPWR _7574_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4458_ _3838_/Y _4458_/A1 _4462_/S VGND VGND VPWR VPWR _7154_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7246_ _7679_/CLK _7246_/D fanout635/X VGND VGND VPWR VPWR _7246_/Q sky130_fd_sc_hd__dfrtp_4
Xhold276 hold276/A VGND VGND VPWR VPWR hold276/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 _5719_/X VGND VGND VPWR VPWR _7326_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold298 hold298/A VGND VGND VPWR VPWR hold298/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7177_ _7255_/CLK _7177_/D fanout616/X VGND VGND VPWR VPWR _7177_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4389_ _6862_/A1 _4389_/A1 _4393_/S VGND VGND VPWR VPWR _4389_/X sky130_fd_sc_hd__mux2_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6128_ _7330_/Q _6309_/C _6127_/X _7370_/Q _6125_/X VGND VGND VPWR VPWR _6128_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6059_ _7620_/Q _7621_/Q _6063_/D VGND VGND VPWR VPWR _6061_/B sky130_fd_sc_hd__nand3_1
XTAP_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_105 _6309_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_116 _6138_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 _6226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 _6450_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_149 _6474_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_650 _6145_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_661 _6465_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_672 _7222_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_683 input80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_694 _4187_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3760_ _7542_/Q _3530_/X _3562_/X _7502_/Q _3759_/X VGND VGND VPWR VPWR _3760_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_60_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3691_ _3691_/A _3691_/B _3691_/C _3691_/D VGND VGND VPWR VPWR _3691_/Y sky130_fd_sc_hd__nor4_1
X_5430_ _4756_/Y _5611_/A2 _4960_/Y _5514_/B VGND VGND VPWR VPWR _5566_/B sky130_fd_sc_hd__o31a_1
XFILLER_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput304 _3658_/X VGND VGND VPWR VPWR serial_data_1 sky130_fd_sc_hd__buf_12
XFILLER_161_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5361_ _4714_/X _5595_/C _5597_/A VGND VGND VPWR VPWR _5361_/X sky130_fd_sc_hd__a21bo_1
Xoutput315 hold630/X VGND VGND VPWR VPWR hold631/A sky130_fd_sc_hd__buf_12
XFILLER_114_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput326 hold784/X VGND VGND VPWR VPWR hold785/A sky130_fd_sc_hd__buf_12
Xoutput337 hold632/X VGND VGND VPWR VPWR hold633/A sky130_fd_sc_hd__buf_12
X_4312_ hold102/X _4312_/A1 _4312_/S VGND VGND VPWR VPWR _4312_/X sky130_fd_sc_hd__mux2_1
X_7100_ _7238_/CLK _7100_/D fanout602/X VGND VGND VPWR VPWR _7100_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5292_ _5108_/B _5131_/B _5291_/C _5311_/A VGND VGND VPWR VPWR _5292_/X sky130_fd_sc_hd__o211a_1
XFILLER_114_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7031_ _7553_/CLK _7031_/D fanout622/X VGND VGND VPWR VPWR _7031_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4243_ hold405/X _6003_/A1 _4257_/S VGND VGND VPWR VPWR _4243_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4174_ _6913_/Q _4174_/B _6912_/Q VGND VGND VPWR VPWR _4174_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_95_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6815_ _6815_/A _6962_/Q VGND VGND VPWR VPWR _6823_/S sky130_fd_sc_hd__nand2_4
XFILLER_51_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6746_ _7073_/Q _6447_/X _6474_/C _7058_/Q _6745_/X VGND VGND VPWR VPWR _6746_/X
+ sky130_fd_sc_hd__a221o_1
X_3958_ _7230_/Q _4547_/A _5678_/B _3957_/X VGND VGND VPWR VPWR _3958_/X sky130_fd_sc_hd__a31o_1
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3889_ _6974_/Q _3560_/X _3695_/X _7048_/Q _3888_/X VGND VGND VPWR VPWR _3889_/X
+ sky130_fd_sc_hd__a221o_1
X_6677_ _7337_/Q _6469_/X _6474_/C _7377_/Q _6676_/X VGND VGND VPWR VPWR _6684_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_109_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5628_ _5628_/A _5661_/B _5659_/C _6861_/C VGND VGND VPWR VPWR _5633_/S sky130_fd_sc_hd__nand4_4
XFILLER_164_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5559_ _4948_/B _5146_/B _5313_/B _5093_/C _5105_/Y VGND VGND VPWR VPWR _5560_/B
+ sky130_fd_sc_hd__a41oi_1
XFILLER_117_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7229_ _7294_/CLK _7229_/D fanout599/X VGND VGND VPWR VPWR _7229_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_132_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout520 hold19/X VGND VGND VPWR VPWR _6043_/A1 sky130_fd_sc_hd__buf_8
XFILLER_132_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout531 hold81/X VGND VGND VPWR VPWR _6041_/A1 sky130_fd_sc_hd__buf_6
XFILLER_120_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout542 hold5/X VGND VGND VPWR VPWR _5761_/A1 sky130_fd_sc_hd__buf_8
XFILLER_59_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout553 hold28/X VGND VGND VPWR VPWR hold29/A sky130_fd_sc_hd__buf_12
XFILLER_59_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout564 _7626_/Q VGND VGND VPWR VPWR _6231_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_58_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout597 fanout600/X VGND VGND VPWR VPWR fanout597/X sky130_fd_sc_hd__clkbuf_8
XFILLER_74_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4930_ _4930_/A _4930_/B _4930_/C VGND VGND VPWR VPWR _4933_/C sky130_fd_sc_hd__nand3_1
XFILLER_33_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_480 _7232_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4861_ _4633_/Y _4777_/Y _4836_/Y _5014_/D _4907_/A VGND VGND VPWR VPWR _5389_/B
+ sky130_fd_sc_hd__o221a_4
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_491 _7202_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6600_ _7350_/Q _6465_/X _6593_/X _6597_/X _6599_/X VGND VGND VPWR VPWR _6600_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_177_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3812_ _7124_/Q _3516_/X _4535_/B _3811_/X VGND VGND VPWR VPWR _3815_/C sky130_fd_sc_hd__a31o_1
XFILLER_178_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7580_ _7580_/CLK _7580_/D fanout605/X VGND VGND VPWR VPWR _7580_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_16 _3516_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4792_ _4783_/X _4786_/Y _4884_/A _4572_/X VGND VGND VPWR VPWR _4969_/B sky130_fd_sc_hd__a211oi_4
XFILLER_177_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_27 _3529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_38 _3544_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3743_ _7045_/Q _4529_/B _5680_/B _7494_/Q _3519_/X VGND VGND VPWR VPWR _3743_/X
+ sky130_fd_sc_hd__a32o_1
X_6531_ _7531_/Q _6480_/X _6528_/X _6530_/X VGND VGND VPWR VPWR _6532_/C sky130_fd_sc_hd__a211o_1
XANTENNA_49 _3555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3674_ _5686_/A _5686_/B hold98/A VGND VGND VPWR VPWR _3674_/X sky130_fd_sc_hd__and3_2
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6462_ _6791_/B _6720_/C _6645_/C VGND VGND VPWR VPWR _6474_/B sky130_fd_sc_hd__and3_4
X_5413_ _5285_/X _4993_/Y _4960_/Y _5604_/B1 _4998_/Y VGND VGND VPWR VPWR _5413_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_146_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6393_ _7069_/Q _6231_/D _6146_/C _6114_/X _7227_/Q VGND VGND VPWR VPWR _6393_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_161_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5344_ _5616_/A _5616_/C _5617_/A _5344_/D VGND VGND VPWR VPWR _5346_/C sky130_fd_sc_hd__and4bb_1
XFILLER_0_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput178 _3447_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[12] sky130_fd_sc_hd__buf_12
Xoutput189 _3437_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[22] sky130_fd_sc_hd__buf_12
XFILLER_102_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5275_ _4629_/Y _5011_/C _5407_/C _4854_/X VGND VGND VPWR VPWR _5279_/B sky130_fd_sc_hd__a211o_1
XFILLER_114_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7014_ _7549_/CLK _7014_/D fanout626/X VGND VGND VPWR VPWR _7706_/A sky130_fd_sc_hd__dfrtp_1
X_4226_ hold117/X hold85/X _4230_/S VGND VGND VPWR VPWR _6977_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4157_ _7010_/Q input77/X _4195_/B VGND VGND VPWR VPWR _4157_/X sky130_fd_sc_hd__mux2_4
XFILLER_110_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4088_ _6914_/Q _6912_/Q _6913_/Q VGND VGND VPWR VPWR _4104_/D sky130_fd_sc_hd__nor3_4
XFILLER_43_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6729_ _7683_/Q _6464_/X _6484_/X _7092_/Q _6728_/X VGND VGND VPWR VPWR _6734_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_52_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7584_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_192_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_67_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7558_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_78_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout383 _4475_/A VGND VGND VPWR VPWR _5759_/B sky130_fd_sc_hd__buf_8
XFILLER_46_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput14 mask_rev_in[19] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__clkbuf_1
Xinput25 mask_rev_in[29] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__clkbuf_1
XFILLER_168_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput36 mgmt_gpio_in[0] VGND VGND VPWR VPWR _4197_/A sky130_fd_sc_hd__clkbuf_4
Xinput47 mgmt_gpio_in[1] VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__buf_2
Xmax_cap506 _5490_/B VGND VGND VPWR VPWR _5186_/B sky130_fd_sc_hd__buf_6
Xinput58 mgmt_gpio_in[2] VGND VGND VPWR VPWR input58/X sky130_fd_sc_hd__buf_8
XFILLER_183_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput69 mgmt_gpio_in[6] VGND VGND VPWR VPWR input69/X sky130_fd_sc_hd__clkbuf_1
Xhold809 hold809/A VGND VGND VPWR VPWR wb_dat_o[12] sky130_fd_sc_hd__buf_12
XFILLER_128_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5060_ _4984_/Y _4987_/Y _5030_/Y _5059_/Y VGND VGND VPWR VPWR _5060_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1509 _7050_/Q VGND VGND VPWR VPWR hold213/A sky130_fd_sc_hd__dlygate4sd3_1
X_4011_ _7076_/Q _4541_/A _4487_/A _5813_/A _7410_/Q VGND VGND VPWR VPWR _4011_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_38_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5962_ _5962_/A0 hold2/X _5965_/S VGND VGND VPWR VPWR hold3/A sky130_fd_sc_hd__mux2_1
X_7701_ _7701_/A VGND VGND VPWR VPWR _7701_/X sky130_fd_sc_hd__clkbuf_2
X_4913_ _5452_/A _5389_/C _4925_/C VGND VGND VPWR VPWR _4915_/A sky130_fd_sc_hd__and3_1
X_5893_ hold888/X _6028_/A1 _5893_/S VGND VGND VPWR VPWR _5893_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7632_ _4167_/A1 _7632_/D fanout620/X VGND VGND VPWR VPWR _7632_/Q sky130_fd_sc_hd__dfstp_1
X_4844_ _4948_/A _5074_/A VGND VGND VPWR VPWR _5112_/B sky130_fd_sc_hd__and2b_4
XFILLER_138_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7563_ _7569_/CLK _7563_/D fanout614/X VGND VGND VPWR VPWR _7563_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_159_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4775_ _4775_/A _4775_/B _5180_/C _4775_/D VGND VGND VPWR VPWR _4775_/Y sky130_fd_sc_hd__nand4_1
XFILLER_165_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6514_ _7411_/Q _6450_/X _6474_/B _7595_/Q VGND VGND VPWR VPWR _6514_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3726_ _4199_/B _5984_/B _6038_/B _3725_/X VGND VGND VPWR VPWR _3726_/X sky130_fd_sc_hd__a31o_1
X_7494_ _7614_/CLK _7494_/D fanout605/X VGND VGND VPWR VPWR _7494_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6445_ _6791_/C _6469_/A _6445_/C VGND VGND VPWR VPWR _6445_/X sky130_fd_sc_hd__and3_4
X_3657_ _3693_/A1 _3656_/X _3904_/S VGND VGND VPWR VPWR _3657_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3588_ _7473_/Q _5903_/A _6020_/A hold56/A _7138_/Q VGND VGND VPWR VPWR _3588_/X
+ sky130_fd_sc_hd__a32o_4
X_6376_ _7063_/Q _6432_/A3 _6427_/B1 _7113_/Q VGND VGND VPWR VPWR _6376_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5327_ _5327_/A _5327_/B _5082_/Y VGND VGND VPWR VPWR _5544_/C sky130_fd_sc_hd__nor3b_2
XFILLER_130_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5258_ _5245_/X _5384_/A _5524_/A _5258_/D VGND VGND VPWR VPWR _5259_/C sky130_fd_sc_hd__and4bb_1
X_4209_ _6965_/Q _6962_/Q VGND VGND VPWR VPWR _4209_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5189_ _5189_/A _5375_/A _5189_/C _5189_/D VGND VGND VPWR VPWR _5189_/Y sky130_fd_sc_hd__nand4_1
XFILLER_96_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_532 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_587 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4560_ _4560_/A0 _6862_/A1 _4564_/S VGND VGND VPWR VPWR _4560_/X sky130_fd_sc_hd__mux2_1
X_3511_ _4229_/S hold22/X _3509_/Y VGND VGND VPWR VPWR hold23/A sky130_fd_sc_hd__o21ai_4
Xhold606 hold606/A VGND VGND VPWR VPWR hold606/X sky130_fd_sc_hd__dlygate4sd3_1
X_4491_ _4491_/A0 _6865_/A1 _4492_/S VGND VGND VPWR VPWR _4491_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold617 _7392_/Q VGND VGND VPWR VPWR hold617/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 hold628/A VGND VGND VPWR VPWR hold628/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold639 _4266_/X VGND VGND VPWR VPWR _6998_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6230_ _7382_/Q _6161_/D _6146_/C _6119_/X _7414_/Q VGND VGND VPWR VPWR _6230_/X
+ sky130_fd_sc_hd__a32o_1
X_3442_ _7453_/Q VGND VGND VPWR VPWR _3442_/Y sky130_fd_sc_hd__inv_2
Xmax_cap369 _5591_/C VGND VGND VPWR VPWR _5549_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_170_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6161_ _6213_/B _6231_/B _6416_/B _6161_/D VGND VGND VPWR VPWR _6161_/X sky130_fd_sc_hd__and4bb_2
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _5316_/A _5112_/B _5311_/C _5249_/C VGND VGND VPWR VPWR _5112_/Y sky130_fd_sc_hd__nand4_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ _6109_/B _7629_/Q _7628_/Q VGND VGND VPWR VPWR _6092_/X sky130_fd_sc_hd__and3_1
XFILLER_112_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1306 _7486_/Q VGND VGND VPWR VPWR hold233/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1317 _7581_/Q VGND VGND VPWR VPWR hold1317/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _5614_/A _5043_/B _5197_/B _5311_/A VGND VGND VPWR VPWR _5043_/Y sky130_fd_sc_hd__nand4_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1328 _7382_/Q VGND VGND VPWR VPWR hold281/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1339 _5655_/X VGND VGND VPWR VPWR _7276_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0_wbbd_sck _7680_/Q VGND VGND VPWR VPWR clkbuf_0_wbbd_sck/X sky130_fd_sc_hd__clkbuf_16
XFILLER_93_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6994_ _7583_/CLK _6994_/D fanout629/X VGND VGND VPWR VPWR _7702_/A sky130_fd_sc_hd__dfrtp_1
X_5945_ hold839/X _5999_/A1 _5947_/S VGND VGND VPWR VPWR _5945_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5876_ _5903_/A _6020_/A _6038_/C VGND VGND VPWR VPWR _5884_/S sky130_fd_sc_hd__and3_4
XFILLER_178_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7615_ _7617_/CLK _7615_/D fanout624/X VGND VGND VPWR VPWR _7615_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_139_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4827_ _4827_/A _4827_/B _4827_/C VGND VGND VPWR VPWR _4827_/Y sky130_fd_sc_hd__nand3_1
XFILLER_178_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7546_ _7613_/CLK _7546_/D fanout626/X VGND VGND VPWR VPWR _7546_/Q sky130_fd_sc_hd__dfstp_1
X_4758_ _5015_/C _5025_/C _5030_/D VGND VGND VPWR VPWR _4758_/X sky130_fd_sc_hd__and3_1
XFILLER_193_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3709_ _5661_/B _5682_/B _4511_/C VGND VGND VPWR VPWR _4358_/A sky130_fd_sc_hd__and3_2
XFILLER_146_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7477_ _7597_/CLK _7477_/D fanout626/X VGND VGND VPWR VPWR _7477_/Q sky130_fd_sc_hd__dfrtp_4
X_4689_ _4747_/B _5490_/C _5614_/C _5595_/B VGND VGND VPWR VPWR _5466_/C sky130_fd_sc_hd__nand4_2
XFILLER_107_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6428_ _7095_/Q _6428_/A2 _6428_/B1 _7223_/Q _6427_/X VGND VGND VPWR VPWR _6428_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_122_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6359_ _7252_/Q _6359_/B VGND VGND VPWR VPWR _6359_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_161_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3 hold3/A VGND VGND VPWR VPWR hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_82_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3991_ _7450_/Q _3516_/X _6002_/A _3990_/X VGND VGND VPWR VPWR _3991_/X sky130_fd_sc_hd__a31o_1
XFILLER_62_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5730_ hold767/X _5991_/A1 _5731_/S VGND VGND VPWR VPWR _5730_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5661_ _5661_/A _5661_/B _6038_/B hold29/X VGND VGND VPWR VPWR hold30/A sky130_fd_sc_hd__nand4_4
XFILLER_31_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7400_ _7445_/CLK _7400_/D fanout628/X VGND VGND VPWR VPWR _7400_/Q sky130_fd_sc_hd__dfrtp_1
X_4612_ _5186_/B _4760_/D _4760_/C _4760_/B VGND VGND VPWR VPWR _5189_/C sky130_fd_sc_hd__and4_1
X_5592_ _4629_/Y _4709_/Y _4811_/Y _4681_/Y _4691_/X VGND VGND VPWR VPWR _5592_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_129_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7331_ _7515_/CLK _7331_/D fanout621/X VGND VGND VPWR VPWR _7331_/Q sky130_fd_sc_hd__dfstp_1
X_4543_ hold585/X _5761_/A1 _4546_/S VGND VGND VPWR VPWR _4543_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold403 _7117_/Q VGND VGND VPWR VPWR hold403/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold414 _4516_/X VGND VGND VPWR VPWR _7203_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold425 _4477_/X VGND VGND VPWR VPWR _7170_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 _7703_/A VGND VGND VPWR VPWR hold436/X sky130_fd_sc_hd__dlygate4sd3_1
X_7262_ _7307_/CLK _7262_/D _6886_/A VGND VGND VPWR VPWR _7262_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_143_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4474_ hold387/X _5926_/A0 _4474_/S VGND VGND VPWR VPWR _4474_/X sky130_fd_sc_hd__mux2_1
Xhold447 _4513_/X VGND VGND VPWR VPWR _7200_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold458 _7252_/Q VGND VGND VPWR VPWR hold458/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 _7536_/Q VGND VGND VPWR VPWR hold469/X sky130_fd_sc_hd__dlygate4sd3_1
X_6213_ _7461_/Q _6213_/B _6309_/C VGND VGND VPWR VPWR _6213_/X sky130_fd_sc_hd__and3_1
X_3425_ _7589_/Q VGND VGND VPWR VPWR _3425_/Y sky130_fd_sc_hd__inv_2
X_7193_ _7207_/CLK _7193_/D fanout616/X VGND VGND VPWR VPWR _7193_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_171_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6144_ _6158_/D _6231_/B _6392_/B _6161_/D VGND VGND VPWR VPWR _6144_/X sky130_fd_sc_hd__and4_4
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1103 _7352_/Q VGND VGND VPWR VPWR _5748_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1114 _7429_/Q VGND VGND VPWR VPWR _5835_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6075_ _6416_/C _6126_/D _6151_/B VGND VGND VPWR VPWR _6075_/X sky130_fd_sc_hd__a21o_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1125 _7167_/Q VGND VGND VPWR VPWR _4473_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1136 _4398_/X VGND VGND VPWR VPWR _7099_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1147 _7064_/Q VGND VGND VPWR VPWR _4356_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1158 hold1592/X VGND VGND VPWR VPWR _4538_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5026_ _5297_/A _5195_/B _5476_/B _5233_/C VGND VGND VPWR VPWR _5026_/Y sky130_fd_sc_hd__nand4_1
Xhold1169 hold1389/X VGND VGND VPWR VPWR _5635_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_309 _4293_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6977_ _7289_/CLK _6977_/D fanout598/X VGND VGND VPWR VPWR _6977_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_41_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5928_ _6045_/A1 hold556/X hold76/A VGND VGND VPWR VPWR _7512_/D sky130_fd_sc_hd__mux2_1
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5859_ hold266/X _6039_/A1 _5866_/S VGND VGND VPWR VPWR _5859_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7529_ _7545_/CLK _7529_/D fanout613/X VGND VGND VPWR VPWR _7529_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_175_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold970 hold970/A VGND VGND VPWR VPWR hold970/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_134_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold981 hold981/A VGND VGND VPWR VPWR hold981/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold992 _4282_/X VGND VGND VPWR VPWR _7005_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4190_ _6923_/Q _4190_/B VGND VGND VPWR VPWR _4190_/X sky130_fd_sc_hd__and2b_4
XFILLER_69_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6900_ _6903_/A _6907_/B VGND VGND VPWR VPWR _6900_/X sky130_fd_sc_hd__and2_1
XFILLER_48_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6831_ _6971_/Q _6831_/A2 _6831_/B1 wire537/X _6830_/X VGND VGND VPWR VPWR _6831_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6762_ _6761_/X _6786_/A1 _6812_/S VGND VGND VPWR VPWR _7660_/D sky130_fd_sc_hd__mux2_1
X_3974_ _6958_/Q _5678_/C _6002_/A VGND VGND VPWR VPWR _3974_/X sky130_fd_sc_hd__and3_1
XFILLER_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5713_ _6028_/A1 hold577/X hold38/X VGND VGND VPWR VPWR _5713_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6693_ _7229_/Q _6720_/C _6536_/C _6471_/X _7046_/Q VGND VGND VPWR VPWR _6693_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_149_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5644_ _5644_/A0 _5697_/A0 _5649_/S VGND VGND VPWR VPWR _7266_/D sky130_fd_sc_hd__mux2_1
XFILLER_191_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5575_ _5400_/X _5454_/B _5575_/C _5575_/D VGND VGND VPWR VPWR _5575_/Y sky130_fd_sc_hd__nand4bb_1
XFILLER_156_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold200 _4507_/X VGND VGND VPWR VPWR _7195_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7314_ _7614_/CLK _7314_/D fanout605/X VGND VGND VPWR VPWR _7314_/Q sky130_fd_sc_hd__dfstp_2
Xhold211 _7414_/Q VGND VGND VPWR VPWR hold211/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_191_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4526_ _5789_/A1 hold343/X _4528_/S VGND VGND VPWR VPWR _4526_/X sky130_fd_sc_hd__mux2_1
Xhold222 hold222/A VGND VGND VPWR VPWR hold222/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 hold233/A VGND VGND VPWR VPWR hold233/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 _4561_/X VGND VGND VPWR VPWR _7240_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold255 _4345_/X VGND VGND VPWR VPWR _7055_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7245_ _7679_/CLK _7245_/D fanout635/X VGND VGND VPWR VPWR _7245_/Q sky130_fd_sc_hd__dfrtp_4
Xhold266 _7450_/Q VGND VGND VPWR VPWR hold266/X sky130_fd_sc_hd__dlygate4sd3_1
X_4457_ _3902_/Y _4457_/A1 _4462_/S VGND VGND VPWR VPWR _7153_/D sky130_fd_sc_hd__mux2_1
XFILLER_171_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold277 hold277/A VGND VGND VPWR VPWR hold277/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold288 hold288/A VGND VGND VPWR VPWR hold288/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 _7529_/Q VGND VGND VPWR VPWR hold299/X sky130_fd_sc_hd__dlygate4sd3_1
X_7176_ _7498_/CLK _7176_/D fanout615/X VGND VGND VPWR VPWR _7176_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_98_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4388_ _4388_/A _5686_/D VGND VGND VPWR VPWR _4393_/S sky130_fd_sc_hd__nand2_4
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6127_ _6231_/B _6392_/B _7624_/Q _7623_/Q VGND VGND VPWR VPWR _6127_/X sky130_fd_sc_hd__and4b_4
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6058_ _4140_/Y _6056_/Y _6057_/X _6053_/A _6058_/B2 VGND VGND VPWR VPWR _7620_/D
+ sky130_fd_sc_hd__a32o_1
XTAP_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5009_ _5108_/B _5094_/D VGND VGND VPWR VPWR _5009_/Y sky130_fd_sc_hd__nand2_4
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_106 _6129_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_117 _6138_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_128 _6297_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_139 _6451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_640 _6131_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_651 _6145_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_662 _6482_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_673 _7222_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_684 input80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_695 _4116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3690_ input57/X _3583_/X _6011_/A _7591_/Q _3689_/X VGND VGND VPWR VPWR _3691_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput305 _3624_/X VGND VGND VPWR VPWR serial_data_2 sky130_fd_sc_hd__buf_12
X_5360_ _4707_/X _4770_/A _5512_/B _4761_/A _5359_/X VGND VGND VPWR VPWR _5597_/A
+ sky130_fd_sc_hd__a221oi_2
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput316 hold608/X VGND VGND VPWR VPWR hold609/A sky130_fd_sc_hd__buf_12
XFILLER_114_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput327 hold642/X VGND VGND VPWR VPWR hold643/A sky130_fd_sc_hd__buf_12
X_4311_ _5991_/A1 hold604/X _4311_/S VGND VGND VPWR VPWR _4311_/X sky130_fd_sc_hd__mux2_1
Xoutput338 hold667/X VGND VGND VPWR VPWR hold668/A sky130_fd_sc_hd__buf_12
X_5291_ _5313_/A _5291_/B _5291_/C VGND VGND VPWR VPWR _5291_/X sky130_fd_sc_hd__and3_1
XFILLER_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7030_ _7617_/CLK _7030_/D fanout624/X VGND VGND VPWR VPWR _7030_/Q sky130_fd_sc_hd__dfrtp_1
X_4242_ _4257_/S _4240_/X _4241_/Y hold29/X VGND VGND VPWR VPWR _4258_/S sky130_fd_sc_hd__o211a_4
XFILLER_113_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4173_ _6920_/Q _6919_/Q VGND VGND VPWR VPWR _4179_/A sky130_fd_sc_hd__nand2b_1
XFILLER_67_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6814_ _6968_/D _4119_/B _6813_/Y _6814_/B2 VGND VGND VPWR VPWR _7663_/D sky130_fd_sc_hd__a22o_1
XFILLER_168_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6745_ _7108_/Q _6099_/B _6694_/C _6474_/A _7171_/Q VGND VGND VPWR VPWR _6745_/X
+ sky130_fd_sc_hd__a32o_1
X_3957_ _7587_/Q _5939_/B _6038_/B _4275_/S input72/X VGND VGND VPWR VPWR _3957_/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_149_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6676_ _7409_/Q _6466_/X _6487_/X _7473_/Q VGND VGND VPWR VPWR _6676_/X sky130_fd_sc_hd__a22o_1
X_3888_ _7289_/Q _5682_/C _5678_/B _3530_/X _7540_/Q VGND VGND VPWR VPWR _3888_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_137_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5627_ _5627_/A1 wire535/X _5626_/X _5624_/X VGND VGND VPWR VPWR _7250_/D sky130_fd_sc_hd__a211o_1
XFILLER_191_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5558_ _5558_/A _5558_/B VGND VGND VPWR VPWR _5558_/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4509_ _4509_/A0 _6865_/A1 _4510_/S VGND VGND VPWR VPWR _4509_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5489_ _5490_/C _4801_/C _5490_/A _5488_/X VGND VGND VPWR VPWR _5493_/B sky130_fd_sc_hd__a31o_1
XFILLER_78_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7228_ _7398_/CLK _7228_/D fanout625/X VGND VGND VPWR VPWR _7228_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout510 hold102/X VGND VGND VPWR VPWR _6046_/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_104_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout521 hold19/X VGND VGND VPWR VPWR _5926_/A0 sky130_fd_sc_hd__buf_8
Xfanout532 hold80/X VGND VGND VPWR VPWR hold81/A sky130_fd_sc_hd__buf_6
XFILLER_132_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout543 _6862_/A1 VGND VGND VPWR VPWR _5697_/A0 sky130_fd_sc_hd__buf_6
X_7159_ _7215_/CLK _7159_/D _6903_/A VGND VGND VPWR VPWR _7159_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout565 _6416_/B VGND VGND VPWR VPWR _6392_/B sky130_fd_sc_hd__buf_6
XFILLER_58_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout587 _5046_/A VGND VGND VPWR VPWR _5297_/A sky130_fd_sc_hd__buf_6
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout598 fanout600/X VGND VGND VPWR VPWR fanout598/X sky130_fd_sc_hd__buf_6
XFILLER_58_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4860_ _4866_/A _4860_/B _4877_/C _4950_/C VGND VGND VPWR VPWR _4935_/C sky130_fd_sc_hd__and4_4
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_470 _7049_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_481 _7232_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_492 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3811_ _7477_/Q _3516_/X _5957_/B _3552_/X _7389_/Q VGND VGND VPWR VPWR _3811_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_60_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4791_ _4781_/Y _4884_/A _4572_/X _4788_/X VGND VGND VPWR VPWR _4791_/Y sky130_fd_sc_hd__a211oi_1
XANTENNA_17 _3516_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 _5661_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_39 _3546_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6530_ _7611_/Q _6451_/X _6466_/X _7403_/Q _6529_/X VGND VGND VPWR VPWR _6530_/X
+ sky130_fd_sc_hd__a221o_1
X_3742_ _7686_/Q _4559_/B hold98/A _3739_/X _3741_/X VGND VGND VPWR VPWR _3753_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_13_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6461_ _7490_/Q _6771_/B _6563_/C VGND VGND VPWR VPWR _6461_/X sky130_fd_sc_hd__and3_1
X_3673_ hold96/X _3673_/B _3673_/C hold69/X VGND VGND VPWR VPWR hold97/A sky130_fd_sc_hd__nor4_4
XFILLER_173_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5412_ _4948_/A _5429_/D _5102_/B _4993_/Y VGND VGND VPWR VPWR _5412_/X sky130_fd_sc_hd__o31a_1
X_6392_ _6231_/B _6392_/B _6416_/C _7182_/Q VGND VGND VPWR VPWR _6392_/X sky130_fd_sc_hd__and4b_1
XFILLER_127_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5343_ _5463_/A _5534_/A _5463_/B _5343_/D VGND VGND VPWR VPWR _5344_/D sky130_fd_sc_hd__and4_1
XFILLER_142_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput179 _3446_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[13] sky130_fd_sc_hd__buf_12
X_5274_ _4629_/Y _5011_/C _5407_/C _4854_/X VGND VGND VPWR VPWR _5274_/X sky130_fd_sc_hd__a211o_1
XFILLER_102_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7013_ _7597_/CLK _7013_/D fanout626/X VGND VGND VPWR VPWR _7705_/A sky130_fd_sc_hd__dfrtp_1
X_4225_ hold83/X hold89/X _4229_/S VGND VGND VPWR VPWR hold90/A sky130_fd_sc_hd__mux2_2
XFILLER_87_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4156_ _6996_/Q _4171_/D _6922_/Q VGND VGND VPWR VPWR _4156_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4087_ _4085_/B hold22/A _4086_/S VGND VGND VPWR VPWR _6924_/D sky130_fd_sc_hd__o21a_1
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4989_ _4992_/D _5195_/B _5476_/B _4989_/D VGND VGND VPWR VPWR _4989_/X sky130_fd_sc_hd__and4b_1
X_6728_ _7072_/Q _6469_/A _6536_/C _6482_/X _7112_/Q VGND VGND VPWR VPWR _6728_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_137_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6659_ _6659_/A _6659_/B _6659_/C _6809_/D VGND VGND VPWR VPWR _6659_/Y sky130_fd_sc_hd__nor4_1
XFILLER_164_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout384 hold70/X VGND VGND VPWR VPWR _4505_/B sky130_fd_sc_hd__buf_12
XFILLER_59_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput15 mask_rev_in[1] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__clkbuf_1
Xinput26 mask_rev_in[2] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput37 mgmt_gpio_in[10] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput48 mgmt_gpio_in[20] VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__clkbuf_4
Xinput59 mgmt_gpio_in[30] VGND VGND VPWR VPWR input59/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4010_ _7546_/Q _3514_/X _3565_/X _7322_/Q _4009_/X VGND VGND VPWR VPWR _4010_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5961_ hold46/X hold9/X _5965_/S VGND VGND VPWR VPWR hold47/A sky130_fd_sc_hd__mux2_1
XFILLER_80_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7700_ _7700_/A VGND VGND VPWR VPWR _7700_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4912_ _5490_/C _4946_/A VGND VGND VPWR VPWR _4912_/Y sky130_fd_sc_hd__nand2_4
X_5892_ hold579/X _6045_/A1 _5893_/S VGND VGND VPWR VPWR _5892_/X sky130_fd_sc_hd__mux2_1
X_7631_ _4167_/A1 _7631_/D fanout620/X VGND VGND VPWR VPWR _7631_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_33_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4843_ _4779_/X _4833_/X _4907_/A _4860_/B _4853_/C VGND VGND VPWR VPWR _4953_/B
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_21_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7562_ _7562_/CLK hold64/X fanout632/X VGND VGND VPWR VPWR _7562_/Q sky130_fd_sc_hd__dfstp_4
X_4774_ _4943_/A _5375_/A _5186_/C _5595_/B _5182_/A VGND VGND VPWR VPWR _4775_/D
+ sky130_fd_sc_hd__a41oi_2
XFILLER_165_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6513_ _7523_/Q _6447_/X _6457_/X _7571_/Q _6512_/X VGND VGND VPWR VPWR _6523_/A
+ sky130_fd_sc_hd__a221o_1
X_3725_ _7188_/Q _5993_/A _5680_/A _3555_/X _7518_/Q VGND VGND VPWR VPWR _3725_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_146_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7493_ _7580_/CLK hold41/X fanout607/X VGND VGND VPWR VPWR hold40/A sky130_fd_sc_hd__dfrtp_4
XFILLER_9_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6444_ _7631_/Q _6485_/B _6469_/A _6771_/C VGND VGND VPWR VPWR _6444_/X sky130_fd_sc_hd__and4_4
X_3656_ _3655_/Y _6948_/Q _3967_/S VGND VGND VPWR VPWR _3656_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6375_ _7221_/Q _7626_/Q _6416_/B _6416_/C VGND VGND VPWR VPWR _6375_/X sky130_fd_sc_hd__and4_1
XFILLER_115_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3587_ _5661_/A _4340_/A _5680_/B VGND VGND VPWR VPWR _6011_/A sky130_fd_sc_hd__and3_4
X_5326_ _5325_/X _5190_/X _6829_/D _5326_/B2 VGND VGND VPWR VPWR _7245_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_161_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5257_ _4867_/X _4889_/Y _5009_/Y _5088_/Y _5256_/X VGND VGND VPWR VPWR _5258_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_87_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4208_ _4208_/A0 _5869_/A1 _4208_/S VGND VGND VPWR VPWR _4208_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5188_ _5188_/A _5555_/D VGND VGND VPWR VPWR _5188_/X sky130_fd_sc_hd__and2_1
XFILLER_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4139_ _6811_/S _4140_/B VGND VGND VPWR VPWR _4139_/X sky130_fd_sc_hd__and2_1
XFILLER_28_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3510_ _4229_/S hold22/X hold128/X VGND VGND VPWR VPWR _3622_/B sky130_fd_sc_hd__o21a_4
XFILLER_128_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4490_ hold359/X _5789_/A1 _4492_/S VGND VGND VPWR VPWR _4490_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold607 hold607/A VGND VGND VPWR VPWR wb_dat_o[15] sky130_fd_sc_hd__buf_12
XFILLER_6_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold618 _5793_/X VGND VGND VPWR VPWR _7392_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold629 hold629/A VGND VGND VPWR VPWR wb_dat_o[13] sky130_fd_sc_hd__buf_12
XFILLER_6_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3441_ _7461_/Q VGND VGND VPWR VPWR _3441_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6160_ _6158_/D _7626_/Q _6416_/B _6160_/D VGND VGND VPWR VPWR _6160_/X sky130_fd_sc_hd__and4bb_4
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5111_ _5316_/A _5112_/B _5311_/C _5111_/D VGND VGND VPWR VPWR _5111_/Y sky130_fd_sc_hd__nand4_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6091_ _7629_/Q _7628_/Q VGND VGND VPWR VPWR _6487_/A sky130_fd_sc_hd__and2_2
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1307 _5899_/X VGND VGND VPWR VPWR _7486_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5042_ _5042_/A _5311_/C _5042_/C VGND VGND VPWR VPWR _5050_/B sky130_fd_sc_hd__and3_1
Xhold1318 _6006_/X VGND VGND VPWR VPWR _7581_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1329 _5782_/X VGND VGND VPWR VPWR _7382_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6993_ _7583_/CLK _6993_/D fanout629/X VGND VGND VPWR VPWR _7701_/A sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_51_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7569_/CLK sky130_fd_sc_hd__clkbuf_16
X_5944_ hold421/X _6043_/A1 _5947_/S VGND VGND VPWR VPWR _5944_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5875_ hold527/X _6028_/A1 _5875_/S VGND VGND VPWR VPWR _5875_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_580 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7614_ _7614_/CLK _7614_/D fanout606/X VGND VGND VPWR VPWR _7614_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4826_ _4597_/Y _4811_/Y _4821_/Y _4825_/Y _4817_/Y VGND VGND VPWR VPWR _4827_/C
+ sky130_fd_sc_hd__o32a_1
Xclkbuf_leaf_66_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7606_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_178_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7545_ _7545_/CLK _7545_/D fanout613/X VGND VGND VPWR VPWR _7545_/Q sky130_fd_sc_hd__dfrtp_1
X_4757_ _4597_/B _4597_/C _4614_/X _4660_/C _4756_/Y VGND VGND VPWR VPWR _4762_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3708_ _4511_/A _5682_/B _4511_/C VGND VGND VPWR VPWR _4346_/A sky130_fd_sc_hd__and3_2
X_7476_ _7603_/CLK _7476_/D fanout606/X VGND VGND VPWR VPWR _7476_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_175_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4688_ _5197_/A _4688_/B _4688_/C VGND VGND VPWR VPWR _5005_/C sky130_fd_sc_hd__and3_1
XFILLER_146_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6427_ _7233_/Q _6160_/D _6427_/A3 _6427_/B1 _7115_/Q VGND VGND VPWR VPWR _6427_/X
+ sky130_fd_sc_hd__a32o_1
X_3639_ hold74/A _5939_/B _5686_/B _5650_/A _7278_/Q VGND VGND VPWR VPWR _3639_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_161_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6358_ _7082_/Q _6146_/X _6151_/X _7215_/Q _6357_/X VGND VGND VPWR VPWR _6358_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5309_ _4825_/Y _4882_/Y _5611_/A2 _4987_/Y VGND VGND VPWR VPWR _5310_/C sky130_fd_sc_hd__a211o_1
XFILLER_130_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6289_ _7552_/Q _6151_/X _6153_/X _7568_/Q _6288_/X VGND VGND VPWR VPWR _6289_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_19_csclk _7202_/CLK VGND VGND VPWR VPWR _7305_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_17_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold4 hold4/A VGND VGND VPWR VPWR hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3990_ _7204_/Q _5984_/A _5666_/B _3702_/X _7061_/Q VGND VGND VPWR VPWR _3990_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_90_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5660_ hold887/X _6862_/A1 _5660_/S VGND VGND VPWR VPWR _7280_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4611_ _4760_/D _4760_/C _4760_/B VGND VGND VPWR VPWR _4704_/D sky130_fd_sc_hd__nand3_2
XFILLER_176_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5591_ _5490_/X _5491_/Y _5591_/C _5591_/D VGND VGND VPWR VPWR _5591_/X sky130_fd_sc_hd__and4bb_1
XFILLER_190_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7330_ _7586_/CLK _7330_/D fanout625/X VGND VGND VPWR VPWR _7330_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_144_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4542_ hold817/X _6003_/A1 _4546_/S VGND VGND VPWR VPWR _4542_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold404 _4420_/X VGND VGND VPWR VPWR _7117_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7261_ _7307_/CLK _7261_/D _6886_/A VGND VGND VPWR VPWR _7261_/Q sky130_fd_sc_hd__dfrtp_4
Xhold415 _7534_/Q VGND VGND VPWR VPWR hold415/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold426 hold426/A VGND VGND VPWR VPWR hold426/X sky130_fd_sc_hd__dlygate4sd3_1
X_4473_ _4473_/A0 _6865_/A1 _4474_/S VGND VGND VPWR VPWR _4473_/X sky130_fd_sc_hd__mux2_1
Xhold437 _4258_/X VGND VGND VPWR VPWR _6995_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 hold448/A VGND VGND VPWR VPWR hold448/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold459 _5630_/X VGND VGND VPWR VPWR _7252_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6212_ _7429_/Q _6432_/A3 _6209_/X _6212_/C1 _6211_/X VGND VGND VPWR VPWR _6212_/X
+ sky130_fd_sc_hd__a2111o_1
X_3424_ _7631_/Q VGND VGND VPWR VPWR _4126_/B sky130_fd_sc_hd__inv_2
XFILLER_131_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7192_ _7192_/CLK _7192_/D fanout619/X VGND VGND VPWR VPWR _7192_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6143_ _7482_/Q _6427_/B1 _6407_/A3 _7490_/Q _6142_/X VGND VGND VPWR VPWR _6143_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1104 _5748_/X VGND VGND VPWR VPWR _7352_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6074_ _6392_/B _6065_/Y _6073_/X _6109_/B VGND VGND VPWR VPWR _7625_/D sky130_fd_sc_hd__a22o_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1115 _5835_/X VGND VGND VPWR VPWR _7429_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1126 _4473_/X VGND VGND VPWR VPWR _7167_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 _7066_/Q VGND VGND VPWR VPWR _4359_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5025_ _5030_/D _5025_/B _5025_/C VGND VGND VPWR VPWR _5233_/C sky130_fd_sc_hd__and3_4
XFILLER_100_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1148 _4356_/X VGND VGND VPWR VPWR _7064_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1159 hold1556/X VGND VGND VPWR VPWR _4532_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6976_ _7289_/CLK _6976_/D fanout598/X VGND VGND VPWR VPWR _6976_/Q sky130_fd_sc_hd__dfstp_2
X_5927_ _5999_/A1 hold810/X hold76/A VGND VGND VPWR VPWR _5927_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5858_ _5903_/A _6002_/A _6038_/C VGND VGND VPWR VPWR _5866_/S sky130_fd_sc_hd__and3_4
XFILLER_166_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4809_ _5311_/A _5071_/B _5071_/C VGND VGND VPWR VPWR _4814_/A sky130_fd_sc_hd__and3_1
X_5789_ hold220/X _5789_/A1 _5794_/S VGND VGND VPWR VPWR _5789_/X sky130_fd_sc_hd__mux2_1
X_7528_ _7608_/CLK _7528_/D fanout611/X VGND VGND VPWR VPWR _7528_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7459_ _7459_/CLK _7459_/D fanout606/X VGND VGND VPWR VPWR _7459_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_135_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold960 _7607_/Q VGND VGND VPWR VPWR hold960/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold971 _7339_/Q VGND VGND VPWR VPWR hold971/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold982 hold982/A VGND VGND VPWR VPWR hold982/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold993 _7188_/Q VGND VGND VPWR VPWR hold993/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6830_ _6969_/Q _6830_/A2 _6830_/B1 _6970_/Q VGND VGND VPWR VPWR _6830_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6761_ _6760_/Y _6759_/X _6761_/B1 _7140_/Q VGND VGND VPWR VPWR _6761_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_62_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3973_ _7474_/Q _6861_/A _3529_/X _3531_/X _7482_/Q VGND VGND VPWR VPWR _3973_/X
+ sky130_fd_sc_hd__a32o_1
X_5712_ _6045_/A1 hold523/X hold38/X VGND VGND VPWR VPWR _5712_/X sky130_fd_sc_hd__mux2_1
X_6692_ _7101_/Q _6486_/X _6487_/X _7126_/Q _6691_/X VGND VGND VPWR VPWR _6692_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5643_ _5678_/C hold98/X _5680_/C VGND VGND VPWR VPWR _5649_/S sky130_fd_sc_hd__and3_2
XFILLER_163_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5574_ _4709_/Y _4960_/Y _4859_/Y _4854_/X VGND VGND VPWR VPWR _5575_/C sky130_fd_sc_hd__a211o_1
X_7313_ _7616_/CLK _7313_/D fanout610/X VGND VGND VPWR VPWR _7313_/Q sky130_fd_sc_hd__dfrtp_1
Xhold201 _7115_/Q VGND VGND VPWR VPWR hold201/X sky130_fd_sc_hd__dlygate4sd3_1
X_4525_ _5761_/A1 hold473/X _4528_/S VGND VGND VPWR VPWR _4525_/X sky130_fd_sc_hd__mux2_1
Xhold212 _5818_/X VGND VGND VPWR VPWR _7414_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 hold223/A VGND VGND VPWR VPWR hold223/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 _7342_/Q VGND VGND VPWR VPWR hold234/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 _7470_/Q VGND VGND VPWR VPWR hold245/X sky130_fd_sc_hd__dlygate4sd3_1
X_7244_ _7679_/CLK _7244_/D fanout635/X VGND VGND VPWR VPWR _7244_/Q sky130_fd_sc_hd__dfrtp_4
X_4456_ _3966_/X _4456_/A1 _4462_/S VGND VGND VPWR VPWR _7152_/D sky130_fd_sc_hd__mux2_1
Xhold256 _7457_/Q VGND VGND VPWR VPWR hold256/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 _7010_/Q VGND VGND VPWR VPWR hold267/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold278 _7198_/Q VGND VGND VPWR VPWR hold278/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold289 _7705_/A VGND VGND VPWR VPWR hold289/X sky130_fd_sc_hd__dlygate4sd3_1
X_7175_ _7197_/CLK _7175_/D fanout615/X VGND VGND VPWR VPWR _7175_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_132_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4387_ _5926_/A0 hold494/X _4387_/S VGND VGND VPWR VPWR _4387_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6126_ _7623_/Q _6151_/B _7624_/Q _6126_/D VGND VGND VPWR VPWR _6309_/C sky130_fd_sc_hd__and4bb_4
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6057_ _7619_/Q _7620_/Q _7142_/Q _6811_/S VGND VGND VPWR VPWR _6057_/X sky130_fd_sc_hd__o22a_1
XTAP_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5008_ _5007_/A _5017_/A _5008_/C _5014_/D VGND VGND VPWR VPWR _5111_/D sky130_fd_sc_hd__and4bb_4
XFILLER_39_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 _6132_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 _6138_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_129 _6329_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6959_ _7286_/CLK _6959_/D fanout604/X VGND VGND VPWR VPWR _6959_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_121_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold790 hold790/A VGND VGND VPWR VPWR hold790/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1490 _4092_/X VGND VGND VPWR VPWR _6922_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_630 _5233_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_641 _6170_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_652 _6145_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_663 _6486_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_674 _7222_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_685 input80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_696 _4116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_0__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _7258_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_60_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput306 _4170_/X VGND VGND VPWR VPWR serial_load sky130_fd_sc_hd__buf_12
Xoutput317 hold808/X VGND VGND VPWR VPWR hold809/A sky130_fd_sc_hd__buf_12
X_4310_ _6044_/A1 hold845/X _4311_/S VGND VGND VPWR VPWR _4310_/X sky130_fd_sc_hd__mux2_1
Xoutput328 hold657/X VGND VGND VPWR VPWR hold658/A sky130_fd_sc_hd__buf_12
XFILLER_114_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput339 hold684/X VGND VGND VPWR VPWR hold685/A sky130_fd_sc_hd__buf_12
X_5290_ _5313_/B _5290_/A2 _5291_/B _5038_/B _5311_/A VGND VGND VPWR VPWR _5290_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_113_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4241_ _7294_/Q _4171_/C _4171_/D _5666_/B VGND VGND VPWR VPWR _4241_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_68_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4172_ hold42/A _4172_/A2 _4171_/Y _4172_/B2 VGND VGND VPWR VPWR _4172_/X sky130_fd_sc_hd__a22o_2
XFILLER_67_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6813_ _6961_/Q _6965_/Q _6962_/Q _6968_/Q _4119_/B VGND VGND VPWR VPWR _6813_/Y
+ sky130_fd_sc_hd__o41ai_1
XFILLER_23_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3956_ _7579_/Q _3584_/X _3952_/X _3954_/X _3955_/X VGND VGND VPWR VPWR _3964_/C
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_149_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6744_ _7078_/Q _6450_/X _6483_/X _7068_/Q _6743_/X VGND VGND VPWR VPWR _6744_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_51_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6675_ _6675_/A _6675_/B _6675_/C _6675_/D VGND VGND VPWR VPWR _6675_/Y sky130_fd_sc_hd__nor4_1
X_3887_ _7564_/Q _3554_/X _3712_/X _7206_/Q _3886_/X VGND VGND VPWR VPWR _3887_/X
+ sky130_fd_sc_hd__a221o_1
X_5626_ _5603_/Y _5625_/Y _5626_/C _5626_/D VGND VGND VPWR VPWR _5626_/X sky130_fd_sc_hd__and4bb_1
X_5557_ _4867_/X _5381_/X _5451_/B _5526_/C _5526_/A VGND VGND VPWR VPWR _5557_/Y
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_117_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4508_ _4508_/A0 _6864_/A1 _4510_/S VGND VGND VPWR VPWR _4508_/X sky130_fd_sc_hd__mux2_1
X_5488_ _5364_/B _5485_/X _5168_/X VGND VGND VPWR VPWR _5488_/X sky130_fd_sc_hd__a21bo_1
XFILLER_117_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4439_ _6864_/A1 _4439_/A1 _4444_/S VGND VGND VPWR VPWR _4439_/X sky130_fd_sc_hd__mux2_1
X_7227_ _7227_/CLK _7227_/D fanout619/X VGND VGND VPWR VPWR _7227_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_104_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout511 hold101/X VGND VGND VPWR VPWR hold102/A sky130_fd_sc_hd__buf_8
XFILLER_132_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout522 hold19/X VGND VGND VPWR VPWR _5935_/A1 sky130_fd_sc_hd__buf_6
Xfanout533 hold80/X VGND VGND VPWR VPWR _5789_/A1 sky130_fd_sc_hd__buf_8
XFILLER_160_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7158_ _7668_/CLK _7158_/D VGND VGND VPWR VPWR _7158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout544 _6039_/A1 VGND VGND VPWR VPWR _6862_/A1 sky130_fd_sc_hd__buf_8
XFILLER_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout555 _6082_/B VGND VGND VPWR VPWR _6159_/B sky130_fd_sc_hd__buf_12
Xfanout566 _7625_/Q VGND VGND VPWR VPWR _6416_/B sky130_fd_sc_hd__buf_4
X_6109_ _6811_/S _6109_/B VGND VGND VPWR VPWR _6109_/X sky130_fd_sc_hd__and2b_4
XFILLER_58_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout577 _5093_/B VGND VGND VPWR VPWR _5452_/B sky130_fd_sc_hd__buf_8
XFILLER_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout588 _3460_/Y VGND VGND VPWR VPWR _5429_/D sky130_fd_sc_hd__clkbuf_16
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7089_ _7254_/CLK _7089_/D fanout617/X VGND VGND VPWR VPWR _7089_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout599 fanout600/X VGND VGND VPWR VPWR fanout599/X sky130_fd_sc_hd__buf_8
XFILLER_58_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_460 _6583_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_471 _7122_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_482 _7232_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3810_ _7469_/Q _3528_/X hold75/A _7509_/Q _3809_/X VGND VGND VPWR VPWR _3815_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA_493 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4790_ _4884_/A _4781_/Y _4788_/X VGND VGND VPWR VPWR _4953_/A sky130_fd_sc_hd__a21o_2
XANTENNA_18 _3516_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_29 _5682_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3741_ _7173_/Q _3700_/X _3713_/X _7100_/Q _3740_/X VGND VGND VPWR VPWR _3741_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_186_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6460_ _6563_/C _6791_/D _6645_/C VGND VGND VPWR VPWR _6460_/X sky130_fd_sc_hd__and3_4
X_3672_ _7495_/Q _5903_/A _5975_/B _3531_/X _7487_/Q VGND VGND VPWR VPWR _3672_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_173_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5411_ _5285_/X _4993_/Y _4960_/Y _5604_/B1 _4987_/Y VGND VGND VPWR VPWR _5605_/B
+ sky130_fd_sc_hd__a311o_1
X_6391_ _6391_/A1 _4139_/X _6109_/X _6390_/X VGND VGND VPWR VPWR _7647_/D sky130_fd_sc_hd__o31a_1
X_5342_ _5339_/X _5011_/A _5201_/D _5341_/X VGND VGND VPWR VPWR _5343_/D sky130_fd_sc_hd__o211a_1
XFILLER_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5273_ _5273_/A _5273_/B _5273_/C VGND VGND VPWR VPWR _5279_/A sky130_fd_sc_hd__and3_1
XFILLER_114_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7012_ _7597_/CLK _7012_/D fanout626/X VGND VGND VPWR VPWR _7704_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_101_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4224_ hold222/X _6866_/A1 _4230_/S VGND VGND VPWR VPWR _6976_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4155_ _6997_/Q _4172_/B2 _6954_/Q VGND VGND VPWR VPWR _4155_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4086_ _3505_/Y _3506_/X _4086_/S VGND VGND VPWR VPWR _6925_/D sky130_fd_sc_hd__mux2_1
XFILLER_71_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4988_ _5094_/A _5131_/A _5512_/C VGND VGND VPWR VPWR _4989_/D sky130_fd_sc_hd__and3_1
XFILLER_168_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6727_ _7170_/Q _6474_/A _6456_/X _7160_/Q _6726_/X VGND VGND VPWR VPWR _6734_/A
+ sky130_fd_sc_hd__a221o_1
X_3939_ _7225_/Q _4541_/A _4469_/B _3697_/X _7165_/Q VGND VGND VPWR VPWR _3946_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_177_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6658_ _7456_/Q _6459_/X _6460_/X _7448_/Q _6657_/X VGND VGND VPWR VPWR _6659_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_192_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5609_ _5311_/A _5131_/B _5291_/C _5094_/D _5432_/X VGND VGND VPWR VPWR _5610_/D
+ sky130_fd_sc_hd__a41o_1
X_6589_ _7606_/Q _6791_/B _6791_/C _6791_/D VGND VGND VPWR VPWR _6589_/X sky130_fd_sc_hd__and4_1
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout385 hold107/X VGND VGND VPWR VPWR _5984_/B sky130_fd_sc_hd__buf_12
XFILLER_143_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput16 mask_rev_in[20] VGND VGND VPWR VPWR input16/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput27 mask_rev_in[30] VGND VGND VPWR VPWR input27/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput38 mgmt_gpio_in[11] VGND VGND VPWR VPWR input38/X sky130_fd_sc_hd__buf_4
XFILLER_167_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput49 mgmt_gpio_in[21] VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__clkbuf_2
XFILLER_182_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5960_ hold769/X _6041_/A1 _5965_/S VGND VGND VPWR VPWR _5960_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4911_ _4935_/B _5007_/D _4946_/A VGND VGND VPWR VPWR _4925_/C sky130_fd_sc_hd__and3_1
X_5891_ hold804/X _5999_/A1 _5893_/S VGND VGND VPWR VPWR _5891_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7630_ _4167_/A1 _7630_/D fanout620/X VGND VGND VPWR VPWR _7630_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_290 _7713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4842_ _4907_/C _4935_/B VGND VGND VPWR VPWR _4957_/B sky130_fd_sc_hd__nor2_2
XFILLER_60_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7561_ _7569_/CLK _7561_/D fanout614/X VGND VGND VPWR VPWR _7561_/Q sky130_fd_sc_hd__dfrtp_1
X_4773_ _5375_/A _5429_/A _5313_/C VGND VGND VPWR VPWR _5182_/A sky130_fd_sc_hd__and3_1
XFILLER_158_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3724_ _7130_/Q _4559_/B _5678_/B _3701_/X _7243_/Q VGND VGND VPWR VPWR _3724_/X
+ sky130_fd_sc_hd__a32o_1
X_6512_ _7395_/Q _6463_/X _6486_/X _7499_/Q _6511_/X VGND VGND VPWR VPWR _6512_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7492_ _7541_/CLK _7492_/D fanout609/X VGND VGND VPWR VPWR _7492_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_119_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6443_ _6771_/C VGND VGND VPWR VPWR _6443_/Y sky130_fd_sc_hd__inv_2
X_3655_ _3655_/A _3655_/B VGND VGND VPWR VPWR _3655_/Y sky130_fd_sc_hd__nand2_4
XFILLER_173_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6374_ _7171_/Q _6131_/C _6371_/X _6373_/X VGND VGND VPWR VPWR _6374_/X sky130_fd_sc_hd__a211o_1
XFILLER_173_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3586_ _3586_/A _5661_/B _5680_/B VGND VGND VPWR VPWR _4275_/S sky130_fd_sc_hd__and3_4
XFILLER_115_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5325_ _5282_/X _5325_/B _5325_/C _6829_/D VGND VGND VPWR VPWR _5325_/X sky130_fd_sc_hd__and4b_1
XFILLER_130_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5256_ _5256_/A _5256_/B _5256_/C VGND VGND VPWR VPWR _5256_/X sky130_fd_sc_hd__and3_1
X_4207_ hold4/X _6835_/A0 _4229_/S VGND VGND VPWR VPWR hold5/A sky130_fd_sc_hd__mux2_8
XFILLER_87_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5187_ _4597_/Y _4811_/Y _4821_/Y _5186_/Y VGND VGND VPWR VPWR _5187_/X sky130_fd_sc_hd__o31a_1
XFILLER_56_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4138_ _4118_/B _4117_/X _4133_/X _4201_/B VGND VGND VPWR VPWR _6967_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4069_ _4069_/A _4069_/B VGND VGND VPWR VPWR _6931_/D sky130_fd_sc_hd__nor2_1
XFILLER_44_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire572 _5096_/Y VGND VGND VPWR VPWR wire572/X sky130_fd_sc_hd__clkbuf_2
Xhold608 hold608/A VGND VGND VPWR VPWR hold608/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3440_ _7469_/Q VGND VGND VPWR VPWR _3440_/Y sky130_fd_sc_hd__inv_2
Xhold619 _7710_/A VGND VGND VPWR VPWR hold619/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5110_ _5313_/B _5452_/B _5110_/C VGND VGND VPWR VPWR _5110_/X sky130_fd_sc_hd__and3_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6090_ _7139_/Q _6109_/B _6090_/A3 _6645_/B _6089_/Y VGND VGND VPWR VPWR _7629_/D
+ sky130_fd_sc_hd__o32a_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _5322_/C _5311_/C _5042_/C VGND VGND VPWR VPWR _5050_/A sky130_fd_sc_hd__and3_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1308 _7323_/Q VGND VGND VPWR VPWR hold978/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1319 _7487_/Q VGND VGND VPWR VPWR hold783/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_wb_clk_i wb_clk_i VGND VGND VPWR VPWR clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_93_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6992_ _7583_/CLK _6992_/D fanout629/X VGND VGND VPWR VPWR _7700_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_65_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5943_ hold87/X hold9/X _5947_/S VGND VGND VPWR VPWR hold88/A sky130_fd_sc_hd__mux2_1
XFILLER_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5874_ hold467/X _6045_/A1 _5875_/S VGND VGND VPWR VPWR _5874_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7613_ _7613_/CLK _7613_/D fanout626/X VGND VGND VPWR VPWR _7613_/Q sky130_fd_sc_hd__dfrtp_4
X_4825_ _5146_/A _5146_/B VGND VGND VPWR VPWR _4825_/Y sky130_fd_sc_hd__nand2_4
XFILLER_166_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7544_ _7608_/CLK _7544_/D fanout610/X VGND VGND VPWR VPWR _7544_/Q sky130_fd_sc_hd__dfrtp_2
X_4756_ _5131_/A _5131_/B VGND VGND VPWR VPWR _4756_/Y sky130_fd_sc_hd__nand2_4
XFILLER_159_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3707_ _7055_/Q _6038_/B _4553_/B VGND VGND VPWR VPWR _3707_/X sky130_fd_sc_hd__and3_1
XFILLER_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7475_ _7580_/CLK _7475_/D fanout605/X VGND VGND VPWR VPWR _7475_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_107_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4687_ _3460_/Y _5000_/C _4568_/Y _4649_/X _5015_/C VGND VGND VPWR VPWR _5197_/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_174_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6426_ _7686_/Q _6145_/X _6158_/X _7243_/Q _6425_/X VGND VGND VPWR VPWR _6426_/X
+ sky130_fd_sc_hd__a221o_1
X_3638_ _6978_/Q _3560_/X _5849_/A _7448_/Q _3637_/X VGND VGND VPWR VPWR _3654_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3569_ _3905_/B _3717_/B _5680_/B VGND VGND VPWR VPWR _3569_/X sky130_fd_sc_hd__and3_4
X_6357_ _7190_/Q _6138_/X _6157_/X _7102_/Q _6356_/X VGND VGND VPWR VPWR _6357_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5308_ _5322_/C _5401_/A _5291_/C _5012_/X _5017_/B VGND VGND VPWR VPWR _5610_/B
+ sky130_fd_sc_hd__o2111a_1
X_6288_ _7520_/Q _6131_/B _6115_/X _6144_/X _7544_/Q VGND VGND VPWR VPWR _6288_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5239_ _4943_/A _4926_/B _4934_/C _5089_/A _5092_/A VGND VGND VPWR VPWR _5263_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_130_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_586 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold5 hold5/A VGND VGND VPWR VPWR hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_94_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4610_ _5025_/B _4706_/D _4608_/Y _4760_/C _4760_/D VGND VGND VPWR VPWR _5186_/C
+ sky130_fd_sc_hd__o311a_4
XFILLER_175_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5590_ _4704_/D _4680_/X _5484_/Y _5371_/B _5177_/X VGND VGND VPWR VPWR _5591_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_128_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4541_ _4541_/A _4541_/B _6861_/C VGND VGND VPWR VPWR _4546_/S sky130_fd_sc_hd__and3_2
XFILLER_191_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold405 _7020_/Q VGND VGND VPWR VPWR hold405/X sky130_fd_sc_hd__dlygate4sd3_1
X_7260_ _7293_/CLK _7260_/D _6886_/A VGND VGND VPWR VPWR _7260_/Q sky130_fd_sc_hd__dfstp_2
Xhold416 _5953_/X VGND VGND VPWR VPWR _7534_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4472_ hold361/X _5789_/A1 _4474_/S VGND VGND VPWR VPWR _4472_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold427 hold427/A VGND VGND VPWR VPWR hold427/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold438 _7235_/Q VGND VGND VPWR VPWR hold438/X sky130_fd_sc_hd__dlygate4sd3_1
X_3423_ _4171_/C VGND VGND VPWR VPWR _3423_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6211_ _7325_/Q _6170_/C _6309_/C _7333_/Q _6210_/X VGND VGND VPWR VPWR _6211_/X
+ sky130_fd_sc_hd__a221o_1
Xhold449 hold449/A VGND VGND VPWR VPWR hold449/X sky130_fd_sc_hd__dlygate4sd3_1
X_7191_ _7192_/CLK _7191_/D fanout617/X VGND VGND VPWR VPWR _7191_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_143_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6142_ _7530_/Q _6160_/D _6427_/A3 _6127_/X _7498_/Q VGND VGND VPWR VPWR _6142_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6073_ _6392_/B _6416_/C VGND VGND VPWR VPWR _6073_/X sky130_fd_sc_hd__xor2_1
XFILLER_98_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1105 hold1406/X VGND VGND VPWR VPWR _5745_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1116 _7272_/Q VGND VGND VPWR VPWR _5651_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1127 _7207_/Q VGND VGND VPWR VPWR _4521_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5024_ _5046_/B _5024_/B _5024_/C _5024_/D VGND VGND VPWR VPWR _5047_/D sky130_fd_sc_hd__nand4_1
Xhold1138 _4359_/X VGND VGND VPWR VPWR _7066_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1149 hold1587/X VGND VGND VPWR VPWR _5823_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6975_ _7289_/CLK _6975_/D fanout596/X VGND VGND VPWR VPWR _6975_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5926_ _5926_/A0 hold373/X hold76/A VGND VGND VPWR VPWR _5926_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5857_ _6046_/A1 hold831/X _5857_/S VGND VGND VPWR VPWR _5857_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4808_ _4808_/A _4808_/B VGND VGND VPWR VPWR _4814_/C sky130_fd_sc_hd__nand2_1
XFILLER_186_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5788_ hold979/X _6040_/A1 _5794_/S VGND VGND VPWR VPWR _5788_/X sky130_fd_sc_hd__mux2_1
X_7527_ _7608_/CLK _7527_/D fanout611/X VGND VGND VPWR VPWR _7527_/Q sky130_fd_sc_hd__dfrtp_1
X_4739_ _4739_/A _4739_/B _4739_/C _4739_/D VGND VGND VPWR VPWR _4741_/B sky130_fd_sc_hd__nand4_1
XFILLER_147_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7458_ _7614_/CLK _7458_/D fanout604/X VGND VGND VPWR VPWR _7458_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_135_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6409_ _7129_/Q _6130_/X _6132_/X _7119_/Q _6408_/X VGND VGND VPWR VPWR _6409_/X
+ sky130_fd_sc_hd__a221o_1
Xhold950 _4268_/X VGND VGND VPWR VPWR _6999_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold961 _6035_/X VGND VGND VPWR VPWR _7607_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7389_ _7445_/CLK _7389_/D fanout628/X VGND VGND VPWR VPWR _7389_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_89_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold972 _5734_/X VGND VGND VPWR VPWR _7339_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold983 hold983/A VGND VGND VPWR VPWR hold983/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold994 _4498_/X VGND VGND VPWR VPWR _7188_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1650 _7245_/Q VGND VGND VPWR VPWR _5326_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_50_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7609_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_140_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_65_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7612_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6760_ _7038_/Q _6759_/D _7140_/Q VGND VGND VPWR VPWR _6760_/Y sky130_fd_sc_hd__o21bai_1
X_3972_ _7041_/Q _4529_/B _5680_/B _4463_/A _7159_/Q VGND VGND VPWR VPWR _3972_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5711_ _5999_/A1 hold779/X hold38/X VGND VGND VPWR VPWR _5711_/X sky130_fd_sc_hd__mux2_1
X_6691_ _7056_/Q _6474_/C _6481_/X _7209_/Q VGND VGND VPWR VPWR _6691_/X sky130_fd_sc_hd__a22o_1
X_5642_ hold205/X _6866_/A1 _5642_/S VGND VGND VPWR VPWR _5642_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5573_ _5460_/X _5573_/B _5573_/C _5573_/D VGND VGND VPWR VPWR _5573_/X sky130_fd_sc_hd__and4b_1
X_7312_ _7312_/CLK hold59/X _6891_/A VGND VGND VPWR VPWR hold58/A sky130_fd_sc_hd__dfrtp_1
XFILLER_8_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold202 _4417_/X VGND VGND VPWR VPWR _7115_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4524_ _6012_/A0 hold682/X _4528_/S VGND VGND VPWR VPWR _4524_/X sky130_fd_sc_hd__mux2_1
Xhold213 hold213/A VGND VGND VPWR VPWR hold213/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_18_csclk _7202_/CLK VGND VGND VPWR VPWR _7227_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold224 _7583_/Q VGND VGND VPWR VPWR hold224/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 _5737_/X VGND VGND VPWR VPWR _7342_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold246 _5881_/X VGND VGND VPWR VPWR _7470_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7243_ _7682_/CLK _7243_/D fanout603/X VGND VGND VPWR VPWR _7243_/Q sky130_fd_sc_hd__dfrtp_1
X_4455_ _4037_/Y _4455_/A1 _4462_/S VGND VGND VPWR VPWR _7151_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold257 _5866_/X VGND VGND VPWR VPWR _7457_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold268 _4292_/X VGND VGND VPWR VPWR _7010_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold279 _4510_/X VGND VGND VPWR VPWR _7198_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7174_ _7194_/CLK _7174_/D fanout615/X VGND VGND VPWR VPWR _7174_/Q sky130_fd_sc_hd__dfrtp_1
X_4386_ _6865_/A1 _4386_/A1 _4387_/S VGND VGND VPWR VPWR _4386_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6125_ _7402_/Q _6160_/D _6146_/C _6077_/X _7378_/Q VGND VGND VPWR VPWR _6125_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ _7619_/Q _7620_/Q VGND VGND VPWR VPWR _6056_/Y sky130_fd_sc_hd__nand2_1
XFILLER_100_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5007_ _5007_/A _5017_/A _5008_/C _5007_/D VGND VGND VPWR VPWR _5007_/Y sky130_fd_sc_hd__nor4_2
XFILLER_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_108 _6132_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_119 _6144_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6958_ _7286_/CLK _6958_/D fanout604/X VGND VGND VPWR VPWR _6958_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_81_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5909_ hold759/X _5999_/A1 _5911_/S VGND VGND VPWR VPWR _5909_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6889_ _6899_/A _6908_/B VGND VGND VPWR VPWR _6889_/X sky130_fd_sc_hd__and2_1
XFILLER_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold780 _5711_/X VGND VGND VPWR VPWR _7319_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold791 hold791/A VGND VGND VPWR VPWR wb_dat_o[24] sky130_fd_sc_hd__buf_12
XFILLER_89_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_727 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1480 _7154_/Q VGND VGND VPWR VPWR _4458_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1491 _7098_/Q VGND VGND VPWR VPWR hold1491/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_55_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_620 _3529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_631 _5021_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_642 _6170_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_653 _6145_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_664 _6486_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_675 _7222_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_686 input80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_697 _4116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput307 _4169_/X VGND VGND VPWR VPWR serial_resetn sky130_fd_sc_hd__buf_12
XFILLER_160_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput318 hold628/X VGND VGND VPWR VPWR hold629/A sky130_fd_sc_hd__buf_12
XFILLER_126_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput329 hold721/X VGND VGND VPWR VPWR hold722/A sky130_fd_sc_hd__buf_12
XFILLER_154_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4240_ _7294_/Q _4171_/C _4171_/D _5975_/B _6038_/B VGND VGND VPWR VPWR _4240_/X
+ sky130_fd_sc_hd__o311a_4
XFILLER_113_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4171_ _4229_/S _7294_/Q _4171_/C _4171_/D VGND VGND VPWR VPWR _4171_/Y sky130_fd_sc_hd__nor4_1
XFILLER_67_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6812_ _6811_/X _6812_/A1 _6812_/S VGND VGND VPWR VPWR _6812_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6743_ _7201_/Q _6694_/B _6445_/C _6463_/X _7226_/Q VGND VGND VPWR VPWR _6743_/X
+ sky130_fd_sc_hd__a32o_1
X_3955_ _7240_/Q _3701_/X _3702_/X _7062_/Q VGND VGND VPWR VPWR _3955_/X sky130_fd_sc_hd__a22o_1
XFILLER_188_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6674_ _7545_/Q _6479_/X _6672_/X _6673_/X _6671_/X VGND VGND VPWR VPWR _6675_/D
+ sky130_fd_sc_hd__a2111o_1
X_3886_ _7274_/Q _5650_/A _3702_/X _7063_/Q _3841_/X VGND VGND VPWR VPWR _3886_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_149_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5625_ _5625_/A _5625_/B _5625_/C _5625_/D VGND VGND VPWR VPWR _5625_/Y sky130_fd_sc_hd__nor4_1
XFILLER_137_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5556_ _5544_/C _5542_/X _5554_/Y _5497_/X VGND VGND VPWR VPWR _5558_/B sky130_fd_sc_hd__a22oi_2
XFILLER_191_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4507_ hold199/X _5869_/A1 _4510_/S VGND VGND VPWR VPWR _4507_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5487_ _5486_/X _5547_/C _5487_/C _5547_/B VGND VGND VPWR VPWR _5493_/A sky130_fd_sc_hd__nand4b_1
X_7226_ _7304_/CLK _7226_/D fanout620/X VGND VGND VPWR VPWR _7226_/Q sky130_fd_sc_hd__dfstp_2
X_4438_ _5869_/A1 hold145/X _4444_/S VGND VGND VPWR VPWR _4438_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout512 hold50/X VGND VGND VPWR VPWR _6045_/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout523 hold9/X VGND VGND VPWR VPWR _5673_/A1 sky130_fd_sc_hd__buf_8
X_7157_ _7668_/CLK _7157_/D VGND VGND VPWR VPWR _7157_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout534 hold80/X VGND VGND VPWR VPWR _5843_/A1 sky130_fd_sc_hd__buf_4
XFILLER_113_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4369_ hold184/X _6866_/A1 _4369_/S VGND VGND VPWR VPWR _4369_/X sky130_fd_sc_hd__mux2_1
Xfanout545 hold44/A VGND VGND VPWR VPWR _6039_/A1 sky130_fd_sc_hd__buf_12
Xfanout556 _3458_/Y VGND VGND VPWR VPWR _6082_/B sky130_fd_sc_hd__buf_12
Xfanout567 _7141_/Q VGND VGND VPWR VPWR _6109_/B sky130_fd_sc_hd__buf_8
X_6108_ _6108_/A0 _6107_/X _6108_/S VGND VGND VPWR VPWR _7636_/D sky130_fd_sc_hd__mux2_1
Xfanout578 _5313_/B VGND VGND VPWR VPWR _5291_/C sky130_fd_sc_hd__buf_4
Xfanout589 input99/X VGND VGND VPWR VPWR _5074_/A sky130_fd_sc_hd__buf_12
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7088_ _7254_/CLK _7088_/D fanout617/X VGND VGND VPWR VPWR _7088_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_46_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6039_ hold293/X _6039_/A1 _6046_/S VGND VGND VPWR VPWR _7610_/D sky130_fd_sc_hd__mux2_1
XFILLER_58_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_450 _6474_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_461 _6700_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_472 _7483_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_483 _7232_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_494 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_19 _3516_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3740_ _7238_/Q _5628_/A _4553_/B _3715_/X _7110_/Q VGND VGND VPWR VPWR _3740_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_13_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3671_ _7391_/Q _3552_/X _3556_/X _7431_/Q _3670_/X VGND VGND VPWR VPWR _3678_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_185_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5410_ _5316_/C _5146_/A _5143_/X _5149_/X VGND VGND VPWR VPWR _5602_/C sky130_fd_sc_hd__a31o_1
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6390_ _6811_/S _6390_/A2 _6812_/S _6389_/X VGND VGND VPWR VPWR _6390_/X sky130_fd_sc_hd__a211o_1
X_5341_ _4984_/Y _5018_/Y _5196_/Y _5197_/Y _5340_/X VGND VGND VPWR VPWR _5341_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_114_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5272_ _4953_/A _4953_/B _4953_/C _4953_/D _5573_/B VGND VGND VPWR VPWR _5273_/C
+ sky130_fd_sc_hd__o41a_1
X_7011_ _7584_/CLK _7011_/D fanout613/X VGND VGND VPWR VPWR _7693_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_99_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4223_ hold1/X hold17/X hold42/X VGND VGND VPWR VPWR _4223_/X sky130_fd_sc_hd__mux2_8
XFILLER_114_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4154_ _6998_/Q input58/X _6922_/Q VGND VGND VPWR VPWR _4154_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4085_ _4085_/A _4085_/B VGND VGND VPWR VPWR _4086_/S sky130_fd_sc_hd__nand2_1
XFILLER_55_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4987_ _5094_/A _5131_/A VGND VGND VPWR VPWR _4987_/Y sky130_fd_sc_hd__nand2_4
X_6726_ _7230_/Q _6720_/C _6536_/C _6453_/X _7062_/Q VGND VGND VPWR VPWR _6726_/X
+ sky130_fd_sc_hd__a32o_1
X_3938_ _7210_/Q hold70/A _4511_/C _3565_/X _7323_/Q VGND VGND VPWR VPWR _3946_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_177_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6657_ _7536_/Q _6720_/C _6536_/C _6444_/X _7432_/Q VGND VGND VPWR VPWR _6657_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_137_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3869_ _7103_/Q _3706_/X _3865_/X _3866_/X _3868_/X VGND VGND VPWR VPWR _3883_/A
+ sky130_fd_sc_hd__a2111o_1
XFILLER_109_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5608_ _5291_/C _5313_/A _5095_/C _5607_/X _5610_/C VGND VGND VPWR VPWR _5625_/D
+ sky130_fd_sc_hd__a311o_1
XFILLER_137_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6588_ _7454_/Q _6645_/B _6720_/D _6645_/C VGND VGND VPWR VPWR _6588_/X sky130_fd_sc_hd__and4_1
XFILLER_118_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5539_ _5322_/A _5068_/C _5250_/X _5538_/X VGND VGND VPWR VPWR _5539_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_132_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7209_ _7253_/CLK _7209_/D fanout618/X VGND VGND VPWR VPWR _7209_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_132_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout386 _3535_/X VGND VGND VPWR VPWR _5680_/A sky130_fd_sc_hd__buf_12
XFILLER_19_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout397 _4553_/B VGND VGND VPWR VPWR _5678_/B sky130_fd_sc_hd__buf_8
XFILLER_19_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_730 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput17 mask_rev_in[21] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput28 mask_rev_in[31] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput39 mgmt_gpio_in[12] VGND VGND VPWR VPWR _4199_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_109_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4910_ _4935_/B _5007_/D VGND VGND VPWR VPWR _4910_/Y sky130_fd_sc_hd__nand2_1
X_5890_ hold168/X _6043_/A1 _5893_/S VGND VGND VPWR VPWR _5890_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4841_ _5025_/B _4608_/Y _4865_/B _5007_/D _4836_/Y VGND VGND VPWR VPWR _4877_/D
+ sky130_fd_sc_hd__o32ai_2
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_280 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_291 _7713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7560_ _7616_/CLK _7560_/D fanout611/X VGND VGND VPWR VPWR _7560_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_60_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4772_ _5186_/C _5595_/B VGND VGND VPWR VPWR _4772_/Y sky130_fd_sc_hd__nand2_1
XFILLER_193_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6511_ _7563_/Q _6099_/B _6720_/D _6483_/X _7387_/Q VGND VGND VPWR VPWR _6511_/X
+ sky130_fd_sc_hd__a32o_1
X_3723_ _7287_/Q _5678_/C _5678_/B _3704_/X _7198_/Q VGND VGND VPWR VPWR _3723_/X
+ sky130_fd_sc_hd__a32o_1
X_7491_ _7547_/CLK _7491_/D fanout609/X VGND VGND VPWR VPWR _7491_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_159_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6442_ _7632_/Q _7633_/Q VGND VGND VPWR VPWR _6442_/Y sky130_fd_sc_hd__nor2_1
X_3654_ _3654_/A _3654_/B _3654_/C _3654_/D VGND VGND VPWR VPWR _3655_/B sky130_fd_sc_hd__nor4_2
XFILLER_173_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6373_ _7098_/Q _6432_/A3 _6124_/X _7236_/Q _6372_/X VGND VGND VPWR VPWR _6373_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3585_ _5939_/B _5768_/C _5768_/B VGND VGND VPWR VPWR _3585_/X sky130_fd_sc_hd__and3_2
XFILLER_161_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5324_ _5234_/Y _5235_/X _5323_/Y _4975_/Y VGND VGND VPWR VPWR _5325_/B sky130_fd_sc_hd__a31o_1
XFILLER_114_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5255_ _4953_/B _4859_/Y _4949_/Y _4880_/Y _5254_/X VGND VGND VPWR VPWR _5256_/C
+ sky130_fd_sc_hd__o311a_1
XFILLER_130_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4206_ _4206_/A0 _5697_/A0 _4208_/S VGND VGND VPWR VPWR _4206_/X sky130_fd_sc_hd__mux2_1
X_5186_ _5375_/A _5186_/B _5186_/C _5614_/C VGND VGND VPWR VPWR _5186_/Y sky130_fd_sc_hd__nand4_1
X_4137_ _6969_/Q _4133_/X _4210_/B VGND VGND VPWR VPWR _6969_/D sky130_fd_sc_hd__a21o_1
XFILLER_28_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4068_ _4067_/A _4067_/C hold33/A VGND VGND VPWR VPWR _4069_/B sky130_fd_sc_hd__a21oi_1
XFILLER_71_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6709_ _6709_/A _6709_/B _6709_/C _6809_/D VGND VGND VPWR VPWR _6709_/Y sky130_fd_sc_hd__nor4_1
XFILLER_149_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7689_ _7689_/A VGND VGND VPWR VPWR _7689_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold609 hold609/A VGND VGND VPWR VPWR wb_dat_o[11] sky130_fd_sc_hd__buf_12
XFILLER_156_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _5040_/A _5297_/C _5040_/C _5094_/D VGND VGND VPWR VPWR _5051_/B sky130_fd_sc_hd__nand4_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1309 _5716_/X VGND VGND VPWR VPWR _7323_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_93_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6991_ _7421_/CLK _6991_/D fanout630/X VGND VGND VPWR VPWR _7699_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_19_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5942_ hold383/X hold81/X _5947_/S VGND VGND VPWR VPWR _5942_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5873_ hold659/X _5999_/A1 _5875_/S VGND VGND VPWR VPWR _5873_/X sky130_fd_sc_hd__mux2_1
X_7612_ _7612_/CLK _7612_/D fanout612/X VGND VGND VPWR VPWR _7612_/Q sky130_fd_sc_hd__dfrtp_1
X_4824_ _5102_/B _5404_/C VGND VGND VPWR VPWR _5322_/C sky130_fd_sc_hd__nor2_4
XFILLER_138_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7543_ _7559_/CLK _7543_/D fanout613/X VGND VGND VPWR VPWR _7543_/Q sky130_fd_sc_hd__dfrtp_1
X_4755_ _5017_/A _5131_/A _5000_/C VGND VGND VPWR VPWR _5313_/C sky130_fd_sc_hd__and3_4
XFILLER_193_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3706_ _3714_/A hold74/A _5666_/B VGND VGND VPWR VPWR _3706_/X sky130_fd_sc_hd__and3_1
X_7474_ _7614_/CLK _7474_/D fanout605/X VGND VGND VPWR VPWR _7474_/Q sky130_fd_sc_hd__dfstp_2
X_4686_ _4747_/B _5490_/C _5196_/A _5595_/B VGND VGND VPWR VPWR _4735_/C sky130_fd_sc_hd__nand4_1
XFILLER_162_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6425_ _7120_/Q _6359_/B _6170_/C _6424_/X VGND VGND VPWR VPWR _6425_/X sky130_fd_sc_hd__a31o_1
XFILLER_147_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3637_ _7440_/Q _5840_/A _3553_/X _3525_/X _7400_/Q VGND VGND VPWR VPWR _3637_/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_146_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6356_ _7062_/Q _6359_/B _6432_/A3 _6130_/X _7127_/Q VGND VGND VPWR VPWR _6356_/X
+ sky130_fd_sc_hd__a32o_1
X_3568_ _3714_/A hold53/X _3568_/C VGND VGND VPWR VPWR _6002_/B sky130_fd_sc_hd__and3_4
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5307_ _5604_/B1 _4991_/Y _5285_/X _5287_/X _5306_/X VGND VGND VPWR VPWR _5310_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_115_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6287_ _7368_/Q _6082_/B _6141_/X _6160_/X _7376_/Q VGND VGND VPWR VPWR _6287_/X
+ sky130_fd_sc_hd__a32o_2
X_3499_ hold133/X hold68/X _4229_/S VGND VGND VPWR VPWR _3513_/D sky130_fd_sc_hd__mux2_8
XFILLER_124_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5238_ _5061_/A _4951_/A _5089_/A _4933_/B VGND VGND VPWR VPWR _5263_/A sky130_fd_sc_hd__a31o_1
XFILLER_69_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5169_ _4681_/Y _5165_/X _5167_/X _5168_/X VGND VGND VPWR VPWR _5169_/X sky130_fd_sc_hd__o211a_1
XFILLER_84_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold6 hold6/A VGND VGND VPWR VPWR hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_59_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4540_ hold274/X _6866_/A1 _4540_/S VGND VGND VPWR VPWR _4540_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire370 _5548_/Y VGND VGND VPWR VPWR _5591_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_7_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4471_ hold395/X _5761_/A1 _4474_/S VGND VGND VPWR VPWR _4471_/X sky130_fd_sc_hd__mux2_1
Xhold406 _4305_/X VGND VGND VPWR VPWR _7020_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold417 hold417/A VGND VGND VPWR VPWR hold417/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold428 hold428/A VGND VGND VPWR VPWR hold428/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 _4555_/X VGND VGND VPWR VPWR _7235_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6210_ _7397_/Q _6166_/B _6146_/C _6124_/X _7405_/Q VGND VGND VPWR VPWR _6210_/X
+ sky130_fd_sc_hd__a32o_1
X_3422_ _7293_/Q VGND VGND VPWR VPWR _3422_/Y sky130_fd_sc_hd__clkinv_2
X_7190_ _7207_/CLK _7190_/D fanout633/X VGND VGND VPWR VPWR _7190_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6141_ _7623_/Q _6151_/B _6392_/B _7624_/Q VGND VGND VPWR VPWR _6141_/X sky130_fd_sc_hd__and4bb_4
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6072_ _7139_/Q _6109_/B _7624_/Q _6071_/Y VGND VGND VPWR VPWR _7624_/D sky130_fd_sc_hd__o31a_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1106 hold1451/X VGND VGND VPWR VPWR _5718_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1117 _5651_/X VGND VGND VPWR VPWR _7272_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1128 _4521_/X VGND VGND VPWR VPWR _7207_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5023_ _4629_/Y _4657_/Y _4750_/Y _5022_/X VGND VGND VPWR VPWR _5024_/B sky130_fd_sc_hd__o31ai_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1139 hold1440/X VGND VGND VPWR VPWR _5724_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6974_ _7291_/CLK _6974_/D fanout596/X VGND VGND VPWR VPWR _6974_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5925_ _6042_/A1 _5925_/A1 hold76/A VGND VGND VPWR VPWR _5925_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5856_ hold50/X hold180/X _5857_/S VGND VGND VPWR VPWR _5856_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4807_ _4943_/A _5318_/B _4806_/X VGND VGND VPWR VPWR _4808_/B sky130_fd_sc_hd__a21oi_1
XFILLER_186_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5787_ hold428/X _6003_/A1 _5794_/S VGND VGND VPWR VPWR _5787_/X sky130_fd_sc_hd__mux2_1
X_7526_ _7602_/CLK _7526_/D fanout615/X VGND VGND VPWR VPWR _7526_/Q sky130_fd_sc_hd__dfrtp_4
X_4738_ _4738_/A _4738_/B _5476_/A _4740_/D VGND VGND VPWR VPWR _4739_/B sky130_fd_sc_hd__nand4_1
XFILLER_147_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7457_ _7569_/CLK _7457_/D fanout614/X VGND VGND VPWR VPWR _7457_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_162_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4669_ _4747_/B _5364_/B VGND VGND VPWR VPWR _4669_/Y sky130_fd_sc_hd__nand2_1
XFILLER_174_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6408_ _7074_/Q _6158_/D _6334_/C _6407_/X VGND VGND VPWR VPWR _6408_/X sky130_fd_sc_hd__a31o_1
Xhold940 _5888_/X VGND VGND VPWR VPWR _7476_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7388_ _7430_/CLK _7388_/D fanout627/X VGND VGND VPWR VPWR _7388_/Q sky130_fd_sc_hd__dfrtp_1
Xhold951 _7615_/Q VGND VGND VPWR VPWR hold951/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold962 hold962/A VGND VGND VPWR VPWR hold962/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold973 _7411_/Q VGND VGND VPWR VPWR hold973/X sky130_fd_sc_hd__dlygate4sd3_1
X_6339_ _7081_/Q _6146_/X _6332_/X _6333_/X _6338_/X VGND VGND VPWR VPWR _6339_/X
+ sky130_fd_sc_hd__a2111o_1
Xhold984 hold984/A VGND VGND VPWR VPWR hold984/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 hold995/A VGND VGND VPWR VPWR hold995/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_532 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1640 _6974_/Q VGND VGND VPWR VPWR hold1640/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1651 hold21/A VGND VGND VPWR VPWR _4085_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3971_ _7426_/Q _5975_/B _4541_/A VGND VGND VPWR VPWR _3971_/X sky130_fd_sc_hd__and3_1
XFILLER_16_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5710_ _6043_/A1 hold271/X hold38/X VGND VGND VPWR VPWR _5710_/X sky130_fd_sc_hd__mux2_1
XFILLER_188_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6690_ _7071_/Q _6447_/X _6483_/X _7066_/Q _6689_/X VGND VGND VPWR VPWR _6700_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5641_ hold510/X _5673_/A1 _5642_/S VGND VGND VPWR VPWR _7264_/D sky130_fd_sc_hd__mux2_1
XFILLER_191_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5572_ _5572_/A _5572_/B _5572_/C _5572_/D VGND VGND VPWR VPWR _5573_/D sky130_fd_sc_hd__nor4_1
XFILLER_157_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7311_ _7616_/CLK _7311_/D fanout610/X VGND VGND VPWR VPWR _7311_/Q sky130_fd_sc_hd__dfrtp_1
X_4523_ _5768_/C hold70/X _6861_/C _5768_/B VGND VGND VPWR VPWR _4528_/S sky130_fd_sc_hd__nand4_4
XFILLER_144_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold203 _7459_/Q VGND VGND VPWR VPWR hold203/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold214 _7021_/Q VGND VGND VPWR VPWR hold214/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7242_ _7242_/CLK _7242_/D fanout616/X VGND VGND VPWR VPWR _7242_/Q sky130_fd_sc_hd__dfrtp_2
Xhold225 _6008_/X VGND VGND VPWR VPWR _7583_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 hold236/A VGND VGND VPWR VPWR hold236/X sky130_fd_sc_hd__dlygate4sd3_1
X_4454_ _6815_/A _4454_/B VGND VGND VPWR VPWR _4462_/S sky130_fd_sc_hd__nand2_4
Xhold247 hold247/A VGND VGND VPWR VPWR hold247/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 _7706_/A VGND VGND VPWR VPWR hold258/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold269 _7428_/Q VGND VGND VPWR VPWR hold269/X sky130_fd_sc_hd__dlygate4sd3_1
X_7173_ _7238_/CLK _7173_/D fanout602/X VGND VGND VPWR VPWR _7173_/Q sky130_fd_sc_hd__dfrtp_1
X_4385_ _5789_/A1 hold349/X _4387_/S VGND VGND VPWR VPWR _4385_/X sky130_fd_sc_hd__mux2_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6124_ _6151_/B _6157_/C _6126_/D VGND VGND VPWR VPWR _6124_/X sky130_fd_sc_hd__and3_4
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _6052_/Y _6053_/X _6064_/A VGND VGND VPWR VPWR _7619_/D sky130_fd_sc_hd__o21a_1
XFILLER_85_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _4990_/A _5014_/D VGND VGND VPWR VPWR _5094_/D sky130_fd_sc_hd__and2b_4
XFILLER_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_109 _6133_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6957_ _6957_/D _4193_/X VGND VGND VPWR VPWR _6957_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_121_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5908_ hold170/X _6043_/A1 _5911_/S VGND VGND VPWR VPWR _5908_/X sky130_fd_sc_hd__mux2_1
X_6888_ _6899_/A _6908_/B VGND VGND VPWR VPWR _6888_/X sky130_fd_sc_hd__and2_1
XFILLER_14_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5839_ hold910/X _6046_/A1 _5839_/S VGND VGND VPWR VPWR _5839_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7509_ _7597_/CLK _7509_/D fanout626/X VGND VGND VPWR VPWR _7509_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_108_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold770 _5960_/X VGND VGND VPWR VPWR _7540_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 _7267_/Q VGND VGND VPWR VPWR hold781/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold792 _7410_/Q VGND VGND VPWR VPWR hold792/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1470 _5778_/X VGND VGND VPWR VPWR _7378_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1481 _7662_/Q VGND VGND VPWR VPWR _6812_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1492 _4397_/X VGND VGND VPWR VPWR _7098_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_610 _6003_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_621 _3562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_632 _5021_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_643 _6127_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_654 _6153_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_665 _7438_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_676 _7189_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_687 input80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_698 _4116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput308 _4196_/X VGND VGND VPWR VPWR spi_sdi sky130_fd_sc_hd__buf_12
Xoutput319 hold594/X VGND VGND VPWR VPWR hold595/A sky130_fd_sc_hd__buf_12
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4170_ _7636_/Q _7288_/Q _7292_/Q VGND VGND VPWR VPWR _4170_/X sky130_fd_sc_hd__mux2_4
XFILLER_68_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6811_ _6810_/X _7661_/Q _6811_/S VGND VGND VPWR VPWR _6811_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6742_ _7191_/Q _6454_/X _6469_/X _7166_/Q _6741_/X VGND VGND VPWR VPWR _6742_/X
+ sky130_fd_sc_hd__a221o_2
X_3954_ input15/X _5669_/B _4529_/B _3953_/X VGND VGND VPWR VPWR _3954_/X sky130_fd_sc_hd__a31o_1
X_6673_ _7521_/Q _6645_/B _6536_/C _6457_/X _7577_/Q VGND VGND VPWR VPWR _6673_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_149_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3885_ _7452_/Q _6861_/A _6002_/A _3558_/X _7556_/Q VGND VGND VPWR VPWR _3901_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_176_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5624_ _5618_/Y _5580_/X _5623_/Y _5622_/X VGND VGND VPWR VPWR _5624_/X sky130_fd_sc_hd__a211o_1
XFILLER_176_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5555_ _5496_/X _5555_/B _5555_/C _5555_/D VGND VGND VPWR VPWR _5589_/B sky130_fd_sc_hd__and4b_1
X_4506_ _4506_/A0 _6862_/A1 _4510_/S VGND VGND VPWR VPWR _4506_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5486_ _5595_/B _5485_/X _5358_/X _5163_/Y VGND VGND VPWR VPWR _5486_/X sky130_fd_sc_hd__a211o_1
X_7225_ _7304_/CLK _7225_/D fanout620/X VGND VGND VPWR VPWR _7225_/Q sky130_fd_sc_hd__dfrtp_4
X_4437_ _5697_/A0 _4437_/A1 _4444_/S VGND VGND VPWR VPWR _7131_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout513 hold50/X VGND VGND VPWR VPWR _5991_/A1 sky130_fd_sc_hd__clkbuf_8
X_7156_ _7668_/CLK _7156_/D VGND VGND VPWR VPWR _7156_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout524 _5988_/A1 VGND VGND VPWR VPWR _6865_/A1 sky130_fd_sc_hd__buf_6
X_4368_ hold465/X _5673_/A1 _4369_/S VGND VGND VPWR VPWR _7074_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout546 _6003_/A1 VGND VGND VPWR VPWR _6012_/A0 sky130_fd_sc_hd__buf_6
XFILLER_98_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6107_ _7620_/Q _7142_/Q _6107_/C _7619_/Q VGND VGND VPWR VPWR _6107_/X sky130_fd_sc_hd__and4b_1
XFILLER_86_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout557 _7630_/Q VGND VGND VPWR VPWR _6485_/B sky130_fd_sc_hd__buf_4
Xfanout568 _7140_/Q VGND VGND VPWR VPWR _6811_/S sky130_fd_sc_hd__buf_6
XFILLER_100_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7087_ _7210_/CLK _7087_/D fanout621/X VGND VGND VPWR VPWR _7087_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout579 _5311_/C VGND VGND VPWR VPWR _5313_/B sky130_fd_sc_hd__buf_6
X_4299_ _4299_/A0 _6042_/A1 _4303_/S VGND VGND VPWR VPWR _4299_/X sky130_fd_sc_hd__mux2_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6038_ hold24/X _6038_/B _6038_/C VGND VGND VPWR VPWR _6046_/S sky130_fd_sc_hd__and3_4
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_64_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7590_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_41_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_79_csclk _7095_/CLK VGND VGND VPWR VPWR _7293_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_173_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_440 _6444_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_451 _6464_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_462 _6700_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_473 _7516_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_484 _7221_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_495 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3670_ _7439_/Q _5840_/A _5984_/B _3555_/X _7519_/Q VGND VGND VPWR VPWR _3670_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_185_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5340_ _5585_/A1 _4825_/Y _5018_/Y _5197_/Y _4976_/Y VGND VGND VPWR VPWR _5340_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5271_ _4953_/C _4949_/Y _4858_/A _4953_/D _5407_/D VGND VGND VPWR VPWR _5573_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_114_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7010_ _7312_/CLK _7010_/D _6891_/A VGND VGND VPWR VPWR _7010_/Q sky130_fd_sc_hd__dfrtp_1
X_4222_ hold455/X _5673_/A1 _4230_/S VGND VGND VPWR VPWR _6975_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4153_ _7303_/Q input81/X _4196_/B VGND VGND VPWR VPWR _4153_/X sky130_fd_sc_hd__mux2_2
XFILLER_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4084_ _4084_/A1 _3508_/S _4043_/Y _4083_/X VGND VGND VPWR VPWR _6926_/D sky130_fd_sc_hd__a31o_1
XFILLER_55_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4986_ _5017_/A _5017_/B _5131_/A VGND VGND VPWR VPWR _5452_/C sky130_fd_sc_hd__and3_2
X_3937_ _7523_/Q _5993_/A _5939_/B _3933_/X _3936_/X VGND VGND VPWR VPWR _3937_/X
+ sky130_fd_sc_hd__a311o_1
X_6725_ _6725_/A _6725_/B _6725_/C _6725_/D VGND VGND VPWR VPWR _6725_/Y sky130_fd_sc_hd__nor4_1
XFILLER_149_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6656_ _7464_/Q _6464_/X _6481_/X _7384_/Q _6655_/X VGND VGND VPWR VPWR _6659_/B
+ sky130_fd_sc_hd__a221o_1
X_3868_ _7604_/Q _5957_/B _6038_/B _3867_/X VGND VGND VPWR VPWR _3868_/X sky130_fd_sc_hd__a31o_1
XFILLER_127_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5607_ _5021_/B _5291_/C _5249_/C _5095_/X _5606_/X VGND VGND VPWR VPWR _5607_/X
+ sky130_fd_sc_hd__a311o_1
X_6587_ _7478_/Q _6791_/C _6720_/D _6791_/D VGND VGND VPWR VPWR _6587_/X sky130_fd_sc_hd__and4_1
X_3799_ _7217_/Q _5993_/A _4529_/B _3557_/X _7573_/Q VGND VGND VPWR VPWR _3799_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_191_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5538_ _5375_/A _5196_/A _5068_/C _5069_/X VGND VGND VPWR VPWR _5538_/X sky130_fd_sc_hd__a31o_1
XFILLER_192_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5469_ _5614_/C _4702_/X _4758_/X _5614_/A VGND VGND VPWR VPWR _5469_/X sky130_fd_sc_hd__o211a_1
XFILLER_133_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7208_ _7686_/CLK _7208_/D _6907_/A VGND VGND VPWR VPWR _7208_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_59_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7139_ _7680_/CLK _7139_/D _6886_/A VGND VGND VPWR VPWR _7139_/Q sky130_fd_sc_hd__dfstp_4
Xfanout387 _3550_/B VGND VGND VPWR VPWR _5628_/A sky130_fd_sc_hd__buf_8
Xfanout398 _3622_/X VGND VGND VPWR VPWR _4553_/B sky130_fd_sc_hd__buf_6
XFILLER_74_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput18 mask_rev_in[22] VGND VGND VPWR VPWR input18/X sky130_fd_sc_hd__clkbuf_1
Xinput29 mask_rev_in[3] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__clkbuf_1
XFILLER_182_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4840_ _4633_/Y _4777_/Y _4836_/Y _5014_/D VGND VGND VPWR VPWR _4853_/C sky130_fd_sc_hd__o22ai_2
XANTENNA_270 input71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_281 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_292 _7713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4771_ _4943_/A _5595_/A _5490_/B _5186_/C VGND VGND VPWR VPWR _5180_/C sky130_fd_sc_hd__nand4_1
XFILLER_193_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6510_ _6510_/A1 _6812_/S _6508_/X _6509_/X VGND VGND VPWR VPWR _7650_/D sky130_fd_sc_hd__a22o_1
X_3722_ _7382_/Q _5993_/B _4511_/C _3718_/X _3721_/X VGND VGND VPWR VPWR _3722_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_119_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7490_ _7580_/CLK _7490_/D fanout605/X VGND VGND VPWR VPWR _7490_/Q sky130_fd_sc_hd__dfstp_4
X_6441_ _6791_/C _6563_/C _6791_/D VGND VGND VPWR VPWR _6441_/X sky130_fd_sc_hd__and3_4
X_3653_ _7552_/Q _3514_/X _3646_/X _3649_/X _3652_/X VGND VGND VPWR VPWR _3654_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_173_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6372_ _7226_/Q _6166_/B _6427_/A3 _6170_/C _7048_/Q VGND VGND VPWR VPWR _6372_/X
+ sky130_fd_sc_hd__a32o_1
X_3584_ _3905_/B _4340_/A _5680_/B VGND VGND VPWR VPWR _3584_/X sky130_fd_sc_hd__and3_2
XFILLER_127_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5323_ _5196_/A _5322_/A _5476_/C _5327_/B VGND VGND VPWR VPWR _5323_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_142_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5254_ _4871_/X _4889_/Y _5015_/Y _5088_/Y _5392_/C VGND VGND VPWR VPWR _5254_/X
+ sky130_fd_sc_hd__o221a_1
X_4205_ input58/X hold14/X hold42/X VGND VGND VPWR VPWR hold43/A sky130_fd_sc_hd__mux2_8
X_5185_ _4597_/Y _4811_/Y _4821_/Y _4817_/Y _4674_/Y VGND VGND VPWR VPWR _5555_/D
+ sky130_fd_sc_hd__o32a_1
Xclkbuf_3_6_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR _7352_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4136_ _6970_/Q _4133_/X _4210_/C VGND VGND VPWR VPWR _6970_/D sky130_fd_sc_hd__a21o_1
XFILLER_83_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4067_ _4067_/A hold33/A _4067_/C VGND VGND VPWR VPWR _4069_/A sky130_fd_sc_hd__and3_1
XFILLER_71_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4969_ _5131_/A _4969_/B _5040_/A _5452_/B VGND VGND VPWR VPWR _4969_/Y sky130_fd_sc_hd__nand4_1
XFILLER_184_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6708_ _7251_/Q _6460_/X _6705_/X _6707_/X VGND VGND VPWR VPWR _6709_/C sky130_fd_sc_hd__a211o_1
XFILLER_177_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7688_ _7688_/A VGND VGND VPWR VPWR _7688_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_177_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6639_ _7440_/Q _6097_/X _6445_/C _6474_/A _7344_/Q VGND VGND VPWR VPWR _6639_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_165_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6990_ _7421_/CLK _6990_/D fanout630/X VGND VGND VPWR VPWR _7698_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_65_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5941_ hold307/X _6031_/A0 _5947_/S VGND VGND VPWR VPWR _5941_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5872_ hold237/X _6866_/A1 _5875_/S VGND VGND VPWR VPWR _5872_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7611_ _7611_/CLK _7611_/D fanout624/X VGND VGND VPWR VPWR _7611_/Q sky130_fd_sc_hd__dfstp_1
X_4823_ _4822_/A _5146_/B VGND VGND VPWR VPWR _4823_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_178_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7542_ _7606_/CLK hold3/X fanout615/X VGND VGND VPWR VPWR _7542_/Q sky130_fd_sc_hd__dfrtp_1
X_4754_ _5017_/B _5025_/B VGND VGND VPWR VPWR _5131_/B sky130_fd_sc_hd__nor2_4
X_3705_ _3714_/A hold74/A _4505_/B VGND VGND VPWR VPWR _4388_/A sky130_fd_sc_hd__and3_2
XFILLER_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7473_ _7547_/CLK _7473_/D fanout607/X VGND VGND VPWR VPWR _7473_/Q sky130_fd_sc_hd__dfrtp_4
X_4685_ _4747_/B _5595_/B VGND VGND VPWR VPWR _4685_/Y sky130_fd_sc_hd__nand2_2
XFILLER_119_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3636_ _7544_/Q _3530_/X _3563_/X _7480_/Q _3635_/X VGND VGND VPWR VPWR _3654_/A
+ sky130_fd_sc_hd__a221o_1
X_6424_ _7255_/Q _6082_/B _6416_/C _6166_/C VGND VGND VPWR VPWR _6424_/X sky130_fd_sc_hd__o211a_1
XFILLER_161_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6355_ _7220_/Q _6428_/B1 _6352_/X _6354_/X VGND VGND VPWR VPWR _6355_/X sky130_fd_sc_hd__a211o_1
XFILLER_115_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3567_ _5768_/C _6020_/A _5768_/B VGND VGND VPWR VPWR _3567_/X sky130_fd_sc_hd__and3_4
X_5306_ _5604_/B1 _4998_/Y _5285_/X _5305_/X VGND VGND VPWR VPWR _5306_/X sky130_fd_sc_hd__o31a_1
X_6286_ _7480_/Q _6309_/B _6286_/C VGND VGND VPWR VPWR _6286_/X sky130_fd_sc_hd__and3_1
XFILLER_170_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3498_ hold94/X hold132/X _3508_/S VGND VGND VPWR VPWR _3498_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5237_ _5322_/A _5512_/B _5452_/B _4975_/Y VGND VGND VPWR VPWR _5327_/A sky130_fd_sc_hd__a31o_1
X_5168_ _4619_/Y _4660_/C _4681_/Y _4912_/Y _4669_/Y VGND VGND VPWR VPWR _5168_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_130_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4119_ hold1638/X _4119_/B VGND VGND VPWR VPWR _6961_/D sky130_fd_sc_hd__nand2b_1
XFILLER_29_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5099_ _4570_/Y _4821_/Y _5097_/Y VGND VGND VPWR VPWR _5099_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_56_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold7 hold7/A VGND VGND VPWR VPWR hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire360 _5696_/Y VGND VGND VPWR VPWR _5703_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_116_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4470_ _4470_/A0 _6012_/A0 _4474_/S VGND VGND VPWR VPWR _4470_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold407 _7566_/Q VGND VGND VPWR VPWR hold407/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold418 _7107_/Q VGND VGND VPWR VPWR hold418/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold429 _7598_/Q VGND VGND VPWR VPWR hold429/X sky130_fd_sc_hd__dlygate4sd3_1
X_3421_ _7142_/Q VGND VGND VPWR VPWR _3421_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6140_ _7450_/Q _6132_/X _6134_/X _6131_/X _6139_/X VGND VGND VPWR VPWR _6140_/X
+ sky130_fd_sc_hd__a2111o_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _6231_/D _6166_/B _6109_/B VGND VGND VPWR VPWR _6071_/Y sky130_fd_sc_hd__o21ai_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1107 _7300_/Q VGND VGND VPWR VPWR _5690_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _4825_/Y _5018_/Y _5021_/Y _5019_/X VGND VGND VPWR VPWR _5022_/X sky130_fd_sc_hd__o211a_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1118 _7274_/Q VGND VGND VPWR VPWR _5653_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1129 _7237_/Q VGND VGND VPWR VPWR _4557_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6973_ _7291_/CLK _6973_/D fanout596/X VGND VGND VPWR VPWR _6973_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_81_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5924_ _6041_/A1 hold800/X hold76/A VGND VGND VPWR VPWR _5924_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5855_ _5999_/A1 hold945/X _5857_/S VGND VGND VPWR VPWR _5855_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4806_ _5375_/A _5186_/C _5364_/B _4946_/A VGND VGND VPWR VPWR _4806_/X sky130_fd_sc_hd__and4_1
XFILLER_166_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5786_ _5840_/A _5786_/B _6029_/B VGND VGND VPWR VPWR _5794_/S sky130_fd_sc_hd__and3_4
XFILLER_119_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7525_ _7603_/CLK hold88/X fanout606/X VGND VGND VPWR VPWR hold87/A sky130_fd_sc_hd__dfrtp_4
X_4737_ _4737_/A _4737_/B VGND VGND VPWR VPWR _4739_/A sky130_fd_sc_hd__nor2_1
XFILLER_147_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4668_ _4747_/B _4684_/A _4668_/C VGND VGND VPWR VPWR _4743_/C sky130_fd_sc_hd__and3_2
X_7456_ _7616_/CLK _7456_/D fanout610/X VGND VGND VPWR VPWR _7456_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3619_ _6917_/Q _4192_/B VGND VGND VPWR VPWR _3967_/S sky130_fd_sc_hd__nand2_4
X_6407_ _7242_/Q _6158_/D _6407_/A3 _6145_/X _7685_/Q VGND VGND VPWR VPWR _6407_/X
+ sky130_fd_sc_hd__a32o_1
Xhold930 _5738_/X VGND VGND VPWR VPWR _7343_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4599_ _5015_/C _5017_/B VGND VGND VPWR VPWR _4599_/Y sky130_fd_sc_hd__nand2_8
XFILLER_190_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold941 hold941/A VGND VGND VPWR VPWR hold941/X sky130_fd_sc_hd__dlygate4sd3_1
X_7387_ _7515_/CLK _7387_/D fanout621/X VGND VGND VPWR VPWR _7387_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_162_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold952 _6044_/X VGND VGND VPWR VPWR _7615_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold963 _7535_/Q VGND VGND VPWR VPWR hold963/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6338_ _7091_/Q _6136_/X _6334_/X _6335_/X _6337_/X VGND VGND VPWR VPWR _6338_/X
+ sky130_fd_sc_hd__a2111o_1
Xhold974 _5815_/X VGND VGND VPWR VPWR _7411_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 _7254_/Q VGND VGND VPWR VPWR hold985/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold996 hold996/A VGND VGND VPWR VPWR hold996/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6269_ _7447_/Q _6082_/B _6416_/C _6166_/C VGND VGND VPWR VPWR _6269_/X sky130_fd_sc_hd__o211a_1
XFILLER_130_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1630 _7141_/Q VGND VGND VPWR VPWR _6103_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1641 _6954_/Q VGND VGND VPWR VPWR hold1641/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1652 _6927_/Q VGND VGND VPWR VPWR _4079_/B1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3970_ _3970_/A VGND VGND VPWR VPWR _3970_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5640_ _5640_/A0 _6864_/A1 _5642_/S VGND VGND VPWR VPWR _5640_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5571_ _5021_/B _5404_/B _5571_/B1 _5074_/A _5278_/X VGND VGND VPWR VPWR _5572_/D
+ sky130_fd_sc_hd__a221o_1
X_7310_ _7616_/CLK _7310_/D fanout610/X VGND VGND VPWR VPWR _7310_/Q sky130_fd_sc_hd__dfrtp_1
X_4522_ hold195/X _6866_/A1 _4522_/S VGND VGND VPWR VPWR _4522_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold204 _5869_/X VGND VGND VPWR VPWR _7459_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold215 _4306_/X VGND VGND VPWR VPWR _7021_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7241_ _7686_/CLK _7241_/D fanout600/X VGND VGND VPWR VPWR _7241_/Q sky130_fd_sc_hd__dfstp_1
X_4453_ _3618_/Y _4453_/A1 _4453_/S VGND VGND VPWR VPWR _7150_/D sky130_fd_sc_hd__mux2_1
Xhold226 _7422_/Q VGND VGND VPWR VPWR hold226/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 _7462_/Q VGND VGND VPWR VPWR hold237/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 hold248/A VGND VGND VPWR VPWR hold248/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold259 _4298_/X VGND VGND VPWR VPWR _7014_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7172_ _7242_/CLK _7172_/D fanout616/X VGND VGND VPWR VPWR _7172_/Q sky130_fd_sc_hd__dfstp_2
X_4384_ _5761_/A1 hold490/X _4387_/S VGND VGND VPWR VPWR _4384_/X sky130_fd_sc_hd__mux2_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6123_ _7410_/Q _6231_/B _6416_/B _6416_/C _6122_/X VGND VGND VPWR VPWR _6123_/X
+ sky130_fd_sc_hd__a41o_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6054_ _7142_/Q _6811_/S _6109_/B _7619_/Q _4140_/Y VGND VGND VPWR VPWR _6063_/D
+ sky130_fd_sc_hd__o311a_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5005_ _5195_/B _5476_/B _5005_/C _5311_/A VGND VGND VPWR VPWR _5466_/B sky130_fd_sc_hd__nand4_2
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6956_ _6956_/D _4193_/X VGND VGND VPWR VPWR _6956_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_54_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5907_ hold40/X hold9/X _5911_/S VGND VGND VPWR VPWR hold41/A sky130_fd_sc_hd__mux2_1
X_6887_ _6899_/A _6908_/B VGND VGND VPWR VPWR _6887_/X sky130_fd_sc_hd__and2_1
XFILLER_22_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5838_ hold680/X _5991_/A1 _5839_/S VGND VGND VPWR VPWR _5838_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5769_ _6003_/A1 hold422/X _5776_/S VGND VGND VPWR VPWR _5769_/X sky130_fd_sc_hd__mux2_1
X_7508_ _7541_/CLK _7508_/D fanout605/X VGND VGND VPWR VPWR _7508_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_108_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7439_ _7445_/CLK _7439_/D fanout631/X VGND VGND VPWR VPWR _7439_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_123_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold760 _5909_/X VGND VGND VPWR VPWR _7495_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 _7596_/Q VGND VGND VPWR VPWR hold771/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold782 _5645_/X VGND VGND VPWR VPWR _7267_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap490 _5093_/C VGND VGND VPWR VPWR _5523_/A3 sky130_fd_sc_hd__clkbuf_2
XFILLER_122_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold793 _5814_/X VGND VGND VPWR VPWR _7410_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1460 _7638_/Q VGND VGND VPWR VPWR _6206_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1471 _7426_/Q VGND VGND VPWR VPWR hold420/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1482 _6812_/X VGND VGND VPWR VPWR _7662_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_600 _5669_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1493 _7394_/Q VGND VGND VPWR VPWR hold1493/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_611 _6003_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_622 _5666_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_633 _5021_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_644 _6137_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_655 _6153_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_666 _7121_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_677 _7382_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_688 input80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_699 _4116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput309 _4190_/X VGND VGND VPWR VPWR spimemio_flash_io0_di sky130_fd_sc_hd__buf_12
XFILLER_181_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6810_ wire372/X _6809_/Y _7040_/Q _6759_/D VGND VGND VPWR VPWR _6810_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6741_ _7083_/Q _6645_/B _6562_/C _6458_/X _7088_/Q VGND VGND VPWR VPWR _6741_/X
+ sky130_fd_sc_hd__a32o_1
X_3953_ input12/X _5669_/B _4535_/B _5650_/A _7273_/Q VGND VGND VPWR VPWR _3953_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_149_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3884_ _7231_/Q _4547_/A _4553_/B _3584_/X _7580_/Q VGND VGND VPWR VPWR _3901_/A
+ sky130_fd_sc_hd__a32o_1
X_6672_ _7481_/Q _6791_/C _6720_/D _6791_/D VGND VGND VPWR VPWR _6672_/X sky130_fd_sc_hd__and4_1
XFILLER_31_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5623_ _5549_/A _5594_/Y _5597_/X _5589_/Y VGND VGND VPWR VPWR _5623_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_164_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5554_ _4805_/Y _4953_/C _5553_/Y VGND VGND VPWR VPWR _5554_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_129_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4505_ _4547_/A _4505_/B _5686_/D VGND VGND VPWR VPWR _4510_/S sky130_fd_sc_hd__and3_2
X_5485_ _5476_/A _5375_/C _4738_/A _5490_/C VGND VGND VPWR VPWR _5485_/X sky130_fd_sc_hd__o211a_1
XFILLER_160_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4436_ hold56/X _5680_/C VGND VGND VPWR VPWR _4444_/S sky130_fd_sc_hd__nand2_4
XFILLER_104_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7224_ _7304_/CLK _7224_/D fanout619/X VGND VGND VPWR VPWR _7224_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_160_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout503 _4702_/X VGND VGND VPWR VPWR _5311_/A sky130_fd_sc_hd__buf_8
XFILLER_160_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout514 hold49/X VGND VGND VPWR VPWR hold50/A sky130_fd_sc_hd__buf_8
X_4367_ _4367_/A0 _6864_/A1 _4369_/S VGND VGND VPWR VPWR _7073_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7155_ _7668_/CLK _7155_/D VGND VGND VPWR VPWR _7155_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout525 _5988_/A1 VGND VGND VPWR VPWR _6042_/A1 sky130_fd_sc_hd__buf_6
Xfanout547 hold44/A VGND VGND VPWR VPWR _6003_/A1 sky130_fd_sc_hd__buf_8
XFILLER_113_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6106_ _6106_/A0 _4129_/X _6108_/S VGND VGND VPWR VPWR _7635_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout558 _6131_/B VGND VGND VPWR VPWR _6309_/B sky130_fd_sc_hd__buf_6
XFILLER_98_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7086_ _7254_/CLK _7086_/D fanout617/X VGND VGND VPWR VPWR _7086_/Q sky130_fd_sc_hd__dfrtp_2
X_4298_ hold258/X _5789_/A1 _4303_/S VGND VGND VPWR VPWR _4298_/X sky130_fd_sc_hd__mux2_1
Xfanout569 _7140_/Q VGND VGND VPWR VPWR _6686_/S sky130_fd_sc_hd__buf_4
XFILLER_86_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6037_ hold102/X hold282/X _6037_/S VGND VGND VPWR VPWR _6037_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6939_ _4183_/A1 _6939_/D _6894_/X VGND VGND VPWR VPWR _6939_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_csclk _4172_/X VGND VGND VPWR VPWR clkbuf_0_csclk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_157_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold590 _5739_/X VGND VGND VPWR VPWR _7344_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1290 _5933_/X VGND VGND VPWR VPWR _7516_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_430 _6192_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_441 _6444_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_452 _6465_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_463 _6700_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_474 _7516_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_485 _7570_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_496 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5270_ _5407_/A _5429_/D _4704_/A _4949_/Y VGND VGND VPWR VPWR _5270_/X sky130_fd_sc_hd__o31a_1
XFILLER_142_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4221_ hold7/X hold11/X _4221_/S VGND VGND VPWR VPWR hold12/A sky130_fd_sc_hd__mux2_1
XFILLER_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4152_ _7301_/Q input78/X _4196_/B VGND VGND VPWR VPWR _4152_/X sky130_fd_sc_hd__mux2_2
XFILLER_110_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4083_ _4085_/B _4062_/Y _4082_/X _3500_/X VGND VGND VPWR VPWR _4083_/X sky130_fd_sc_hd__a31o_1
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4985_ _5313_/C _4985_/B VGND VGND VPWR VPWR _4985_/Y sky130_fd_sc_hd__nand2_1
XFILLER_189_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6724_ _7057_/Q _6474_/C _6720_/X _6721_/X _6723_/X VGND VGND VPWR VPWR _6725_/D
+ sky130_fd_sc_hd__a2111o_1
X_3936_ _7170_/Q _4475_/A _5678_/B _3935_/X VGND VGND VPWR VPWR _3936_/X sky130_fd_sc_hd__a31o_1
Xclkbuf_3_2_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_2_0_csclk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_176_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6655_ _7496_/Q _6694_/B _6720_/D _6452_/X _7584_/Q VGND VGND VPWR VPWR _6655_/X
+ sky130_fd_sc_hd__a32o_1
X_3867_ _7283_/Q _5993_/B _6038_/B _7492_/Q _3519_/X VGND VGND VPWR VPWR _3867_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_137_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5606_ _4948_/B _5146_/B _5291_/C _5249_/C _5423_/X VGND VGND VPWR VPWR _5606_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_192_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6586_ _6585_/X _6610_/A1 _6611_/S VGND VGND VPWR VPWR _6586_/X sky130_fd_sc_hd__mux2_1
X_3798_ _7222_/Q _5984_/A _4535_/B _3797_/X VGND VGND VPWR VPWR _3798_/X sky130_fd_sc_hd__a31o_1
XFILLER_118_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5537_ _5537_/A _5537_/B _5537_/C VGND VGND VPWR VPWR _5583_/C sky130_fd_sc_hd__and3_1
XFILLER_145_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5468_ _5537_/A _5537_/B _5468_/C VGND VGND VPWR VPWR _5473_/A sky130_fd_sc_hd__and3_1
XFILLER_172_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7207_ _7207_/CLK _7207_/D fanout616/X VGND VGND VPWR VPWR _7207_/Q sky130_fd_sc_hd__dfrtp_4
X_4419_ _6012_/A0 _4419_/A1 _4423_/S VGND VGND VPWR VPWR _4419_/X sky130_fd_sc_hd__mux2_1
X_5399_ _5382_/X _5399_/B _5399_/C _5399_/D VGND VGND VPWR VPWR _5403_/C sky130_fd_sc_hd__and4b_1
XFILLER_99_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7138_ _7614_/CLK _7138_/D fanout604/X VGND VGND VPWR VPWR _7138_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_86_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout388 _5840_/A VGND VGND VPWR VPWR _4541_/A sky130_fd_sc_hd__buf_6
Xfanout399 _3551_/Y VGND VGND VPWR VPWR _6002_/A sky130_fd_sc_hd__buf_12
XFILLER_47_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7069_ _7212_/CLK _7069_/D fanout619/X VGND VGND VPWR VPWR _7069_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_74_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput19 mask_rev_in[23] VGND VGND VPWR VPWR input19/X sky130_fd_sc_hd__clkbuf_2
XFILLER_168_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_260 input61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_271 input78/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_282 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_293 input95/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4770_ _4770_/A _5490_/B _5186_/C _5181_/C VGND VGND VPWR VPWR _4775_/B sky130_fd_sc_hd__nand4_1
XFILLER_14_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3721_ _7213_/Q _4505_/B _4511_/C _3720_/X VGND VGND VPWR VPWR _3721_/X sky130_fd_sc_hd__a31o_1
XFILLER_158_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6440_ _7629_/Q _7628_/Q VGND VGND VPWR VPWR _6562_/B sky130_fd_sc_hd__nor2_2
X_3652_ _7432_/Q _3556_/X _4257_/S input50/X _3651_/X VGND VGND VPWR VPWR _3652_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3583_ _3713_/A _5661_/A _4481_/A VGND VGND VPWR VPWR _3583_/X sky130_fd_sc_hd__and3_4
X_6371_ _7166_/Q _6166_/B _6145_/C _6428_/A2 _7211_/Q VGND VGND VPWR VPWR _6371_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_127_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5322_ _5322_/A _5512_/B _5322_/C VGND VGND VPWR VPWR _5327_/B sky130_fd_sc_hd__and3_1
X_5253_ _4859_/Y _4949_/Y _5018_/Y _4873_/Y _4889_/Y VGND VGND VPWR VPWR _5392_/C
+ sky130_fd_sc_hd__o32a_1
XFILLER_142_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4204_ _5678_/C _6002_/A _5686_/D VGND VGND VPWR VPWR _4208_/S sky130_fd_sc_hd__and3_1
X_5184_ _4813_/X _5184_/B _5184_/C VGND VGND VPWR VPWR _5188_/A sky130_fd_sc_hd__and3b_1
XFILLER_68_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4135_ _6971_/Q _4133_/X _4210_/A VGND VGND VPWR VPWR _6971_/D sky130_fd_sc_hd__a21o_1
XFILLER_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_63_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7614_/CLK sky130_fd_sc_hd__clkbuf_16
X_4066_ _6929_/Q _4085_/B _4064_/X _3478_/X VGND VGND VPWR VPWR _4067_/C sky130_fd_sc_hd__a31o_1
XFILLER_56_559 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_78_csclk _7095_/CLK VGND VGND VPWR VPWR _7291_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_52_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4968_ _4968_/A _4968_/B _4968_/C VGND VGND VPWR VPWR _4971_/A sky130_fd_sc_hd__nor3_1
X_6707_ _7051_/Q _6474_/B _6482_/X _7111_/Q _6706_/X VGND VGND VPWR VPWR _6707_/X
+ sky130_fd_sc_hd__a221o_1
X_3919_ input44/X _6002_/B _5666_/B _3714_/X _7220_/Q VGND VGND VPWR VPWR _3919_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_137_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4899_ _4901_/B _5021_/B _4899_/C _4950_/C VGND VGND VPWR VPWR _4900_/D sky130_fd_sc_hd__nand4_1
X_6638_ _7600_/Q _6791_/B _6720_/C _6645_/C VGND VGND VPWR VPWR _6638_/X sky130_fd_sc_hd__and4_1
XFILLER_106_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6569_ _7413_/Q _6450_/X _6483_/X _7389_/Q _6568_/X VGND VGND VPWR VPWR _6569_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_16_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7192_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_133_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire575 _5191_/C VGND VGND VPWR VPWR _5137_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_109_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5940_ hold399/X _6039_/A1 _5947_/S VGND VGND VPWR VPWR _7522_/D sky130_fd_sc_hd__mux2_1
XFILLER_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5871_ _5871_/A0 hold9/X _5875_/S VGND VGND VPWR VPWR hold13/A sky130_fd_sc_hd__mux2_1
XFILLER_179_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7610_ _7614_/CLK _7610_/D fanout606/X VGND VGND VPWR VPWR _7610_/Q sky130_fd_sc_hd__dfstp_2
X_4822_ _4822_/A _5404_/C VGND VGND VPWR VPWR _5512_/C sky130_fd_sc_hd__nor2_2
XFILLER_33_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7541_ _7541_/CLK hold47/X fanout605/X VGND VGND VPWR VPWR hold46/A sky130_fd_sc_hd__dfrtp_4
X_4753_ _4990_/A _5014_/D VGND VGND VPWR VPWR _5131_/A sky130_fd_sc_hd__nor2_8
XFILLER_147_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3704_ _4547_/A _5661_/B _5659_/C VGND VGND VPWR VPWR _3704_/X sky130_fd_sc_hd__and3_2
X_7472_ _7616_/CLK _7472_/D fanout610/X VGND VGND VPWR VPWR _7472_/Q sky130_fd_sc_hd__dfrtp_1
X_4684_ _4684_/A _5015_/C _4706_/D VGND VGND VPWR VPWR _5595_/B sky130_fd_sc_hd__and3_4
X_6423_ _6416_/X _6418_/X _6422_/X _6082_/B VGND VGND VPWR VPWR _6423_/X sky130_fd_sc_hd__o31a_2
X_3635_ _7456_/Q _5903_/A _6002_/A _3580_/X _7616_/Q VGND VGND VPWR VPWR _3635_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_147_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6354_ _7092_/Q _6428_/A2 _6427_/B1 _7112_/Q _6353_/X VGND VGND VPWR VPWR _6354_/X
+ sky130_fd_sc_hd__a221o_1
X_3566_ _5661_/A _3717_/B _4511_/C VGND VGND VPWR VPWR _5741_/A sky130_fd_sc_hd__and3_4
XFILLER_115_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5305_ _5604_/B1 _5001_/Y _5285_/X _5288_/X _5304_/Y VGND VGND VPWR VPWR _5305_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_161_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3497_ hold34/X hold53/X hold61/X hold73/A VGND VGND VPWR VPWR hold62/A sky130_fd_sc_hd__and4bb_1
X_6285_ _7560_/Q _6309_/B _6432_/A3 _6145_/X _7464_/Q VGND VGND VPWR VPWR _6285_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_170_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5236_ _4800_/Y _4816_/Y _4821_/Y _5080_/Y VGND VGND VPWR VPWR _5236_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_69_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5167_ _4685_/Y _5165_/X _5166_/X _5164_/X VGND VGND VPWR VPWR _5167_/X sky130_fd_sc_hd__o211a_1
XFILLER_29_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4118_ _4117_/X _4118_/B VGND VGND VPWR VPWR _4119_/B sky130_fd_sc_hd__nand2b_1
XFILLER_68_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5098_ _5071_/C _5137_/C wire572/X _5311_/C VGND VGND VPWR VPWR _5098_/X sky130_fd_sc_hd__a31o_1
X_4049_ _6915_/Q _4049_/B VGND VGND VPWR VPWR _4049_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold8 hold8/A VGND VGND VPWR VPWR hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_87_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire350 _3617_/Y VGND VGND VPWR VPWR _3618_/C sky130_fd_sc_hd__clkbuf_1
Xwire361 _5696_/Y VGND VGND VPWR VPWR _5704_/S sky130_fd_sc_hd__clkbuf_2
Xwire372 _6800_/Y VGND VGND VPWR VPWR wire372/X sky130_fd_sc_hd__clkbuf_1
XFILLER_156_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold408 _5989_/X VGND VGND VPWR VPWR _7566_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold419 _4408_/X VGND VGND VPWR VPWR _7107_/D sky130_fd_sc_hd__dlygate4sd3_1
Xwire394 _4469_/B VGND VGND VPWR VPWR _4541_/B sky130_fd_sc_hd__clkbuf_2
X_3420_ _5096_/A VGND VGND VPWR VPWR _4794_/D sky130_fd_sc_hd__inv_2
XFILLER_109_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6070_ _7624_/Q _7623_/Q VGND VGND VPWR VPWR _6157_/C sky130_fd_sc_hd__and2_4
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1108 _5690_/X VGND VGND VPWR VPWR _7300_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5021_ _5021_/A _5021_/B VGND VGND VPWR VPWR _5021_/Y sky130_fd_sc_hd__nand2_1
Xhold1119 _5653_/X VGND VGND VPWR VPWR _7274_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6972_ _7291_/CLK _6972_/D fanout596/X VGND VGND VPWR VPWR _6972_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_53_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5923_ _6031_/A0 hold149/X hold76/A VGND VGND VPWR VPWR _5923_/X sky130_fd_sc_hd__mux2_1
X_5854_ hold19/X _5854_/A1 _5857_/S VGND VGND VPWR VPWR hold20/A sky130_fd_sc_hd__mux2_1
XFILLER_110_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4805_ _5071_/B _5071_/C VGND VGND VPWR VPWR _4805_/Y sky130_fd_sc_hd__nand2_1
XFILLER_167_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5785_ _6046_/A1 hold855/X _5785_/S VGND VGND VPWR VPWR _5785_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7524_ _7545_/CLK _7524_/D fanout613/X VGND VGND VPWR VPWR _7524_/Q sky130_fd_sc_hd__dfrtp_4
X_4736_ _4738_/A _4738_/B _5297_/A _5595_/B VGND VGND VPWR VPWR _4737_/A sky130_fd_sc_hd__and4_1
XFILLER_175_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7455_ _7584_/CLK _7455_/D fanout613/X VGND VGND VPWR VPWR _7455_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4667_ _5025_/B _4706_/D _4684_/A VGND VGND VPWR VPWR _5364_/B sky130_fd_sc_hd__and3_2
XFILLER_147_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6406_ _7094_/Q _6136_/X _6144_/X _7222_/Q _6401_/X VGND VGND VPWR VPWR _6406_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_190_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3618_ _3592_/X _3618_/B _3618_/C VGND VGND VPWR VPWR _3618_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_134_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold920 _7069_/Q VGND VGND VPWR VPWR hold920/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold931 _7003_/Q VGND VGND VPWR VPWR hold931/X sky130_fd_sc_hd__dlygate4sd3_1
X_7386_ _7518_/CLK _7386_/D fanout625/X VGND VGND VPWR VPWR _7386_/Q sky130_fd_sc_hd__dfstp_1
X_4598_ _5015_/C _5017_/B VGND VGND VPWR VPWR _5094_/A sky130_fd_sc_hd__and2_4
Xhold942 hold942/A VGND VGND VPWR VPWR wb_ack_o sky130_fd_sc_hd__buf_12
XFILLER_122_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold953 _7689_/A VGND VGND VPWR VPWR hold953/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold964 _5954_/X VGND VGND VPWR VPWR _7535_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6337_ _7126_/Q _6130_/X _6159_/X _7106_/Q _6336_/X VGND VGND VPWR VPWR _6337_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3549_ _3714_/A hold74/A _5939_/B VGND VGND VPWR VPWR _3549_/X sky130_fd_sc_hd__and3_4
Xhold975 _7379_/Q VGND VGND VPWR VPWR hold975/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold986 _5632_/X VGND VGND VPWR VPWR _7254_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold997 _7543_/Q VGND VGND VPWR VPWR hold997/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6268_ _7455_/Q _6213_/B _6170_/C _6159_/X _7439_/Q VGND VGND VPWR VPWR _6268_/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_76_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5219_ _4625_/Y _5585_/A1 _4677_/Y _4984_/Y _4998_/Y VGND VGND VPWR VPWR _5221_/B
+ sky130_fd_sc_hd__o32a_1
X_6199_ _7524_/Q _6309_/B _6334_/C _6132_/X _7452_/Q VGND VGND VPWR VPWR _6199_/X
+ sky130_fd_sc_hd__a32o_1
Xhold1620 _7294_/Q VGND VGND VPWR VPWR hold1620/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1631 _6100_/Y VGND VGND VPWR VPWR _7632_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1642 _7049_/Q VGND VGND VPWR VPWR hold452/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1653 _4079_/X VGND VGND VPWR VPWR _4081_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_532 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5570_ _5570_/A _5570_/B _5570_/C _5570_/D VGND VGND VPWR VPWR _5572_/C sky130_fd_sc_hd__nand4_1
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4521_ _4521_/A0 _6865_/A1 _4522_/S VGND VGND VPWR VPWR _4521_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold205 _7265_/Q VGND VGND VPWR VPWR hold205/X sky130_fd_sc_hd__dlygate4sd3_1
X_7240_ _7240_/CLK _7240_/D fanout603/X VGND VGND VPWR VPWR _7240_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_117_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4452_ _3655_/Y _4452_/A1 _4453_/S VGND VGND VPWR VPWR _7149_/D sky130_fd_sc_hd__mux2_1
Xhold216 _7350_/Q VGND VGND VPWR VPWR hold216/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 _5827_/X VGND VGND VPWR VPWR _7422_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 _5872_/X VGND VGND VPWR VPWR _7462_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 _7606_/Q VGND VGND VPWR VPWR hold249/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7171_ _7238_/CLK _7171_/D fanout602/X VGND VGND VPWR VPWR _7171_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_171_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4383_ _6012_/A0 _4383_/A1 _4387_/S VGND VGND VPWR VPWR _4383_/X sky130_fd_sc_hd__mux2_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6122_ _7434_/Q _6416_/B _6159_/A _6170_/C _7322_/Q VGND VGND VPWR VPWR _6122_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _6053_/A _6053_/B VGND VGND VPWR VPWR _6053_/X sky130_fd_sc_hd__and2_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _5094_/A _5109_/A VGND VGND VPWR VPWR _5004_/Y sky130_fd_sc_hd__nand2_2
XFILLER_66_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6955_ _6955_/D _4193_/X VGND VGND VPWR VPWR _6955_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5906_ hold806/X _6041_/A1 _5911_/S VGND VGND VPWR VPWR _5906_/X sky130_fd_sc_hd__mux2_1
X_6886_ _6886_/A _6911_/B VGND VGND VPWR VPWR _6886_/X sky130_fd_sc_hd__and2_1
X_5837_ hold924/X _6044_/A1 _5839_/S VGND VGND VPWR VPWR _5837_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5768_ _5984_/B _5768_/B _5768_/C _6861_/C VGND VGND VPWR VPWR _5776_/S sky130_fd_sc_hd__nand4_4
XFILLER_6_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7507_ _7601_/CLK _7507_/D fanout611/X VGND VGND VPWR VPWR _7507_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_147_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4719_ _5143_/B _4706_/D _4580_/Y _4950_/D _4718_/X VGND VGND VPWR VPWR _4770_/A
+ sky130_fd_sc_hd__o311a_2
X_5699_ _6041_/A1 hold727/X _5704_/S VGND VGND VPWR VPWR _5699_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7438_ _7586_/CLK _7438_/D fanout625/X VGND VGND VPWR VPWR _7438_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_190_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold750 _7220_/Q VGND VGND VPWR VPWR hold750/X sky130_fd_sc_hd__dlygate4sd3_1
X_7369_ _7445_/CLK _7369_/D fanout628/X VGND VGND VPWR VPWR _7369_/Q sky130_fd_sc_hd__dfrtp_2
Xhold761 _7580_/Q VGND VGND VPWR VPWR hold761/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold772 _6023_/X VGND VGND VPWR VPWR _7596_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap480 _6363_/A1 VGND VGND VPWR VPWR _6082_/A sky130_fd_sc_hd__clkbuf_2
Xhold783 hold783/A VGND VGND VPWR VPWR hold783/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap491 _5291_/B VGND VGND VPWR VPWR _5093_/C sky130_fd_sc_hd__clkbuf_2
Xhold794 _7471_/Q VGND VGND VPWR VPWR hold794/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1450 _7158_/Q VGND VGND VPWR VPWR _4462_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1461 _6185_/X VGND VGND VPWR VPWR _7638_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_55_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1472 _5832_/X VGND VGND VPWR VPWR _7426_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1483 _7145_/Q VGND VGND VPWR VPWR _4448_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_601 _6428_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1494 _5796_/X VGND VGND VPWR VPWR _7394_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_612 _4172_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_623 _5666_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_634 _5021_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_645 _6137_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_656 _6153_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_667 _7122_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_678 _7703_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_689 input80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6740_ _7128_/Q _6487_/X _6738_/X _6739_/X VGND VGND VPWR VPWR _6740_/X sky130_fd_sc_hd__a211o_1
X_3952_ input96/X _3780_/X _3947_/X _3948_/X _3951_/X VGND VGND VPWR VPWR _3952_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_189_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6671_ _7433_/Q _6444_/X _6465_/X _7353_/Q _6670_/X VGND VGND VPWR VPWR _6671_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_31_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3883_ _3883_/A _3883_/B _3883_/C _3883_/D VGND VGND VPWR VPWR _3883_/Y sky130_fd_sc_hd__nor4_1
X_5622_ _5577_/X _5621_/Y _5573_/X VGND VGND VPWR VPWR _5622_/X sky130_fd_sc_hd__o21a_1
XFILLER_176_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5553_ _5553_/A _5553_/B VGND VGND VPWR VPWR _5553_/Y sky130_fd_sc_hd__nor2_1
XFILLER_191_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4504_ _5926_/A0 hold391/X _4504_/S VGND VGND VPWR VPWR _4504_/X sky130_fd_sc_hd__mux2_1
X_5484_ _5476_/A _5375_/C _4747_/B VGND VGND VPWR VPWR _5484_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_144_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7223_ _7294_/CLK _7223_/D fanout599/X VGND VGND VPWR VPWR _7223_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_105_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4435_ hold550/X _4564_/A1 _4435_/S VGND VGND VPWR VPWR _4435_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7154_ _7668_/CLK _7154_/D VGND VGND VPWR VPWR _7154_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout504 _4673_/X VGND VGND VPWR VPWR _5614_/C sky130_fd_sc_hd__buf_6
X_4366_ hold649/X _6863_/A1 _4369_/S VGND VGND VPWR VPWR _4366_/X sky130_fd_sc_hd__mux2_1
Xfanout515 hold85/X VGND VGND VPWR VPWR _5999_/A1 sky130_fd_sc_hd__buf_6
XFILLER_59_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout526 _5988_/A1 VGND VGND VPWR VPWR _6006_/A1 sky130_fd_sc_hd__clkbuf_4
X_6105_ _7142_/Q _7139_/Q _6811_/S _6109_/B _6104_/X VGND VGND VPWR VPWR _6108_/S
+ sky130_fd_sc_hd__o41a_1
XFILLER_98_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout548 _5686_/D VGND VGND VPWR VPWR _5680_/C sky130_fd_sc_hd__buf_6
XFILLER_100_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7085_ _7130_/CLK _7085_/D fanout602/X VGND VGND VPWR VPWR _7085_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout559 _6359_/B VGND VGND VPWR VPWR _6131_/B sky130_fd_sc_hd__buf_6
X_4297_ hold289/X _5761_/A1 _4303_/S VGND VGND VPWR VPWR _4297_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6036_ _6045_/A1 hold573/X _6037_/S VGND VGND VPWR VPWR _6036_/X sky130_fd_sc_hd__mux2_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6938_ _4172_/B2 _6938_/D _6893_/X VGND VGND VPWR VPWR _6938_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6869_ _6899_/A _6911_/B VGND VGND VPWR VPWR _6869_/X sky130_fd_sc_hd__and2_1
XFILLER_22_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold580 _5892_/X VGND VGND VPWR VPWR _7480_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold591 _7416_/Q VGND VGND VPWR VPWR hold591/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_106_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1280 _7438_/Q VGND VGND VPWR VPWR hold552/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1291 _7681_/Q VGND VGND VPWR VPWR _4203_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_420 _6124_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_431 _6192_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_442 _6645_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_453 _6465_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_464 _6700_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_475 _7071_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_486 _7570_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_497 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4220_ _4220_/A0 _6864_/A1 _4230_/S VGND VGND VPWR VPWR _6974_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4151_ _7300_/Q input80/X _4196_/B VGND VGND VPWR VPWR _4151_/X sky130_fd_sc_hd__mux2_2
XFILLER_68_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4082_ _6925_/Q hold21/A hold94/A VGND VGND VPWR VPWR _4082_/X sky130_fd_sc_hd__a21o_1
XFILLER_83_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4984_ _5042_/A _5297_/C VGND VGND VPWR VPWR _4984_/Y sky130_fd_sc_hd__nand2_2
XFILLER_51_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6723_ _7180_/Q _6465_/X _6479_/X _7220_/Q _6722_/X VGND VGND VPWR VPWR _6723_/X
+ sky130_fd_sc_hd__a221o_1
X_3935_ _7459_/Q _3549_/X _3716_/X _7262_/Q _3934_/X VGND VGND VPWR VPWR _3935_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_32_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6654_ _7544_/Q _6479_/X _6486_/X _7504_/Q _6653_/X VGND VGND VPWR VPWR _6659_/A
+ sky130_fd_sc_hd__a221o_1
X_3866_ _7468_/Q _5903_/A _6020_/A _3703_/X _7113_/Q VGND VGND VPWR VPWR _3866_/X
+ sky130_fd_sc_hd__a32o_1
X_5605_ _5314_/B _5605_/B _5605_/C _5605_/D VGND VGND VPWR VPWR _5626_/C sky130_fd_sc_hd__and4b_1
XFILLER_176_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6585_ _6686_/S _7652_/Q _6583_/X _6584_/X VGND VGND VPWR VPWR _6585_/X sky130_fd_sc_hd__a22o_1
X_3797_ _7104_/Q _3516_/X _5666_/B _4257_/S input46/X VGND VGND VPWR VPWR _3797_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_176_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5536_ _5536_/A _5536_/B _5536_/C VGND VGND VPWR VPWR _5537_/C sky130_fd_sc_hd__and3_1
X_5467_ _5617_/A _5534_/B _5586_/B _5617_/B VGND VGND VPWR VPWR _5468_/C sky130_fd_sc_hd__and4_1
X_7206_ _7217_/CLK _7206_/D _6903_/A VGND VGND VPWR VPWR _7206_/Q sky130_fd_sc_hd__dfstp_2
X_4418_ _4541_/A _5661_/B _4493_/C _6861_/C VGND VGND VPWR VPWR _4423_/S sky130_fd_sc_hd__nand4_4
X_5398_ _5017_/A _4877_/C _4859_/Y _5381_/X _5526_/A VGND VGND VPWR VPWR _5399_/D
+ sky130_fd_sc_hd__o41a_1
XFILLER_99_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7137_ _7462_/CLK hold57/X fanout604/X VGND VGND VPWR VPWR _7137_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_113_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4349_ _5789_/A1 hold357/X _4351_/S VGND VGND VPWR VPWR _4349_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout378 _6038_/B VGND VGND VPWR VPWR _5680_/B sky130_fd_sc_hd__buf_6
XFILLER_47_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout389 _3550_/B VGND VGND VPWR VPWR _5840_/A sky130_fd_sc_hd__buf_8
X_7068_ _7212_/CLK _7068_/D fanout619/X VGND VGND VPWR VPWR _7068_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_86_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6019_ _6046_/A1 hold918/X _6019_/S VGND VGND VPWR VPWR _6019_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_250 input38/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_261 input62/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_272 input80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_283 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_294 input95/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3720_ _7203_/Q _3696_/X _4499_/A _7193_/Q _3719_/X VGND VGND VPWR VPWR _3720_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3651_ input9/X _5957_/B _3573_/C _3650_/X VGND VGND VPWR VPWR _3651_/X sky130_fd_sc_hd__a31o_1
XFILLER_158_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6370_ _7078_/Q _6119_/X _6213_/B _6369_/X VGND VGND VPWR VPWR _6370_/X sky130_fd_sc_hd__a211o_2
X_3582_ _5661_/A _3717_/B _4481_/A VGND VGND VPWR VPWR _6029_/A sky130_fd_sc_hd__and3_4
X_5321_ _5319_/Y _5320_/X _5149_/X VGND VGND VPWR VPWR _5325_/C sky130_fd_sc_hd__a21o_1
XFILLER_161_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5252_ _4882_/Y _5604_/B1 _5015_/Y _5251_/X _4874_/Y VGND VGND VPWR VPWR _5256_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_142_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4203_ hold27/X _4203_/A1 _4229_/S VGND VGND VPWR VPWR hold28/A sky130_fd_sc_hd__mux2_1
XFILLER_114_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5183_ _4597_/Y _4629_/Y _4706_/Y _4805_/Y _5011_/C VGND VGND VPWR VPWR _5184_/C
+ sky130_fd_sc_hd__o32a_1
X_4134_ _6950_/Q hold27/A _6907_/B VGND VGND VPWR VPWR _4202_/A sky130_fd_sc_hd__o21ai_1
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4065_ _6929_/Q _4064_/X _3478_/X VGND VGND VPWR VPWR _4065_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_37_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4967_ _5021_/B _5404_/B VGND VGND VPWR VPWR _4971_/D sky130_fd_sc_hd__nand2_1
X_3918_ _7547_/Q _3514_/X _3569_/X _7595_/Q _3917_/X VGND VGND VPWR VPWR _3918_/X
+ sky130_fd_sc_hd__a221o_1
X_6706_ _7106_/Q _6099_/B _6694_/C _6469_/X _7164_/Q VGND VGND VPWR VPWR _6706_/X
+ sky130_fd_sc_hd__a32o_1
X_7686_ _7686_/CLK _7686_/D fanout600/X VGND VGND VPWR VPWR _7686_/Q sky130_fd_sc_hd__dfrtp_2
X_4898_ _4946_/A _4901_/B _4901_/C _4950_/C VGND VGND VPWR VPWR _4900_/C sky130_fd_sc_hd__nand4_1
XFILLER_165_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6637_ _7608_/Q _6791_/B _6791_/C _6791_/D VGND VGND VPWR VPWR _6637_/X sky130_fd_sc_hd__and4_1
X_3849_ _7128_/Q _4559_/B _4553_/B _3846_/X _3848_/X VGND VGND VPWR VPWR _3849_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_164_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6568_ _7365_/Q _6694_/B _6445_/C _6463_/X _7397_/Q VGND VGND VPWR VPWR _6568_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_152_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5519_ _5602_/D _5316_/X _5516_/X _5501_/Y VGND VGND VPWR VPWR _5519_/X sky130_fd_sc_hd__o31a_1
X_6499_ _7402_/Q _6466_/X _6485_/X _7546_/Q _6461_/X VGND VGND VPWR VPWR _6499_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_106_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire576 _5002_/B VGND VGND VPWR VPWR _5191_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_109_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5870_ hold647/X _6041_/A1 _5875_/S VGND VGND VPWR VPWR _5870_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4821_ _5131_/A _5040_/A VGND VGND VPWR VPWR _4821_/Y sky130_fd_sc_hd__nand2_8
XFILLER_21_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7540_ _7580_/CLK _7540_/D fanout605/X VGND VGND VPWR VPWR _7540_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4752_ _5233_/A _4748_/B _4751_/Y VGND VGND VPWR VPWR _4762_/A sky130_fd_sc_hd__a21oi_1
X_3703_ _3714_/A hold74/A _4529_/B VGND VGND VPWR VPWR _3703_/X sky130_fd_sc_hd__and3_1
X_7471_ _7512_/CLK _7471_/D fanout610/X VGND VGND VPWR VPWR _7471_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_174_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4683_ _4738_/A _4738_/B _5614_/C _4740_/D VGND VGND VPWR VPWR _4739_/D sky130_fd_sc_hd__nand4_1
XFILLER_119_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6422_ _7090_/Q _6149_/X _6420_/X _6421_/X VGND VGND VPWR VPWR _6422_/X sky130_fd_sc_hd__a211o_1
XFILLER_147_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3634_ _7368_/Q _3581_/X _3626_/X _3628_/X _3633_/X VGND VGND VPWR VPWR _3634_/Y
+ sky130_fd_sc_hd__a2111oi_4
XFILLER_162_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6353_ _7683_/Q _6166_/B _6166_/C _6082_/B VGND VGND VPWR VPWR _6353_/X sky130_fd_sc_hd__a31o_1
XFILLER_162_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3565_ _5768_/C _6002_/A _5768_/B VGND VGND VPWR VPWR _3565_/X sky130_fd_sc_hd__and3_4
XFILLER_108_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5304_ _5038_/B _5313_/A _5289_/X _5303_/X VGND VGND VPWR VPWR _5304_/Y sky130_fd_sc_hd__a211oi_1
X_6284_ _7536_/Q _6160_/D _6427_/A3 _6137_/X _7488_/Q VGND VGND VPWR VPWR _6284_/X
+ sky130_fd_sc_hd__a32o_1
X_3496_ hold53/X _3568_/C VGND VGND VPWR VPWR _5686_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5235_ _4800_/Y _4816_/Y _4821_/Y _5080_/Y VGND VGND VPWR VPWR _5235_/X sky130_fd_sc_hd__o31a_1
XFILLER_69_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5166_ _4619_/Y _4660_/C _4685_/Y _4912_/Y _4681_/Y VGND VGND VPWR VPWR _5166_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_69_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4117_ input123/X input122/X _4117_/C _4117_/D VGND VGND VPWR VPWR _4117_/X sky130_fd_sc_hd__and4bb_4
X_5097_ _5189_/D _5108_/B _5146_/B _5131_/A VGND VGND VPWR VPWR _5097_/Y sky130_fd_sc_hd__nand4_1
XFILLER_56_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4048_ _4049_/B _4048_/B VGND VGND VPWR VPWR _4048_/Y sky130_fd_sc_hd__nor2_1
XFILLER_71_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5999_ hold827/X _5999_/A1 _6001_/S VGND VGND VPWR VPWR _5999_/X sky130_fd_sc_hd__mux2_1
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7669_ _7672_/CLK _7669_/D VGND VGND VPWR VPWR _7669_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_149_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput290 _6975_/Q VGND VGND VPWR VPWR pll_trim[3] sky130_fd_sc_hd__buf_12
XFILLER_160_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold9 hold9/A VGND VGND VPWR VPWR hold9/X sky130_fd_sc_hd__buf_6
XFILLER_87_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire351 _4005_/Y VGND VGND VPWR VPWR _4037_/B sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_62_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7580_/CLK sky130_fd_sc_hd__clkbuf_16
Xwire373 _6775_/Y VGND VGND VPWR VPWR wire373/X sky130_fd_sc_hd__clkbuf_1
XFILLER_156_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold409 _7082_/Q VGND VGND VPWR VPWR hold409/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire395 wire396/X VGND VGND VPWR VPWR _4469_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_171_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_77_csclk _7095_/CLK VGND VGND VPWR VPWR _7294_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _5316_/A _5512_/B _5112_/B VGND VGND VPWR VPWR _5020_/X sky130_fd_sc_hd__and3_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1109 hold1595/X VGND VGND VPWR VPWR _4367_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6971_ _7680_/CLK _6971_/D _6815_/A VGND VGND VPWR VPWR _6971_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5922_ hold44/X _5922_/A1 hold76/A VGND VGND VPWR VPWR hold77/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_15_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7207_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5853_ _6006_/A1 _5853_/A1 _5857_/S VGND VGND VPWR VPWR _7445_/D sky130_fd_sc_hd__mux2_1
XFILLER_21_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4804_ _5108_/B _5131_/A _5146_/C VGND VGND VPWR VPWR _5318_/B sky130_fd_sc_hd__and3_2
XFILLER_179_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5784_ hold50/X hold111/X _5785_/S VGND VGND VPWR VPWR _5784_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4735_ _4735_/A _4735_/B _4735_/C _5466_/C VGND VGND VPWR VPWR _4737_/B sky130_fd_sc_hd__nand4_1
X_7523_ _7602_/CLK _7523_/D fanout615/X VGND VGND VPWR VPWR _7523_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_159_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7454_ _7601_/CLK _7454_/D fanout611/X VGND VGND VPWR VPWR _7454_/Q sky130_fd_sc_hd__dfrtp_4
X_4666_ _5000_/C _4568_/Y _5015_/C VGND VGND VPWR VPWR _4706_/B sky130_fd_sc_hd__a21oi_1
XFILLER_175_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6405_ _7109_/Q _6159_/X _6402_/X _6404_/X VGND VGND VPWR VPWR _6405_/X sky130_fd_sc_hd__a211o_1
XFILLER_190_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3617_ _3617_/A _3617_/B _3617_/C _3617_/D VGND VGND VPWR VPWR _3617_/Y sky130_fd_sc_hd__nor4_1
XFILLER_134_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7385_ _7568_/CLK _7385_/D fanout622/X VGND VGND VPWR VPWR _7385_/Q sky130_fd_sc_hd__dfrtp_2
Xhold910 _7433_/Q VGND VGND VPWR VPWR hold910/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 _4362_/X VGND VGND VPWR VPWR _7069_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4597_ _4884_/A _4597_/B _4597_/C _5143_/A VGND VGND VPWR VPWR _4597_/Y sky130_fd_sc_hd__nand4b_4
Xhold932 _4276_/X VGND VGND VPWR VPWR _7003_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold943 _7567_/Q VGND VGND VPWR VPWR hold943/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold954 _4284_/X VGND VGND VPWR VPWR _7006_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6336_ _7189_/Q _6082_/B _6427_/B1 _6157_/X _7101_/Q VGND VGND VPWR VPWR _6336_/X
+ sky130_fd_sc_hd__a32o_1
X_3548_ _5661_/A _5661_/B _5682_/C VGND VGND VPWR VPWR hold37/A sky130_fd_sc_hd__and3_2
Xhold965 _7419_/Q VGND VGND VPWR VPWR hold965/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold976 hold976/A VGND VGND VPWR VPWR hold976/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 hold987/A VGND VGND VPWR VPWR hold987/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold998 _5963_/X VGND VGND VPWR VPWR _7543_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6267_ _7567_/Q _6153_/X _6157_/X _7503_/Q _6266_/X VGND VGND VPWR VPWR _6267_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3479_ _6912_/Q _3500_/C VGND VGND VPWR VPWR _3508_/S sky130_fd_sc_hd__nand2_4
X_5218_ _5217_/X _5002_/X _5218_/C _5218_/D VGND VGND VPWR VPWR _5221_/A sky130_fd_sc_hd__and4bb_1
XFILLER_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6198_ _7516_/Q _6146_/X _6160_/X _7372_/Q _6197_/X VGND VGND VPWR VPWR _6198_/X
+ sky130_fd_sc_hd__a221o_1
Xhold1610 hold94/A VGND VGND VPWR VPWR _4084_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1621 _7256_/Q VGND VGND VPWR VPWR _3470_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1632 _7578_/Q VGND VGND VPWR VPWR hold818/A sky130_fd_sc_hd__dlygate4sd3_1
X_5149_ _5517_/A2 _5143_/X _6969_/Q _6971_/Q _6970_/Q VGND VGND VPWR VPWR _5149_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_185_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1643 _7499_/Q VGND VGND VPWR VPWR _5914_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1654 _7147_/Q VGND VGND VPWR VPWR _4450_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4520_ _4520_/A0 _4556_/A1 _4522_/S VGND VGND VPWR VPWR _4520_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold206 _5642_/X VGND VGND VPWR VPWR _7265_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4451_ _3692_/Y _4451_/A1 _4453_/S VGND VGND VPWR VPWR _7148_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold217 _5746_/X VGND VGND VPWR VPWR _7350_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 hold228/A VGND VGND VPWR VPWR hold228/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold239 _7125_/Q VGND VGND VPWR VPWR hold239/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7170_ _7238_/CLK _7170_/D fanout602/X VGND VGND VPWR VPWR _7170_/Q sky130_fd_sc_hd__dfrtp_2
X_4382_ _4382_/A _6861_/C VGND VGND VPWR VPWR _4387_/S sky130_fd_sc_hd__nand2_2
XFILLER_98_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6121_ _7624_/Q _6151_/B _6126_/D _7623_/Q VGND VGND VPWR VPWR _6170_/C sky130_fd_sc_hd__and4bb_4
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6052_ _6053_/B _6053_/A VGND VGND VPWR VPWR _6052_/Y sky130_fd_sc_hd__nor2_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _5007_/A _5094_/A _5007_/D VGND VGND VPWR VPWR _5110_/C sky130_fd_sc_hd__and3_4
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6954_ _4183_/A1 _6954_/D _6908_/X VGND VGND VPWR VPWR _6954_/Q sky130_fd_sc_hd__dfrtp_4
X_5905_ hold143/X _6031_/A0 _5911_/S VGND VGND VPWR VPWR _5905_/X sky130_fd_sc_hd__mux2_1
X_6885_ _6911_/A _6911_/B VGND VGND VPWR VPWR _6885_/X sky130_fd_sc_hd__and2_1
XFILLER_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5836_ hold284/X _5935_/A1 _5839_/S VGND VGND VPWR VPWR _5836_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5767_ hold109/X hold102/X _5767_/S VGND VGND VPWR VPWR _5767_/X sky130_fd_sc_hd__mux2_1
X_7506_ _7566_/CLK hold77/X fanout621/X VGND VGND VPWR VPWR _7506_/Q sky130_fd_sc_hd__dfstp_1
X_4718_ _4781_/B _4781_/C _4581_/X _4595_/B VGND VGND VPWR VPWR _4718_/X sky130_fd_sc_hd__a31o_1
X_5698_ _6863_/A1 hold736/X _5703_/S VGND VGND VPWR VPWR _5698_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7437_ _7445_/CLK _7437_/D fanout628/X VGND VGND VPWR VPWR _7437_/Q sky130_fd_sc_hd__dfrtp_4
X_4649_ _5189_/A _4992_/B _4822_/A _4992_/D _5008_/C VGND VGND VPWR VPWR _4649_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_107_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold740 _6973_/Q VGND VGND VPWR VPWR hold740/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 _4537_/X VGND VGND VPWR VPWR _7220_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7368_ _7445_/CLK _7368_/D fanout628/X VGND VGND VPWR VPWR _7368_/Q sky130_fd_sc_hd__dfrtp_2
Xhold762 _6005_/X VGND VGND VPWR VPWR _7580_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap481 _6180_/A2 VGND VGND VPWR VPWR _6363_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_116_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold773 _7360_/Q VGND VGND VPWR VPWR hold773/X sky130_fd_sc_hd__dlygate4sd3_1
X_6319_ _7321_/Q _6082_/Y _6686_/S VGND VGND VPWR VPWR _6319_/X sky130_fd_sc_hd__o21ba_1
Xhold784 hold784/A VGND VGND VPWR VPWR hold784/X sky130_fd_sc_hd__dlygate4sd3_1
X_7299_ _7462_/CLK _7299_/D fanout604/X VGND VGND VPWR VPWR _7299_/Q sky130_fd_sc_hd__dfrtp_1
Xhold795 _5882_/X VGND VGND VPWR VPWR _7471_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1440 _7330_/Q VGND VGND VPWR VPWR hold1440/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1451 _7325_/Q VGND VGND VPWR VPWR hold1451/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1462 _7354_/Q VGND VGND VPWR VPWR hold449/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1473 _6918_/Q VGND VGND VPWR VPWR _4099_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1484 _7157_/Q VGND VGND VPWR VPWR _4461_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_176_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1495 _7151_/Q VGND VGND VPWR VPWR _4455_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_602 _6302_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_613 hold85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_624 _5666_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_635 _5884_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_646 _6137_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_657 _6645_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_668 _7114_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_679 input38/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3951_ _7127_/Q _4559_/B _5678_/B _3949_/X _3950_/X VGND VGND VPWR VPWR _3951_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_63_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6670_ _7529_/Q _6469_/A _6562_/C _6474_/A _7345_/Q VGND VGND VPWR VPWR _6670_/X
+ sky130_fd_sc_hd__a32o_1
X_3882_ _7596_/Q _3569_/X _3875_/X _3876_/X _3881_/X VGND VGND VPWR VPWR _3883_/D
+ sky130_fd_sc_hd__a2111o_1
X_5621_ _5621_/A _5621_/B _5621_/C VGND VGND VPWR VPWR _5621_/Y sky130_fd_sc_hd__nand3_1
XFILLER_188_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5552_ _5552_/A _5552_/B _5552_/C VGND VGND VPWR VPWR _5553_/B sky130_fd_sc_hd__nand3_1
X_4503_ _5988_/A1 hold786/X _4504_/S VGND VGND VPWR VPWR _4503_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5483_ _5597_/A _5597_/C _5597_/D VGND VGND VPWR VPWR _5487_/C sky130_fd_sc_hd__and3_1
XFILLER_145_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7222_ _7231_/CLK _7222_/D fanout599/X VGND VGND VPWR VPWR _7222_/Q sky130_fd_sc_hd__dfrtp_4
X_4434_ hold640/X _5673_/A1 _4435_/S VGND VGND VPWR VPWR _4434_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7153_ _7668_/CLK _7153_/D VGND VGND VPWR VPWR _7153_/Q sky130_fd_sc_hd__dfxtp_1
X_4365_ _4365_/A0 _5697_/A0 _4369_/S VGND VGND VPWR VPWR _7071_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout505 _5068_/A VGND VGND VPWR VPWR _5476_/A sky130_fd_sc_hd__buf_6
XFILLER_116_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout516 hold85/X VGND VGND VPWR VPWR _6044_/A1 sky130_fd_sc_hd__buf_6
X_6104_ _6107_/C _6056_/Y _3421_/Y VGND VGND VPWR VPWR _6104_/X sky130_fd_sc_hd__a21o_1
Xfanout527 hold9/X VGND VGND VPWR VPWR _5988_/A1 sky130_fd_sc_hd__buf_6
Xfanout538 _5869_/A1 VGND VGND VPWR VPWR _6863_/A1 sky130_fd_sc_hd__buf_6
X_7084_ _7192_/CLK _7084_/D fanout619/X VGND VGND VPWR VPWR _7084_/Q sky130_fd_sc_hd__dfrtp_1
X_4296_ hold453/X _6003_/A1 _4303_/S VGND VGND VPWR VPWR _4296_/X sky130_fd_sc_hd__mux2_1
Xfanout549 hold29/X VGND VGND VPWR VPWR _5686_/D sky130_fd_sc_hd__buf_6
XFILLER_112_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6035_ _6044_/A1 hold960/X _6037_/S VGND VGND VPWR VPWR _6035_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6937_ _4172_/B2 _6937_/D _6892_/X VGND VGND VPWR VPWR hold48/A sky130_fd_sc_hd__dfrtp_1
XFILLER_54_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6868_ _6899_/A _6911_/B VGND VGND VPWR VPWR _6868_/X sky130_fd_sc_hd__and2_1
X_5819_ hold85/X hold262/X _5821_/S VGND VGND VPWR VPWR _5819_/X sky130_fd_sc_hd__mux2_1
XFILLER_167_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6799_ _7090_/Q _6458_/X _6481_/X _7213_/Q _6798_/X VGND VGND VPWR VPWR _6800_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_167_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold570 hold570/A VGND VGND VPWR VPWR hold570/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 _7304_/Q VGND VGND VPWR VPWR hold581/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold592 _5820_/X VGND VGND VPWR VPWR _7416_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1270 _7477_/Q VGND VGND VPWR VPWR hold1270/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1281 _5845_/X VGND VGND VPWR VPWR _7438_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1292 _5779_/X VGND VGND VPWR VPWR _7379_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_410 _5884_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_421 _6153_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_432 _6192_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_443 _6645_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_454 _6465_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_465 _6754_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_476 _7071_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_487 _7579_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_498 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4150_ _7597_/Q _4196_/B _4149_/Y VGND VGND VPWR VPWR _4150_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4081_ _4081_/A1 _4080_/X _3498_/X _4043_/Y VGND VGND VPWR VPWR _6927_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4983_ _5143_/A _5042_/A _4983_/C VGND VGND VPWR VPWR _4985_/B sky130_fd_sc_hd__and3_2
XFILLER_189_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6722_ _7240_/Q _6694_/B _6720_/D _6485_/X _7215_/Q VGND VGND VPWR VPWR _6722_/X
+ sky130_fd_sc_hd__a32o_1
X_3934_ _7683_/Q _4559_/B hold98/A _3710_/X _7072_/Q VGND VGND VPWR VPWR _3934_/X
+ sky130_fd_sc_hd__a32o_1
X_6653_ _7480_/Q _6441_/X _6482_/X _7488_/Q _6652_/X VGND VGND VPWR VPWR _6653_/X
+ sky130_fd_sc_hd__a221o_1
X_3865_ input45/X _4257_/S _3583_/X input54/X _3864_/X VGND VGND VPWR VPWR _3865_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_31_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5604_ _4816_/Y _4953_/C _5604_/B1 _4756_/Y VGND VGND VPWR VPWR _5605_/D sky130_fd_sc_hd__a211o_1
XFILLER_164_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6584_ _7317_/Q _6759_/D _6686_/S VGND VGND VPWR VPWR _6584_/X sky130_fd_sc_hd__o21ba_1
X_3796_ _7581_/Q _3584_/X _3784_/X _3788_/X _3795_/X VGND VGND VPWR VPWR _3796_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_191_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5535_ _5614_/C _4702_/X _5614_/A _5043_/B _5614_/B VGND VGND VPWR VPWR _5536_/C
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_127_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5466_ _5209_/C _5466_/B _5466_/C VGND VGND VPWR VPWR _5617_/B sky130_fd_sc_hd__and3b_1
XFILLER_127_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4417_ hold201/X _6866_/A1 _4417_/S VGND VGND VPWR VPWR _4417_/X sky130_fd_sc_hd__mux2_1
X_7205_ _7217_/CLK _7205_/D _6903_/A VGND VGND VPWR VPWR _7205_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_105_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5397_ _4769_/Y _4953_/C _4867_/X _4910_/Y VGND VGND VPWR VPWR _5526_/B sky130_fd_sc_hd__a211o_1
X_7136_ _7614_/CLK hold91/X fanout604/X VGND VGND VPWR VPWR _7136_/Q sky130_fd_sc_hd__dfstp_2
X_4348_ _5761_/A1 hold385/X _4351_/S VGND VGND VPWR VPWR _4348_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7067_ _7210_/CLK _7067_/D fanout621/X VGND VGND VPWR VPWR _7067_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout379 _6002_/B VGND VGND VPWR VPWR _6038_/B sky130_fd_sc_hd__buf_12
X_4279_ _5697_/A1 _5697_/A0 _4291_/S VGND VGND VPWR VPWR _4279_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6018_ _6045_/A1 hold553/X _6019_/S VGND VGND VPWR VPWR _6018_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_240 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_251 input38/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_262 _4196_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_273 input80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_284 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_295 input95/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3650_ _7496_/Q _5903_/A _5975_/B hold75/A _7512_/Q VGND VGND VPWR VPWR _3650_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_9_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3581_ _3713_/A _3581_/B _5759_/B VGND VGND VPWR VPWR _3581_/X sky130_fd_sc_hd__and3_4
XFILLER_161_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5320_ _5407_/B _5102_/B _4821_/Y _4948_/A _4795_/Y VGND VGND VPWR VPWR _5320_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5251_ _4629_/Y _5011_/C _4953_/B _4859_/Y VGND VGND VPWR VPWR _5251_/X sky130_fd_sc_hd__a211o_1
X_4202_ _4202_/A _6969_/Q VGND VGND VPWR VPWR _6966_/D sky130_fd_sc_hd__and2_1
XFILLER_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5182_ _5182_/A _5182_/B _5182_/C VGND VGND VPWR VPWR _5184_/B sky130_fd_sc_hd__nor3_1
X_4133_ _6950_/Q hold27/A _6907_/B VGND VGND VPWR VPWR _4133_/X sky130_fd_sc_hd__o21a_1
XFILLER_110_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4064_ _6928_/Q _4064_/B VGND VGND VPWR VPWR _4064_/X sky130_fd_sc_hd__and2_1
XFILLER_113_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4966_ _4966_/A _4966_/B _5452_/B VGND VGND VPWR VPWR _4968_/B sky130_fd_sc_hd__and3_1
XFILLER_189_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6705_ _7239_/Q _6694_/B _6720_/D _6451_/X _7041_/Q VGND VGND VPWR VPWR _6705_/X
+ sky130_fd_sc_hd__a32o_1
X_3917_ _7411_/Q _5628_/A _3529_/X _3916_/X VGND VGND VPWR VPWR _3917_/X sky130_fd_sc_hd__a31o_1
XFILLER_149_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7685_ _7685_/CLK _7685_/D fanout617/X VGND VGND VPWR VPWR _7685_/Q sky130_fd_sc_hd__dfrtp_2
X_4897_ _4779_/X _4833_/X _4892_/B _4907_/C _4907_/A VGND VGND VPWR VPWR _4901_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6636_ _6635_/X _6661_/A1 _6812_/S VGND VGND VPWR VPWR _6636_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3848_ _7484_/Q _3531_/X _4388_/A _7093_/Q _3847_/X VGND VGND VPWR VPWR _3848_/X
+ sky130_fd_sc_hd__a221o_1
X_3779_ _7044_/Q _4529_/B _4481_/A VGND VGND VPWR VPWR _3779_/X sky130_fd_sc_hd__and3_1
XFILLER_164_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6567_ _7357_/Q _6454_/X _6469_/X _7333_/Q VGND VGND VPWR VPWR _6567_/X sky130_fd_sc_hd__a22o_1
XFILLER_192_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5518_ _5042_/A _5084_/X _5319_/A _5517_/X VGND VGND VPWR VPWR _5602_/D sky130_fd_sc_hd__a211o_1
XFILLER_105_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6498_ _7410_/Q _6450_/X _6481_/X _7378_/Q _6488_/X VGND VGND VPWR VPWR _6498_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_145_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5449_ _5604_/B1 _4960_/Y _4998_/Y _4912_/Y _4867_/X VGND VGND VPWR VPWR _5449_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_160_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7119_ _7685_/CLK _7119_/D fanout617/X VGND VGND VPWR VPWR _7119_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_86_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_wbbd_sck clkbuf_0_wbbd_sck/X VGND VGND VPWR VPWR _4172_/A2 sky130_fd_sc_hd__clkbuf_16
XFILLER_42_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4820_ _4990_/A _5014_/D _5015_/C _5017_/B VGND VGND VPWR VPWR _5021_/A sky130_fd_sc_hd__nor4_4
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751_ _4751_/A _4751_/B _4751_/C VGND VGND VPWR VPWR _4751_/Y sky130_fd_sc_hd__nand3_1
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3702_ _5993_/A _5682_/A _5659_/C VGND VGND VPWR VPWR _3702_/X sky130_fd_sc_hd__and3_4
XFILLER_119_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4682_ _4747_/B _4738_/B _5196_/A _4740_/D VGND VGND VPWR VPWR _4739_/C sky130_fd_sc_hd__nand4_1
X_7470_ _7606_/CLK _7470_/D fanout606/X VGND VGND VPWR VPWR _7470_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_147_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6421_ _7050_/Q _6231_/D _6166_/C _6432_/A3 _7100_/Q VGND VGND VPWR VPWR _6421_/X
+ sky130_fd_sc_hd__a32o_1
X_3633_ input59/X _5975_/B _4481_/A _3630_/X _3632_/X VGND VGND VPWR VPWR _3633_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_146_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3564_ _5686_/B _3568_/C hold53/X VGND VGND VPWR VPWR _4475_/A sky130_fd_sc_hd__and3_4
X_6352_ _7230_/Q _6160_/D _6427_/A3 _6429_/A3 _7122_/Q VGND VGND VPWR VPWR _6352_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_174_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5303_ _5311_/A _5038_/B _5091_/B _5093_/C _5302_/X VGND VGND VPWR VPWR _5303_/X
+ sky130_fd_sc_hd__a221o_1
X_6283_ _7456_/Q _6132_/X _6158_/X _7496_/Q _6282_/X VGND VGND VPWR VPWR _6283_/X
+ sky130_fd_sc_hd__a221o_1
X_3495_ _3494_/X hold52/X _4229_/S VGND VGND VPWR VPWR hold53/A sky130_fd_sc_hd__mux2_8
XFILLER_142_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5234_ _5429_/A _5318_/B _5233_/X _5232_/X VGND VGND VPWR VPWR _5234_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_130_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5165_ _4674_/Y _4769_/Y _5015_/D _4760_/D VGND VGND VPWR VPWR _5165_/X sky130_fd_sc_hd__a211o_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4116_ _4116_/A _4116_/B _4116_/C _4116_/D VGND VGND VPWR VPWR _4117_/D sky130_fd_sc_hd__and4_1
XFILLER_29_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5096_ _5096_/A _5096_/B _5096_/C _4884_/A VGND VGND VPWR VPWR _5096_/Y sky130_fd_sc_hd__nor4b_1
XFILLER_83_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4047_ _6941_/Q _6940_/Q _6939_/Q _4192_/B _4192_/C VGND VGND VPWR VPWR _4048_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5998_ hold264/X _6043_/A1 _6001_/S VGND VGND VPWR VPWR _5998_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4949_ _5189_/D _5112_/B VGND VGND VPWR VPWR _4949_/Y sky130_fd_sc_hd__nand2_4
XFILLER_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7668_ _7668_/CLK _7668_/D VGND VGND VPWR VPWR _7668_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6619_ _7519_/Q _6455_/C _6562_/C _6466_/X _7407_/Q VGND VGND VPWR VPWR _6619_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_193_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7599_ _7599_/CLK _7599_/D fanout629/X VGND VGND VPWR VPWR _7599_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_193_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput280 _7274_/Q VGND VGND VPWR VPWR pll_trim[18] sky130_fd_sc_hd__buf_12
XFILLER_160_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput291 _6976_/Q VGND VGND VPWR VPWR pll_trim[4] sky130_fd_sc_hd__buf_12
XFILLER_94_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire352 _3932_/Y VGND VGND VPWR VPWR _3965_/C sky130_fd_sc_hd__clkbuf_2
Xwire363 _4304_/Y VGND VGND VPWR VPWR _4311_/S sky130_fd_sc_hd__clkbuf_2
Xwire374 _6725_/Y VGND VGND VPWR VPWR wire374/X sky130_fd_sc_hd__clkbuf_1
XFILLER_156_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire396 hold97/X VGND VGND VPWR VPWR wire396/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6970_ _7680_/CLK _6970_/D _6815_/A VGND VGND VPWR VPWR _6970_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_66_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5921_ hold75/X _6038_/C VGND VGND VPWR VPWR hold76/A sky130_fd_sc_hd__nand2_8
XFILLER_80_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5852_ hold81/X hold311/X _5857_/S VGND VGND VPWR VPWR _5852_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4803_ _5131_/A _5025_/B _5017_/B VGND VGND VPWR VPWR _5071_/C sky130_fd_sc_hd__and3_2
XFILLER_167_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5783_ _6044_/A1 hold813/X _5785_/S VGND VGND VPWR VPWR _5783_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7522_ _7590_/CLK _7522_/D fanout605/X VGND VGND VPWR VPWR _7522_/Q sky130_fd_sc_hd__dfstp_2
X_4734_ _4747_/B _5490_/C _5476_/A _5595_/B VGND VGND VPWR VPWR _4735_/B sky130_fd_sc_hd__nand4_1
XFILLER_119_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7453_ _7553_/CLK _7453_/D fanout622/X VGND VGND VPWR VPWR _7453_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_190_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4665_ _5358_/A _5490_/C _5476_/A VGND VGND VPWR VPWR _4744_/A sky130_fd_sc_hd__and3_1
XFILLER_135_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6404_ _7192_/Q _6138_/X _6152_/X _7202_/Q _6403_/X VGND VGND VPWR VPWR _6404_/X
+ sky130_fd_sc_hd__a221o_1
X_3616_ _7441_/Q _3579_/X _3612_/X _3614_/X _3615_/X VGND VGND VPWR VPWR _3617_/D
+ sky130_fd_sc_hd__a2111o_1
Xhold900 _7345_/Q VGND VGND VPWR VPWR hold900/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold911 _5839_/X VGND VGND VPWR VPWR _7433_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7384_ _7568_/CLK _7384_/D fanout622/X VGND VGND VPWR VPWR _7384_/Q sky130_fd_sc_hd__dfrtp_4
Xhold922 _7184_/Q VGND VGND VPWR VPWR hold922/X sky130_fd_sc_hd__dlygate4sd3_1
X_4596_ _4884_/A _4597_/B _4597_/C _5143_/A VGND VGND VPWR VPWR _5375_/A sky130_fd_sc_hd__and4b_4
Xhold933 hold933/A VGND VGND VPWR VPWR hold933/X sky130_fd_sc_hd__dlygate4sd3_1
X_6335_ _7239_/Q _6359_/B _6407_/A3 _6133_/X _7121_/Q VGND VGND VPWR VPWR _6335_/X
+ sky130_fd_sc_hd__a32o_1
Xhold944 _5990_/X VGND VGND VPWR VPWR _7567_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3547_ hold34/X hold61/A hold53/A _3547_/D VGND VGND VPWR VPWR hold35/A sky130_fd_sc_hd__nor4_1
Xhold955 _7503_/Q VGND VGND VPWR VPWR hold955/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 hold966/A VGND VGND VPWR VPWR hold966/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold977 hold977/A VGND VGND VPWR VPWR hold977/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold988 hold988/A VGND VGND VPWR VPWR hold988/X sky130_fd_sc_hd__dlygate4sd3_1
X_3478_ _6912_/Q _3500_/C VGND VGND VPWR VPWR _3478_/X sky130_fd_sc_hd__and2_1
Xhold999 _7001_/Q VGND VGND VPWR VPWR hold999/X sky130_fd_sc_hd__dlygate4sd3_1
X_6266_ _7495_/Q _6309_/B _6407_/A3 _6145_/X _7463_/Q VGND VGND VPWR VPWR _6266_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_142_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5217_ _5614_/B _5614_/D _5195_/X _4985_/B _5092_/B VGND VGND VPWR VPWR _5217_/X
+ sky130_fd_sc_hd__a32o_1
Xhold1600 _6964_/Q VGND VGND VPWR VPWR _4210_/C sky130_fd_sc_hd__dlygate4sd3_1
X_6197_ _7556_/Q _6309_/B _6432_/A3 _6157_/X _7500_/Q VGND VGND VPWR VPWR _6197_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_130_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1611 _6923_/Q VGND VGND VPWR VPWR _4090_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1622 _7644_/Q VGND VGND VPWR VPWR _6321_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1633 _6916_/Q VGND VGND VPWR VPWR hold1633/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5148_ _4795_/Y _4821_/Y _4993_/Y _6858_/C VGND VGND VPWR VPWR _5148_/X sky130_fd_sc_hd__o31a_1
Xhold1644 _6984_/Q VGND VGND VPWR VPWR _4236_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1655 _7619_/Q VGND VGND VPWR VPWR _6053_/B sky130_fd_sc_hd__dlygate4sd3_1
X_5079_ _5079_/A _5079_/B VGND VGND VPWR VPWR _5079_/Y sky130_fd_sc_hd__nor2_1
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4450_ _6820_/A0 _4450_/A1 _4453_/S VGND VGND VPWR VPWR _7147_/D sky130_fd_sc_hd__mux2_1
Xhold207 _7324_/Q VGND VGND VPWR VPWR hold207/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_156_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold218 _7390_/Q VGND VGND VPWR VPWR hold218/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold229 _7334_/Q VGND VGND VPWR VPWR hold229/X sky130_fd_sc_hd__dlygate4sd3_1
X_4381_ hold561/X _4564_/A1 _4381_/S VGND VGND VPWR VPWR _4381_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6120_ _7624_/Q _7623_/Q _6231_/B VGND VGND VPWR VPWR _6159_/A sky130_fd_sc_hd__and3_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6051_ _6811_/S _4130_/B _7142_/Q _6053_/A VGND VGND VPWR VPWR _6064_/A sky130_fd_sc_hd__a211o_1
XFILLER_140_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _5311_/C _5002_/B _5092_/B VGND VGND VPWR VPWR _5002_/X sky130_fd_sc_hd__and3_1
XFILLER_66_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6953_ _6953_/CLK _6953_/D _3473_/X VGND VGND VPWR VPWR _6953_/Q sky130_fd_sc_hd__dfstp_2
X_5904_ hold368/X _6039_/A1 _5911_/S VGND VGND VPWR VPWR _5904_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6884_ _6899_/A _6907_/B VGND VGND VPWR VPWR _6884_/X sky130_fd_sc_hd__and2_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5835_ _5835_/A0 _6006_/A1 _5839_/S VGND VGND VPWR VPWR _5835_/X sky130_fd_sc_hd__mux2_1
XFILLER_167_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5766_ hold621/X _5991_/A1 _5767_/S VGND VGND VPWR VPWR _5766_/X sky130_fd_sc_hd__mux2_1
X_7505_ _7617_/CLK _7505_/D fanout624/X VGND VGND VPWR VPWR _7505_/Q sky130_fd_sc_hd__dfrtp_2
X_4717_ _4747_/B _5297_/A _5595_/B _5358_/B VGND VGND VPWR VPWR _5156_/A sky130_fd_sc_hd__nand4_1
XFILLER_175_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5697_ _5697_/A0 _5697_/A1 _5703_/S VGND VGND VPWR VPWR _5697_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7436_ _7566_/CLK _7436_/D fanout621/X VGND VGND VPWR VPWR _7436_/Q sky130_fd_sc_hd__dfrtp_4
X_4648_ _5595_/A _5476_/A VGND VGND VPWR VPWR _4648_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold730 _4390_/X VGND VGND VPWR VPWR _7092_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 _4218_/X VGND VGND VPWR VPWR _6973_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7367_ _7599_/CLK _7367_/D fanout630/X VGND VGND VPWR VPWR _7367_/Q sky130_fd_sc_hd__dfrtp_1
X_4579_ _4579_/A _4579_/B VGND VGND VPWR VPWR _4781_/C sky130_fd_sc_hd__nor2_2
XFILLER_190_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold752 hold752/A VGND VGND VPWR VPWR hold752/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold763 _7600_/Q VGND VGND VPWR VPWR hold763/X sky130_fd_sc_hd__dlygate4sd3_1
X_6318_ _6082_/B _6304_/X _6317_/X VGND VGND VPWR VPWR _6318_/X sky130_fd_sc_hd__a21o_1
Xmax_cap482 _6212_/C1 VGND VGND VPWR VPWR _6180_/A2 sky130_fd_sc_hd__clkbuf_2
Xhold774 _5757_/X VGND VGND VPWR VPWR _7360_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 hold785/A VGND VGND VPWR VPWR wb_dat_o[20] sky130_fd_sc_hd__buf_12
Xmax_cap493 _5007_/Y VGND VGND VPWR VPWR _5042_/C sky130_fd_sc_hd__clkbuf_2
X_7298_ _7462_/CLK _7298_/D fanout604/X VGND VGND VPWR VPWR _7298_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold796 _7102_/Q VGND VGND VPWR VPWR hold796/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6249_ _6309_/B _6238_/X _6244_/X _6248_/X VGND VGND VPWR VPWR _6249_/X sky130_fd_sc_hd__a211o_1
XFILLER_77_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1430 _7453_/Q VGND VGND VPWR VPWR hold644/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1441 _5724_/X VGND VGND VPWR VPWR _7330_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1452 _5718_/X VGND VGND VPWR VPWR _7325_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1463 _5751_/X VGND VGND VPWR VPWR _7354_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1474 _7637_/Q VGND VGND VPWR VPWR _6163_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_61_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7541_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1485 _7206_/Q VGND VGND VPWR VPWR hold1485/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1496 _7153_/Q VGND VGND VPWR VPWR _4457_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_603 _6427_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_614 _4493_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_625 _3589_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_636 _5884_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_647 _6137_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_658 _6454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_669 _7232_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_76_csclk _7095_/CLK VGND VGND VPWR VPWR _7233_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_14_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7242_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_136_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold90 hold90/A VGND VGND VPWR VPWR hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_29_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7430_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_152_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3950_ _7052_/Q _5680_/B _5678_/B _7475_/Q _3563_/X VGND VGND VPWR VPWR _3950_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_51_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3881_ _7295_/Q _3843_/X _3878_/X _3879_/X _3880_/X VGND VGND VPWR VPWR _3881_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_189_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5620_ _4873_/Y _5381_/X _5619_/X _5259_/A _5259_/B VGND VGND VPWR VPWR _5621_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5551_ _5551_/A1 _5318_/B _5182_/B _4797_/X _5550_/Y VGND VGND VPWR VPWR _5552_/C
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_157_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4502_ _5789_/A1 hold369/X _4504_/S VGND VGND VPWR VPWR _4502_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5482_ _5297_/A _5595_/C _4801_/C _5595_/A _5595_/D VGND VGND VPWR VPWR _5547_/B
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7221_ _7686_/CLK _7221_/D fanout599/X VGND VGND VPWR VPWR _7221_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_105_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4433_ _4433_/A0 _6864_/A1 _4435_/S VGND VGND VPWR VPWR _7128_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7152_ _7668_/CLK _7152_/D VGND VGND VPWR VPWR _7152_/Q sky130_fd_sc_hd__dfxtp_1
X_4364_ _4547_/A hold98/X _5680_/C VGND VGND VPWR VPWR _4369_/S sky130_fd_sc_hd__and3_2
XFILLER_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout517 hold84/X VGND VGND VPWR VPWR hold85/A sky130_fd_sc_hd__buf_8
X_6103_ _6103_/A1 _6065_/Y _6102_/X _6103_/B2 VGND VGND VPWR VPWR _7633_/D sky130_fd_sc_hd__a22o_1
Xfanout528 hold8/X VGND VGND VPWR VPWR hold9/A sky130_fd_sc_hd__buf_6
XFILLER_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout539 hold5/X VGND VGND VPWR VPWR _5869_/A1 sky130_fd_sc_hd__buf_8
XFILLER_59_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7083_ _7207_/CLK _7083_/D fanout616/X VGND VGND VPWR VPWR _7083_/Q sky130_fd_sc_hd__dfstp_2
X_4295_ _4295_/A _4481_/A _6029_/B VGND VGND VPWR VPWR _4303_/S sky130_fd_sc_hd__and3_4
XFILLER_113_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6034_ _6043_/A1 hold249/X _6037_/S VGND VGND VPWR VPWR _6034_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6936_ _4172_/B2 _6936_/D _6891_/X VGND VGND VPWR VPWR hold83/A sky130_fd_sc_hd__dfrtp_1
XFILLER_35_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6867_ _6899_/A _6911_/B VGND VGND VPWR VPWR _6867_/X sky130_fd_sc_hd__and2_1
XFILLER_179_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5818_ _5935_/A1 hold211/X _5821_/S VGND VGND VPWR VPWR _5818_/X sky130_fd_sc_hd__mux2_1
X_6798_ _7125_/Q _6441_/X _6482_/X _7115_/Q VGND VGND VPWR VPWR _6798_/X sky130_fd_sc_hd__a22o_1
XFILLER_41_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5749_ _6046_/A1 hold916/X _5749_/S VGND VGND VPWR VPWR _5749_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7419_ _7553_/CLK _7419_/D fanout624/X VGND VGND VPWR VPWR _7419_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_163_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold560 _6000_/X VGND VGND VPWR VPWR _7576_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold571 _7035_/Q VGND VGND VPWR VPWR hold571/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold582 _5694_/X VGND VGND VPWR VPWR _7304_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_173_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold593 hold593/A VGND VGND VPWR VPWR hold593/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1260 _7366_/Q VGND VGND VPWR VPWR hold288/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1271 _5889_/X VGND VGND VPWR VPWR _7477_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1282 _7673_/Q VGND VGND VPWR VPWR _6835_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1293 _7105_/Q VGND VGND VPWR VPWR hold549/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_400 _3838_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_411 _5938_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_422 _6158_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_433 _6192_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_444 _6451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_455 _6468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_466 _7040_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_477 _7232_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_488 _7162_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_499 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4080_ _4064_/B _4192_/C _4193_/B _6913_/Q VGND VGND VPWR VPWR _4080_/X sky130_fd_sc_hd__and4b_1
XFILLER_110_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4982_ _5322_/C _4995_/A VGND VGND VPWR VPWR _4982_/Y sky130_fd_sc_hd__nand2_2
X_6721_ _7205_/Q _6099_/B _6720_/D _6452_/X _7185_/Q VGND VGND VPWR VPWR _6721_/X
+ sky130_fd_sc_hd__a32o_1
X_3933_ _7235_/Q _5628_/A _4553_/B _3715_/X _7107_/Q VGND VGND VPWR VPWR _3933_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_189_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6652_ _7560_/Q _6453_/X _6485_/X _7552_/Q _6638_/X VGND VGND VPWR VPWR _6652_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3864_ _7043_/Q _4529_/B _6038_/B _3574_/X input22/X VGND VGND VPWR VPWR _3864_/X
+ sky130_fd_sc_hd__a32o_4
X_5603_ _5603_/A _5603_/B _5603_/C _5603_/D VGND VGND VPWR VPWR _5603_/Y sky130_fd_sc_hd__nand4_1
XFILLER_118_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6583_ _7325_/Q _6471_/X _6565_/X _6574_/X _6582_/X VGND VGND VPWR VPWR _6583_/X
+ sky130_fd_sc_hd__a2111o_4
X_3795_ _7405_/Q _3545_/X _3790_/X _3791_/X _3794_/X VGND VGND VPWR VPWR _3795_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_117_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5534_ _5534_/A _5534_/B _5534_/C VGND VGND VPWR VPWR _5618_/A sky130_fd_sc_hd__and3_1
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5465_ _5339_/X _5011_/A _5202_/Y _5464_/X VGND VGND VPWR VPWR _5586_/B sky130_fd_sc_hd__o211a_1
XFILLER_172_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7204_ _7207_/CLK _7204_/D fanout616/X VGND VGND VPWR VPWR _7204_/Q sky130_fd_sc_hd__dfrtp_1
X_4416_ hold426/X _5673_/A1 _4417_/S VGND VGND VPWR VPWR _4416_/X sky130_fd_sc_hd__mux2_1
X_5396_ _4811_/Y _4871_/X _4910_/Y _5121_/D _5527_/B VGND VGND VPWR VPWR _5399_/C
+ sky130_fd_sc_hd__o311a_1
X_7135_ _7286_/CLK _7135_/D fanout598/X VGND VGND VPWR VPWR _7135_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_99_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4347_ _6012_/A0 _4347_/A1 _4351_/S VGND VGND VPWR VPWR _4347_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7066_ _7212_/CLK _7066_/D fanout619/X VGND VGND VPWR VPWR _7066_/Q sky130_fd_sc_hd__dfrtp_2
X_4278_ _4293_/S _4240_/X _4277_/Y _6038_/C VGND VGND VPWR VPWR _4294_/S sky130_fd_sc_hd__o211ai_4
XFILLER_101_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6017_ _6044_/A1 hold871/X _6019_/S VGND VGND VPWR VPWR _6017_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_wbbd_sck clkbuf_0_wbbd_sck/X VGND VGND VPWR VPWR _6854_/A sky130_fd_sc_hd__clkbuf_16
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6919_ _7258_/CLK _6919_/D _6874_/X VGND VGND VPWR VPWR _6919_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold390 _4492_/X VGND VGND VPWR VPWR _7183_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1090 _5952_/X VGND VGND VPWR VPWR _7533_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_230 _6922_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_241 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_252 _4199_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_263 _4196_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_274 input81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_285 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_296 input95/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3580_ _3713_/A _3905_/B _4481_/A VGND VGND VPWR VPWR _3580_/X sky130_fd_sc_hd__and3_4
XFILLER_173_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_586 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5250_ _5189_/A _4992_/B _5404_/A _5311_/A VGND VGND VPWR VPWR _5250_/X sky130_fd_sc_hd__a31o_1
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4201_ _4202_/A _4201_/B VGND VGND VPWR VPWR _6964_/D sky130_fd_sc_hd__and2_1
XFILLER_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5181_ _5375_/A _5375_/B _5181_/C VGND VGND VPWR VPWR _5182_/B sky130_fd_sc_hd__and3_1
X_4132_ _6791_/B _6694_/B _4130_/Y _4121_/Y _4132_/B2 VGND VGND VPWR VPWR _7142_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_96_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4063_ _6927_/Q hold94/A _6925_/Q hold21/A VGND VGND VPWR VPWR _4064_/B sky130_fd_sc_hd__and4_1
XFILLER_96_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4965_ _5476_/A _4966_/A _4966_/B VGND VGND VPWR VPWR _4968_/A sky130_fd_sc_hd__and3_1
X_6704_ _7061_/Q _6453_/X _6484_/X _7091_/Q _6703_/X VGND VGND VPWR VPWR _6709_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3916_ _7531_/Q _5984_/A _6020_/A _3573_/C _5723_/A VGND VGND VPWR VPWR _3916_/X
+ sky130_fd_sc_hd__a32o_1
X_7684_ _7686_/CLK _7684_/D fanout600/X VGND VGND VPWR VPWR _7684_/Q sky130_fd_sc_hd__dfstp_1
X_4896_ _4943_/A _4901_/B _4896_/C _4950_/C VGND VGND VPWR VPWR _4900_/B sky130_fd_sc_hd__nand4_1
X_6635_ _6634_/Y _6633_/X _7654_/Q _6686_/S VGND VGND VPWR VPWR _6635_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_137_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3847_ _7083_/Q _4559_/B _5680_/A _3562_/X _7500_/Q VGND VGND VPWR VPWR _3847_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_22_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6566_ hold87/A _6447_/X _6474_/C _7373_/Q _6564_/X VGND VGND VPWR VPWR _6566_/X
+ sky130_fd_sc_hd__a221o_1
X_3778_ _6945_/Q _3777_/X _3904_/S VGND VGND VPWR VPWR _6946_/D sky130_fd_sc_hd__mux2_1
XFILLER_138_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5517_ _5318_/B _5517_/A2 _5143_/X _5311_/A VGND VGND VPWR VPWR _5517_/X sky130_fd_sc_hd__a22o_1
XFILLER_145_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6497_ _7338_/Q _6474_/A _6494_/X _6496_/X VGND VGND VPWR VPWR _6497_/X sky130_fd_sc_hd__a211o_1
XFILLER_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5448_ _4867_/X _4912_/Y _4998_/Y _5440_/Y _5260_/B VGND VGND VPWR VPWR _5527_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_154_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5379_ _5102_/B _5404_/C _4817_/Y _5189_/Y _4613_/X VGND VGND VPWR VPWR _5555_/B
+ sky130_fd_sc_hd__o311a_1
X_7118_ _7242_/CLK _7118_/D fanout616/X VGND VGND VPWR VPWR _7118_/Q sky130_fd_sc_hd__dfstp_2
X_7049_ _7289_/CLK _7049_/D fanout598/X VGND VGND VPWR VPWR _7049_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_87_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4750_ _4836_/A _4694_/Y _4693_/Y _5027_/C VGND VGND VPWR VPWR _4750_/Y sky130_fd_sc_hd__o211ai_4
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3701_ _3713_/A _6861_/A _5659_/C VGND VGND VPWR VPWR _3701_/X sky130_fd_sc_hd__and3_4
XFILLER_119_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4681_ _4747_/B _4801_/C VGND VGND VPWR VPWR _4681_/Y sky130_fd_sc_hd__nand2_2
X_6420_ _7173_/Q _6160_/D _6166_/C _6419_/X VGND VGND VPWR VPWR _6420_/X sky130_fd_sc_hd__a31o_1
X_3632_ _7600_/Q _3569_/X _6029_/A _7608_/Q _3631_/X VGND VGND VPWR VPWR _3632_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_146_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6351_ _7180_/Q wire452/X _6346_/X _6359_/B _6350_/X VGND VGND VPWR VPWR _6351_/X
+ sky130_fd_sc_hd__a2111o_1
X_3563_ _3714_/A hold74/A _5957_/B VGND VGND VPWR VPWR _3563_/X sky130_fd_sc_hd__and3_1
XFILLER_127_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5302_ _5094_/D _5293_/X _5291_/X _5301_/X VGND VGND VPWR VPWR _5302_/X sky130_fd_sc_hd__a211o_1
X_6282_ _7528_/Q _6309_/B _6334_/C _6136_/X _7512_/Q VGND VGND VPWR VPWR _6282_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_142_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3494_ hold153/X _6929_/Q _3508_/S VGND VGND VPWR VPWR _3494_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5233_ _5233_/A _5233_/B _5233_/C VGND VGND VPWR VPWR _5233_/X sky130_fd_sc_hd__and3_1
XFILLER_130_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5164_ _4660_/C _4728_/Y _4912_/Y _4685_/Y _5162_/Y VGND VGND VPWR VPWR _5164_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_124_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4115_ _5143_/A _4115_/B _4115_/C _4115_/D VGND VGND VPWR VPWR _4117_/C sky130_fd_sc_hd__and4_1
XFILLER_69_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5095_ _5291_/C _5130_/B _5095_/C VGND VGND VPWR VPWR _5095_/X sky130_fd_sc_hd__and3_1
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4046_ _4046_/A0 _4099_/A0 _4049_/B VGND VGND VPWR VPWR _6941_/D sky130_fd_sc_hd__mux2_1
XFILLER_24_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5997_ _5997_/A0 _6042_/A1 _6001_/S VGND VGND VPWR VPWR _7573_/D sky130_fd_sc_hd__mux2_1
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4948_ _4948_/A _4948_/B _4959_/C _5429_/D VGND VGND VPWR VPWR _4948_/Y sky130_fd_sc_hd__nor4_2
X_7667_ _7672_/CLK _7667_/D VGND VGND VPWR VPWR _7667_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4879_ _4953_/A _4953_/C _4953_/D _4878_/X _4900_/A VGND VGND VPWR VPWR _4879_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_177_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6618_ _7615_/Q _6451_/X _6482_/X _7487_/Q _6617_/X VGND VGND VPWR VPWR _6623_/B
+ sky130_fd_sc_hd__a221o_1
X_7598_ _7603_/CLK _7598_/D fanout612/X VGND VGND VPWR VPWR _7598_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6549_ _7532_/Q _6720_/C _6536_/C _6460_/X _7444_/Q VGND VGND VPWR VPWR _6549_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput270 _7268_/Q VGND VGND VPWR VPWR pll_sel[2] sky130_fd_sc_hd__buf_12
Xoutput281 _7275_/Q VGND VGND VPWR VPWR pll_trim[19] sky130_fd_sc_hd__buf_12
Xoutput292 _6977_/Q VGND VGND VPWR VPWR pll_trim[5] sky130_fd_sc_hd__buf_12
XFILLER_181_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire353 _3816_/Y VGND VGND VPWR VPWR _3838_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_128_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire375 _6478_/Y VGND VGND VPWR VPWR _6759_/D sky130_fd_sc_hd__buf_8
XFILLER_109_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5920_ hold906/X _6046_/A1 _5920_/S VGND VGND VPWR VPWR _5920_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5851_ _6040_/A1 hold983/X _5857_/S VGND VGND VPWR VPWR _7443_/D sky130_fd_sc_hd__mux2_1
XFILLER_34_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4802_ _4775_/Y _4798_/Y _4801_/X VGND VGND VPWR VPWR _4808_/A sky130_fd_sc_hd__a21oi_1
X_5782_ _5926_/A0 hold281/X _5785_/S VGND VGND VPWR VPWR _5782_/X sky130_fd_sc_hd__mux2_1
X_7521_ _7609_/CLK _7521_/D fanout614/X VGND VGND VPWR VPWR _7521_/Q sky130_fd_sc_hd__dfrtp_1
X_4733_ _4733_/A _4733_/B _4733_/C VGND VGND VPWR VPWR _4735_/A sky130_fd_sc_hd__nor3_1
XFILLER_159_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7452_ _7616_/CLK hold82/X fanout610/X VGND VGND VPWR VPWR _7452_/Q sky130_fd_sc_hd__dfrtp_2
X_4664_ _5000_/C _4836_/A _4660_/C _4688_/B _5007_/D VGND VGND VPWR VPWR _5614_/B
+ sky130_fd_sc_hd__o311a_4
XFILLER_174_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6403_ _7064_/Q _6158_/D _6432_/A3 _6146_/X _7084_/Q VGND VGND VPWR VPWR _6403_/X
+ sky130_fd_sc_hd__a32o_1
X_3615_ _7337_/Q _5939_/B _5759_/B _3571_/X _7361_/Q VGND VGND VPWR VPWR _3615_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_175_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7383_ _7421_/CLK _7383_/D fanout630/X VGND VGND VPWR VPWR _7383_/Q sky130_fd_sc_hd__dfrtp_1
Xhold901 _5740_/X VGND VGND VPWR VPWR _7345_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4595_ _5143_/B _4595_/B VGND VGND VPWR VPWR _4595_/Y sky130_fd_sc_hd__nor2_2
Xhold912 _7585_/Q VGND VGND VPWR VPWR hold912/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold923 _4494_/X VGND VGND VPWR VPWR _7184_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6334_ _7071_/Q _6359_/B _6334_/C VGND VGND VPWR VPWR _6334_/X sky130_fd_sc_hd__and3_1
Xhold934 hold934/A VGND VGND VPWR VPWR hold934/X sky130_fd_sc_hd__dlygate4sd3_1
X_3546_ _3714_/A _5686_/A _3546_/C VGND VGND VPWR VPWR _3546_/X sky130_fd_sc_hd__and3_4
Xhold945 _7447_/Q VGND VGND VPWR VPWR hold945/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold956 _5918_/X VGND VGND VPWR VPWR _7503_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold967 hold967/A VGND VGND VPWR VPWR hold967/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold978 hold978/A VGND VGND VPWR VPWR hold978/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6265_ _7511_/Q _6428_/A2 _6428_/B1 _7543_/Q _6264_/X VGND VGND VPWR VPWR _6265_/X
+ sky130_fd_sc_hd__a221o_1
Xhold989 _7002_/Q VGND VGND VPWR VPWR hold989/X sky130_fd_sc_hd__dlygate4sd3_1
X_3477_ _6914_/Q _6913_/Q VGND VGND VPWR VPWR _3500_/C sky130_fd_sc_hd__nor2_4
XFILLER_135_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5216_ _4625_/Y _5585_/A1 _5212_/Y _5001_/Y _4984_/Y VGND VGND VPWR VPWR _5216_/X
+ sky130_fd_sc_hd__o32a_1
X_6196_ _7476_/Q _6309_/B _6286_/C _6195_/X VGND VGND VPWR VPWR _6196_/X sky130_fd_sc_hd__a31o_1
Xhold1601 _7618_/Q VGND VGND VPWR VPWR _6049_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1612 _6939_/Q VGND VGND VPWR VPWR _4054_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1623 _7679_/Q VGND VGND VPWR VPWR _6853_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5147_ _5147_/A _5147_/B _5147_/C VGND VGND VPWR VPWR _5147_/Y sky130_fd_sc_hd__nand3_1
Xhold1634 _6972_/Q VGND VGND VPWR VPWR hold1634/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1645 _6967_/Q VGND VGND VPWR VPWR _4201_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1656 _7629_/Q VGND VGND VPWR VPWR _6090_/A3 sky130_fd_sc_hd__dlygate4sd3_1
X_5078_ _5322_/A _5021_/A _5401_/A _5077_/X VGND VGND VPWR VPWR _5079_/B sky130_fd_sc_hd__a31o_1
XFILLER_178_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4029_ _7111_/Q _4559_/B _4529_/B _5678_/B _5669_/B VGND VGND VPWR VPWR _4029_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_44_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold208 _5717_/X VGND VGND VPWR VPWR _7324_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold219 _5791_/X VGND VGND VPWR VPWR _7390_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4380_ hold815/X _5988_/A1 _4381_/S VGND VGND VPWR VPWR _4380_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ _7142_/Q _6811_/S _6109_/B _4140_/Y VGND VGND VPWR VPWR _6053_/A sky130_fd_sc_hd__o31ai_2
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ _5109_/A _5131_/B VGND VGND VPWR VPWR _5001_/Y sky130_fd_sc_hd__nand2_4
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6952_ _4172_/B2 _6952_/D _6907_/X VGND VGND VPWR VPWR hold27/A sky130_fd_sc_hd__dfrtn_1
X_5903_ _5903_/A _5975_/B _6038_/C VGND VGND VPWR VPWR _5911_/S sky130_fd_sc_hd__and3_4
X_6883_ _6899_/A _6908_/B VGND VGND VPWR VPWR _6883_/X sky130_fd_sc_hd__and2_1
XFILLER_179_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5834_ hold269/X _5843_/A1 _5839_/S VGND VGND VPWR VPWR _5834_/X sky130_fd_sc_hd__mux2_1
X_5765_ hold875/X _6044_/A1 _5767_/S VGND VGND VPWR VPWR _5765_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4716_ _4738_/A _5476_/A _4740_/D _5358_/B VGND VGND VPWR VPWR _4721_/B sky130_fd_sc_hd__nand4_1
X_7504_ _7568_/CLK _7504_/D fanout622/X VGND VGND VPWR VPWR _7504_/Q sky130_fd_sc_hd__dfrtp_4
X_5696_ _7294_/Q _4171_/C _4171_/D _4293_/S _6038_/C VGND VGND VPWR VPWR _5696_/Y
+ sky130_fd_sc_hd__o311ai_4
X_7435_ _7435_/CLK _7435_/D fanout623/X VGND VGND VPWR VPWR _7435_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_175_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4647_ _5476_/A _5195_/B _5476_/B VGND VGND VPWR VPWR _4761_/A sky130_fd_sc_hd__and3_4
XFILLER_107_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold720 _4414_/X VGND VGND VPWR VPWR _7112_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7366_ _7597_/CLK _7366_/D fanout626/X VGND VGND VPWR VPWR _7366_/Q sky130_fd_sc_hd__dfrtp_4
X_4578_ _4585_/C _4585_/D _4584_/A _4584_/B VGND VGND VPWR VPWR _4579_/B sky130_fd_sc_hd__nand4_1
Xhold731 _7127_/Q VGND VGND VPWR VPWR hold731/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold742 _7230_/Q VGND VGND VPWR VPWR hold742/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold753 _7548_/Q VGND VGND VPWR VPWR hold753/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 _6027_/X VGND VGND VPWR VPWR _7600_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6317_ _6307_/X _6131_/B _6306_/X _6308_/X _6316_/X VGND VGND VPWR VPWR _6317_/X
+ sky130_fd_sc_hd__a2111o_1
X_3529_ _3622_/A _3717_/B hold23/X VGND VGND VPWR VPWR _3529_/X sky130_fd_sc_hd__and3_4
Xmax_cap483 wire484/X VGND VGND VPWR VPWR _6212_/C1 sky130_fd_sc_hd__clkbuf_2
X_7297_ _7497_/CLK _7297_/D fanout607/X VGND VGND VPWR VPWR _7297_/Q sky130_fd_sc_hd__dfrtp_2
Xhold775 _7095_/Q VGND VGND VPWR VPWR hold775/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap494 _5290_/A2 VGND VGND VPWR VPWR _5088_/B sky130_fd_sc_hd__clkbuf_2
Xhold786 _7192_/Q VGND VGND VPWR VPWR hold786/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 _4402_/X VGND VGND VPWR VPWR _7102_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6248_ _7366_/Q _6152_/X _6153_/X _7566_/Q _6247_/X VGND VGND VPWR VPWR _6248_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6179_ _7555_/Q _6131_/B _6432_/A3 _6160_/X _7371_/Q VGND VGND VPWR VPWR _6179_/X
+ sky130_fd_sc_hd__a32o_1
Xhold1420 _7458_/Q VGND VGND VPWR VPWR hold296/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1431 _7474_/Q VGND VGND VPWR VPWR hold280/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1442 _6987_/Q VGND VGND VPWR VPWR _4239_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1453 _7667_/Q VGND VGND VPWR VPWR _6819_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1464 _7144_/Q VGND VGND VPWR VPWR _4447_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1475 _6981_/Q VGND VGND VPWR VPWR _4233_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1486 _4520_/X VGND VGND VPWR VPWR _7206_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1497 _7490_/Q VGND VGND VPWR VPWR hold368/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_604 _6166_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_615 _4493_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_626 _4019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_637 _6131_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_648 _6137_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_659 _6464_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold80 hold80/A VGND VGND VPWR VPWR hold80/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 hold91/A VGND VGND VPWR VPWR hold91/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3880_ _7508_/Q _5903_/A _5993_/B _3573_/X input5/X VGND VGND VPWR VPWR _3880_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_188_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5550_ _4597_/Y _4769_/Y _4772_/Y _5180_/C _4775_/D VGND VGND VPWR VPWR _5550_/Y
+ sky130_fd_sc_hd__o311ai_1
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4501_ _5761_/A1 hold381/X _4504_/S VGND VGND VPWR VPWR _4501_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5481_ _4629_/Y _4709_/Y _4811_/Y _4692_/Y VGND VGND VPWR VPWR _5547_/C sky130_fd_sc_hd__a31o_1
X_7220_ _7233_/CLK _7220_/D fanout599/X VGND VGND VPWR VPWR _7220_/Q sky130_fd_sc_hd__dfrtp_4
X_4432_ hold731/X _6863_/A1 _4435_/S VGND VGND VPWR VPWR _4432_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7151_ _7668_/CLK _7151_/D VGND VGND VPWR VPWR _7151_/Q sky130_fd_sc_hd__dfxtp_1
X_4363_ _5926_/A0 hold379/X _4363_/S VGND VGND VPWR VPWR _4363_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout507 _4569_/X VGND VGND VPWR VPWR _4943_/A sky130_fd_sc_hd__buf_8
X_6102_ _6099_/B _6563_/C _6099_/Y _7633_/Q VGND VGND VPWR VPWR _6102_/X sky130_fd_sc_hd__a22o_1
Xfanout518 hold19/X VGND VGND VPWR VPWR _6866_/A1 sky130_fd_sc_hd__buf_6
XFILLER_112_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout529 _4556_/A1 VGND VGND VPWR VPWR _6864_/A1 sky130_fd_sc_hd__buf_6
X_7082_ _7130_/CLK _7082_/D fanout602/X VGND VGND VPWR VPWR _7082_/Q sky130_fd_sc_hd__dfrtp_4
X_4294_ _4293_/X _4294_/A1 _4294_/S VGND VGND VPWR VPWR _4294_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6033_ _6042_/A1 _6033_/A1 _6037_/S VGND VGND VPWR VPWR _6033_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6935_ _6950_/CLK _6935_/D _6890_/X VGND VGND VPWR VPWR _6935_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6866_ hold182/X _6866_/A1 _6866_/S VGND VGND VPWR VPWR _6866_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5817_ _6006_/A1 hold892/X _5821_/S VGND VGND VPWR VPWR _5817_/X sky130_fd_sc_hd__mux2_1
X_6797_ _7168_/Q _6469_/X _6485_/X _7218_/Q _6796_/X VGND VGND VPWR VPWR _6800_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_167_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5748_ _5991_/A1 _5748_/A1 _5749_/S VGND VGND VPWR VPWR _5748_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5679_ _5679_/A1 _3623_/X _5680_/C _5678_/Y VGND VGND VPWR VPWR _5679_/X sky130_fd_sc_hd__o211a_1
XFILLER_135_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7418_ _7586_/CLK _7418_/D fanout625/X VGND VGND VPWR VPWR _7418_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_190_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold550 _7130_/Q VGND VGND VPWR VPWR hold550/X sky130_fd_sc_hd__dlygate4sd3_1
X_7349_ _7599_/CLK _7349_/D fanout628/X VGND VGND VPWR VPWR _7349_/Q sky130_fd_sc_hd__dfrtp_4
Xhold561 _7085_/Q VGND VGND VPWR VPWR hold561/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 _4321_/X VGND VGND VPWR VPWR _7035_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold583 _7544_/Q VGND VGND VPWR VPWR hold583/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold594 hold594/A VGND VGND VPWR VPWR hold594/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1250 _7351_/Q VGND VGND VPWR VPWR hold928/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1261 _5764_/X VGND VGND VPWR VPWR _7366_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1272 _7281_/Q VGND VGND VPWR VPWR hold298/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1283 _5824_/X VGND VGND VPWR VPWR _7419_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_401 _3957_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1294 _4405_/X VGND VGND VPWR VPWR _7105_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_412 _5938_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_423 _6158_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_434 _6341_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_445 _6451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_456 _6478_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_467 _7224_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_478 _7232_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_489 _7610_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput170 wb_we_i VGND VGND VPWR VPWR _6827_/A sky130_fd_sc_hd__buf_2
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4981_ _5146_/A _5146_/B _5311_/C VGND VGND VPWR VPWR _4981_/X sky130_fd_sc_hd__and3_2
XFILLER_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6720_ _7102_/Q _6791_/C _6720_/C _6720_/D VGND VGND VPWR VPWR _6720_/X sky130_fd_sc_hd__and4_1
X_3932_ _7371_/Q _3572_/X _3927_/X _3929_/X _3931_/X VGND VGND VPWR VPWR _3932_/Y
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_149_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6651_ _6651_/A _6651_/B _6651_/C VGND VGND VPWR VPWR _6651_/Y sky130_fd_sc_hd__nor3_4
X_3863_ _7548_/Q _3514_/X _3849_/X _3853_/X _3862_/X VGND VGND VPWR VPWR _3863_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_177_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5602_ _5602_/A _5602_/B _5602_/C _5602_/D VGND VGND VPWR VPWR _5603_/D sky130_fd_sc_hd__nor4_1
X_6582_ _7597_/Q _6474_/B _6578_/X _6581_/X _6477_/X VGND VGND VPWR VPWR _6582_/X
+ sky130_fd_sc_hd__a2111o_1
X_3794_ _7429_/Q _3556_/X _3792_/X _3793_/X VGND VGND VPWR VPWR _3794_/X sky130_fd_sc_hd__a211o_1
XFILLER_192_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5533_ _4994_/X _5111_/D _5027_/X _4761_/A _5532_/X VGND VGND VPWR VPWR _5534_/C
+ sky130_fd_sc_hd__a221oi_1
XFILLER_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_60_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7603_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_133_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5464_ _5011_/A _4674_/Y _5197_/Y _5192_/X _5026_/Y VGND VGND VPWR VPWR _5464_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_105_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7203_ _7207_/CLK _7203_/D fanout616/X VGND VGND VPWR VPWR _7203_/Q sky130_fd_sc_hd__dfrtp_2
X_4415_ _4415_/A0 _6864_/A1 _4417_/S VGND VGND VPWR VPWR _4415_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5395_ _4769_/Y _4953_/C _4871_/X _4910_/Y VGND VGND VPWR VPWR _5527_/B sky130_fd_sc_hd__a211o_1
XFILLER_99_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7134_ _7614_/CLK _7134_/D fanout604/X VGND VGND VPWR VPWR _7134_/Q sky130_fd_sc_hd__dfstp_2
X_4346_ _4346_/A _6861_/C VGND VGND VPWR VPWR _4351_/S sky130_fd_sc_hd__nand2_2
XFILLER_59_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_75_csclk _7095_/CLK VGND VGND VPWR VPWR _7231_/CLK sky130_fd_sc_hd__clkbuf_16
X_7065_ _7217_/CLK _7065_/D _6903_/A VGND VGND VPWR VPWR _7065_/Q sky130_fd_sc_hd__dfrtp_2
X_4277_ _7294_/Q _4171_/C _4171_/D _4505_/B VGND VGND VPWR VPWR _4277_/Y sky130_fd_sc_hd__o31ai_2
X_6016_ _6043_/A1 hold294/X _6019_/S VGND VGND VPWR VPWR _6016_/X sky130_fd_sc_hd__mux2_1
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6918_ _4183_/A1 _6918_/D _6873_/X VGND VGND VPWR VPWR _6918_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_13_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7685_/CLK sky130_fd_sc_hd__clkbuf_16
X_6849_ _6969_/Q _6849_/A2 _6849_/B1 wire537/X _6848_/X VGND VGND VPWR VPWR _6849_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_167_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_28_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7557_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold380 _4363_/X VGND VGND VPWR VPWR _7070_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold391 _7193_/Q VGND VGND VPWR VPWR hold391/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1080 hold1379/X VGND VGND VPWR VPWR _5727_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1091 hold1317/X VGND VGND VPWR VPWR _6006_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_93_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_220 _7534_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_231 _6922_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_242 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_253 _4199_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_264 _7714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_275 input81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_286 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_297 input96/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4200_ _4202_/A _6970_/Q VGND VGND VPWR VPWR _6963_/D sky130_fd_sc_hd__and2_1
XFILLER_142_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5180_ _5180_/A _5552_/A _5180_/C VGND VGND VPWR VPWR _5182_/C sky130_fd_sc_hd__nand3_1
XFILLER_123_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4131_ _7139_/Q _7293_/Q _4130_/Y _4127_/Y VGND VGND VPWR VPWR _7141_/D sky130_fd_sc_hd__a22o_1
XFILLER_110_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4062_ hold94/A _6925_/Q hold21/A VGND VGND VPWR VPWR _4062_/Y sky130_fd_sc_hd__nand3_1
XFILLER_95_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4964_ _4964_/A _4964_/B _5570_/A VGND VGND VPWR VPWR _4968_/C sky130_fd_sc_hd__nand3_1
X_6703_ _7194_/Q _6457_/X _6807_/A2 _7234_/Q VGND VGND VPWR VPWR _6703_/X sky130_fd_sc_hd__a22o_1
XFILLER_189_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3915_ _7603_/Q _5957_/B _6038_/B _3914_/X VGND VGND VPWR VPWR _3915_/X sky130_fd_sc_hd__a31o_1
XFILLER_177_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7683_ _7686_/CLK _7683_/D fanout600/X VGND VGND VPWR VPWR _7683_/Q sky130_fd_sc_hd__dfrtp_2
X_4895_ _5014_/D _4836_/Y _4907_/A _5389_/C VGND VGND VPWR VPWR _4896_/C sky130_fd_sc_hd__o211a_1
X_6634_ _7319_/Q _6759_/D _6686_/S VGND VGND VPWR VPWR _6634_/Y sky130_fd_sc_hd__o21bai_1
X_3846_ input58/X _4293_/S _3701_/X _7241_/Q _3844_/X VGND VGND VPWR VPWR _3846_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_165_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3777_ _4459_/A0 _3777_/A1 _3967_/S VGND VGND VPWR VPWR _3777_/X sky130_fd_sc_hd__mux2_1
X_6565_ _7405_/Q _6466_/X _6501_/X _7565_/Q _6562_/X VGND VGND VPWR VPWR _6565_/X
+ sky130_fd_sc_hd__a221o_1
X_5516_ _5429_/A _5313_/C _5137_/A _5515_/Y VGND VGND VPWR VPWR _5516_/X sky130_fd_sc_hd__a31o_1
X_6496_ _7474_/Q _6441_/X _6445_/X _7362_/Q _6495_/X VGND VGND VPWR VPWR _6496_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5447_ _5621_/A _5447_/B _5524_/C VGND VGND VPWR VPWR _5451_/A sky130_fd_sc_hd__and3_1
XFILLER_160_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5378_ _5555_/D _5378_/B _5555_/C VGND VGND VPWR VPWR _5378_/Y sky130_fd_sc_hd__nand3_1
X_4329_ _4329_/A0 _6862_/A1 _4333_/S VGND VGND VPWR VPWR _4329_/X sky130_fd_sc_hd__mux2_1
X_7117_ _7242_/CLK _7117_/D fanout616/X VGND VGND VPWR VPWR _7117_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7048_ _7289_/CLK _7048_/D fanout598/X VGND VGND VPWR VPWR _7048_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire535 wire535/A VGND VGND VPWR VPWR wire535/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3700_ _4340_/A _5682_/B _4475_/A VGND VGND VPWR VPWR _3700_/X sky130_fd_sc_hd__and3_2
XFILLER_186_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4680_ _5015_/C _4684_/A _4668_/C VGND VGND VPWR VPWR _4680_/X sky130_fd_sc_hd__a21o_1
XFILLER_187_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3631_ _7320_/Q _5993_/B _5682_/C hold56/A _7137_/Q VGND VGND VPWR VPWR _3631_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_174_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6350_ _7235_/Q _6124_/X _6347_/X _6349_/X VGND VGND VPWR VPWR _6350_/X sky130_fd_sc_hd__a211o_1
X_3562_ _3714_/A hold74/A _5984_/B VGND VGND VPWR VPWR _3562_/X sky130_fd_sc_hd__and3_4
XFILLER_127_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5301_ _5291_/C _5294_/X _5295_/X _5296_/X _5300_/X VGND VGND VPWR VPWR _5301_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_127_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6281_ _7384_/Q _6077_/X _6276_/X _6278_/X _6280_/X VGND VGND VPWR VPWR _6281_/X
+ sky130_fd_sc_hd__a2111o_4
X_3493_ hold34/X hold61/X VGND VGND VPWR VPWR _3714_/A sky130_fd_sc_hd__and2b_4
XFILLER_142_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5232_ _5196_/A _5322_/A _5068_/C _5231_/X _5230_/Y VGND VGND VPWR VPWR _5232_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_142_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5163_ _4617_/X _4660_/C _4691_/X _4912_/Y _4685_/Y VGND VGND VPWR VPWR _5163_/Y
+ sky130_fd_sc_hd__o32ai_1
X_4114_ _4884_/A _5096_/A _4586_/A _4586_/B VGND VGND VPWR VPWR _4115_/D sky130_fd_sc_hd__a211oi_1
XFILLER_68_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5094_ _5094_/A _5189_/D _5112_/B _5094_/D VGND VGND VPWR VPWR _5094_/Y sky130_fd_sc_hd__nand4_1
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4045_ _6940_/Q _6939_/Q _4043_/Y _4045_/B1 VGND VGND VPWR VPWR _4045_/X sky130_fd_sc_hd__o31a_1
XFILLER_84_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5996_ hold347/X hold81/X _6001_/S VGND VGND VPWR VPWR _5996_/X sky130_fd_sc_hd__mux2_1
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4947_ _4947_/A _4947_/B VGND VGND VPWR VPWR _4947_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7666_ _7676_/CLK _7666_/D VGND VGND VPWR VPWR _7666_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_130_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4878_ _5000_/C _4777_/Y _4830_/Y _4907_/C _4935_/B VGND VGND VPWR VPWR _4878_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_20_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6617_ _7399_/Q _6463_/X _6474_/C _7375_/Q VGND VGND VPWR VPWR _6617_/X sky130_fd_sc_hd__a22o_1
X_3829_ _7373_/Q _3572_/X _4382_/A _7089_/Q _3828_/X VGND VGND VPWR VPWR _3837_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_165_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7597_ _7597_/CLK _7597_/D fanout626/X VGND VGND VPWR VPWR _7597_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6548_ _7364_/Q _6445_/X _6542_/X _6546_/X _6547_/X VGND VGND VPWR VPWR _6548_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_165_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6479_ _7631_/Q _6485_/B _6563_/C _6791_/D VGND VGND VPWR VPWR _6479_/X sky130_fd_sc_hd__and4_4
XFILLER_121_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput260 _7280_/Q VGND VGND VPWR VPWR pll_bypass sky130_fd_sc_hd__buf_12
XFILLER_121_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput271 _6972_/Q VGND VGND VPWR VPWR pll_trim[0] sky130_fd_sc_hd__buf_12
Xoutput282 _6973_/Q VGND VGND VPWR VPWR pll_trim[1] sky130_fd_sc_hd__buf_12
XFILLER_160_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput293 _6978_/Q VGND VGND VPWR VPWR pll_trim[6] sky130_fd_sc_hd__buf_12
XFILLER_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire354 _3691_/Y VGND VGND VPWR VPWR _3692_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_156_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire365 _4276_/S VGND VGND VPWR VPWR _4274_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_144_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5850_ hold44/X _5850_/A1 _5857_/S VGND VGND VPWR VPWR hold45/A sky130_fd_sc_hd__mux2_1
XFILLER_179_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4801_ _5375_/A _5186_/C _4801_/C _4946_/A VGND VGND VPWR VPWR _4801_/X sky130_fd_sc_hd__and4_1
XFILLER_15_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5781_ _6042_/A1 _5781_/A1 _5785_/S VGND VGND VPWR VPWR _5781_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7520_ _7547_/CLK _7520_/D fanout609/X VGND VGND VPWR VPWR _7520_/Q sky130_fd_sc_hd__dfrtp_4
X_4732_ _5153_/A _5297_/A _5595_/D VGND VGND VPWR VPWR _4733_/B sky130_fd_sc_hd__and3_1
XFILLER_30_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4663_ _5000_/C _4836_/A _4631_/Y _4688_/B VGND VGND VPWR VPWR _5027_/C sky130_fd_sc_hd__o31ai_4
X_7451_ _7607_/CLK _7451_/D fanout624/X VGND VGND VPWR VPWR _7451_/Q sky130_fd_sc_hd__dfstp_1
X_3614_ _7585_/Q _6002_/A _4481_/A _3613_/X VGND VGND VPWR VPWR _3614_/X sky130_fd_sc_hd__a31o_1
X_6402_ _7124_/Q _6158_/D _6113_/Y _6153_/X _7207_/Q VGND VGND VPWR VPWR _6402_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_174_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4594_ _5096_/A _4884_/A VGND VGND VPWR VPWR _4595_/B sky130_fd_sc_hd__and2b_2
X_7382_ _7430_/CLK _7382_/D fanout627/X VGND VGND VPWR VPWR _7382_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_162_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold902 _7617_/Q VGND VGND VPWR VPWR hold902/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold913 _6010_/X VGND VGND VPWR VPWR _7585_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6333_ _7219_/Q _6359_/B _6428_/B1 _6151_/X _7214_/Q VGND VGND VPWR VPWR _6333_/X
+ sky130_fd_sc_hd__a32o_1
X_3545_ hold73/A _5768_/C _6020_/A VGND VGND VPWR VPWR _3545_/X sky130_fd_sc_hd__and3_4
XFILLER_127_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold924 _7431_/Q VGND VGND VPWR VPWR hold924/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold935 _7532_/Q VGND VGND VPWR VPWR hold935/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold946 _5855_/X VGND VGND VPWR VPWR _7447_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold957 hold957/A VGND VGND VPWR VPWR hold957/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 _7702_/A VGND VGND VPWR VPWR hold968/X sky130_fd_sc_hd__dlygate4sd3_1
X_6264_ _7535_/Q _6160_/D _6427_/A3 _6137_/X _7487_/Q VGND VGND VPWR VPWR _6264_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3476_ _6913_/Q _4193_/B VGND VGND VPWR VPWR _4192_/B sky130_fd_sc_hd__and2_4
Xhold979 hold979/A VGND VGND VPWR VPWR hold979/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5215_ _5215_/A _5215_/B _5215_/C VGND VGND VPWR VPWR _5218_/D sky130_fd_sc_hd__and3_1
XFILLER_142_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6195_ _7468_/Q _6309_/B _6131_/C _6151_/X _7548_/Q VGND VGND VPWR VPWR _6195_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_69_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5146_ _5146_/A _5146_/B _5146_/C _5512_/B VGND VGND VPWR VPWR _5147_/C sky130_fd_sc_hd__nand4_1
Xhold1602 _7045_/Q VGND VGND VPWR VPWR hold614/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1613 hold89/A VGND VGND VPWR VPWR _6847_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1624 _6912_/Q VGND VGND VPWR VPWR _3474_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1635 _7633_/Q VGND VGND VPWR VPWR _6103_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1646 _7131_/Q VGND VGND VPWR VPWR hold1646/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1657 _7668_/Q VGND VGND VPWR VPWR _6820_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5077_ _5297_/A _5233_/B _5233_/C VGND VGND VPWR VPWR _5077_/X sky130_fd_sc_hd__and3_1
XFILLER_84_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4028_ _7442_/Q _5849_/A _3973_/X _4022_/X _4027_/X VGND VGND VPWR VPWR _4036_/C
+ sky130_fd_sc_hd__a2111o_2
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5979_ _5979_/A0 _6042_/A1 _5983_/S VGND VGND VPWR VPWR _7557_/D sky130_fd_sc_hd__mux2_1
XFILLER_12_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7649_ _7680_/CLK _7649_/D fanout596/X VGND VGND VPWR VPWR _7649_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_138_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold209 _7374_/Q VGND VGND VPWR VPWR hold209/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _5017_/A _5109_/A _5000_/C VGND VGND VPWR VPWR _5092_/B sky130_fd_sc_hd__and3_4
XFILLER_39_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6951_ _4183_/A1 _6951_/D _6906_/X VGND VGND VPWR VPWR _6951_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5902_ hold511/X _6028_/A1 hold25/X VGND VGND VPWR VPWR _5902_/X sky130_fd_sc_hd__mux2_1
X_6882_ _6899_/A _6908_/B VGND VGND VPWR VPWR _6882_/X sky130_fd_sc_hd__and2_1
XFILLER_179_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5833_ hold981/X _6040_/A1 _5839_/S VGND VGND VPWR VPWR _5833_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5764_ hold288/X _5935_/A1 _5767_/S VGND VGND VPWR VPWR _5764_/X sky130_fd_sc_hd__mux2_1
X_7503_ _7584_/CLK _7503_/D fanout613/X VGND VGND VPWR VPWR _7503_/Q sky130_fd_sc_hd__dfrtp_2
X_4715_ _4740_/D _5595_/B _5358_/B _5233_/A _4738_/A VGND VGND VPWR VPWR _4721_/A
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_148_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5695_ hold85/X hold626/X _5695_/S VGND VGND VPWR VPWR _5695_/X sky130_fd_sc_hd__mux2_1
X_7434_ _7586_/CLK _7434_/D fanout625/X VGND VGND VPWR VPWR _7434_/Q sky130_fd_sc_hd__dfstp_1
X_4646_ _4637_/A _4595_/Y _4799_/A _5195_/B VGND VGND VPWR VPWR _5011_/A sky130_fd_sc_hd__o211ai_4
XFILLER_175_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold710 hold710/A VGND VGND VPWR VPWR hold710/X sky130_fd_sc_hd__dlygate4sd3_1
X_4577_ _4584_/C _4584_/D _5015_/C VGND VGND VPWR VPWR _4579_/A sky130_fd_sc_hd__nand3_1
Xhold721 hold721/A VGND VGND VPWR VPWR hold721/X sky130_fd_sc_hd__dlygate4sd3_1
X_7365_ _7445_/CLK _7365_/D fanout628/X VGND VGND VPWR VPWR _7365_/Q sky130_fd_sc_hd__dfrtp_4
Xhold732 _4432_/X VGND VGND VPWR VPWR _7127_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap451 wire452/X VGND VGND VPWR VPWR _6429_/A3 sky130_fd_sc_hd__clkbuf_2
Xhold743 _4549_/X VGND VGND VPWR VPWR _7230_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold754 _5969_/X VGND VGND VPWR VPWR _7548_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6316_ _7481_/Q _6133_/X _6309_/X _6310_/X _6315_/X VGND VGND VPWR VPWR _6316_/X
+ sky130_fd_sc_hd__a2111o_1
Xmax_cap462 _4877_/D VGND VGND VPWR VPWR _4907_/C sky130_fd_sc_hd__clkbuf_2
X_3528_ _3714_/A hold74/A _6020_/A VGND VGND VPWR VPWR _3528_/X sky130_fd_sc_hd__and3_4
Xhold765 _7500_/Q VGND VGND VPWR VPWR hold765/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7296_ _7547_/CLK _7296_/D fanout607/X VGND VGND VPWR VPWR _7296_/Q sky130_fd_sc_hd__dfrtp_2
Xhold776 _4393_/X VGND VGND VPWR VPWR _7095_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 _4503_/X VGND VGND VPWR VPWR _7192_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold798 _7033_/Q VGND VGND VPWR VPWR hold798/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6247_ _7478_/Q _6309_/B _6286_/C _6245_/X _6246_/X VGND VGND VPWR VPWR _6247_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_131_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3459_ _6392_/B VGND VGND VPWR VPWR _6126_/D sky130_fd_sc_hd__clkinv_2
XFILLER_39_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6178_ _7507_/Q _6428_/A2 _6124_/X _7531_/Q _6177_/X VGND VGND VPWR VPWR _6178_/X
+ sky130_fd_sc_hd__a221o_1
Xhold1410 _7146_/Q VGND VGND VPWR VPWR _4449_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1421 _5868_/X VGND VGND VPWR VPWR _7458_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1432 _7665_/Q VGND VGND VPWR VPWR _6817_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1443 _7664_/Q VGND VGND VPWR VPWR _6816_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5129_ _5611_/A2 _4960_/Y _4987_/Y _5128_/Y VGND VGND VPWR VPWR _5129_/Y sky130_fd_sc_hd__o31ai_1
Xhold1454 _7554_/Q VGND VGND VPWR VPWR hold513/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1465 _7103_/Q VGND VGND VPWR VPWR hold1465/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1476 _7498_/Q VGND VGND VPWR VPWR hold534/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1487 _7642_/Q VGND VGND VPWR VPWR _6297_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1498 _5904_/X VGND VGND VPWR VPWR _7490_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_605 _6160_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_616 _7001_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_627 _4522_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_638 _6131_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_649 _6137_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold70 hold70/A VGND VGND VPWR VPWR hold70/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold81 hold81/A VGND VGND VPWR VPWR hold81/X sky130_fd_sc_hd__buf_6
Xhold92 hold92/A VGND VGND VPWR VPWR hold92/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4500_ _6012_/A0 _4500_/A1 _4504_/S VGND VGND VPWR VPWR _4500_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5480_ _5480_/A _5595_/A VGND VGND VPWR VPWR _5597_/C sky130_fd_sc_hd__nand2_1
XFILLER_117_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1 _4276_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4431_ _4431_/A0 _6862_/A1 _4435_/S VGND VGND VPWR VPWR _4431_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7150_ _7672_/CLK _7150_/D VGND VGND VPWR VPWR _7150_/Q sky130_fd_sc_hd__dfxtp_1
X_4362_ _5988_/A1 hold920/X _4363_/S VGND VGND VPWR VPWR _4362_/X sky130_fd_sc_hd__mux2_1
X_6101_ _7633_/Q _7632_/Q VGND VGND VPWR VPWR _6516_/C sky130_fd_sc_hd__and2b_4
X_7081_ _7130_/CLK _7081_/D fanout602/X VGND VGND VPWR VPWR _7081_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout508 _4569_/X VGND VGND VPWR VPWR _5551_/A1 sky130_fd_sc_hd__buf_4
X_4293_ hold508/X _6028_/A1 _4293_/S VGND VGND VPWR VPWR _4293_/X sky130_fd_sc_hd__mux2_1
Xfanout519 hold19/X VGND VGND VPWR VPWR _4564_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_58_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6032_ _6041_/A1 hold744/X _6037_/S VGND VGND VPWR VPWR _6032_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6934_ _6950_/CLK _6934_/D _6889_/X VGND VGND VPWR VPWR hold7/A sky130_fd_sc_hd__dfrtp_1
XFILLER_54_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6865_ _6865_/A0 _6865_/A1 _6866_/S VGND VGND VPWR VPWR _6865_/X sky130_fd_sc_hd__mux2_1
X_5816_ _5843_/A1 hold252/X _5821_/S VGND VGND VPWR VPWR _5816_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6796_ _7208_/Q _6099_/B _6720_/D _6464_/X _7686_/Q VGND VGND VPWR VPWR _6796_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_10_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5747_ _6044_/A1 hold928/X _5749_/S VGND VGND VPWR VPWR _5747_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5678_ _5697_/A0 _5678_/B _5678_/C VGND VGND VPWR VPWR _5678_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_136_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7417_ _7568_/CLK _7417_/D fanout622/X VGND VGND VPWR VPWR _7417_/Q sky130_fd_sc_hd__dfrtp_1
X_4629_ _5407_/A _5074_/A _5404_/A VGND VGND VPWR VPWR _4629_/Y sky130_fd_sc_hd__nand3_4
Xhold540 _4480_/X VGND VGND VPWR VPWR _7173_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold551 _4435_/X VGND VGND VPWR VPWR _7130_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7348_ _7562_/CLK _7348_/D fanout621/X VGND VGND VPWR VPWR _7348_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_190_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold562 _4381_/X VGND VGND VPWR VPWR _7085_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 _7608_/Q VGND VGND VPWR VPWR hold573/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold584 _5964_/X VGND VGND VPWR VPWR _7544_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 hold595/A VGND VGND VPWR VPWR wb_dat_o[14] sky130_fd_sc_hd__buf_12
X_7279_ _7614_/CLK _7279_/D fanout604/X VGND VGND VPWR VPWR _7279_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_89_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1240 _7452_/Q VGND VGND VPWR VPWR _5861_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1251 _5747_/X VGND VGND VPWR VPWR _7351_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1262 _7251_/Q VGND VGND VPWR VPWR hold1262/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1273 _5662_/X VGND VGND VPWR VPWR _7281_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1284 _7549_/Q VGND VGND VPWR VPWR hold1284/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_402 _3975_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1295 _7440_/Q VGND VGND VPWR VPWR hold718/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_413 _5983_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_424 _6158_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_435 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_446 _6451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_457 _6484_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_468 _7428_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_479 _7232_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput160 wb_dat_i[6] VGND VGND VPWR VPWR _6849_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4980_ _5027_/D _5011_/A _5472_/C VGND VGND VPWR VPWR _5066_/A sky130_fd_sc_hd__o21ai_1
XFILLER_63_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3931_ _7395_/Q _3525_/X _4499_/A _7190_/Q _3930_/X VGND VGND VPWR VPWR _3931_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_16_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6650_ _7352_/Q _6465_/X _6644_/X _6647_/X _6649_/X VGND VGND VPWR VPWR _6651_/C
+ sky130_fd_sc_hd__a2111o_1
XFILLER_149_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3862_ _7396_/Q _3525_/X _3855_/X _3856_/X _3861_/X VGND VGND VPWR VPWR _3862_/X
+ sky130_fd_sc_hd__a2111o_2
X_5601_ _5429_/A _5084_/X _5069_/X _5501_/B _5140_/X VGND VGND VPWR VPWR _5601_/Y
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_177_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6581_ hold46/A _6479_/X _6486_/X _7501_/Q _6580_/X VGND VGND VPWR VPWR _6581_/X
+ sky130_fd_sc_hd__a221o_1
X_3793_ _7079_/Q _5840_/A _4535_/B _3602_/X _7421_/Q VGND VGND VPWR VPWR _3793_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_118_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5532_ _5614_/C _4702_/X _5027_/X _5614_/A VGND VGND VPWR VPWR _5532_/X sky130_fd_sc_hd__o211a_1
XFILLER_157_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_9_csclk _7236_/CLK VGND VGND VPWR VPWR _7197_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_117_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5463_ _5463_/A _5463_/B _5463_/C VGND VGND VPWR VPWR _5534_/B sky130_fd_sc_hd__and3_1
XFILLER_172_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7202_ _7202_/CLK _7202_/D fanout619/X VGND VGND VPWR VPWR _7202_/Q sky130_fd_sc_hd__dfrtp_2
X_4414_ hold719/X _6863_/A1 _4417_/S VGND VGND VPWR VPWR _4414_/X sky130_fd_sc_hd__mux2_1
X_5394_ _4873_/Y _5381_/X _5393_/X _5259_/B VGND VGND VPWR VPWR _5399_/B sky130_fd_sc_hd__o211a_1
XFILLER_160_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7133_ _7462_/CLK _7133_/D fanout604/X VGND VGND VPWR VPWR _7133_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_99_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4345_ _6866_/A1 hold254/X _4345_/S VGND VGND VPWR VPWR _4345_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4276_ _4275_/X hold931/X _4276_/S VGND VGND VPWR VPWR _4276_/X sky130_fd_sc_hd__mux2_1
X_7064_ _7192_/CLK _7064_/D fanout617/X VGND VGND VPWR VPWR _7064_/Q sky130_fd_sc_hd__dfrtp_1
X_6015_ _6042_/A1 _6015_/A1 _6019_/S VGND VGND VPWR VPWR _7589_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6917_ _6950_/CLK _6917_/D _6872_/X VGND VGND VPWR VPWR _6917_/Q sky130_fd_sc_hd__dfrtp_2
X_6848_ _6971_/Q _6848_/A2 _6848_/B1 _6970_/Q VGND VGND VPWR VPWR _6848_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6779_ _7099_/Q _6444_/X _6468_/X _7177_/Q _6778_/X VGND VGND VPWR VPWR _6784_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_183_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold370 _4502_/X VGND VGND VPWR VPWR _7191_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 _7190_/Q VGND VGND VPWR VPWR hold381/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold392 _4504_/X VGND VGND VPWR VPWR _7193_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1070 _4476_/X VGND VGND VPWR VPWR _7169_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 hold1300/X VGND VGND VPWR VPWR _5808_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1092 _7684_/Q VGND VGND VPWR VPWR _6864_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_210 _7047_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_221 _7222_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_232 _6953_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_243 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_254 _4199_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_265 _7714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_276 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_287 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_298 input96/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4130_ _4140_/B _4130_/B _6811_/S VGND VGND VPWR VPWR _4130_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_123_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4061_ _4061_/A0 input58/X _4192_/B VGND VGND VPWR VPWR _6932_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4963_ _4948_/B _4966_/A _5112_/B _4966_/B VGND VGND VPWR VPWR _4963_/X sky130_fd_sc_hd__and4b_1
XFILLER_189_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6702_ _7096_/Q _6444_/X _6485_/X _7214_/Q _6701_/X VGND VGND VPWR VPWR _6709_/A
+ sky130_fd_sc_hd__a221o_1
X_3914_ _7215_/Q _5993_/A _4529_/B _3557_/X _7571_/Q VGND VGND VPWR VPWR _3914_/X
+ sky130_fd_sc_hd__a32o_1
X_7682_ _7682_/CLK _7682_/D fanout603/X VGND VGND VPWR VPWR _7682_/Q sky130_fd_sc_hd__dfrtp_4
X_4894_ _4767_/Y _4892_/Y _4893_/Y _4891_/Y VGND VGND VPWR VPWR _4902_/C sky130_fd_sc_hd__o211ai_1
XFILLER_149_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6633_ _6612_/X _6614_/X _6633_/C _6633_/D VGND VGND VPWR VPWR _6633_/X sky130_fd_sc_hd__and4bb_2
X_3845_ _7253_/Q _4541_/A hold70/A VGND VGND VPWR VPWR _3845_/X sky130_fd_sc_hd__and3_1
XFILLER_20_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6564_ _7437_/Q _6097_/X _6445_/C _6474_/A _7341_/Q VGND VGND VPWR VPWR _6564_/X
+ sky130_fd_sc_hd__a32o_1
X_3776_ _7398_/Q _3525_/X _3722_/X _3732_/X _3775_/Y VGND VGND VPWR VPWR _3776_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_118_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5515_ _5605_/C _5515_/B _5515_/C VGND VGND VPWR VPWR _5515_/Y sky130_fd_sc_hd__nand3_1
XFILLER_145_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6495_ _7514_/Q _6645_/B _6536_/C _6447_/X _7522_/Q VGND VGND VPWR VPWR _6495_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_133_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5446_ _4953_/B _5088_/Y _5387_/X _4880_/Y _5445_/X VGND VGND VPWR VPWR _5446_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_172_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5377_ _4597_/Y _4821_/Y _4882_/Y _4816_/Y _4817_/Y VGND VGND VPWR VPWR _5555_/C
+ sky130_fd_sc_hd__o32a_1
XFILLER_114_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7116_ _7685_/CLK _7116_/D fanout617/X VGND VGND VPWR VPWR _7116_/Q sky130_fd_sc_hd__dfrtp_4
X_4328_ _4529_/B _4481_/A _6861_/C VGND VGND VPWR VPWR _4333_/S sky130_fd_sc_hd__and3_4
XFILLER_59_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7047_ _7286_/CLK _7047_/D fanout598/X VGND VGND VPWR VPWR _7047_/Q sky130_fd_sc_hd__dfrtp_4
X_4259_ _7294_/Q _4171_/C _4171_/D _5984_/B VGND VGND VPWR VPWR _4259_/Y sky130_fd_sc_hd__o31ai_2
XFILLER_47_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_606 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_74_csclk _7095_/CLK VGND VGND VPWR VPWR _7289_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_147_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3630_ _7328_/Q _3565_/X _5741_/A _7352_/Q _3629_/X VGND VGND VPWR VPWR _3630_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3561_ _5993_/A _5661_/A _4340_/A VGND VGND VPWR VPWR _3561_/X sky130_fd_sc_hd__and3_2
X_5300_ _5291_/C _5012_/X _5313_/A _5298_/X VGND VGND VPWR VPWR _5300_/X sky130_fd_sc_hd__a31o_1
XFILLER_161_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3492_ _3491_/X hold60/X _4229_/S VGND VGND VPWR VPWR hold61/A sky130_fd_sc_hd__mux2_2
XFILLER_6_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6280_ _7352_/Q wire455/X _6149_/X _7424_/Q _6279_/X VGND VGND VPWR VPWR _6280_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_142_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5231_ _5313_/C _5231_/B _5231_/C _5316_/C VGND VGND VPWR VPWR _5231_/X sky130_fd_sc_hd__and4_1
X_5162_ _5162_/A _5162_/B _5162_/C VGND VGND VPWR VPWR _5162_/Y sky130_fd_sc_hd__nor3_1
XFILLER_123_580 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_12_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7253_/CLK sky130_fd_sc_hd__clkbuf_16
X_4113_ _4584_/C _4584_/D _4113_/C input116/X VGND VGND VPWR VPWR _4116_/D sky130_fd_sc_hd__nor4b_1
X_5093_ _5313_/B _5093_/B _5093_/C VGND VGND VPWR VPWR _5093_/X sky130_fd_sc_hd__and3_1
XFILLER_68_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4044_ _6956_/Q _6957_/Q _6955_/Q VGND VGND VPWR VPWR _4049_/B sky130_fd_sc_hd__nor3b_2
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_27_csclk _7352_/CLK VGND VGND VPWR VPWR _7515_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_52_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5995_ hold351/X _6031_/A0 _6001_/S VGND VGND VPWR VPWR _5995_/X sky130_fd_sc_hd__mux2_1
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4946_ _4946_/A _4946_/B _5261_/D VGND VGND VPWR VPWR _4947_/A sky130_fd_sc_hd__and3_1
XFILLER_33_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7665_ _7676_/CLK _7665_/D VGND VGND VPWR VPWR _7665_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_193_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4877_ _4990_/A _5017_/A _4877_/C _4877_/D VGND VGND VPWR VPWR _4966_/B sky130_fd_sc_hd__nor4_2
XFILLER_177_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6616_ _7431_/Q _6444_/X _6474_/A _7343_/Q _6615_/X VGND VGND VPWR VPWR _6623_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_192_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3828_ _7325_/Q _5786_/B _5759_/B _3571_/X _7357_/Q VGND VGND VPWR VPWR _3828_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_165_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7596_ _7606_/CLK _7596_/D fanout612/X VGND VGND VPWR VPWR _7596_/Q sky130_fd_sc_hd__dfrtp_1
X_6547_ _7572_/Q _6457_/X _6465_/X _7348_/Q _6540_/X VGND VGND VPWR VPWR _6547_/X
+ sky130_fd_sc_hd__a221o_1
X_3759_ _7558_/Q _5993_/A _5975_/B _3758_/X VGND VGND VPWR VPWR _3759_/X sky130_fd_sc_hd__a31o_1
XFILLER_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6478_ _6457_/X _6468_/X _6478_/C _6478_/D VGND VGND VPWR VPWR _6478_/Y sky130_fd_sc_hd__nand4bb_4
XFILLER_106_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5429_ _5429_/A _5512_/B _5512_/D _5429_/D VGND VGND VPWR VPWR _5514_/B sky130_fd_sc_hd__nand4_1
XFILLER_160_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput250 _4182_/Y VGND VGND VPWR VPWR pad_flash_csb_oeb sky130_fd_sc_hd__buf_12
Xoutput261 _7260_/Q VGND VGND VPWR VPWR pll_dco_ena sky130_fd_sc_hd__buf_12
Xoutput272 _7133_/Q VGND VGND VPWR VPWR pll_trim[10] sky130_fd_sc_hd__buf_12
XFILLER_121_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput283 _7276_/Q VGND VGND VPWR VPWR pll_trim[20] sky130_fd_sc_hd__buf_12
Xoutput294 _6979_/Q VGND VGND VPWR VPWR pll_trim[7] sky130_fd_sc_hd__buf_12
XFILLER_58_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_523 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire355 _3634_/Y VGND VGND VPWR VPWR _3655_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_156_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire366 _6684_/Y VGND VGND VPWR VPWR wire366/X sky130_fd_sc_hd__clkbuf_1
Xwire377 _6204_/Y VGND VGND VPWR VPWR wire377/X sky130_fd_sc_hd__clkbuf_1
XFILLER_171_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4800_ _5476_/B _5476_/D VGND VGND VPWR VPWR _4800_/Y sky130_fd_sc_hd__nand2_2
XFILLER_34_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5780_ _5843_/A1 hold313/X _5785_/S VGND VGND VPWR VPWR _5780_/X sky130_fd_sc_hd__mux2_1
X_4731_ _5153_/A _5196_/A _5358_/B VGND VGND VPWR VPWR _4733_/A sky130_fd_sc_hd__and3_1
XFILLER_187_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7450_ _7616_/CLK _7450_/D fanout610/X VGND VGND VPWR VPWR _7450_/Q sky130_fd_sc_hd__dfstp_2
X_4662_ _5000_/C _4836_/A _4660_/C _5007_/D VGND VGND VPWR VPWR _5027_/B sky130_fd_sc_hd__o31ai_4
XFILLER_147_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6401_ _7254_/Q _6159_/B _6416_/C _6166_/C VGND VGND VPWR VPWR _6401_/X sky130_fd_sc_hd__o211a_1
X_3613_ _4198_/B _4505_/B _6002_/B _4275_/S input42/X VGND VGND VPWR VPWR _3613_/X
+ sky130_fd_sc_hd__a32o_1
X_7381_ _7421_/CLK _7381_/D fanout630/X VGND VGND VPWR VPWR _7381_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_190_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4593_ _4884_/A _5096_/A VGND VGND VPWR VPWR _5143_/B sky130_fd_sc_hd__and2b_4
XFILLER_128_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold903 _6046_/X VGND VGND VPWR VPWR _7617_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_127_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6332_ _7251_/Q _6082_/B _6416_/C _6166_/C VGND VGND VPWR VPWR _6332_/X sky130_fd_sc_hd__o211a_1
Xhold914 _7441_/Q VGND VGND VPWR VPWR hold914/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3544_ _3717_/B _3573_/C _5682_/B VGND VGND VPWR VPWR _3544_/X sky130_fd_sc_hd__and3_4
Xhold925 _5837_/X VGND VGND VPWR VPWR _7431_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 _5951_/X VGND VGND VPWR VPWR _7532_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold947 _7551_/Q VGND VGND VPWR VPWR hold947/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_142_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold958 _7327_/Q VGND VGND VPWR VPWR hold958/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold969 _4256_/X VGND VGND VPWR VPWR _6994_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6263_ _7519_/Q _6146_/X _6161_/X _7351_/Q _6262_/X VGND VGND VPWR VPWR _6263_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3475_ _6914_/Q _6912_/Q VGND VGND VPWR VPWR _4193_/B sky130_fd_sc_hd__nor2_2
XFILLER_142_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5214_ _4761_/A _5614_/B _5614_/D _5038_/B _5002_/B VGND VGND VPWR VPWR _5215_/C
+ sky130_fd_sc_hd__a32oi_1
X_6194_ _7532_/Q _6160_/D _6427_/A3 _6427_/B1 _7484_/Q VGND VGND VPWR VPWR _6194_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_97_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1603 hold72/A VGND VGND VPWR VPWR _5569_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5145_ _4811_/Y _4816_/Y _4821_/Y _4795_/Y VGND VGND VPWR VPWR _5147_/B sky130_fd_sc_hd__a211o_1
Xhold1614 _6917_/Q VGND VGND VPWR VPWR _4101_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1625 _6951_/Q VGND VGND VPWR VPWR _3474_/B1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1636 _6961_/Q VGND VGND VPWR VPWR _4118_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1647 _7620_/Q VGND VGND VPWR VPWR _6058_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1658 _6964_/Q VGND VGND VPWR VPWR _4454_/B sky130_fd_sc_hd__dlygate4sd3_1
X_5076_ _5075_/X _5076_/B _5076_/C VGND VGND VPWR VPWR _5079_/A sky130_fd_sc_hd__nand3b_1
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4027_ _7164_/Q _3697_/X _4023_/X _4024_/X _4026_/X VGND VGND VPWR VPWR _4027_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_84_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5978_ hold937/X _6041_/A1 _5983_/S VGND VGND VPWR VPWR _5978_/X sky130_fd_sc_hd__mux2_1
X_4929_ _4943_/A _5261_/D _4957_/C _4934_/C VGND VGND VPWR VPWR _4930_/C sky130_fd_sc_hd__nand4_1
XFILLER_166_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7648_ _7662_/CLK _7648_/D fanout597/X VGND VGND VPWR VPWR _7648_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7579_ _7580_/CLK _7579_/D fanout605/X VGND VGND VPWR VPWR _7579_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_193_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmgmt_gpio_9_buff_inst _4155_/X VGND VGND VPWR VPWR mgmt_gpio_out[9] sky130_fd_sc_hd__clkbuf_8
XFILLER_134_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6950_ _6950_/CLK _6950_/D _6905_/X VGND VGND VPWR VPWR _6950_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_66_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5901_ hold485/X _6045_/A1 hold25/X VGND VGND VPWR VPWR _5901_/X sky130_fd_sc_hd__mux2_1
X_6881_ _6899_/A _6911_/B VGND VGND VPWR VPWR _6881_/X sky130_fd_sc_hd__and2_1
XFILLER_62_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5832_ hold420/X _6003_/A1 _5839_/S VGND VGND VPWR VPWR _5832_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5763_ _5763_/A0 _6042_/A1 _5767_/S VGND VGND VPWR VPWR _5763_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7502_ _7614_/CLK _7502_/D fanout605/X VGND VGND VPWR VPWR _7502_/Q sky130_fd_sc_hd__dfrtp_4
X_4714_ _4801_/C _5595_/B _5595_/D _4738_/A VGND VGND VPWR VPWR _4714_/X sky130_fd_sc_hd__o211a_1
X_5694_ _5926_/A0 hold581/X _5695_/S VGND VGND VPWR VPWR _5694_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7433_ _7435_/CLK _7433_/D fanout623/X VGND VGND VPWR VPWR _7433_/Q sky130_fd_sc_hd__dfrtp_1
X_4645_ _4637_/A _4595_/Y _4799_/A _5195_/B VGND VGND VPWR VPWR _5061_/A sky130_fd_sc_hd__o211a_4
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold700 _7292_/Q VGND VGND VPWR VPWR hold700/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7364_ _7518_/CLK _7364_/D fanout627/X VGND VGND VPWR VPWR _7364_/Q sky130_fd_sc_hd__dfrtp_4
Xhold711 hold711/A VGND VGND VPWR VPWR wb_dat_o[7] sky130_fd_sc_hd__buf_12
XFILLER_116_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4576_ _4576_/A _4576_/B VGND VGND VPWR VPWR _4781_/B sky130_fd_sc_hd__nor2_2
Xhold722 hold722/A VGND VGND VPWR VPWR wb_dat_o[23] sky130_fd_sc_hd__buf_12
Xhold733 hold733/A VGND VGND VPWR VPWR hold733/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 _7604_/Q VGND VGND VPWR VPWR hold744/X sky130_fd_sc_hd__dlygate4sd3_1
X_6315_ _7377_/Q _6160_/X _6311_/X _6312_/X _6314_/X VGND VGND VPWR VPWR _6315_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_190_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap463 _4740_/D VGND VGND VPWR VPWR _4801_/C sky130_fd_sc_hd__buf_4
Xhold755 _7468_/Q VGND VGND VPWR VPWR hold755/X sky130_fd_sc_hd__dlygate4sd3_1
X_3527_ hold69/X _3622_/A hold23/X _3559_/B VGND VGND VPWR VPWR _3546_/C sky130_fd_sc_hd__and4bb_2
X_7295_ _7497_/CLK _7295_/D fanout607/X VGND VGND VPWR VPWR _7295_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_143_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold766 _5915_/X VGND VGND VPWR VPWR _7500_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap474 _6141_/X VGND VGND VPWR VPWR _6407_/A3 sky130_fd_sc_hd__buf_6
Xhold777 _7160_/Q VGND VGND VPWR VPWR hold777/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold788 _7584_/Q VGND VGND VPWR VPWR hold788/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap496 _4948_/Y VGND VGND VPWR VPWR _4951_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_131_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold799 _4319_/X VGND VGND VPWR VPWR _7033_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6246_ _7558_/Q _6309_/B _6432_/A3 _6138_/X _7358_/Q VGND VGND VPWR VPWR _6246_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3458_ _6158_/D VGND VGND VPWR VPWR _3458_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6177_ _7515_/Q _6067_/X _6146_/C _6137_/X _7483_/Q VGND VGND VPWR VPWR _6177_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_190_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1400 _6958_/Q VGND VGND VPWR VPWR hold1400/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1411 _7587_/Q VGND VGND VPWR VPWR _6013_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1422 _7666_/Q VGND VGND VPWR VPWR _6818_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1433 _7074_/Q VGND VGND VPWR VPWR hold465/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5128_ _4948_/B _5090_/B _5452_/C _5127_/Y VGND VGND VPWR VPWR _5128_/Y sky130_fd_sc_hd__a31oi_1
Xhold1444 _7108_/Q VGND VGND VPWR VPWR hold1444/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1455 _7660_/Q VGND VGND VPWR VPWR _6786_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1466 _4403_/X VGND VGND VPWR VPWR _7103_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1477 _5913_/X VGND VGND VPWR VPWR _7498_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1488 _6275_/X VGND VGND VPWR VPWR _7642_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5059_ _5059_/A _5059_/B _5059_/C _5059_/D VGND VGND VPWR VPWR _5059_/Y sky130_fd_sc_hd__nor4_1
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1499 _7054_/Q VGND VGND VPWR VPWR hold450/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_606 _6416_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_617 hold833/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_628 _4522_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_639 _6131_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold60 hold60/A VGND VGND VPWR VPWR hold60/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 hold71/A VGND VGND VPWR VPWR hold71/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 hold82/A VGND VGND VPWR VPWR hold82/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 hold93/A VGND VGND VPWR VPWR hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4430_ _4559_/B _5678_/B _5680_/C VGND VGND VPWR VPWR _4435_/S sky130_fd_sc_hd__and3_2
XANTENNA_2 _4318_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4361_ _5789_/A1 hold506/X _4363_/S VGND VGND VPWR VPWR _4361_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6100_ _6103_/B2 _7632_/Q _6099_/B _6098_/Y VGND VGND VPWR VPWR _6100_/Y sky130_fd_sc_hd__a31oi_1
Xfanout509 hold102/X VGND VGND VPWR VPWR _6028_/A1 sky130_fd_sc_hd__buf_8
X_7080_ _7212_/CLK _7080_/D fanout619/X VGND VGND VPWR VPWR _7080_/Q sky130_fd_sc_hd__dfrtp_4
X_4292_ _4291_/X hold267/X _4292_/S VGND VGND VPWR VPWR _4292_/X sky130_fd_sc_hd__mux2_1
X_6031_ _6031_/A0 hold331/X _6037_/S VGND VGND VPWR VPWR _6031_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6933_ _4172_/B2 _6933_/D _6888_/X VGND VGND VPWR VPWR hold79/A sky130_fd_sc_hd__dfrtp_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6864_ _6864_/A0 _6864_/A1 _6866_/S VGND VGND VPWR VPWR _6864_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5815_ _6040_/A1 hold973/X _5821_/S VGND VGND VPWR VPWR _5815_/X sky130_fd_sc_hd__mux2_1
X_6795_ _7080_/Q _6450_/X _6791_/X _6792_/X _6794_/X VGND VGND VPWR VPWR _6800_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_50_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5746_ _5926_/A0 hold216/X _5749_/S VGND VGND VPWR VPWR _5746_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5677_ hold700/X _6863_/A1 _5677_/S VGND VGND VPWR VPWR _5677_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7416_ _7445_/CLK _7416_/D fanout628/X VGND VGND VPWR VPWR _7416_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_163_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4628_ _5407_/A _5074_/A _5404_/A VGND VGND VPWR VPWR _5068_/A sky130_fd_sc_hd__and3_2
Xhold530 _7226_/Q VGND VGND VPWR VPWR hold530/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7347_ _7611_/CLK _7347_/D fanout621/X VGND VGND VPWR VPWR _7347_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_151_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4559_ _5682_/A _4559_/B _5659_/C _5686_/D VGND VGND VPWR VPWR _4564_/S sky130_fd_sc_hd__and4_4
Xhold541 _7238_/Q VGND VGND VPWR VPWR hold541/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold552 hold552/A VGND VGND VPWR VPWR hold552/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_9_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold563 hold563/A VGND VGND VPWR VPWR hold563/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold574 _6036_/X VGND VGND VPWR VPWR _7608_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7278_ _7462_/CLK hold67/X fanout604/X VGND VGND VPWR VPWR _7278_/Q sky130_fd_sc_hd__dfstp_1
Xhold585 _7225_/Q VGND VGND VPWR VPWR hold585/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 _7178_/Q VGND VGND VPWR VPWR hold596/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_106_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6229_ _6228_/X _6252_/A1 _6812_/S VGND VGND VPWR VPWR _7640_/D sky130_fd_sc_hd__mux2_1
XFILLER_77_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1230 _6823_/A1 VGND VGND VPWR VPWR hold667/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1241 _7446_/Q VGND VGND VPWR VPWR _5854_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1252 _7218_/Q VGND VGND VPWR VPWR hold248/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1263 _5629_/X VGND VGND VPWR VPWR _7251_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1274 _7224_/Q VGND VGND VPWR VPWR hold817/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1285 _7358_/Q VGND VGND VPWR VPWR hold276/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_403 _4033_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1296 _5847_/X VGND VGND VPWR VPWR _7440_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_414 _6157_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_425 _6158_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_436 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_447 _6452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_458 _6486_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_469 _7049_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput150 wb_dat_i[26] VGND VGND VPWR VPWR _6836_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput161 wb_dat_i[7] VGND VGND VPWR VPWR _6852_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3930_ _7347_/Q _5957_/B _4511_/C _4346_/A _7057_/Q VGND VGND VPWR VPWR _3930_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_32_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3861_ _7324_/Q _5786_/B _4487_/B _3858_/X _3860_/X VGND VGND VPWR VPWR _3861_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_149_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5600_ _4821_/Y _5611_/A2 _4993_/Y _5566_/D VGND VGND VPWR VPWR _5603_/B sky130_fd_sc_hd__o31a_1
X_6580_ _7581_/Q _6452_/X _6485_/X _7549_/Q _6579_/X VGND VGND VPWR VPWR _6580_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_32_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3792_ _7557_/Q _5984_/A _5975_/B _3696_/X _7202_/Q VGND VGND VPWR VPWR _3792_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_192_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5531_ _5530_/X _5570_/C _5409_/X _5522_/X VGND VGND VPWR VPWR _5558_/A sky130_fd_sc_hd__a211o_1
XFILLER_191_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5462_ _5462_/A1 _5585_/A1 _4823_/Y _5015_/Y _5461_/X VGND VGND VPWR VPWR _5463_/C
+ sky130_fd_sc_hd__o41a_1
XFILLER_117_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7201_ _7212_/CLK _7201_/D fanout619/X VGND VGND VPWR VPWR _7201_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_172_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4413_ _4413_/A0 _5697_/A0 _4417_/S VGND VGND VPWR VPWR _4413_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5393_ _5442_/B _5524_/B _5393_/C VGND VGND VPWR VPWR _5393_/X sky130_fd_sc_hd__and3_1
XFILLER_126_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7132_ _7286_/CLK _7132_/D fanout598/X VGND VGND VPWR VPWR _7132_/Q sky130_fd_sc_hd__dfstp_2
X_4344_ _5673_/A1 hold450/X _4345_/S VGND VGND VPWR VPWR _7054_/D sky130_fd_sc_hd__mux2_1
XFILLER_125_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7063_ _7686_/CLK _7063_/D fanout599/X VGND VGND VPWR VPWR _7063_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_59_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4275_ hold571/X _6028_/A1 _4275_/S VGND VGND VPWR VPWR _4275_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6014_ _6041_/A1 hold829/X _6019_/S VGND VGND VPWR VPWR _6014_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6916_ _6950_/CLK _6916_/D _6871_/X VGND VGND VPWR VPWR _6916_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_54_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6847_ _6847_/A0 _6846_/X _6853_/S VGND VGND VPWR VPWR _7677_/D sky130_fd_sc_hd__mux2_1
XFILLER_22_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6778_ _7207_/Q _6099_/B _6563_/C _6487_/X _7129_/Q VGND VGND VPWR VPWR _6778_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5729_ hold877/X _6044_/A1 _5731_/S VGND VGND VPWR VPWR _5729_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold360 _4490_/X VGND VGND VPWR VPWR _7181_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 _7436_/Q VGND VGND VPWR VPWR hold371/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold382 _4501_/X VGND VGND VPWR VPWR _7190_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 _7180_/Q VGND VGND VPWR VPWR hold393/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1060 hold1256/X VGND VGND VPWR VPWR _6862_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_93_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1071 hold1276/X VGND VGND VPWR VPWR _6024_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_532 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1082 hold1313/X VGND VGND VPWR VPWR _5853_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_200 _6846_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1093 hold1353/X VGND VGND VPWR VPWR _5736_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_211 _7047_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_222 _7163_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_233 mgmt_gpio_in[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_244 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_255 _4199_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_266 _7714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_277 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_288 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_299 input96/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4060_ _4060_/A0 _4061_/A0 _4192_/B VGND VGND VPWR VPWR _6933_/D sky130_fd_sc_hd__mux2_1
XFILLER_49_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4962_ _5311_/A _5404_/B VGND VGND VPWR VPWR _5570_/C sky130_fd_sc_hd__nand2_1
X_3913_ _7491_/Q _3519_/X _3908_/X _3910_/X _3912_/X VGND VGND VPWR VPWR _3913_/X
+ sky130_fd_sc_hd__a2111o_1
X_6701_ _7224_/Q _6463_/X _6468_/X _7174_/Q VGND VGND VPWR VPWR _6701_/X sky130_fd_sc_hd__a22o_1
XFILLER_32_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7681_ _4167_/A1 _7681_/D fanout635/X VGND VGND VPWR VPWR _7681_/Q sky130_fd_sc_hd__dfrtp_4
X_4893_ _4953_/D _4953_/A _5021_/B _4899_/C VGND VGND VPWR VPWR _4893_/Y sky130_fd_sc_hd__nand4b_1
X_6632_ _6632_/A _6632_/B _6632_/C _6809_/D VGND VGND VPWR VPWR _6633_/D sky130_fd_sc_hd__nor4_1
X_3844_ _7476_/Q _5903_/A _5957_/B VGND VGND VPWR VPWR _3844_/X sky130_fd_sc_hd__and3_1
XFILLER_177_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6563_ _7477_/Q _6791_/C _6563_/C _6791_/D VGND VGND VPWR VPWR _6563_/X sky130_fd_sc_hd__and4_1
XFILLER_158_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3775_ _3775_/A _3775_/B _3775_/C VGND VGND VPWR VPWR _3775_/Y sky130_fd_sc_hd__nand3_2
XFILLER_118_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5514_ _5314_/A _5514_/B _5514_/C _5514_/D VGND VGND VPWR VPWR _5515_/C sky130_fd_sc_hd__and4b_1
XFILLER_157_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6494_ _7530_/Q _6720_/C _6536_/C _6464_/X _7458_/Q VGND VGND VPWR VPWR _6494_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_173_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5445_ _4859_/Y _4960_/Y _5018_/Y _5261_/Y _4890_/X VGND VGND VPWR VPWR _5445_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_118_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5376_ _5376_/A _5376_/B _5376_/C VGND VGND VPWR VPWR _5378_/B sky130_fd_sc_hd__nor3_1
X_7115_ _7686_/CLK _7115_/D fanout599/X VGND VGND VPWR VPWR _7115_/Q sky130_fd_sc_hd__dfrtp_2
X_4327_ hold228/X _6866_/A1 _4327_/S VGND VGND VPWR VPWR _7040_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7046_ _7291_/CLK _7046_/D fanout596/X VGND VGND VPWR VPWR _7046_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4258_ hold436/X _4257_/X _4258_/S VGND VGND VPWR VPWR _4258_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4189_ input85/X input58/X _6923_/Q VGND VGND VPWR VPWR _4189_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire537 _6858_/C VGND VGND VPWR VPWR wire537/X sky130_fd_sc_hd__buf_2
XFILLER_7_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold190 _4208_/X VGND VGND VPWR VPWR _6959_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_120_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3560_ hold74/A _5686_/B _4505_/B VGND VGND VPWR VPWR _3560_/X sky130_fd_sc_hd__and3_4
XFILLER_155_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3491_ _6929_/Q _6912_/Q _3500_/C _3490_/X VGND VGND VPWR VPWR _3491_/X sky130_fd_sc_hd__a31o_1
XFILLER_6_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5230_ _5066_/A _5230_/B _5230_/C _5472_/B VGND VGND VPWR VPWR _5230_/Y sky130_fd_sc_hd__nand4b_1
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5161_ _4743_/C _5153_/C _5358_/B _5160_/X _5159_/X VGND VGND VPWR VPWR _5162_/C
+ sky130_fd_sc_hd__a311o_1
XFILLER_96_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4112_ _4585_/C _4585_/D _4584_/A _4584_/B VGND VGND VPWR VPWR _4115_/C sky130_fd_sc_hd__nor4_1
X_5092_ _5092_/A _5092_/B VGND VGND VPWR VPWR _5121_/C sky130_fd_sc_hd__nand2_1
XFILLER_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4043_ _4192_/B _4192_/C VGND VGND VPWR VPWR _4043_/Y sky130_fd_sc_hd__nand2_2
XFILLER_84_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5994_ hold448/X _6003_/A1 _6001_/S VGND VGND VPWR VPWR _7570_/D sky130_fd_sc_hd__mux2_1
X_4945_ _4946_/B _5261_/D VGND VGND VPWR VPWR _4945_/Y sky130_fd_sc_hd__nand2_1
XFILLER_177_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7664_ _7668_/CLK _7664_/D VGND VGND VPWR VPWR _7664_/Q sky130_fd_sc_hd__dfxtp_2
X_4876_ _4629_/Y _4953_/B _4950_/C _4901_/B VGND VGND VPWR VPWR _4900_/A sky130_fd_sc_hd__nand4bb_1
XFILLER_165_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3827_ _7589_/Q _6011_/A _3821_/X _3824_/X _3826_/X VGND VGND VPWR VPWR _3837_/A
+ sky130_fd_sc_hd__a2111o_1
X_6615_ _7335_/Q _6469_/X _6481_/X _7383_/Q VGND VGND VPWR VPWR _6615_/X sky130_fd_sc_hd__a22o_1
X_7595_ _7603_/CLK _7595_/D fanout611/X VGND VGND VPWR VPWR _7595_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_193_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6546_ _7396_/Q _6463_/X _6543_/X _6545_/X VGND VGND VPWR VPWR _6546_/X sky130_fd_sc_hd__a211o_1
XFILLER_146_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3758_ _7178_/Q _6038_/B hold98/A _4388_/A _7095_/Q VGND VGND VPWR VPWR _3758_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_165_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6477_ _6457_/X _6468_/X _6478_/C _6478_/D VGND VGND VPWR VPWR _6477_/X sky130_fd_sc_hd__and4bb_2
X_3689_ _7583_/Q _6002_/A _4481_/A _3567_/X _7343_/Q VGND VGND VPWR VPWR _3689_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_133_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5428_ _5605_/B _5428_/B _5428_/C VGND VGND VPWR VPWR _5428_/X sky130_fd_sc_hd__and3_1
Xoutput240 _4144_/X VGND VGND VPWR VPWR mgmt_gpio_out[36] sky130_fd_sc_hd__buf_12
Xoutput251 _4189_/X VGND VGND VPWR VPWR pad_flash_io0_do sky130_fd_sc_hd__buf_12
Xoutput262 _7261_/Q VGND VGND VPWR VPWR pll_div[0] sky130_fd_sc_hd__buf_12
XFILLER_160_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput273 _7134_/Q VGND VGND VPWR VPWR pll_trim[11] sky130_fd_sc_hd__buf_12
XFILLER_160_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput284 _7277_/Q VGND VGND VPWR VPWR pll_trim[21] sky130_fd_sc_hd__buf_12
XFILLER_59_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5359_ _4708_/X _5181_/C _5186_/B _5186_/C _5595_/A VGND VGND VPWR VPWR _5359_/X
+ sky130_fd_sc_hd__o2111a_1
Xoutput295 _7131_/Q VGND VGND VPWR VPWR pll_trim[8] sky130_fd_sc_hd__buf_12
XFILLER_58_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7029_ _7584_/CLK _7029_/D fanout613/X VGND VGND VPWR VPWR _7029_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_74_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire356 _3963_/Y VGND VGND VPWR VPWR _3964_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire367 _6659_/Y VGND VGND VPWR VPWR wire367/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4730_ _4629_/Y _4728_/Y _4729_/Y _4727_/Y VGND VGND VPWR VPWR _4733_/C sky130_fd_sc_hd__o211ai_1
XFILLER_21_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4661_ _5000_/C _4836_/A _4660_/C _5007_/D VGND VGND VPWR VPWR _4688_/C sky130_fd_sc_hd__o31a_2
X_6400_ _7232_/Q _6160_/D _6146_/C _6427_/B1 _7114_/Q VGND VGND VPWR VPWR _6400_/X
+ sky130_fd_sc_hd__a32o_1
X_3612_ input33/X _3544_/X _3565_/X _7329_/Q _3611_/X VGND VGND VPWR VPWR _3612_/X
+ sky130_fd_sc_hd__a221o_1
X_7380_ _7515_/CLK _7380_/D fanout621/X VGND VGND VPWR VPWR _7380_/Q sky130_fd_sc_hd__dfrtp_4
X_4592_ _5096_/A _4785_/C _4785_/A _4592_/D VGND VGND VPWR VPWR _4597_/C sky130_fd_sc_hd__nand4_4
XFILLER_128_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold904 _7688_/A VGND VGND VPWR VPWR hold904/X sky130_fd_sc_hd__dlygate4sd3_1
X_6331_ _7199_/Q _6159_/B _6407_/A3 _6145_/X _7682_/Q VGND VGND VPWR VPWR _6331_/X
+ sky130_fd_sc_hd__a32o_1
X_3543_ _3622_/A _3622_/B _3717_/B VGND VGND VPWR VPWR _3543_/X sky130_fd_sc_hd__and3_4
Xhold915 _5848_/X VGND VGND VPWR VPWR _7441_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold926 _7391_/Q VGND VGND VPWR VPWR hold926/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold937 _7556_/Q VGND VGND VPWR VPWR hold937/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold948 _5972_/X VGND VGND VPWR VPWR _7551_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6262_ _7527_/Q _6309_/B _6334_/C _6130_/X _7471_/Q VGND VGND VPWR VPWR _6262_/X
+ sky130_fd_sc_hd__a32o_1
Xhold959 _5720_/X VGND VGND VPWR VPWR _7327_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3474_ _3474_/A1 _3464_/X _3474_/B1 VGND VGND VPWR VPWR _6951_/D sky130_fd_sc_hd__a21o_1
XFILLER_115_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5213_ _4761_/A _5614_/B _5614_/D _5110_/C _4994_/X VGND VGND VPWR VPWR _5616_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_88_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6193_ _7444_/Q _6082_/B _6416_/C _6166_/C VGND VGND VPWR VPWR _6193_/X sky130_fd_sc_hd__o211a_1
XFILLER_142_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5144_ _4946_/A _5143_/X _5142_/Y VGND VGND VPWR VPWR _5147_/A sky130_fd_sc_hd__a21oi_1
Xhold1604 hold52/A VGND VGND VPWR VPWR _5613_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1615 _6940_/Q VGND VGND VPWR VPWR _4052_/B1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1626 _7562_/Q VGND VGND VPWR VPWR _5985_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1637 _4215_/Y VGND VGND VPWR VPWR _6960_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5075_ _5614_/C _5322_/A _5233_/C VGND VGND VPWR VPWR _5075_/X sky130_fd_sc_hd__and3_1
Xhold1648 _6978_/Q VGND VGND VPWR VPWR _4228_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_4026_ _7251_/Q _4541_/A hold70/A _3971_/X _4025_/X VGND VGND VPWR VPWR _4026_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_25_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5977_ hold341/X _6031_/A0 _5983_/S VGND VGND VPWR VPWR _5977_/X sky130_fd_sc_hd__mux2_1
X_4928_ _5181_/C _5452_/A _4957_/C _4934_/C VGND VGND VPWR VPWR _4930_/B sky130_fd_sc_hd__nand4_1
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7647_ _7662_/CLK _7647_/D _6911_/A VGND VGND VPWR VPWR _7647_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4859_ _4866_/A _4950_/C VGND VGND VPWR VPWR _4859_/Y sky130_fd_sc_hd__nand2_8
XFILLER_165_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7578_ _7586_/CLK _7578_/D fanout625/X VGND VGND VPWR VPWR _7578_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_153_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6529_ _7427_/Q _6444_/X _6452_/X _7579_/Q VGND VGND VPWR VPWR _6529_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_73_csclk _7095_/CLK VGND VGND VPWR VPWR _7286_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_87_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_11_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7252_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_157_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_26_csclk _7352_/CLK VGND VGND VPWR VPWR _7562_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_166_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5900_ hold783/X _5999_/A1 hold25/X VGND VGND VPWR VPWR _7487_/D sky130_fd_sc_hd__mux2_1
XFILLER_46_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6880_ _6891_/A _6911_/B VGND VGND VPWR VPWR _6880_/X sky130_fd_sc_hd__and2_1
XFILLER_74_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5831_ _5975_/B _5840_/A _6029_/B VGND VGND VPWR VPWR _5839_/S sky130_fd_sc_hd__and3_4
XFILLER_34_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5762_ hold164/X _5789_/A1 _5767_/S VGND VGND VPWR VPWR _5762_/X sky130_fd_sc_hd__mux2_1
X_7501_ _7557_/CLK _7501_/D fanout627/X VGND VGND VPWR VPWR _7501_/Q sky130_fd_sc_hd__dfrtp_4
X_4713_ _4712_/Y wire428/X _5595_/A VGND VGND VPWR VPWR _4722_/B sky130_fd_sc_hd__o21a_1
X_5693_ _6865_/A1 _5693_/A1 _5695_/S VGND VGND VPWR VPWR _5693_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7432_ _7432_/CLK _7432_/D fanout631/X VGND VGND VPWR VPWR _7432_/Q sky130_fd_sc_hd__dfrtp_4
X_4644_ _4637_/A _4595_/Y _4950_/D _5024_/C VGND VGND VPWR VPWR _5476_/B sky130_fd_sc_hd__o211a_4
XFILLER_190_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4575_ _4586_/A _4586_/B _4990_/A _5014_/D VGND VGND VPWR VPWR _4576_/B sky130_fd_sc_hd__nand4_1
Xhold701 _5677_/X VGND VGND VPWR VPWR _7292_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7363_ _7557_/CLK _7363_/D fanout631/X VGND VGND VPWR VPWR _7363_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_162_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold712 hold712/A VGND VGND VPWR VPWR hold712/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap420 _5407_/Y VGND VGND VPWR VPWR _5571_/B1 sky130_fd_sc_hd__clkbuf_1
Xmax_cap431 hold23/X VGND VGND VPWR VPWR _3673_/B sky130_fd_sc_hd__buf_4
Xhold723 _7177_/Q VGND VGND VPWR VPWR hold723/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3526_ hold69/X _3559_/B VGND VGND VPWR VPWR _3717_/B sky130_fd_sc_hd__and2b_4
X_6314_ _7369_/Q _6152_/X _6158_/X _7497_/Q _6313_/X VGND VGND VPWR VPWR _6314_/X
+ sky130_fd_sc_hd__a221o_1
Xhold734 _7034_/Q VGND VGND VPWR VPWR hold734/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 _6032_/X VGND VGND VPWR VPWR _7604_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7294_ _7294_/CLK _7294_/D fanout597/X VGND VGND VPWR VPWR _7294_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_89_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap453 _6113_/Y VGND VGND VPWR VPWR wire452/A sky130_fd_sc_hd__clkbuf_2
Xhold756 _5879_/X VGND VGND VPWR VPWR _7468_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap464 _4619_/Y VGND VGND VPWR VPWR _5244_/A1 sky130_fd_sc_hd__buf_2
Xhold767 _7336_/Q VGND VGND VPWR VPWR hold767/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap475 _6137_/X VGND VGND VPWR VPWR _6427_/B1 sky130_fd_sc_hd__buf_12
Xhold778 _4465_/X VGND VGND VPWR VPWR _7160_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6245_ _7494_/Q _6309_/B _6407_/A3 _6145_/X _7462_/Q VGND VGND VPWR VPWR _6245_/X
+ sky130_fd_sc_hd__a32o_1
Xhold789 _6009_/X VGND VGND VPWR VPWR _7584_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap497 _4948_/Y VGND VGND VPWR VPWR _5290_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6176_ _7419_/Q _6150_/X _6153_/X _7563_/Q _6175_/X VGND VGND VPWR VPWR _6176_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1401 _4206_/X VGND VGND VPWR VPWR _6958_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1412 _7264_/Q VGND VGND VPWR VPWR hold510/A sky130_fd_sc_hd__dlygate4sd3_1
X_5127_ _5127_/A _5127_/B _5127_/C VGND VGND VPWR VPWR _5127_/Y sky130_fd_sc_hd__nand3_1
Xhold1423 _6980_/Q VGND VGND VPWR VPWR _4232_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1434 _7266_/Q VGND VGND VPWR VPWR hold1434/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1445 _4409_/X VGND VGND VPWR VPWR _7108_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1456 hold11/A VGND VGND VPWR VPWR _6841_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1467 _7148_/Q VGND VGND VPWR VPWR _4451_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5058_ _5322_/C _5311_/C _5089_/A VGND VGND VPWR VPWR _5059_/C sky130_fd_sc_hd__and3_1
Xhold1478 _6941_/Q VGND VGND VPWR VPWR _4045_/B1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1489 _6919_/Q VGND VGND VPWR VPWR _4097_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_607 _5935_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4009_ _7184_/Q _4547_/A _5680_/A _3905_/X _7259_/Q VGND VGND VPWR VPWR _4009_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_44_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_618 _6853_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_629 _5233_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold50 hold50/A VGND VGND VPWR VPWR hold50/X sky130_fd_sc_hd__buf_8
Xhold61 hold61/A VGND VGND VPWR VPWR hold61/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold72 hold72/A VGND VGND VPWR VPWR hold72/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold83/A VGND VGND VPWR VPWR hold83/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 hold94/A VGND VGND VPWR VPWR hold94/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_3 _4319_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4360_ _5761_/A1 hold501/X _4363_/S VGND VGND VPWR VPWR _4360_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4291_ hold58/X hold50/X _4291_/S VGND VGND VPWR VPWR _4291_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6030_ _6039_/A1 hold503/X _6037_/S VGND VGND VPWR VPWR _7602_/D sky130_fd_sc_hd__mux2_1
XFILLER_140_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6932_ _4172_/B2 _6932_/D _6887_/X VGND VGND VPWR VPWR hold4/A sky130_fd_sc_hd__dfrtp_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6863_ hold678/X _6863_/A1 _6866_/S VGND VGND VPWR VPWR _6863_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5814_ _6003_/A1 hold792/X _5821_/S VGND VGND VPWR VPWR _5814_/X sky130_fd_sc_hd__mux2_1
X_6794_ _7255_/Q _6460_/X _6486_/X _7105_/Q _6793_/X VGND VGND VPWR VPWR _6794_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_179_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5745_ _6006_/A1 _5745_/A1 _5749_/S VGND VGND VPWR VPWR _7349_/D sky130_fd_sc_hd__mux2_1
XFILLER_157_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5676_ _5676_/A0 hold50/X _5677_/S VGND VGND VPWR VPWR hold51/A sky130_fd_sc_hd__mux2_1
XFILLER_175_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7415_ _7599_/CLK _7415_/D fanout629/X VGND VGND VPWR VPWR _7415_/Q sky130_fd_sc_hd__dfrtp_4
X_4627_ _4959_/C _4948_/B VGND VGND VPWR VPWR _5407_/B sky130_fd_sc_hd__nand2b_2
XFILLER_135_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold520 hold520/A VGND VGND VPWR VPWR hold520/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4558_ hold541/X _4564_/A1 _4558_/S VGND VGND VPWR VPWR _4558_/X sky130_fd_sc_hd__mux2_1
X_7346_ _7518_/CLK _7346_/D fanout627/X VGND VGND VPWR VPWR _7346_/Q sky130_fd_sc_hd__dfstp_1
Xhold531 _4544_/X VGND VGND VPWR VPWR _7226_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold542 _4558_/X VGND VGND VPWR VPWR _7238_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold553 _7592_/Q VGND VGND VPWR VPWR hold553/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 _7077_/Q VGND VGND VPWR VPWR hold564/X sky130_fd_sc_hd__dlygate4sd3_1
X_3509_ hold127/X _4229_/S VGND VGND VPWR VPWR _3509_/Y sky130_fd_sc_hd__nand2b_2
Xhold575 _7528_/Q VGND VGND VPWR VPWR hold575/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7277_ _7614_/CLK hold86/X fanout604/X VGND VGND VPWR VPWR _7277_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_103_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4489_ hold393/X _5761_/A1 _4492_/S VGND VGND VPWR VPWR _4489_/X sky130_fd_sc_hd__mux2_1
Xhold586 _4543_/X VGND VGND VPWR VPWR _7225_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 _4486_/X VGND VGND VPWR VPWR _7178_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6228_ _6686_/S _6228_/A2 _6226_/X _6227_/X VGND VGND VPWR VPWR _6228_/X sky130_fd_sc_hd__a22o_1
XFILLER_103_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6159_ _6159_/A _6159_/B _6392_/B VGND VGND VPWR VPWR _6159_/X sky130_fd_sc_hd__and3_4
Xhold1220 _4448_/A1 VGND VGND VPWR VPWR hold698/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1231 _4446_/A1 VGND VGND VPWR VPWR hold843/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1242 _7542_/Q VGND VGND VPWR VPWR _5962_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1253 _4534_/X VGND VGND VPWR VPWR _7218_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1264 _7605_/Q VGND VGND VPWR VPWR hold1264/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1275 _4542_/X VGND VGND VPWR VPWR _7224_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1286 _5755_/X VGND VGND VPWR VPWR _7358_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_404 _6469_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1297 _7398_/Q VGND VGND VPWR VPWR hold625/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_415 _6157_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_426 _6158_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_437 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_448 _6452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_459 _6486_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput140 wb_dat_i[17] VGND VGND VPWR VPWR _6834_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_95_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput151 wb_dat_i[27] VGND VGND VPWR VPWR _6839_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput162 wb_dat_i[8] VGND VGND VPWR VPWR _6830_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3860_ _7412_/Q _5813_/A _4358_/A _7068_/Q _3859_/X VGND VGND VPWR VPWR _3860_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_177_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3791_ _7413_/Q _5840_/A _5957_/B _3525_/X _7397_/Q VGND VGND VPWR VPWR _3791_/X
+ sky130_fd_sc_hd__a32o_1
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5530_ _5621_/B _5530_/B _5530_/C _5530_/D VGND VGND VPWR VPWR _5530_/X sky130_fd_sc_hd__and4_1
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5461_ _4629_/Y _4674_/Y _5011_/C _5011_/B _5585_/A1 VGND VGND VPWR VPWR _5461_/X
+ sky130_fd_sc_hd__a311o_1
X_4412_ _4559_/B _4529_/B _5680_/C VGND VGND VPWR VPWR _4417_/S sky130_fd_sc_hd__and3_2
X_7200_ _7255_/CLK _7200_/D fanout618/X VGND VGND VPWR VPWR _7200_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_145_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5392_ _5389_/X _5392_/B _5392_/C _5392_/D VGND VGND VPWR VPWR _5393_/C sky130_fd_sc_hd__and4b_1
XFILLER_126_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4343_ _4556_/A1 hold525/X _4345_/S VGND VGND VPWR VPWR _4343_/X sky130_fd_sc_hd__mux2_1
X_7131_ _7289_/CLK _7131_/D fanout598/X VGND VGND VPWR VPWR _7131_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7062_ _7686_/CLK _7062_/D _6891_/A VGND VGND VPWR VPWR _7062_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_86_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4274_ _4273_/X hold989/X _4274_/S VGND VGND VPWR VPWR _4274_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6013_ hold5/X _6013_/A1 _6019_/S VGND VGND VPWR VPWR hold6/A sky130_fd_sc_hd__mux2_1
XFILLER_39_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6915_ _4183_/A1 _6915_/D _6870_/X VGND VGND VPWR VPWR _6915_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_63_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6846_ _6971_/Q _6846_/A2 _6846_/B1 wire537/X _6845_/X VGND VGND VPWR VPWR _6846_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_50_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6777_ _7162_/Q _6456_/X _6486_/X _7104_/Q _6776_/X VGND VGND VPWR VPWR _6784_/A
+ sky130_fd_sc_hd__a221o_1
X_3989_ _7194_/Q _3704_/X _3986_/X _3987_/X _3988_/X VGND VGND VPWR VPWR _3989_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_183_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5728_ hold229/X _5935_/A1 _5731_/S VGND VGND VPWR VPWR _5728_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5659_ _5682_/A _5669_/B _5659_/C _5686_/D VGND VGND VPWR VPWR _5660_/S sky130_fd_sc_hd__and4_1
XFILLER_136_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold350 _4385_/X VGND VGND VPWR VPWR _7088_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold361 _7166_/Q VGND VGND VPWR VPWR hold361/X sky130_fd_sc_hd__dlygate4sd3_1
X_7329_ _7435_/CLK _7329_/D fanout623/X VGND VGND VPWR VPWR _7329_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_104_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold372 _5843_/X VGND VGND VPWR VPWR _7436_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold383 _7524_/Q VGND VGND VPWR VPWR hold383/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold394 _4489_/X VGND VGND VPWR VPWR _7180_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1050 _7204_/Q VGND VGND VPWR VPWR _4518_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1061 _7061_/Q VGND VGND VPWR VPWR _4353_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1072 _7707_/A VGND VGND VPWR VPWR _4299_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1083 _7397_/Q VGND VGND VPWR VPWR _5799_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1094 _7234_/Q VGND VGND VPWR VPWR _4554_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_201 _7295_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_212 _7482_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_223 _7160_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_234 hold92/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_245 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_256 _4199_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_267 _7714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_278 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_289 _7713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4961_ _4961_/A _5452_/B VGND VGND VPWR VPWR _5570_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6700_ _6700_/A _6700_/B _6700_/C _6700_/D VGND VGND VPWR VPWR _6700_/Y sky130_fd_sc_hd__nor4_2
X_3912_ input35/X _3573_/X _3713_/X _7097_/Q _3911_/X VGND VGND VPWR VPWR _3912_/X
+ sky130_fd_sc_hd__a221o_1
X_7680_ _7680_/CLK _7680_/D _6815_/A VGND VGND VPWR VPWR _7680_/Q sky130_fd_sc_hd__dfrtp_2
X_4892_ _4901_/B _4892_/B _5389_/B _4950_/C VGND VGND VPWR VPWR _4892_/Y sky130_fd_sc_hd__nand4_1
XFILLER_189_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6631_ _7503_/Q _6486_/X _6628_/X _6630_/X VGND VGND VPWR VPWR _6632_/C sky130_fd_sc_hd__a211o_1
X_3843_ _5682_/A _5682_/B _5682_/C VGND VGND VPWR VPWR _3843_/X sky130_fd_sc_hd__and3_1
XFILLER_32_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3774_ _3774_/A _3774_/B _3774_/C _3774_/D VGND VGND VPWR VPWR _3774_/Y sky130_fd_sc_hd__nor4_1
X_6562_ _7509_/Q _6562_/B _6562_/C VGND VGND VPWR VPWR _6562_/X sky130_fd_sc_hd__and3_1
XFILLER_9_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5513_ _4756_/Y _5611_/A2 _5285_/X _5514_/B _5514_/D VGND VGND VPWR VPWR _5603_/A
+ sky130_fd_sc_hd__o311a_1
X_6493_ _7594_/Q _6474_/B _6474_/C _7370_/Q _6492_/X VGND VGND VPWR VPWR _6493_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_157_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5444_ _5009_/Y _5440_/Y _5256_/A _4904_/D _5392_/B VGND VGND VPWR VPWR _5524_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_105_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5375_ _5375_/A _5375_/B _5375_/C VGND VGND VPWR VPWR _5376_/A sky130_fd_sc_hd__and3_1
XFILLER_114_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7114_ _7686_/CLK _7114_/D fanout599/X VGND VGND VPWR VPWR _7114_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_113_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4326_ hold505/X _5673_/A1 _4327_/S VGND VGND VPWR VPWR _7039_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4257_ _4312_/A1 hold102/X _4257_/S VGND VGND VPWR VPWR _4257_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7045_ _7398_/CLK _7045_/D fanout619/X VGND VGND VPWR VPWR _7045_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_86_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4188_ _4188_/A VGND VGND VPWR VPWR _4188_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6829_ _6828_/X _6858_/D _6829_/C _6829_/D VGND VGND VPWR VPWR _6853_/S sky130_fd_sc_hd__and4b_4
XFILLER_10_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold180 _7448_/Q VGND VGND VPWR VPWR hold180/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 _7135_/Q VGND VGND VPWR VPWR hold191/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3490_ _3508_/S _4067_/A VGND VGND VPWR VPWR _3490_/X sky130_fd_sc_hd__and2_1
XFILLER_155_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5160_ _4743_/C _5358_/B _4946_/A _4722_/A VGND VGND VPWR VPWR _5160_/X sky130_fd_sc_hd__a31o_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4111_ _4586_/C _4586_/D _4585_/A _4585_/B VGND VGND VPWR VPWR _4115_/B sky130_fd_sc_hd__nor4_1
XFILLER_96_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5091_ _5092_/B _5091_/B VGND VGND VPWR VPWR _5121_/D sky130_fd_sc_hd__nand2_1
XFILLER_96_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4042_ _6913_/Q _4193_/B _4192_/C VGND VGND VPWR VPWR _4085_/B sky130_fd_sc_hd__and3_2
XFILLER_110_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5993_ _5993_/A _5993_/B _6038_/C VGND VGND VPWR VPWR _6001_/S sky130_fd_sc_hd__and3_4
XFILLER_18_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4944_ _4767_/Y _4939_/Y _4943_/Y _4941_/Y VGND VGND VPWR VPWR _4947_/B sky130_fd_sc_hd__o211ai_1
XFILLER_33_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7663_ _7668_/CLK _7663_/D _6815_/A VGND VGND VPWR VPWR _7663_/Q sky130_fd_sc_hd__dfrtp_1
X_4875_ _4709_/Y _4862_/Y _4871_/X _4874_/Y VGND VGND VPWR VPWR _4875_/X sky130_fd_sc_hd__o31a_1
X_6614_ _7447_/Q _6460_/X _6465_/X _7351_/Q _6613_/X VGND VGND VPWR VPWR _6614_/X
+ sky130_fd_sc_hd__a221o_1
X_3826_ _7613_/Q _3580_/X _3704_/X _7197_/Q _3825_/X VGND VGND VPWR VPWR _3826_/X
+ sky130_fd_sc_hd__a221o_1
X_7594_ _7602_/CLK _7594_/D fanout615/X VGND VGND VPWR VPWR _7594_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_193_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6545_ _7356_/Q _6454_/X _6469_/X _7332_/Q _6544_/X VGND VGND VPWR VPWR _6545_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3757_ _7566_/Q _3554_/X _4293_/S _4172_/B2 _3756_/X VGND VGND VPWR VPWR _3757_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_192_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6476_ _6444_/X _6454_/X _6476_/C _6476_/D VGND VGND VPWR VPWR _6478_/D sky130_fd_sc_hd__and4bb_1
X_3688_ _7383_/Q _5777_/A _3581_/X _7367_/Q _3687_/X VGND VGND VPWR VPWR _3691_/C
+ sky130_fd_sc_hd__a221o_1
Xoutput230 _7707_/X VGND VGND VPWR VPWR mgmt_gpio_out[27] sky130_fd_sc_hd__buf_12
X_5427_ _5285_/X _4993_/Y _4960_/Y _5604_/B1 _4991_/Y VGND VGND VPWR VPWR _5428_/C
+ sky130_fd_sc_hd__a311o_1
Xoutput241 _4143_/X VGND VGND VPWR VPWR mgmt_gpio_out[37] sky130_fd_sc_hd__buf_12
Xoutput252 _4186_/A VGND VGND VPWR VPWR pad_flash_io0_ieb sky130_fd_sc_hd__buf_12
Xoutput263 _7262_/Q VGND VGND VPWR VPWR pll_div[1] sky130_fd_sc_hd__buf_12
Xoutput274 _7135_/Q VGND VGND VPWR VPWR pll_trim[12] sky130_fd_sc_hd__buf_12
XFILLER_160_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput285 _7278_/Q VGND VGND VPWR VPWR pll_trim[22] sky130_fd_sc_hd__buf_12
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5358_ _5358_/A _5358_/B _5595_/C VGND VGND VPWR VPWR _5358_/X sky130_fd_sc_hd__and3_1
Xoutput296 _7132_/Q VGND VGND VPWR VPWR pll_trim[9] sky130_fd_sc_hd__buf_12
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4309_ _5935_/A1 hold241/X _4312_/S VGND VGND VPWR VPWR _4309_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5289_ _5311_/A _5313_/B _5092_/B _5110_/C _5091_/B VGND VGND VPWR VPWR _5289_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7028_ _7569_/CLK _7028_/D fanout613/X VGND VGND VPWR VPWR _7028_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire346 _3901_/Y VGND VGND VPWR VPWR _3902_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_183_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire357 _3815_/Y VGND VGND VPWR VPWR wire357/X sky130_fd_sc_hd__clkbuf_1
Xwire368 _6532_/Y VGND VGND VPWR VPWR wire368/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4660_ _5000_/C _4836_/A _4660_/C VGND VGND VPWR VPWR _4660_/Y sky130_fd_sc_hd__nor3_2
XFILLER_187_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3611_ _7369_/Q _5975_/B _5759_/B _3610_/X VGND VGND VPWR VPWR _3611_/X sky130_fd_sc_hd__a31o_1
XFILLER_175_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4591_ _4785_/C _4785_/A _4592_/D _5096_/A VGND VGND VPWR VPWR _4597_/B sky130_fd_sc_hd__a31o_2
X_6330_ _7229_/Q _6160_/D _6427_/A3 _6427_/B1 _7111_/Q VGND VGND VPWR VPWR _6330_/X
+ sky130_fd_sc_hd__a32o_1
X_3542_ hold74/A _5686_/B _4535_/B VGND VGND VPWR VPWR _3542_/X sky130_fd_sc_hd__and3_2
Xhold905 _5670_/X VGND VGND VPWR VPWR _7286_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold916 _7353_/Q VGND VGND VPWR VPWR hold916/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold927 _5792_/X VGND VGND VPWR VPWR _7391_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold938 _5978_/X VGND VGND VPWR VPWR _7556_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3473_ _6886_/A _6911_/B VGND VGND VPWR VPWR _3473_/X sky130_fd_sc_hd__and2_1
X_6261_ _7479_/Q _6133_/X _6138_/X _7359_/Q _6260_/X VGND VGND VPWR VPWR _6261_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold949 _7694_/A VGND VGND VPWR VPWR hold949/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5212_ _5614_/B _5614_/D VGND VGND VPWR VPWR _5212_/Y sky130_fd_sc_hd__nand2_1
XFILLER_170_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6192_ _6187_/X _6189_/X _6191_/X _6159_/B VGND VGND VPWR VPWR _6192_/Y sky130_fd_sc_hd__o31ai_4
X_5143_ _5143_/A _5143_/B _5512_/B VGND VGND VPWR VPWR _5143_/X sky130_fd_sc_hd__and3_1
XFILLER_111_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1605 _7039_/Q VGND VGND VPWR VPWR hold505/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1616 _6928_/Q VGND VGND VPWR VPWR _4078_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5074_ _5074_/A _5074_/B VGND VGND VPWR VPWR _5076_/C sky130_fd_sc_hd__nand2_1
Xhold1627 _7628_/Q VGND VGND VPWR VPWR _6086_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold1638 _6965_/Q VGND VGND VPWR VPWR hold1638/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1649 _7142_/Q VGND VGND VPWR VPWR _4132_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4025_ _7179_/Q _4487_/A _4511_/C _3567_/X _7338_/Q VGND VGND VPWR VPWR _4025_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_56_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5976_ hold513/X _6039_/A1 _5983_/S VGND VGND VPWR VPWR _7554_/D sky130_fd_sc_hd__mux2_1
XFILLER_52_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7715_ _7715_/A VGND VGND VPWR VPWR _7715_/X sky130_fd_sc_hd__buf_2
X_4927_ _4927_/A _4927_/B _4927_/C VGND VGND VPWR VPWR _4930_/A sky130_fd_sc_hd__nor3_1
XFILLER_100_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7646_ _7662_/CLK _7646_/D fanout597/X VGND VGND VPWR VPWR _7646_/Q sky130_fd_sc_hd__dfrtp_1
X_4858_ _4858_/A _4950_/C _4950_/D VGND VGND VPWR VPWR _5261_/D sky130_fd_sc_hd__and3_4
XFILLER_193_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3809_ _7597_/Q _6020_/A _4481_/A _3546_/X _7533_/Q VGND VGND VPWR VPWR _3809_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_20_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7577_ _7609_/CLK _7577_/D fanout614/X VGND VGND VPWR VPWR _7577_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4789_ _4781_/Y _4884_/A _4788_/X VGND VGND VPWR VPWR _4858_/A sky130_fd_sc_hd__a21oi_2
XFILLER_180_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6528_ _7355_/Q _6454_/X _6459_/X _7451_/Q VGND VGND VPWR VPWR _6528_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6459_ _6645_/B _6563_/C _6645_/C VGND VGND VPWR VPWR _6459_/X sky130_fd_sc_hd__and3_4
XFILLER_69_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5830_ hold869/X _6046_/A1 _5830_/S VGND VGND VPWR VPWR _5830_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5761_ hold305/X _5761_/A1 _5767_/S VGND VGND VPWR VPWR _5761_/X sky130_fd_sc_hd__mux2_1
X_7500_ _7580_/CLK _7500_/D fanout607/X VGND VGND VPWR VPWR _7500_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_91_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4712_ _4570_/Y _4706_/Y _4710_/Y _4704_/C VGND VGND VPWR VPWR _4712_/Y sky130_fd_sc_hd__o22ai_1
X_5692_ _5789_/A1 hold483/X _5695_/S VGND VGND VPWR VPWR _5692_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7431_ _7432_/CLK _7431_/D fanout631/X VGND VGND VPWR VPWR _7431_/Q sky130_fd_sc_hd__dfrtp_1
X_4643_ _4637_/A _4884_/A _4572_/X VGND VGND VPWR VPWR _4799_/A sky130_fd_sc_hd__a21oi_2
XFILLER_147_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7362_ _7518_/CLK hold16/X fanout626/X VGND VGND VPWR VPWR _7362_/Q sky130_fd_sc_hd__dfstp_1
X_4574_ _4586_/C _4586_/D _4585_/A _4585_/B VGND VGND VPWR VPWR _4576_/A sky130_fd_sc_hd__nand4_1
Xhold702 _7260_/Q VGND VGND VPWR VPWR hold702/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 hold713/A VGND VGND VPWR VPWR wb_dat_o[5] sky130_fd_sc_hd__buf_12
Xmax_cap432 hold96/X VGND VGND VPWR VPWR _3559_/B sky130_fd_sc_hd__buf_4
X_6313_ _7561_/Q _6131_/B _6432_/A3 _6153_/X _7569_/Q VGND VGND VPWR VPWR _6313_/X
+ sky130_fd_sc_hd__a32o_1
Xhold724 _4485_/X VGND VGND VPWR VPWR _7177_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap443 _5358_/A VGND VGND VPWR VPWR _5153_/A sky130_fd_sc_hd__clkbuf_2
X_3525_ hold73/A _5939_/B _5768_/C VGND VGND VPWR VPWR _3525_/X sky130_fd_sc_hd__and3_4
Xhold735 _4320_/X VGND VGND VPWR VPWR _7034_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7293_ _7293_/CLK _7293_/D fanout597/X VGND VGND VPWR VPWR _7293_/Q sky130_fd_sc_hd__dfrtp_1
Xhold746 _7316_/Q VGND VGND VPWR VPWR hold746/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap454 wire455/X VGND VGND VPWR VPWR _6302_/B1 sky130_fd_sc_hd__clkbuf_2
Xhold757 _7122_/Q VGND VGND VPWR VPWR hold757/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold768 _5730_/X VGND VGND VPWR VPWR _7336_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold779 _7319_/Q VGND VGND VPWR VPWR hold779/X sky130_fd_sc_hd__dlygate4sd3_1
X_6244_ _7510_/Q _6136_/X _6144_/X _7542_/Q _6239_/X VGND VGND VPWR VPWR _6244_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3456_ _7333_/Q VGND VGND VPWR VPWR _3456_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6175_ _7499_/Q _6131_/B _6127_/X _6130_/X _7467_/Q VGND VGND VPWR VPWR _6175_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_97_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1402 _7669_/Q VGND VGND VPWR VPWR _6821_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1413 _7670_/Q VGND VGND VPWR VPWR _6822_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5126_ _5401_/A _5107_/B _5124_/Y _5125_/X VGND VGND VPWR VPWR _5127_/A sky130_fd_sc_hd__a22oi_1
Xhold1424 _7284_/Q VGND VGND VPWR VPWR _5665_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1435 _7386_/Q VGND VGND VPWR VPWR hold428/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1446 _7150_/Q VGND VGND VPWR VPWR _4453_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1457 _7655_/Q VGND VGND VPWR VPWR _6661_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1468 _6921_/Q VGND VGND VPWR VPWR _4053_/A sky130_fd_sc_hd__dlygate4sd3_1
X_5057_ _5011_/A _4823_/Y _4998_/Y _4996_/Y _5056_/Y VGND VGND VPWR VPWR _5059_/D
+ sky130_fd_sc_hd__o311ai_1
Xhold1479 _4045_/X VGND VGND VPWR VPWR _4046_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_608 _6039_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4008_ _7066_/Q _5680_/A _4487_/B _5777_/A _7378_/Q VGND VGND VPWR VPWR _4008_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_619 _5007_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5959_ hold197/X _6031_/A0 _5965_/S VGND VGND VPWR VPWR _5959_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7629_ _4167_/A1 _7629_/D fanout620/X VGND VGND VPWR VPWR _7629_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold40 hold40/A VGND VGND VPWR VPWR hold40/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A VGND VGND VPWR VPWR hold51/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A VGND VGND VPWR VPWR hold62/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hold73/A VGND VGND VPWR VPWR hold73/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 hold90/X VGND VGND VPWR VPWR hold84/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 hold95/A VGND VGND VPWR VPWR hold95/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_4 _4474_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4290_ _4289_/X _4290_/A1 _4294_/S VGND VGND VPWR VPWR _4290_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6931_ _7258_/CLK _6931_/D _6886_/X VGND VGND VPWR VPWR hold32/A sky130_fd_sc_hd__dfrtp_1
XFILLER_19_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6862_ _6862_/A0 _6862_/A1 _6866_/S VGND VGND VPWR VPWR _6862_/X sky130_fd_sc_hd__mux2_1
XFILLER_81_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5813_ _5813_/A hold29/X VGND VGND VPWR VPWR _5821_/S sky130_fd_sc_hd__nand2_8
XFILLER_50_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6793_ _7203_/Q _6694_/B _6694_/C _6474_/C _7060_/Q VGND VGND VPWR VPWR _6793_/X
+ sky130_fd_sc_hd__a32o_1
X_5744_ _5843_/A1 hold319/X _5749_/S VGND VGND VPWR VPWR _5744_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5675_ hold92/X hold85/X _5677_/S VGND VGND VPWR VPWR hold93/A sky130_fd_sc_hd__mux2_1
XFILLER_148_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_72_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7462_/CLK sky130_fd_sc_hd__clkbuf_16
X_7414_ _7518_/CLK _7414_/D fanout625/X VGND VGND VPWR VPWR _7414_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_175_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4626_ _4959_/C _4948_/B VGND VGND VPWR VPWR _5404_/A sky130_fd_sc_hd__and2b_4
XFILLER_190_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold510 hold510/A VGND VGND VPWR VPWR hold510/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7345_ _7435_/CLK _7345_/D fanout623/X VGND VGND VPWR VPWR _7345_/Q sky130_fd_sc_hd__dfrtp_1
Xhold521 _7513_/Q VGND VGND VPWR VPWR hold521/X sky130_fd_sc_hd__dlygate4sd3_1
X_4557_ _4557_/A0 _6865_/A1 _4558_/S VGND VGND VPWR VPWR _4557_/X sky130_fd_sc_hd__mux2_1
Xhold532 _7279_/Q VGND VGND VPWR VPWR hold532/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 _7110_/Q VGND VGND VPWR VPWR hold543/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold554 _6018_/X VGND VGND VPWR VPWR _7592_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3508_ input58/X hold21/X _3508_/S VGND VGND VPWR VPWR hold22/A sky130_fd_sc_hd__mux2_2
XFILLER_104_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold565 _4372_/X VGND VGND VPWR VPWR _7077_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7276_ _7286_/CLK _7276_/D fanout598/X VGND VGND VPWR VPWR _7276_/Q sky130_fd_sc_hd__dfstp_1
Xhold576 _5946_/X VGND VGND VPWR VPWR _7528_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4488_ _4488_/A0 _6012_/A0 _4492_/S VGND VGND VPWR VPWR _4488_/X sky130_fd_sc_hd__mux2_1
Xhold587 _7473_/Q VGND VGND VPWR VPWR hold587/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold598 _7243_/Q VGND VGND VPWR VPWR hold598/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6227_ _7317_/Q _6082_/Y _6686_/S VGND VGND VPWR VPWR _6227_/X sky130_fd_sc_hd__o21ba_1
XFILLER_104_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3439_ _7477_/Q VGND VGND VPWR VPWR _3439_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6158_ _6151_/B _6392_/B _6166_/B _6158_/D VGND VGND VPWR VPWR _6158_/X sky130_fd_sc_hd__and4b_4
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1210 _4456_/A1 VGND VGND VPWR VPWR hold651/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1221 _4460_/A1 VGND VGND VPWR VPWR hold712/A sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_10_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7255_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1232 _4450_/A1 VGND VGND VPWR VPWR hold784/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1243 _7185_/Q VGND VGND VPWR VPWR _4495_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5109_ _5109_/A _5131_/B _5291_/C _5452_/B VGND VGND VPWR VPWR _5121_/B sky130_fd_sc_hd__nand4_1
Xhold1254 _7052_/Q VGND VGND VPWR VPWR _4342_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_6089_ _6469_/A _6109_/B VGND VGND VPWR VPWR _6089_/Y sky130_fd_sc_hd__nand2b_1
Xhold1265 _6033_/X VGND VGND VPWR VPWR _7605_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1276 _7597_/Q VGND VGND VPWR VPWR hold1276/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1287 _7233_/Q VGND VGND VPWR VPWR hold247/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1298 _7395_/Q VGND VGND VPWR VPWR hold976/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_405 _6469_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_416 _6516_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_427 _6158_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_438 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7210_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_449 _6454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput130 wb_adr_i[9] VGND VGND VPWR VPWR _4586_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput141 wb_dat_i[18] VGND VGND VPWR VPWR _6837_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput152 wb_dat_i[28] VGND VGND VPWR VPWR _6843_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput163 wb_dat_i[9] VGND VGND VPWR VPWR _6833_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_726 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3790_ _7349_/Q _5741_/A _4358_/A _7069_/Q _3789_/X VGND VGND VPWR VPWR _3790_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_188_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5460_ _5429_/D _5407_/Y _4850_/X _5280_/X _5409_/X VGND VGND VPWR VPWR _5460_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4411_ hold543/X _4564_/A1 _4411_/S VGND VGND VPWR VPWR _4411_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5391_ _4871_/X _4889_/Y _5015_/Y _5088_/Y _5390_/X VGND VGND VPWR VPWR _5392_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_132_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7130_ _7130_/CLK _7130_/D _6903_/A VGND VGND VPWR VPWR _7130_/Q sky130_fd_sc_hd__dfrtp_1
X_4342_ _5869_/A1 _4342_/A1 _4345_/S VGND VGND VPWR VPWR _4342_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7061_ _7242_/CLK _7061_/D fanout616/X VGND VGND VPWR VPWR _7061_/Q sky130_fd_sc_hd__dfrtp_2
X_4273_ hold734/X _5991_/A1 _4275_/S VGND VGND VPWR VPWR _4273_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6012_ _6012_/A0 _6012_/A1 _6019_/S VGND VGND VPWR VPWR _7586_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
.ends

