magic
tech sky130A
magscale 1 2
timestamp 1637704106
<< error_p >>
rect 111554 1006757 112632 1006758
rect 111554 1006005 111555 1006757
rect 112631 1006005 112632 1006757
rect 111554 1006004 112632 1006005
rect 162954 1006757 164032 1006758
rect 162954 1006005 162955 1006757
rect 164031 1006005 164032 1006757
rect 162954 1006004 164032 1006005
rect 214354 1006757 215432 1006758
rect 214354 1006005 214355 1006757
rect 215431 1006005 215432 1006757
rect 214354 1006004 215432 1006005
rect 265754 1006757 266832 1006758
rect 265754 1006005 265755 1006757
rect 266831 1006005 266832 1006757
rect 265754 1006004 266832 1006005
rect 317354 1006757 318432 1006758
rect 317354 1006005 317355 1006757
rect 318431 1006005 318432 1006757
rect 317354 1006004 318432 1006005
rect 367754 1006757 368832 1006758
rect 367754 1006005 367755 1006757
rect 368831 1006005 368832 1006757
rect 367754 1006004 368832 1006005
rect 435154 1006757 436232 1006758
rect 435154 1006005 435155 1006757
rect 436231 1006005 436232 1006757
rect 435154 1006004 436232 1006005
rect 512154 1006757 513232 1006758
rect 512154 1006005 512155 1006757
rect 513231 1006005 513232 1006757
rect 512154 1006004 513232 1006005
rect 563554 1006757 564632 1006758
rect 563554 1006005 563555 1006757
rect 564631 1006005 564632 1006757
rect 563554 1006004 564632 1006005
rect 109980 1000219 111064 1000220
rect 109980 999459 109981 1000219
rect 111063 999459 111064 1000219
rect 109980 999458 111064 999459
rect 161380 1000219 162464 1000220
rect 161380 999459 161381 1000219
rect 162463 999459 162464 1000219
rect 161380 999458 162464 999459
rect 212780 1000219 213864 1000220
rect 212780 999459 212781 1000219
rect 213863 999459 213864 1000219
rect 212780 999458 213864 999459
rect 264180 1000219 265264 1000220
rect 264180 999459 264181 1000219
rect 265263 999459 265264 1000219
rect 264180 999458 265264 999459
rect 315780 1000219 316864 1000220
rect 315780 999459 315781 1000219
rect 316863 999459 316864 1000219
rect 315780 999458 316864 999459
rect 366180 1000219 367264 1000220
rect 366180 999459 366181 1000219
rect 367263 999459 367264 1000219
rect 366180 999458 367264 999459
rect 433580 1000219 434664 1000220
rect 433580 999459 433581 1000219
rect 434663 999459 434664 1000219
rect 433580 999458 434664 999459
rect 510580 1000219 511664 1000220
rect 510580 999459 510581 1000219
rect 511663 999459 511664 1000219
rect 510580 999458 511664 999459
rect 561980 1000219 563064 1000220
rect 561980 999459 561981 1000219
rect 563063 999459 563064 1000219
rect 561980 999458 563064 999459
rect 670976 992506 673264 992530
rect 670976 990378 671000 992506
rect 673240 990378 673264 992506
rect 670976 990354 673264 990378
rect 41034 986424 43574 986448
rect 41034 985902 41058 986424
rect 43550 985902 43574 986424
rect 41034 985878 43574 985902
rect 44242 985474 46772 985498
rect 44242 984942 44266 985474
rect 46748 984942 46772 985474
rect 44242 984918 46772 984942
rect 670858 984512 673384 984536
rect 670858 983974 670882 984512
rect 673360 983974 673384 984512
rect 670858 983950 673384 983974
rect 674056 983550 676582 983574
rect 674056 983012 674080 983550
rect 676558 983012 676582 983550
rect 674056 982988 676582 983012
rect 61424 953079 61962 953080
rect 44278 953006 46734 953030
rect 44278 952000 44302 953006
rect 46710 952000 46734 953006
rect 44278 951976 46734 952000
rect 61424 951961 61425 953079
rect 61961 951961 61962 953079
rect 61424 951960 61962 951961
rect 60460 951487 60998 951488
rect 41068 951424 43524 951448
rect 41068 951330 41092 951424
rect 43500 951330 43524 951424
rect 60460 950369 60461 951487
rect 60997 950369 60998 951487
rect 60460 950368 60998 950369
rect 63350 949631 63872 949632
rect 63350 948523 63351 949631
rect 63871 948523 63872 949631
rect 63350 948522 63872 948523
rect 62382 948123 62904 948124
rect 62382 947015 62383 948123
rect 62903 947015 62904 948123
rect 62382 947014 62904 947015
rect 30820 946631 31574 946632
rect 30820 945555 30821 946631
rect 31573 945555 31574 946631
rect 30820 945554 31574 945555
rect 650654 946345 651202 946346
rect 650654 945225 650655 946345
rect 651201 945225 651202 946345
rect 650654 945224 651202 945225
rect 37358 945063 38120 945064
rect 37358 943981 37359 945063
rect 38119 943981 38120 945063
rect 37358 943980 38120 943981
rect 651602 944749 652170 944750
rect 651602 943613 651603 944749
rect 652169 943613 652170 944749
rect 651602 943612 652170 943613
rect 686002 943031 686756 943032
rect 686002 941955 686003 943031
rect 686755 941955 686756 943031
rect 686002 941954 686756 941955
rect 679456 941463 680218 941464
rect 679456 940381 679457 941463
rect 680217 940381 680218 941463
rect 679456 940380 680218 940381
rect 650654 901145 651202 901146
rect 650654 900025 650655 901145
rect 651201 900025 651202 901145
rect 674734 901088 675740 901112
rect 674734 900098 674758 901088
rect 675716 900098 675740 901088
rect 674734 900074 675740 900098
rect 650654 900024 651202 900025
rect 651602 899549 652170 899550
rect 651602 898413 651603 899549
rect 652169 898413 652170 899549
rect 671566 899480 672596 899504
rect 671566 898490 671590 899480
rect 672572 898490 672596 899480
rect 671566 898466 672596 898490
rect 651602 898412 652170 898413
rect 650654 856145 651202 856146
rect 650654 855025 650655 856145
rect 651201 855025 651202 856145
rect 674116 856092 675180 856116
rect 674116 855076 674140 856092
rect 675156 855076 675180 856092
rect 674116 855052 675180 855076
rect 650654 855024 651202 855025
rect 651602 854549 652170 854550
rect 651602 853413 651603 854549
rect 652169 853413 652170 854549
rect 671570 854498 672638 854522
rect 671570 853466 671594 854498
rect 672614 853466 672638 854498
rect 671570 853442 672638 853466
rect 651602 853412 652170 853413
rect 61424 827279 61962 827280
rect 44278 827206 46734 827230
rect 44278 826200 44302 827206
rect 46710 826200 46734 827206
rect 44278 826176 46734 826200
rect 61424 826161 61425 827279
rect 61961 826161 61962 827279
rect 61424 826160 61962 826161
rect 60460 825687 60998 825688
rect 41068 825624 43524 825648
rect 41068 825530 41092 825624
rect 43500 825530 43524 825624
rect 60460 824569 60461 825687
rect 60997 824569 60998 825687
rect 60460 824568 60998 824569
rect 63350 824131 63872 824132
rect 63350 823023 63351 824131
rect 63871 823023 63872 824131
rect 63350 823022 63872 823023
rect 62382 822523 62904 822524
rect 62382 821415 62383 822523
rect 62903 821415 62904 822523
rect 62382 821414 62904 821415
rect 30820 820831 31574 820832
rect 30820 819755 30821 820831
rect 31573 819755 31574 820831
rect 30820 819754 31574 819755
rect 37358 819263 38120 819264
rect 37358 818181 37359 819263
rect 38119 818181 38120 819263
rect 37358 818180 38120 818181
rect 61424 785679 61962 785680
rect 44278 785606 46734 785630
rect 44278 784600 44302 785606
rect 46710 784600 46734 785606
rect 44278 784576 46734 784600
rect 61424 784561 61425 785679
rect 61961 784561 61962 785679
rect 61424 784560 61962 784561
rect 60460 784087 60998 784088
rect 41068 784024 43524 784048
rect 41068 783018 41092 784024
rect 43500 783018 43524 784024
rect 41068 782994 43524 783018
rect 60460 782969 60461 784087
rect 60997 782969 60998 784087
rect 60460 782968 60998 782969
rect 63350 782131 63872 782132
rect 63350 781023 63351 782131
rect 63871 781023 63872 782131
rect 63350 781022 63872 781023
rect 62382 779323 62904 779324
rect 62382 778215 62383 779323
rect 62903 778215 62904 779323
rect 62382 778214 62904 778215
rect 30820 777631 31574 777632
rect 30820 776555 30821 777631
rect 31573 776555 31574 777631
rect 30820 776554 31574 776555
rect 37358 776063 38120 776064
rect 37358 774981 37359 776063
rect 38119 774981 38120 776063
rect 37358 774980 38120 774981
rect 650654 767945 651202 767946
rect 650654 766825 650655 767945
rect 651201 766825 651202 767945
rect 650654 766824 651202 766825
rect 651602 766349 652170 766350
rect 651602 765213 651603 766349
rect 652169 765213 652170 766349
rect 651602 765212 652170 765213
rect 686012 764631 686766 764632
rect 686012 763555 686013 764631
rect 686765 763555 686766 764631
rect 686012 763554 686766 763555
rect 679466 763063 680228 763064
rect 679466 761981 679467 763063
rect 680227 761981 680228 763063
rect 679466 761980 680228 761981
rect 61424 740879 61962 740880
rect 44278 740806 46734 740830
rect 44278 739800 44302 740806
rect 46710 739800 46734 740806
rect 44278 739776 46734 739800
rect 61424 739761 61425 740879
rect 61961 739761 61962 740879
rect 61424 739760 61962 739761
rect 60460 739287 60998 739288
rect 41068 739224 43524 739248
rect 41068 739130 41092 739224
rect 43500 739130 43524 739224
rect 60460 738169 60461 739287
rect 60997 738169 60998 739287
rect 60460 738168 60998 738169
rect 63350 737731 63872 737732
rect 63350 736623 63351 737731
rect 63871 736623 63872 737731
rect 63350 736622 63872 736623
rect 62382 736123 62904 736124
rect 62382 735015 62383 736123
rect 62903 735015 62904 736123
rect 62382 735014 62904 735015
rect 30820 734431 31574 734432
rect 30820 733355 30821 734431
rect 31573 733355 31574 734431
rect 30820 733354 31574 733355
rect 37358 732863 38120 732864
rect 37358 731781 37359 732863
rect 38119 731781 38120 732863
rect 37358 731780 38120 731781
rect 650654 722945 651202 722946
rect 650654 721825 650655 722945
rect 651201 721825 651202 722945
rect 650654 721824 651202 721825
rect 651602 721349 652170 721350
rect 651602 720213 651603 721349
rect 652169 720213 652170 721349
rect 651602 720212 652170 720213
rect 686012 719631 686766 719632
rect 686012 718555 686013 719631
rect 686765 718555 686766 719631
rect 686012 718554 686766 718555
rect 679466 718063 680228 718064
rect 679466 716981 679467 718063
rect 680227 716981 680228 718063
rect 679466 716980 680228 716981
rect 61424 697679 61962 697680
rect 44278 697606 46734 697630
rect 44278 696600 44302 697606
rect 46710 696600 46734 697606
rect 44278 696576 46734 696600
rect 61424 696561 61425 697679
rect 61961 696561 61962 697679
rect 61424 696560 61962 696561
rect 60460 696087 60998 696088
rect 41068 696024 43524 696048
rect 41068 695930 41092 696024
rect 43500 695930 43524 696024
rect 60460 694969 60461 696087
rect 60997 694969 60998 696087
rect 60460 694968 60998 694969
rect 63350 694531 63872 694532
rect 63350 693423 63351 694531
rect 63871 693423 63872 694531
rect 63350 693422 63872 693423
rect 62382 692923 62904 692924
rect 62382 691815 62383 692923
rect 62903 691815 62904 692923
rect 62382 691814 62904 691815
rect 30820 691231 31574 691232
rect 30820 690155 30821 691231
rect 31573 690155 31574 691231
rect 30820 690154 31574 690155
rect 37358 689663 38120 689664
rect 37358 688581 37359 689663
rect 38119 688581 38120 689663
rect 37358 688580 38120 688581
rect 650654 677745 651202 677746
rect 650654 676625 650655 677745
rect 651201 676625 651202 677745
rect 650654 676624 651202 676625
rect 651602 676149 652170 676150
rect 651602 675013 651603 676149
rect 652169 675013 652170 676149
rect 651602 675012 652170 675013
rect 686012 674431 686766 674432
rect 686012 673355 686013 674431
rect 686765 673355 686766 674431
rect 686012 673354 686766 673355
rect 679466 672863 680228 672864
rect 679466 671781 679467 672863
rect 680227 671781 680228 672863
rect 679466 671780 680228 671781
rect 61424 654479 61962 654480
rect 44278 654406 46734 654430
rect 44278 653400 44302 654406
rect 46710 653400 46734 654406
rect 44278 653376 46734 653400
rect 61424 653361 61425 654479
rect 61961 653361 61962 654479
rect 61424 653360 61962 653361
rect 60460 652887 60998 652888
rect 41068 652824 43524 652848
rect 41068 652730 41092 652824
rect 43500 652730 43524 652824
rect 60460 651769 60461 652887
rect 60997 651769 60998 652887
rect 60460 651768 60998 651769
rect 63350 651331 63872 651332
rect 63350 650223 63351 651331
rect 63871 650223 63872 651331
rect 63350 650222 63872 650223
rect 62382 649723 62904 649724
rect 62382 648615 62383 649723
rect 62903 648615 62904 649723
rect 62382 648614 62904 648615
rect 30820 648031 31574 648032
rect 30820 646955 30821 648031
rect 31573 646955 31574 648031
rect 30820 646954 31574 646955
rect 37358 646463 38120 646464
rect 37358 645381 37359 646463
rect 38119 645381 38120 646463
rect 37358 645380 38120 645381
rect 650654 632745 651202 632746
rect 650654 631625 650655 632745
rect 651201 631625 651202 632745
rect 650654 631624 651202 631625
rect 651602 629949 652170 629950
rect 651602 628813 651603 629949
rect 652169 628813 652170 629949
rect 651602 628812 652170 628813
rect 686012 629431 686766 629432
rect 686012 628355 686013 629431
rect 686765 628355 686766 629431
rect 686012 628354 686766 628355
rect 679466 627863 680228 627864
rect 679466 626781 679467 627863
rect 680227 626781 680228 627863
rect 679466 626780 680228 626781
rect 61424 612339 61962 612340
rect 44278 612266 46734 612290
rect 44278 611260 44302 612266
rect 46710 611260 46734 612266
rect 44278 611236 46734 611260
rect 61424 611221 61425 612339
rect 61961 611221 61962 612339
rect 61424 611220 61962 611221
rect 60460 610747 60998 610748
rect 41068 610684 43524 610708
rect 41068 609678 41092 610684
rect 43500 609678 43524 610684
rect 41068 609654 43524 609678
rect 60460 609629 60461 610747
rect 60997 609629 60998 610747
rect 60460 609628 60998 609629
rect 63350 608131 63872 608132
rect 63350 607023 63351 608131
rect 63871 607023 63872 608131
rect 63350 607022 63872 607023
rect 62382 606523 62904 606524
rect 62382 605415 62383 606523
rect 62903 605415 62904 606523
rect 62382 605414 62904 605415
rect 30820 604831 31574 604832
rect 30820 603755 30821 604831
rect 31573 603755 31574 604831
rect 30820 603754 31574 603755
rect 37358 603263 38120 603264
rect 37358 602181 37359 603263
rect 38119 602181 38120 603263
rect 37358 602180 38120 602181
rect 650654 587545 651202 587546
rect 650654 586425 650655 587545
rect 651201 586425 651202 587545
rect 650654 586424 651202 586425
rect 651602 585949 652170 585950
rect 651602 584813 651603 585949
rect 652169 584813 652170 585949
rect 651602 584812 652170 584813
rect 686012 584231 686766 584232
rect 686012 583155 686013 584231
rect 686765 583155 686766 584231
rect 686012 583154 686766 583155
rect 679466 582663 680228 582664
rect 679466 581581 679467 582663
rect 680227 581581 680228 582663
rect 679466 581580 680228 581581
rect 61424 568079 61962 568080
rect 44278 568006 46734 568030
rect 44278 567000 44302 568006
rect 46710 567000 46734 568006
rect 44278 566976 46734 567000
rect 61424 566961 61425 568079
rect 61961 566961 61962 568079
rect 61424 566960 61962 566961
rect 60460 566487 60998 566488
rect 41068 566424 43524 566448
rect 41068 566330 41092 566424
rect 43500 566330 43524 566424
rect 60460 565369 60461 566487
rect 60997 565369 60998 566487
rect 60460 565368 60998 565369
rect 63350 564931 63872 564932
rect 63350 563823 63351 564931
rect 63871 563823 63872 564931
rect 63350 563822 63872 563823
rect 62382 563323 62904 563324
rect 62382 562215 62383 563323
rect 62903 562215 62904 563323
rect 62382 562214 62904 562215
rect 30820 561631 31574 561632
rect 30820 560555 30821 561631
rect 31573 560555 31574 561631
rect 30820 560554 31574 560555
rect 37358 560063 38120 560064
rect 37358 558981 37359 560063
rect 38119 558981 38120 560063
rect 37358 558980 38120 558981
rect 650654 542545 651202 542546
rect 650654 541425 650655 542545
rect 651201 541425 651202 542545
rect 650654 541424 651202 541425
rect 651602 540949 652170 540950
rect 651602 539813 651603 540949
rect 652169 539813 652170 540949
rect 651602 539812 652170 539813
rect 686012 539231 686766 539232
rect 686012 538155 686013 539231
rect 686765 538155 686766 539231
rect 686012 538154 686766 538155
rect 679466 537663 680228 537664
rect 679466 536581 679467 537663
rect 680227 536581 680228 537663
rect 679466 536580 680228 536581
rect 650654 499145 651202 499146
rect 650654 498025 650655 499145
rect 651201 498025 651202 499145
rect 650654 498024 651202 498025
rect 651602 496949 652170 496950
rect 651602 495813 651603 496949
rect 652169 495813 652170 496949
rect 651602 495812 652170 495813
rect 686012 495231 686766 495232
rect 686012 494155 686013 495231
rect 686765 494155 686766 495231
rect 686012 494154 686766 494155
rect 679466 493663 680228 493664
rect 679466 492581 679467 493663
rect 680227 492581 680228 493663
rect 679466 492580 680228 492581
rect 61424 440479 61962 440480
rect 44278 440406 46734 440430
rect 44278 439400 44302 440406
rect 46710 439400 46734 440406
rect 44278 439376 46734 439400
rect 61424 439361 61425 440479
rect 61961 439361 61962 440479
rect 61424 439360 61962 439361
rect 60460 438887 60998 438888
rect 41068 438824 43524 438848
rect 41068 438730 41092 438824
rect 43500 438730 43524 438824
rect 60460 437769 60461 438887
rect 60997 437769 60998 438887
rect 60460 437768 60998 437769
rect 63350 437331 63872 437332
rect 63350 436223 63351 437331
rect 63871 436223 63872 437331
rect 63350 436222 63872 436223
rect 62382 435723 62904 435724
rect 62382 434615 62383 435723
rect 62903 434615 62904 435723
rect 62382 434614 62904 434615
rect 30820 434031 31574 434032
rect 30820 432955 30821 434031
rect 31573 432955 31574 434031
rect 30820 432954 31574 432955
rect 37358 432463 38120 432464
rect 37358 431381 37359 432463
rect 38119 431381 38120 432463
rect 37358 431380 38120 431381
rect 650654 410345 651202 410346
rect 650654 409225 650655 410345
rect 651201 409225 651202 410345
rect 650654 409224 651202 409225
rect 651602 408749 652170 408750
rect 651602 407613 651603 408749
rect 652169 407613 652170 408749
rect 651602 407612 652170 407613
rect 686012 407031 686766 407032
rect 686012 405955 686013 407031
rect 686765 405955 686766 407031
rect 686012 405954 686766 405955
rect 679466 405463 680228 405464
rect 679466 404381 679467 405463
rect 680227 404381 680228 405463
rect 679466 404380 680228 404381
rect 61424 397279 61962 397280
rect 44278 397206 46734 397230
rect 44278 396200 44302 397206
rect 46710 396200 46734 397206
rect 44278 396176 46734 396200
rect 61424 396161 61425 397279
rect 61961 396161 61962 397279
rect 61424 396160 61962 396161
rect 60460 395687 60998 395688
rect 41068 395624 43524 395648
rect 41068 395530 41092 395624
rect 43500 395530 43524 395624
rect 60460 394569 60461 395687
rect 60997 394569 60998 395687
rect 60460 394568 60998 394569
rect 63350 394131 63872 394132
rect 63350 393023 63351 394131
rect 63871 393023 63872 394131
rect 63350 393022 63872 393023
rect 62382 392523 62904 392524
rect 62382 391415 62383 392523
rect 62903 391415 62904 392523
rect 62382 391414 62904 391415
rect 30820 390831 31574 390832
rect 30820 389755 30821 390831
rect 31573 389755 31574 390831
rect 30820 389754 31574 389755
rect 37358 389263 38120 389264
rect 37358 388181 37359 389263
rect 38119 388181 38120 389263
rect 37358 388180 38120 388181
rect 650654 366545 651202 366546
rect 650654 365425 650655 366545
rect 651201 365425 651202 366545
rect 650654 365424 651202 365425
rect 651602 363549 652170 363550
rect 651602 362413 651603 363549
rect 652169 362413 652170 363549
rect 651602 362412 652170 362413
rect 686012 361831 686766 361832
rect 686012 360755 686013 361831
rect 686765 360755 686766 361831
rect 686012 360754 686766 360755
rect 679466 360263 680228 360264
rect 679466 359181 679467 360263
rect 680227 359181 680228 360263
rect 679466 359180 680228 359181
rect 61424 355079 61962 355080
rect 44278 355006 46734 355030
rect 44278 354000 44302 355006
rect 46710 354000 46734 355006
rect 44278 353976 46734 354000
rect 61424 353961 61425 355079
rect 61961 353961 61962 355079
rect 61424 353960 61962 353961
rect 60460 353487 60998 353488
rect 41068 353424 43524 353448
rect 41068 352418 41092 353424
rect 43500 352418 43524 353424
rect 41068 352394 43524 352418
rect 60460 352369 60461 353487
rect 60997 352369 60998 353487
rect 60460 352368 60998 352369
rect 63350 351731 63872 351732
rect 63350 350623 63351 351731
rect 63871 350623 63872 351731
rect 63350 350622 63872 350623
rect 62382 349323 62904 349324
rect 62382 348215 62383 349323
rect 62903 348215 62904 349323
rect 62382 348214 62904 348215
rect 30820 347631 31574 347632
rect 30820 346555 30821 347631
rect 31573 346555 31574 347631
rect 30820 346554 31574 346555
rect 37358 346063 38120 346064
rect 37358 344981 37359 346063
rect 38119 344981 38120 346063
rect 37358 344980 38120 344981
rect 650654 320145 651202 320146
rect 650654 319025 650655 320145
rect 651201 319025 651202 320145
rect 650654 319024 651202 319025
rect 651602 318549 652170 318550
rect 651602 317413 651603 318549
rect 652169 317413 652170 318549
rect 651602 317412 652170 317413
rect 686012 316831 686766 316832
rect 686012 315755 686013 316831
rect 686765 315755 686766 316831
rect 686012 315754 686766 315755
rect 679466 315263 680228 315264
rect 679466 314181 679467 315263
rect 680227 314181 680228 315263
rect 679466 314180 680228 314181
rect 61424 310879 61962 310880
rect 44278 310806 46734 310830
rect 44278 309800 44302 310806
rect 46710 309800 46734 310806
rect 44278 309776 46734 309800
rect 61424 309761 61425 310879
rect 61961 309761 61962 310879
rect 61424 309760 61962 309761
rect 60460 309287 60998 309288
rect 41068 309224 43524 309248
rect 41068 309130 41092 309224
rect 43500 309130 43524 309224
rect 60460 308169 60461 309287
rect 60997 308169 60998 309287
rect 60460 308168 60998 308169
rect 63350 307731 63872 307732
rect 63350 306623 63351 307731
rect 63871 306623 63872 307731
rect 63350 306622 63872 306623
rect 62382 306123 62904 306124
rect 62382 305015 62383 306123
rect 62903 305015 62904 306123
rect 62382 305014 62904 305015
rect 30820 304431 31574 304432
rect 30820 303355 30821 304431
rect 31573 303355 31574 304431
rect 30820 303354 31574 303355
rect 37358 302863 38120 302864
rect 37358 301781 37359 302863
rect 38119 301781 38120 302863
rect 37358 301780 38120 301781
rect 674084 278332 676564 278356
rect 670884 277386 673364 277410
rect 44228 277238 46762 277262
rect 44228 275912 44252 277238
rect 46738 275912 46762 277238
rect 670884 276530 670908 277386
rect 673340 276530 673364 277386
rect 674084 276844 674108 278332
rect 676540 276844 676564 278332
rect 674084 276820 676564 276844
rect 670884 276098 670908 276504
rect 673340 276098 673364 276504
rect 670884 276074 673364 276098
rect 44228 275888 46762 275912
rect 42830 275434 43528 275458
rect 42830 269402 42854 275434
rect 43504 269402 43528 275434
rect 675408 275122 676490 275146
rect 675408 274072 675432 275122
rect 676466 274072 676490 275122
rect 675408 274048 676490 274072
rect 671702 273504 672784 273528
rect 671702 272454 671726 273504
rect 672760 272454 672784 273504
rect 671702 272430 672784 272454
rect 686012 271831 686766 271832
rect 56616 271082 56632 271118
rect 686012 270755 686013 271831
rect 686765 270755 686766 271831
rect 686012 270754 686766 270755
rect 42830 269378 43528 269402
rect 679466 270263 680228 270264
rect 679466 269181 679467 270263
rect 680227 269181 680228 270263
rect 679466 269180 680228 269181
rect 30820 261231 31574 261232
rect 30820 260155 30821 261231
rect 31573 260155 31574 261231
rect 30820 260154 31574 260155
rect 37358 259663 38120 259664
rect 37358 258581 37359 259663
rect 38119 258581 38120 259663
rect 37358 258580 38120 258581
rect 674156 249272 676452 249296
rect 674156 246640 674180 249272
rect 676428 246640 676452 249272
rect 674156 246616 676452 246640
rect 41066 245364 43530 245388
rect 41066 238386 41090 245364
rect 43506 238386 43530 245364
rect 41066 238362 43530 238386
rect 44254 241334 46718 241358
rect 44254 234556 44278 241334
rect 46694 234556 46718 241334
rect 44254 234532 46718 234556
rect 675408 229922 676490 229946
rect 675408 228872 675432 229922
rect 676466 228872 676490 229922
rect 675408 228848 676490 228872
rect 671702 228304 672784 228328
rect 671702 227254 671726 228304
rect 672760 227254 672784 228304
rect 671702 227230 672784 227254
rect 686012 226631 686766 226632
rect 686012 225555 686013 226631
rect 686765 225555 686766 226631
rect 686012 225554 686766 225555
rect 679466 225063 680228 225064
rect 679466 223981 679467 225063
rect 680227 223981 680228 225063
rect 679466 223980 680228 223981
rect 30820 218031 31574 218032
rect 30820 216955 30821 218031
rect 31573 216955 31574 218031
rect 30820 216954 31574 216955
rect 37358 216463 38120 216464
rect 37358 215381 37359 216463
rect 38119 215381 38120 216463
rect 37358 215380 38120 215381
rect 675408 184922 676490 184946
rect 675408 183872 675432 184922
rect 676466 183872 676490 184922
rect 675408 183848 676490 183872
rect 671702 183304 672784 183328
rect 671702 182254 671726 183304
rect 672760 182254 672784 183304
rect 671702 182230 672784 182254
rect 686012 181631 686766 181632
rect 686012 180555 686013 181631
rect 686765 180555 686766 181631
rect 686012 180554 686766 180555
rect 679466 180063 680228 180064
rect 679466 178981 679467 180063
rect 680227 178981 680228 180063
rect 679466 178980 680228 178981
rect 675408 139722 676490 139746
rect 675408 138672 675432 139722
rect 676466 138672 676490 139722
rect 675408 138648 676490 138672
rect 671702 138104 672784 138128
rect 671702 137054 671726 138104
rect 672760 137054 672784 138104
rect 671702 137030 672784 137054
rect 686012 136431 686766 136432
rect 686012 135355 686013 136431
rect 686765 135355 686766 136431
rect 686012 135354 686766 135355
rect 679466 134863 680228 134864
rect 679466 133781 679467 134863
rect 680227 133781 680228 134863
rect 679466 133780 680228 133781
rect 234842 38177 237788 38178
rect 234842 37337 234843 38177
rect 237787 37337 237788 38177
rect 234842 37336 237788 37337
rect 149632 35995 150436 35996
rect 149632 35167 149633 35995
rect 150435 35167 150436 35995
rect 149632 35166 150436 35167
rect 148098 34787 148902 34788
rect 148098 33959 148099 34787
rect 148901 33959 148902 34787
rect 642026 34759 643634 34760
rect 642026 33989 642027 34759
rect 643633 33989 643634 34759
rect 642026 33988 643634 33989
rect 148098 33958 148902 33959
rect 204996 31645 207928 31646
rect 204996 30787 204997 31645
rect 207927 30787 207928 31645
rect 204996 30786 207928 30787
<< error_s >>
rect 41068 950418 41092 951330
rect 43500 950418 43524 951330
rect 41068 950394 43524 950418
rect 675398 946322 676480 946346
rect 675398 945272 675422 946322
rect 676456 945272 676480 946322
rect 675398 945248 676480 945272
rect 671692 944704 672774 944728
rect 671692 943654 671716 944704
rect 672750 943654 672774 944704
rect 671692 943630 672774 943654
rect 41068 824618 41092 825530
rect 43500 824618 43524 825530
rect 41068 824594 43524 824618
rect 675408 767922 676490 767946
rect 675408 766872 675432 767922
rect 676466 766872 676490 767922
rect 675408 766848 676490 766872
rect 671702 766304 672784 766328
rect 671702 765254 671726 766304
rect 672760 765254 672784 766304
rect 671702 765230 672784 765254
rect 41068 738218 41092 739130
rect 43500 738218 43524 739130
rect 41068 738194 43524 738218
rect 675408 722922 676490 722946
rect 675408 721872 675432 722922
rect 676466 721872 676490 722922
rect 675408 721848 676490 721872
rect 671702 721304 672784 721328
rect 671702 720254 671726 721304
rect 672760 720254 672784 721304
rect 671702 720230 672784 720254
rect 41068 695018 41092 695930
rect 43500 695018 43524 695930
rect 41068 694994 43524 695018
rect 675408 677722 676490 677746
rect 675408 676672 675432 677722
rect 676466 676672 676490 677722
rect 675408 676648 676490 676672
rect 671702 676104 672784 676128
rect 671702 675054 671726 676104
rect 672760 675054 672784 676104
rect 671702 675030 672784 675054
rect 41068 651818 41092 652730
rect 43500 651818 43524 652730
rect 41068 651794 43524 651818
rect 675408 632722 676490 632746
rect 675408 631672 675432 632722
rect 676466 631672 676490 632722
rect 675408 631648 676490 631672
rect 671702 631104 672784 631128
rect 671702 630054 671726 631104
rect 672760 630054 672784 631104
rect 671702 630030 672784 630054
rect 675408 587522 676490 587546
rect 675408 586472 675432 587522
rect 676466 586472 676490 587522
rect 675408 586448 676490 586472
rect 671702 585904 672784 585928
rect 671702 584854 671726 585904
rect 672760 584854 672784 585904
rect 671702 584830 672784 584854
rect 41068 565418 41092 566330
rect 43500 565418 43524 566330
rect 41068 565394 43524 565418
rect 675408 542522 676490 542546
rect 675408 541472 675432 542522
rect 676466 541472 676490 542522
rect 675408 541448 676490 541472
rect 671702 540904 672784 540928
rect 671702 539854 671726 540904
rect 672760 539854 672784 540904
rect 671702 539830 672784 539854
rect 675408 498522 676490 498546
rect 675408 497472 675432 498522
rect 676466 497472 676490 498522
rect 675408 497448 676490 497472
rect 671702 496904 672784 496928
rect 671702 495854 671726 496904
rect 672760 495854 672784 496904
rect 671702 495830 672784 495854
rect 41068 437818 41092 438730
rect 43500 437818 43524 438730
rect 41068 437794 43524 437818
rect 675408 410322 676490 410346
rect 675408 409272 675432 410322
rect 676466 409272 676490 410322
rect 675408 409248 676490 409272
rect 671702 408704 672784 408728
rect 671702 407654 671726 408704
rect 672760 407654 672784 408704
rect 671702 407630 672784 407654
rect 41068 394618 41092 395530
rect 43500 394618 43524 395530
rect 41068 394594 43524 394618
rect 675408 365122 676490 365146
rect 675408 364072 675432 365122
rect 676466 364072 676490 365122
rect 675408 364048 676490 364072
rect 671702 363504 672784 363528
rect 671702 362454 671726 363504
rect 672760 362454 672784 363504
rect 671702 362430 672784 362454
rect 675408 320122 676490 320146
rect 675408 319072 675432 320122
rect 676466 319072 676490 320122
rect 675408 319048 676490 319072
rect 671702 318504 672784 318528
rect 671702 317454 671726 318504
rect 672760 317454 672784 318504
rect 671702 317430 672784 317454
rect 41068 308218 41092 309130
rect 43500 308218 43524 309130
rect 41068 308194 43524 308218
<< metal1 >>
rect 648104 47124 649670 47188
rect 648104 46660 648166 47124
rect 649608 46738 649670 47124
rect 649608 46660 650160 46738
rect 648104 46598 650160 46660
rect 648104 46590 649670 46598
<< via1 >>
rect 648166 46660 649608 47124
<< metal2 >>
rect 648104 47124 649670 47188
rect 648104 46660 648166 47124
rect 649608 46660 649670 47124
rect 648104 46590 649670 46660
<< via2 >>
rect 648166 46660 649608 47124
<< metal3 >>
rect 575700 997056 580479 997678
rect 575700 995134 575788 997056
rect 580384 995134 580479 997056
rect 575700 995032 580479 995134
rect 585678 997062 590458 997678
rect 585678 995140 585758 997062
rect 590354 995140 590458 997062
rect 585678 995032 590458 995140
rect 44198 953080 61996 953124
rect 44198 953030 61424 953080
rect 44198 951976 44278 953030
rect 46734 951976 61424 953030
rect 44198 951960 61424 951976
rect 61962 951960 61996 953080
rect 44198 951924 61996 951960
rect 40984 951488 61032 951524
rect 40984 951448 60460 951488
rect 40984 950394 41068 951448
rect 43524 950394 60460 951448
rect 40984 950368 60460 950394
rect 60998 950368 61032 951488
rect 40984 950324 61032 950368
rect 55372 949682 58218 949982
rect 55372 949632 63922 949682
rect 55372 948782 63350 949632
rect 57038 948522 63350 948782
rect 63872 948522 63922 949632
rect 57038 948482 63922 948522
rect 53768 948182 56610 948382
rect 53768 948124 62944 948182
rect 53768 947182 62382 948124
rect 55432 947014 62382 947182
rect 62904 947014 62944 948124
rect 55432 946982 62944 947014
rect 650616 946346 675364 946382
rect 650616 945224 650654 946346
rect 651202 945224 675364 946346
rect 650616 945182 675364 945224
rect 651580 944750 671668 944782
rect 651580 943612 651602 944750
rect 652170 943612 671668 944750
rect 651580 943582 671668 943612
rect 650616 901146 675830 901182
rect 650616 900024 650654 901146
rect 651202 901112 675830 901146
rect 651202 900074 674734 901112
rect 675740 900074 675830 901112
rect 651202 900024 675830 900074
rect 650616 899982 675830 900024
rect 651580 899550 672676 899582
rect 651580 898412 651602 899550
rect 652170 899504 672676 899550
rect 652170 898466 671566 899504
rect 672596 898466 672676 899504
rect 652170 898412 672676 898466
rect 651580 898382 672676 898412
rect 650616 856146 675264 856182
rect 650616 855024 650654 856146
rect 651202 856116 675264 856146
rect 651202 855052 674116 856116
rect 675180 855052 675264 856116
rect 651202 855024 675264 855052
rect 650616 854982 675264 855024
rect 651580 854550 672708 854582
rect 651580 853412 651602 854550
rect 652170 854522 672708 854550
rect 652170 853442 671570 854522
rect 672638 853442 672708 854522
rect 652170 853412 672708 853442
rect 651580 853382 672708 853412
rect 39852 842324 50002 842458
rect 39852 837800 47908 842324
rect 49694 837800 50002 842324
rect 39852 837678 50002 837800
rect 667172 833206 677818 833301
rect 39852 832392 50002 832479
rect 39852 827868 47908 832392
rect 49694 827868 50002 832392
rect 667172 828630 667284 833206
rect 669732 828630 677818 833206
rect 667172 828521 677818 828630
rect 39852 827699 50002 827868
rect 44198 827280 61996 827324
rect 44198 827230 61424 827280
rect 44198 826176 44278 827230
rect 46734 826176 61424 827230
rect 44198 826160 61424 826176
rect 61962 826160 61996 827280
rect 44198 826124 61996 826160
rect 40984 825688 61032 825724
rect 40984 825648 60460 825688
rect 40984 824594 41068 825648
rect 43524 824594 60460 825648
rect 40984 824568 60460 824594
rect 60998 824568 61032 825688
rect 40984 824524 61032 824568
rect 55372 824132 63922 824182
rect 55372 823022 63350 824132
rect 63872 823022 63922 824132
rect 55372 822982 63922 823022
rect 667172 823212 677818 823322
rect 53768 822524 62944 822582
rect 53768 821414 62382 822524
rect 62904 821414 62944 822524
rect 53768 821382 62944 821414
rect 667172 818636 667270 823212
rect 669718 818636 677818 823212
rect 667172 818542 677818 818636
rect 44198 785680 61996 785724
rect 44198 785630 61424 785680
rect 44198 784576 44278 785630
rect 46734 784576 61424 785630
rect 44198 784560 61424 784576
rect 61962 784560 61996 785680
rect 44198 784524 61996 784560
rect 40984 784088 61032 784124
rect 40984 784048 60460 784088
rect 40984 782994 41068 784048
rect 43524 782994 60460 784048
rect 40984 782968 60460 782994
rect 60998 782968 61032 784088
rect 40984 782924 61032 782968
rect 56078 782132 63922 782182
rect 56078 781022 63350 782132
rect 63872 781022 63922 782132
rect 56078 780982 63922 781022
rect 55372 779782 57370 780982
rect 53768 779324 62944 779382
rect 53768 778214 62382 779324
rect 62904 778214 62944 779324
rect 53768 778182 62944 778214
rect 650616 767946 675364 767982
rect 650616 766824 650654 767946
rect 651202 766824 675364 767946
rect 650616 766782 675364 766824
rect 651580 766350 671668 766382
rect 651580 765212 651602 766350
rect 652170 765212 671668 766350
rect 651580 765182 671668 765212
rect 44198 740880 61996 740924
rect 44198 740830 61424 740880
rect 44198 739776 44278 740830
rect 46734 739776 61424 740830
rect 44198 739760 61424 739776
rect 61962 739760 61996 740880
rect 44198 739724 61996 739760
rect 40984 739288 61032 739324
rect 40984 739248 60460 739288
rect 40984 738194 41068 739248
rect 43524 738194 60460 739248
rect 40984 738168 60460 738194
rect 60998 738168 61032 739288
rect 40984 738124 61032 738168
rect 55372 737732 63922 737782
rect 55372 736622 63350 737732
rect 63872 736622 63922 737732
rect 55372 736582 63922 736622
rect 53768 736124 62944 736182
rect 53768 735014 62382 736124
rect 62904 735014 62944 736124
rect 53768 734982 62944 735014
rect 650616 722946 675364 722982
rect 650616 721824 650654 722946
rect 651202 721824 675364 722946
rect 650616 721782 675364 721824
rect 651580 721350 671668 721382
rect 651580 720212 651602 721350
rect 652170 720212 671668 721350
rect 651580 720182 671668 720212
rect 44198 697680 61996 697724
rect 44198 697630 61424 697680
rect 44198 696576 44278 697630
rect 46734 696576 61424 697630
rect 44198 696560 61424 696576
rect 61962 696560 61996 697680
rect 44198 696524 61996 696560
rect 40984 696088 61032 696124
rect 40984 696048 60460 696088
rect 40984 694994 41068 696048
rect 43524 694994 60460 696048
rect 40984 694968 60460 694994
rect 60998 694968 61032 696088
rect 40984 694924 61032 694968
rect 55372 694532 63922 694582
rect 55372 693422 63350 694532
rect 63872 693422 63922 694532
rect 55372 693382 63922 693422
rect 53768 692924 62944 692982
rect 53768 691814 62382 692924
rect 62904 691814 62944 692924
rect 53768 691782 62944 691814
rect 650616 677746 675364 677782
rect 650616 676624 650654 677746
rect 651202 676624 675364 677746
rect 650616 676582 675364 676624
rect 651580 676150 671668 676182
rect 651580 675012 651602 676150
rect 652170 675012 671668 676150
rect 651580 674982 671668 675012
rect 44198 654480 61996 654524
rect 44198 654430 61424 654480
rect 44198 653376 44278 654430
rect 46734 653376 61424 654430
rect 44198 653360 61424 653376
rect 61962 653360 61996 654480
rect 44198 653324 61996 653360
rect 40984 652888 61032 652924
rect 40984 652848 60460 652888
rect 40984 651794 41068 652848
rect 43524 651794 60460 652848
rect 40984 651768 60460 651794
rect 60998 651768 61032 652888
rect 40984 651724 61032 651768
rect 55372 651332 63922 651382
rect 55372 650222 63350 651332
rect 63872 650222 63922 651332
rect 55372 650182 63922 650222
rect 53768 649724 62944 649782
rect 53768 648614 62382 649724
rect 62904 648614 62944 649724
rect 53768 648582 62944 648614
rect 650616 632746 675364 632782
rect 650616 631624 650654 632746
rect 651202 631624 675364 632746
rect 650616 631582 675364 631624
rect 659310 629982 671668 631182
rect 651580 629950 660600 629982
rect 651580 628812 651602 629950
rect 652170 628812 660600 629950
rect 651580 628782 660600 628812
rect 44198 612340 61996 612384
rect 44198 612290 61424 612340
rect 44198 611236 44278 612290
rect 46734 611236 61424 612290
rect 44198 611220 61424 611236
rect 61962 611220 61996 612340
rect 44198 611184 61996 611220
rect 40984 610748 61032 610784
rect 40984 610708 60460 610748
rect 40984 609654 41068 610708
rect 43524 609654 60460 610708
rect 40984 609628 60460 609654
rect 60998 609628 61032 610748
rect 40984 609584 61032 609628
rect 55372 608132 63922 608182
rect 55372 607022 63350 608132
rect 63872 607022 63922 608132
rect 55372 606982 63922 607022
rect 53768 606524 62944 606582
rect 53768 605414 62382 606524
rect 62904 605414 62944 606524
rect 53768 605382 62944 605414
rect 650616 587546 675364 587582
rect 650616 586424 650654 587546
rect 651202 586424 675364 587546
rect 650616 586382 675364 586424
rect 651580 585950 671668 585982
rect 651580 584812 651602 585950
rect 652170 584812 671668 585950
rect 651580 584782 671668 584812
rect 44198 568080 61996 568124
rect 44198 568030 61424 568080
rect 44198 566976 44278 568030
rect 46734 566976 61424 568030
rect 44198 566960 61424 566976
rect 61962 566960 61996 568080
rect 44198 566924 61996 566960
rect 40984 566488 61032 566524
rect 40984 566448 60460 566488
rect 40984 565394 41068 566448
rect 43524 565394 60460 566448
rect 40984 565368 60460 565394
rect 60998 565368 61032 566488
rect 40984 565324 61032 565368
rect 55372 564932 63922 564982
rect 55372 563822 63350 564932
rect 63872 563822 63922 564932
rect 55372 563782 63922 563822
rect 53768 563324 62944 563382
rect 53768 562214 62382 563324
rect 62904 562214 62944 563324
rect 53768 562182 62944 562214
rect 650616 542546 675364 542582
rect 650616 541424 650654 542546
rect 651202 541424 675364 542546
rect 650616 541382 675364 541424
rect 651580 540950 671668 540982
rect 651580 539812 651602 540950
rect 652170 539812 671668 540950
rect 651580 539782 671668 539812
rect 667062 518582 677700 518701
rect 667062 514056 667336 518582
rect 669706 514056 677700 518582
rect 667062 513921 677700 514056
rect 667062 508592 677700 508722
rect 667062 504066 667350 508592
rect 669720 504066 677700 508592
rect 667062 503942 677700 504066
rect 650616 499146 659758 499182
rect 650616 498024 650654 499146
rect 651202 498582 659758 499146
rect 651202 498024 675364 498582
rect 650616 497982 675364 498024
rect 39924 497732 52292 497858
rect 39924 493250 50364 497732
rect 52092 493250 52292 497732
rect 658568 497382 675364 497982
rect 651580 496950 671668 496982
rect 651580 495812 651602 496950
rect 652170 495812 671668 496950
rect 651580 495782 671668 495812
rect 39924 493078 52292 493250
rect 39924 487742 52292 487879
rect 39924 483260 50352 487742
rect 52080 483260 52292 487742
rect 39924 483099 52292 483260
rect 44198 440480 61996 440524
rect 44198 440430 61424 440480
rect 44198 439376 44278 440430
rect 46734 439376 61424 440430
rect 44198 439360 61424 439376
rect 61962 439360 61996 440480
rect 44198 439324 61996 439360
rect 40984 438888 61032 438924
rect 40984 438848 60460 438888
rect 40984 437794 41068 438848
rect 43524 437794 60460 438848
rect 40984 437768 60460 437794
rect 60998 437768 61032 438888
rect 40984 437724 61032 437768
rect 55372 437332 63922 437382
rect 55372 436222 63350 437332
rect 63872 436222 63922 437332
rect 55372 436182 63922 436222
rect 53768 435724 62944 435782
rect 53768 434614 62382 435724
rect 62904 434614 62944 435724
rect 53768 434582 62944 434614
rect 663914 430390 677712 430501
rect 663914 425684 664134 430390
rect 666540 425748 677712 430390
rect 666540 425684 667110 425748
rect 663914 425562 667110 425684
rect 663914 420462 677712 420522
rect 663914 415856 664112 420462
rect 666528 415856 677712 420462
rect 663914 415742 677712 415856
rect 650616 410346 675364 410382
rect 650616 409224 650654 410346
rect 651202 409224 675364 410346
rect 650616 409182 675364 409224
rect 651580 408750 671668 408782
rect 651580 407612 651602 408750
rect 652170 407612 671668 408750
rect 651580 407582 671668 407612
rect 44198 397280 61996 397324
rect 44198 397230 61424 397280
rect 44198 396176 44278 397230
rect 46734 396176 61424 397230
rect 44198 396160 61424 396176
rect 61962 396160 61996 397280
rect 44198 396124 61996 396160
rect 40984 395688 61032 395724
rect 40984 395648 60460 395688
rect 40984 394594 41068 395648
rect 43524 394594 60460 395648
rect 40984 394568 60460 394594
rect 60998 394568 61032 395688
rect 40984 394524 61032 394568
rect 55372 394132 63922 394182
rect 55372 393022 63350 394132
rect 63872 393022 63922 394132
rect 55372 392982 63922 393022
rect 53768 392524 62944 392582
rect 53768 391414 62382 392524
rect 62904 391414 62944 392524
rect 53768 391382 62944 391414
rect 650616 366546 665664 366582
rect 650616 365424 650654 366546
rect 651202 365424 665664 366546
rect 650616 365382 665664 365424
rect 664464 365182 665664 365382
rect 664464 363982 675364 365182
rect 651580 363550 671668 363582
rect 651580 362412 651602 363550
rect 652170 362412 671668 363550
rect 651580 362382 671668 362412
rect 44198 355080 61996 355124
rect 44198 355030 61424 355080
rect 44198 353976 44278 355030
rect 46734 353976 61424 355030
rect 44198 353960 61424 353976
rect 61962 353960 61996 355080
rect 44198 353924 61996 353960
rect 40984 353488 61032 353524
rect 40984 353448 60460 353488
rect 40984 352394 41068 353448
rect 43524 352394 60460 353448
rect 40984 352368 60460 352394
rect 60998 352368 61032 353488
rect 40984 352324 61032 352368
rect 55968 351732 63922 351782
rect 55968 350982 63350 351732
rect 55372 350622 63350 350982
rect 63872 350622 63922 351732
rect 55372 350582 63922 350622
rect 55372 349782 57264 350582
rect 53768 349324 62944 349382
rect 53768 348214 62382 349324
rect 62904 348214 62944 349324
rect 53768 348182 62944 348214
rect 650616 320146 676922 320182
rect 650616 319024 650654 320146
rect 651202 319024 676922 320146
rect 650616 318982 676922 319024
rect 651580 318550 673726 318582
rect 651580 317412 651602 318550
rect 652170 317412 673726 318550
rect 651580 317382 673726 317412
rect 44198 310880 61996 310924
rect 44198 310830 61424 310880
rect 44198 309776 44278 310830
rect 46734 309776 61424 310830
rect 44198 309760 61424 309776
rect 61962 309760 61996 310880
rect 44198 309724 61996 309760
rect 40984 309288 61032 309324
rect 40984 309248 60460 309288
rect 40984 308194 41068 309248
rect 43524 308194 60460 309248
rect 40984 308168 60460 308194
rect 60998 308168 61032 309288
rect 40984 308124 61032 308168
rect 55432 307732 63922 307782
rect 55432 306622 63350 307732
rect 63872 306622 63922 307732
rect 55432 306582 63922 306622
rect 53790 306124 62944 306182
rect 53790 305014 62382 306124
rect 62904 305014 62944 306124
rect 53790 304982 62944 305014
rect 39456 82706 45844 82744
rect 39456 78242 41946 82706
rect 45672 78242 45844 82706
rect 39456 78151 45844 78242
rect 39456 72802 45844 72900
rect 39456 68338 41922 72802
rect 45648 68338 45844 72802
rect 39456 68256 45844 68338
rect 648104 47124 649670 47188
rect 241690 46616 246049 46686
rect 241690 42842 241740 46616
rect 245986 42842 246049 46616
rect 149600 41148 150458 41207
rect 149600 40988 149618 41148
rect 150440 40988 150458 41148
rect 148068 40752 148926 40782
rect 148068 40592 148086 40752
rect 148908 40592 148926 40752
rect 148068 34788 148926 40592
rect 149600 35996 150458 40988
rect 241690 39426 246049 42842
rect 251300 46630 255702 46686
rect 251300 42856 251392 46630
rect 255638 42856 255702 46630
rect 648104 46660 648166 47124
rect 649608 46660 649670 47124
rect 648104 46590 649670 46660
rect 653462 45026 656910 45156
rect 251300 39426 255702 42856
rect 641954 43988 643694 44026
rect 641954 42198 641994 43988
rect 643660 42198 643694 43988
rect 149600 35166 149632 35996
rect 150436 35166 150458 35996
rect 149600 35114 150458 35166
rect 234814 38178 237814 38242
rect 234814 37336 234842 38178
rect 237788 37336 237814 38178
rect 148068 33958 148098 34788
rect 148902 33958 148926 34788
rect 148068 33900 148926 33958
rect 204958 31646 207958 31734
rect 204958 30786 204996 31646
rect 207928 30786 207958 31646
rect 204958 18004 207958 30786
rect 234814 19380 237814 37336
rect 641954 34760 643694 42198
rect 653462 42634 653578 45026
rect 656772 42634 656910 45026
rect 653462 35808 656910 42634
rect 641954 33988 642026 34760
rect 643634 33988 643694 34760
rect 641954 33920 643694 33988
rect 234814 18544 234884 19380
rect 237754 18544 237814 19380
rect 234814 18466 237814 18544
rect 204958 17128 205020 18004
rect 207872 17128 207958 18004
rect 204958 17038 207958 17128
<< via3 >>
rect 575788 995134 580384 997056
rect 585758 995140 590354 997062
rect 44278 951976 46734 953030
rect 61424 951960 61962 953080
rect 41068 950394 43524 951448
rect 60460 950368 60998 951488
rect 63350 948522 63872 949632
rect 62382 947014 62904 948124
rect 650654 945224 651202 946346
rect 651602 943612 652170 944750
rect 650654 900024 651202 901146
rect 674734 900074 675740 901112
rect 651602 898412 652170 899550
rect 671566 898466 672596 899504
rect 650654 855024 651202 856146
rect 674116 855052 675180 856116
rect 651602 853412 652170 854550
rect 671570 853442 672638 854522
rect 47908 837800 49694 842324
rect 47908 827868 49694 832392
rect 667284 828630 669732 833206
rect 44278 826176 46734 827230
rect 61424 826160 61962 827280
rect 41068 824594 43524 825648
rect 60460 824568 60998 825688
rect 63350 823022 63872 824132
rect 62382 821414 62904 822524
rect 667270 818636 669718 823212
rect 44278 784576 46734 785630
rect 61424 784560 61962 785680
rect 41068 782994 43524 784048
rect 60460 782968 60998 784088
rect 63350 781022 63872 782132
rect 62382 778214 62904 779324
rect 650654 766824 651202 767946
rect 651602 765212 652170 766350
rect 44278 739776 46734 740830
rect 61424 739760 61962 740880
rect 41068 738194 43524 739248
rect 60460 738168 60998 739288
rect 63350 736622 63872 737732
rect 62382 735014 62904 736124
rect 650654 721824 651202 722946
rect 651602 720212 652170 721350
rect 44278 696576 46734 697630
rect 61424 696560 61962 697680
rect 41068 694994 43524 696048
rect 60460 694968 60998 696088
rect 63350 693422 63872 694532
rect 62382 691814 62904 692924
rect 650654 676624 651202 677746
rect 651602 675012 652170 676150
rect 44278 653376 46734 654430
rect 61424 653360 61962 654480
rect 41068 651794 43524 652848
rect 60460 651768 60998 652888
rect 63350 650222 63872 651332
rect 62382 648614 62904 649724
rect 650654 631624 651202 632746
rect 651602 628812 652170 629950
rect 44278 611236 46734 612290
rect 61424 611220 61962 612340
rect 41068 609654 43524 610708
rect 60460 609628 60998 610748
rect 63350 607022 63872 608132
rect 62382 605414 62904 606524
rect 650654 586424 651202 587546
rect 651602 584812 652170 585950
rect 44278 566976 46734 568030
rect 61424 566960 61962 568080
rect 41068 565394 43524 566448
rect 60460 565368 60998 566488
rect 63350 563822 63872 564932
rect 62382 562214 62904 563324
rect 650654 541424 651202 542546
rect 651602 539812 652170 540950
rect 667336 514056 669706 518582
rect 667350 504066 669720 508592
rect 650654 498024 651202 499146
rect 50364 493250 52092 497732
rect 651602 495812 652170 496950
rect 50352 483260 52080 487742
rect 44278 439376 46734 440430
rect 61424 439360 61962 440480
rect 41068 437794 43524 438848
rect 60460 437768 60998 438888
rect 63350 436222 63872 437332
rect 62382 434614 62904 435724
rect 664134 425684 666540 430390
rect 664112 415856 666528 420462
rect 650654 409224 651202 410346
rect 651602 407612 652170 408750
rect 44278 396176 46734 397230
rect 61424 396160 61962 397280
rect 41068 394594 43524 395648
rect 60460 394568 60998 395688
rect 63350 393022 63872 394132
rect 62382 391414 62904 392524
rect 650654 365424 651202 366546
rect 651602 362412 652170 363550
rect 44278 353976 46734 355030
rect 61424 353960 61962 355080
rect 41068 352394 43524 353448
rect 60460 352368 60998 353488
rect 63350 350622 63872 351732
rect 62382 348214 62904 349324
rect 650654 319024 651202 320146
rect 651602 317412 652170 318550
rect 44278 309776 46734 310830
rect 61424 309760 61962 310880
rect 41068 308194 43524 309248
rect 60460 308168 60998 309288
rect 63350 306622 63872 307732
rect 62382 305014 62904 306124
rect 41946 78242 45672 82706
rect 41922 68338 45648 72802
rect 241740 42842 245986 46616
rect 149618 40988 150440 41148
rect 148086 40592 148908 40752
rect 251392 42856 255638 46630
rect 648166 46660 649608 47124
rect 641994 42198 643660 43988
rect 149632 35166 150436 35996
rect 234842 37336 237788 38178
rect 148098 33958 148902 34788
rect 204996 30786 207928 31646
rect 653578 42634 656772 45026
rect 642026 33988 643634 34760
rect 234884 18544 237754 19380
rect 205020 17128 207872 18004
<< metal4 >>
rect 575680 997056 580478 997130
rect 575680 995134 575788 997056
rect 580384 995134 580478 997056
rect 575680 993314 580478 995134
rect 575680 990884 575762 993314
rect 580384 990884 580478 993314
rect 575680 990788 580478 990884
rect 585670 997062 590468 997144
rect 585670 995140 585758 997062
rect 590354 995140 590468 997062
rect 670816 996692 673426 996696
rect 670808 996584 676654 996692
rect 670808 995628 670928 996584
rect 676500 995628 676654 996584
rect 670808 995492 676654 995628
rect 585670 993328 590468 995140
rect 585670 990898 585758 993328
rect 590380 990898 590468 993328
rect 585670 990802 590468 990898
rect 670816 992530 673426 995492
rect 670816 990354 670976 992530
rect 673264 990354 673426 992530
rect 47796 990278 56582 990310
rect 47796 990276 55820 990278
rect 47796 989738 47836 990276
rect 49748 989738 55820 990276
rect 56394 989738 56582 990278
rect 670816 990200 673426 990354
rect 47796 989692 56582 989738
rect 50194 989318 56434 989348
rect 50194 989312 55824 989318
rect 50194 988774 50242 989312
rect 52154 988778 55824 989312
rect 56398 988778 56434 989318
rect 52154 988774 56434 988778
rect 50194 988736 56434 988774
rect 658380 987386 669826 987436
rect 658380 987376 667268 987386
rect 658380 986872 658430 987376
rect 663120 986872 667268 987376
rect 669770 986872 669826 987386
rect 658380 986812 669826 986872
rect 40993 986448 56414 986468
rect 40993 985878 41034 986448
rect 43574 986436 56414 986448
rect 43574 985886 55804 986436
rect 56378 985886 56414 986436
rect 43574 985878 56414 985886
rect 40993 985854 56414 985878
rect 44200 985498 56440 985526
rect 44200 984918 44242 985498
rect 46772 985478 56440 985498
rect 46772 984918 55804 985478
rect 44200 984916 55804 984918
rect 56408 984916 56440 985478
rect 44200 984874 56440 984916
rect 52596 984520 56404 984548
rect 52596 984510 55802 984520
rect 52596 983968 52628 984510
rect 53766 983968 55802 984510
rect 52596 983958 55802 983968
rect 56376 983958 56404 984520
rect 52596 983928 56404 983958
rect 658316 984536 673430 984570
rect 658316 984492 670858 984536
rect 658316 983984 658380 984492
rect 663118 983984 670858 984492
rect 658316 983950 670858 983984
rect 673384 983950 673430 984536
rect 658316 983928 673430 983950
rect 658288 983574 676624 983602
rect 658288 983536 674056 983574
rect 658288 983028 658362 983536
rect 663100 983028 674056 983536
rect 658288 982988 674056 983028
rect 676582 982988 676624 983574
rect 658288 982960 676624 982988
rect 44200 953030 46792 953126
rect 44200 951976 44278 953030
rect 46734 951976 46792 953030
rect 44200 951922 46792 951976
rect 40994 951448 43588 951522
rect 40994 950394 41068 951448
rect 43524 950394 43588 951448
rect 40994 950326 43588 950394
rect 674630 901112 675830 901182
rect 674630 900074 674734 901112
rect 675740 900074 675830 901112
rect 674630 899982 675830 900074
rect 671476 899504 672676 899582
rect 671476 898466 671566 899504
rect 672596 898466 672676 899504
rect 671476 898382 672676 898466
rect 674054 856116 675254 856182
rect 674054 855052 674116 856116
rect 675180 855052 675254 856116
rect 674054 854982 675254 855052
rect 671508 854522 672708 854582
rect 671508 853442 671570 854522
rect 672638 853442 672708 854522
rect 671508 853382 672708 853442
rect 47792 842324 49822 842462
rect 47792 837800 47908 842324
rect 49694 837800 49822 842324
rect 47792 837658 49822 837800
rect 667202 833206 669802 833310
rect 47792 832392 49822 832506
rect 47792 827868 47908 832392
rect 49694 827868 49822 832392
rect 667202 828630 667284 833206
rect 669732 828630 669802 833206
rect 667202 828520 669802 828630
rect 47792 827702 49822 827868
rect 44200 827230 46792 827326
rect 44200 826176 44278 827230
rect 46734 826176 46792 827230
rect 44200 826122 46792 826176
rect 40994 825648 43588 825722
rect 40994 824594 41068 825648
rect 43524 824594 43588 825648
rect 40994 824526 43588 824594
rect 667214 823212 669814 823336
rect 667214 818636 667270 823212
rect 669718 818636 669814 823212
rect 667214 818546 669814 818636
rect 44200 785630 46792 785726
rect 44200 784576 44278 785630
rect 46734 784576 46792 785630
rect 44200 784522 46792 784576
rect 40994 784048 43588 784122
rect 40994 782994 41068 784048
rect 43524 782994 43588 784048
rect 40994 782926 43588 782994
rect 44200 740830 46792 740926
rect 44200 739776 44278 740830
rect 46734 739776 46792 740830
rect 44200 739722 46792 739776
rect 40994 739248 43588 739322
rect 40994 738194 41068 739248
rect 43524 738194 43588 739248
rect 40994 738126 43588 738194
rect 44200 697630 46792 697726
rect 44200 696576 44278 697630
rect 46734 696576 46792 697630
rect 44200 696522 46792 696576
rect 40994 696048 43588 696122
rect 40994 694994 41068 696048
rect 43524 694994 43588 696048
rect 40994 694926 43588 694994
rect 44200 654430 46792 654526
rect 44200 653376 44278 654430
rect 46734 653376 46792 654430
rect 44200 653322 46792 653376
rect 40994 652848 43588 652922
rect 40994 651794 41068 652848
rect 43524 651794 43588 652848
rect 40994 651726 43588 651794
rect 44200 612290 46792 612386
rect 44200 611236 44278 612290
rect 46734 611236 46792 612290
rect 44200 611182 46792 611236
rect 40994 610708 43588 610782
rect 40994 609654 41068 610708
rect 43524 609654 43588 610708
rect 40994 609586 43588 609654
rect 44200 568030 46792 568126
rect 44200 566976 44278 568030
rect 46734 566976 46792 568030
rect 44200 566922 46792 566976
rect 40994 566448 43588 566522
rect 40994 565394 41068 566448
rect 43524 565394 43588 566448
rect 40994 565326 43588 565394
rect 667206 518582 669814 518696
rect 667206 514056 667336 518582
rect 669706 514056 669814 518582
rect 667206 513920 669814 514056
rect 667218 508592 669826 508726
rect 667218 504066 667350 508592
rect 669720 504066 669826 508592
rect 667218 503950 669826 504066
rect 50172 497732 52196 497874
rect 50172 493250 50364 497732
rect 52092 493250 52196 497732
rect 50172 493084 52196 493250
rect 50198 487742 52222 487884
rect 50198 483260 50352 487742
rect 52080 483260 52222 487742
rect 50198 483094 52222 483260
rect 44200 440430 46792 440526
rect 44200 439376 44278 440430
rect 46734 439376 46792 440430
rect 44200 439322 46792 439376
rect 40994 438848 43588 438922
rect 40994 437794 41068 438848
rect 43524 437794 43588 438848
rect 40994 437726 43588 437794
rect 664008 430390 666612 430490
rect 664008 425684 664134 430390
rect 666540 425684 666612 430390
rect 664008 425572 666612 425684
rect 664018 420462 666634 420524
rect 664018 415856 664112 420462
rect 666528 415856 666634 420462
rect 664018 415760 666634 415856
rect 44200 397230 46792 397326
rect 44200 396176 44278 397230
rect 46734 396176 46792 397230
rect 44200 396122 46792 396176
rect 40994 395648 43588 395722
rect 40994 394594 41068 395648
rect 43524 394594 43588 395648
rect 40994 394526 43588 394594
rect 44200 355030 46792 355126
rect 44200 353976 44278 355030
rect 46734 353976 46792 355030
rect 44200 353922 46792 353976
rect 40994 353448 43588 353522
rect 40994 352394 41068 353448
rect 43524 352394 43588 353448
rect 40994 352326 43588 352394
rect 44200 310830 46792 310926
rect 44200 309776 44278 310830
rect 46734 309776 46792 310830
rect 44200 309722 46792 309776
rect 40994 309248 43588 309322
rect 40994 308194 41068 309248
rect 43524 308194 43588 309248
rect 40994 308126 43588 308194
rect 658882 278356 676628 278406
rect 658882 278344 674084 278356
rect 52582 278014 53800 278046
rect 44195 277262 46802 277284
rect 44195 275888 44228 277262
rect 46762 276484 46802 277262
rect 52582 276882 52652 278014
rect 53730 277446 53800 278014
rect 658882 277842 658950 278344
rect 663094 277842 674084 278344
rect 53730 277420 56416 277446
rect 53730 276882 55790 277420
rect 52582 276854 55790 276882
rect 56378 276854 56416 277420
rect 52582 276822 56416 276854
rect 46762 276442 56432 276484
rect 46762 275898 55782 276442
rect 56406 275898 56432 276442
rect 46762 275888 56432 275898
rect 44195 275858 56432 275888
rect 42746 275488 56448 275532
rect 42746 275458 55790 275488
rect 42746 269378 42830 275458
rect 43528 274944 55790 275458
rect 56414 274944 56448 275488
rect 43528 274906 56448 274944
rect 43528 269378 43610 274906
rect 50186 273390 52198 273438
rect 50186 272078 50248 273390
rect 52134 272638 52198 273390
rect 52134 272618 56406 272638
rect 52134 272078 55782 272618
rect 50186 272052 55782 272078
rect 56378 272052 56406 272618
rect 50186 272026 56406 272052
rect 47792 271656 56616 271688
rect 47792 271652 55782 271656
rect 47792 270310 47848 271652
rect 49746 271088 55782 271652
rect 56486 271088 56616 271656
rect 49746 271082 56616 271088
rect 49746 271058 57202 271082
rect 49746 270310 49802 271058
rect 47792 270258 49802 270310
rect 42746 269278 43610 269378
rect 56572 261466 57202 271058
rect 57542 264698 58162 272042
rect 58502 269428 59122 272992
rect 58502 266504 58532 269428
rect 59082 266504 59122 269428
rect 58502 266408 59122 266504
rect 59462 266618 60082 273952
rect 60422 267578 61042 274922
rect 61382 268538 62002 275876
rect 62342 269498 62962 276834
rect 63302 270458 63922 277792
rect 63302 269838 67172 270458
rect 62342 268878 66212 269498
rect 61382 267918 65252 268538
rect 60422 266958 64292 267578
rect 59462 265998 63332 266618
rect 62712 265424 63332 265998
rect 57542 264078 61412 264698
rect 47770 261338 59470 261466
rect 47770 258676 48050 261338
rect 49608 261232 59470 261338
rect 49608 258676 56554 261232
rect 47770 258660 56554 258676
rect 59352 258660 59470 261232
rect 47770 258466 59470 258660
rect 60792 257466 61412 264078
rect 62712 262500 62740 265424
rect 63290 262500 63332 265424
rect 62712 262402 63332 262500
rect 50170 257424 61412 257466
rect 50170 257338 60826 257424
rect 50170 254676 50450 257338
rect 52008 257232 60826 257338
rect 52008 254676 56554 257232
rect 50170 254660 56554 254676
rect 60330 254660 60826 257232
rect 50170 254504 60826 254660
rect 61370 254504 61412 257424
rect 50170 254466 61412 254504
rect 60792 254422 61412 254466
rect 52578 253402 63292 253466
rect 52578 250538 52654 253402
rect 53746 253396 63292 253402
rect 53746 250548 56204 253396
rect 63216 250548 63292 253396
rect 53746 250538 63292 250548
rect 52578 250466 63292 250538
rect 63672 245466 64292 266958
rect 40984 245434 64292 245466
rect 40984 245388 63706 245434
rect 40984 238362 41066 245388
rect 43530 245296 63706 245388
rect 43530 242590 56394 245296
rect 63344 242590 63706 245296
rect 43530 242510 63706 242590
rect 64256 242510 64292 245434
rect 43530 242466 64292 242510
rect 43530 238362 43612 242466
rect 63672 242358 64292 242466
rect 64632 241466 65252 267918
rect 65592 253422 66212 268878
rect 65592 250498 65618 253422
rect 66168 250498 66212 253422
rect 65592 250386 66212 250498
rect 66552 249434 67172 269838
rect 393442 269370 394228 269470
rect 393442 266556 393536 269370
rect 394142 266556 394228 269370
rect 393442 266474 394228 266556
rect 394044 262208 394224 266474
rect 409094 265462 409274 265476
rect 408466 265334 409274 265462
rect 408466 262926 408538 265334
rect 409192 262926 409274 265334
rect 408466 262854 409274 262926
rect 409094 262244 409274 262854
rect 394504 261336 395406 261450
rect 394504 258566 394590 261336
rect 395320 258566 395406 261336
rect 394504 258468 395406 258566
rect 409686 257378 410808 257470
rect 409686 254558 409786 257378
rect 410720 254558 410808 257378
rect 409686 254452 410808 254558
rect 211712 253384 212610 253472
rect 211712 250572 211800 253384
rect 212518 250572 212610 253384
rect 211712 250470 212610 250572
rect 241812 253384 242710 253472
rect 241812 250572 241900 253384
rect 242618 250572 242710 253384
rect 241812 250470 242710 250572
rect 272232 253384 272620 253472
rect 272232 250470 272620 250572
rect 302162 253384 302714 253472
rect 302162 250470 302714 250572
rect 332112 253384 333010 253472
rect 332112 250572 332200 253384
rect 332918 250572 333010 253384
rect 332112 250470 333010 250572
rect 362212 253384 363110 253472
rect 362212 250572 362300 253384
rect 363018 250572 363110 253384
rect 362212 250470 363110 250572
rect 392572 253384 393110 253472
rect 393018 250572 393110 253384
rect 392572 250470 393110 250572
rect 66552 246510 66582 249434
rect 67132 246510 67172 249434
rect 66552 246348 67172 246510
rect 196676 249384 197618 249464
rect 196676 246554 196766 249384
rect 197520 246554 197618 249384
rect 196676 246468 197618 246554
rect 226776 249384 227718 249464
rect 226776 246554 226866 249384
rect 227620 246554 227718 249384
rect 226776 246468 227718 246554
rect 256876 249384 257818 249464
rect 256876 246554 256966 249384
rect 257720 246554 257818 249384
rect 287156 249384 287658 249464
rect 347176 249384 348118 249464
rect 256876 246468 257818 246554
rect 317354 246468 317802 246554
rect 347176 246554 347266 249384
rect 348020 246554 348118 249384
rect 347176 246468 348118 246554
rect 377176 249384 378118 249464
rect 377176 246554 377266 249384
rect 378020 246554 378118 249384
rect 377176 246468 378118 246554
rect 407176 249384 408118 249464
rect 407176 246554 407266 249384
rect 408020 246554 408118 249384
rect 407176 246468 408118 246554
rect 650618 249440 651238 277798
rect 658882 277774 674084 277842
rect 658856 277410 673450 277456
rect 658856 277396 670884 277410
rect 658856 276900 658916 277396
rect 663090 276900 670884 277396
rect 651578 253422 652198 276844
rect 658856 276816 670884 276900
rect 670818 276074 670884 276816
rect 673364 276074 673450 277410
rect 674016 276820 674084 277774
rect 676564 276820 676628 278356
rect 674016 276774 676628 276820
rect 670818 276016 673450 276074
rect 651578 250496 651612 253422
rect 652172 250496 652198 253422
rect 651578 250392 652198 250496
rect 650618 246514 650646 249440
rect 651206 246514 651238 249440
rect 650618 246296 651238 246514
rect 212568 245420 213540 245462
rect 212568 242526 212622 245420
rect 213464 242526 213540 245420
rect 212568 242464 213540 242526
rect 242668 245420 243640 245462
rect 242668 242526 242722 245420
rect 243564 242526 243640 245420
rect 242668 242464 243640 242526
rect 272982 245420 273314 245462
rect 272982 242464 273314 242526
rect 303168 245420 303460 245462
rect 303168 242464 303460 242526
rect 332968 245420 333940 245462
rect 332968 242526 333022 245420
rect 333864 242526 333940 245420
rect 332968 242464 333940 242526
rect 363068 245420 364040 245462
rect 363068 242526 363122 245420
rect 363964 242526 364040 245420
rect 363068 242464 364040 242526
rect 393210 245420 393800 245462
rect 393210 242464 393800 242526
rect 40984 238266 43612 238362
rect 44196 241430 65252 241466
rect 44196 241358 64656 241430
rect 44196 234532 44254 241358
rect 46718 241330 64656 241358
rect 46718 238624 56424 241330
rect 63344 238624 64656 241330
rect 46718 238506 64656 238624
rect 65206 238506 65252 241430
rect 46718 238466 65252 238506
rect 197542 241402 198398 241470
rect 197542 238534 197632 241402
rect 198322 238534 198398 241402
rect 197542 238480 198398 238534
rect 227642 241402 228498 241470
rect 227642 238534 227732 241402
rect 228422 238534 228498 241402
rect 227642 238480 228498 238534
rect 257742 241402 258598 241470
rect 257742 238534 257832 241402
rect 258522 238534 258598 241402
rect 257742 238480 258598 238534
rect 288068 241402 288566 241470
rect 288068 238480 288566 238534
rect 318226 241402 318574 241470
rect 318226 238480 318574 238534
rect 348042 241402 348898 241470
rect 348042 238534 348132 241402
rect 348822 238534 348898 241402
rect 348042 238480 348898 238534
rect 378042 241402 378898 241470
rect 378042 238534 378132 241402
rect 378822 238534 378898 241402
rect 378042 238480 378898 238534
rect 408410 241402 408734 241470
rect 408410 238480 408734 238534
rect 652538 241428 653158 275876
rect 653498 245430 654118 274916
rect 658950 274502 669812 274574
rect 658950 274494 667296 274502
rect 658950 274000 659050 274494
rect 663076 274000 667296 274494
rect 654458 265422 655078 273956
rect 658950 273938 667296 274000
rect 667216 273206 667296 273938
rect 669756 273206 669812 274502
rect 667216 273138 669812 273206
rect 655418 269424 656038 273004
rect 655418 266502 655458 269424
rect 655992 266502 656038 269424
rect 655418 266386 656038 266502
rect 654458 262500 654500 265422
rect 655034 262500 655078 265422
rect 654458 262362 655078 262500
rect 656378 257418 656998 272036
rect 657338 261436 657958 271082
rect 657338 258514 657374 261436
rect 657908 258514 657958 261436
rect 657338 258390 657958 258514
rect 656378 254496 656412 257418
rect 656946 254496 656998 257418
rect 656378 254386 656998 254496
rect 666890 249296 676670 249476
rect 666890 249288 674156 249296
rect 666890 246662 667058 249288
rect 669642 246662 674156 249288
rect 666890 246616 674156 246662
rect 676452 246616 676670 249296
rect 666890 246466 676670 246616
rect 653498 242520 653536 245430
rect 654058 242520 654118 245430
rect 653498 242362 654118 242520
rect 652538 238518 652578 241428
rect 653100 238518 653158 241428
rect 46718 234532 46802 238466
rect 64632 238400 65252 238466
rect 652538 238266 653158 238518
rect 44196 234466 46802 234532
rect 47786 237372 63250 237466
rect 47786 237366 56424 237372
rect 47786 234588 47980 237366
rect 50678 234594 56424 237366
rect 63122 234594 63250 237372
rect 50678 234588 63250 234594
rect 47786 234466 63250 234588
rect 210866 237386 211814 237474
rect 210866 234540 210958 237386
rect 211722 234540 211814 237386
rect 210866 234448 211814 234540
rect 240966 237386 241914 237474
rect 240966 234540 241058 237386
rect 241822 234540 241914 237386
rect 240966 234448 241914 234540
rect 271344 237386 272014 237474
rect 271922 234540 272014 237386
rect 331414 237386 332214 237474
rect 271344 234448 272014 234540
rect 302022 234540 302114 237290
rect 301514 234448 302114 234540
rect 332122 234540 332214 237386
rect 331414 234448 332214 234540
rect 361366 237386 362314 237474
rect 361366 234540 361458 237386
rect 362222 234540 362314 237386
rect 361366 234448 362314 234540
rect 391834 237386 392314 237474
rect 392222 234540 392314 237386
rect 391834 234448 392314 234540
rect 44186 233340 63160 233466
rect 44186 230606 56406 233340
rect 63018 230606 63160 233340
rect 44186 230466 63160 230606
rect 195988 233390 196616 233464
rect 195988 230538 196058 233390
rect 196556 230538 196616 233390
rect 195988 230466 196616 230538
rect 226088 233390 226716 233464
rect 226088 230538 226158 233390
rect 226656 230538 226716 233390
rect 226088 230466 226716 230538
rect 256188 233390 256816 233464
rect 256188 230538 256258 233390
rect 256756 230538 256816 233390
rect 256188 230466 256816 230538
rect 286288 233390 286916 233464
rect 286288 230538 286358 233390
rect 286856 230538 286916 233390
rect 286288 230466 286916 230538
rect 316388 233390 317016 233464
rect 316388 230538 316458 233390
rect 316956 230538 317016 233390
rect 316388 230466 317016 230538
rect 346488 233390 347116 233464
rect 346488 230538 346558 233390
rect 347056 230538 347116 233390
rect 346488 230466 347116 230538
rect 376488 233390 377116 233464
rect 376488 230538 376558 233390
rect 377056 230538 377116 233390
rect 376488 230466 377116 230538
rect 406660 233390 407116 233464
rect 407056 230538 407116 233390
rect 406660 230466 407116 230538
rect 44198 197498 46798 230466
rect 598368 212326 610962 212504
rect 598368 209740 598598 212326
rect 601098 209740 607452 212326
rect 609952 209740 610962 212326
rect 598368 209504 610962 209740
rect 641044 212352 642108 212460
rect 641044 209640 641152 212352
rect 642010 209640 642108 212352
rect 641044 209528 642108 209640
rect 596262 208442 605388 208502
rect 596262 207926 596332 208442
rect 597664 208434 605388 208442
rect 597664 207934 602456 208434
rect 605326 207934 605388 208434
rect 597664 207926 605388 207934
rect 596262 207862 605388 207926
rect 610642 207692 610962 209504
rect 641362 207684 641682 209528
rect 598496 197778 601174 197876
rect 44198 197454 52344 197498
rect 44198 196934 51420 197454
rect 52282 196934 52344 197454
rect 598496 197108 598684 197778
rect 601038 197528 601174 197778
rect 601038 197492 606976 197528
rect 601038 197238 606016 197492
rect 606936 197238 606976 197492
rect 601038 197208 606976 197238
rect 601038 197108 601174 197208
rect 598496 196992 601174 197108
rect 44198 196858 52344 196934
rect 44198 176742 46798 196858
rect 596072 184442 605388 184502
rect 596072 183902 596116 184442
rect 596848 184418 605388 184442
rect 596848 183918 602456 184418
rect 605326 183918 605388 184418
rect 596848 183902 605388 183918
rect 596072 183862 605388 183902
rect 41864 176610 46798 176742
rect 41864 173284 42002 176610
rect 45608 173284 46798 176610
rect 41864 173126 46798 173284
rect 42646 171444 52246 171498
rect 42646 170908 42828 171444
rect 45682 171440 52246 171444
rect 45682 170920 51312 171440
rect 52174 170920 52246 171440
rect 45682 170908 52246 170920
rect 42646 170858 52246 170908
rect 598496 167138 601174 167236
rect 598496 166468 598684 167138
rect 601038 166892 601174 167138
rect 601038 166866 606976 166892
rect 601038 166608 605986 166866
rect 606932 166608 606976 166866
rect 601038 166572 606976 166608
rect 601038 166468 601174 166572
rect 598496 166352 601174 166468
rect 594072 158446 605388 158502
rect 594072 157906 594114 158446
rect 596846 158430 605388 158446
rect 596846 157930 602430 158430
rect 605300 157930 605388 158430
rect 596846 157906 605388 157930
rect 594072 157862 605388 157906
rect 42578 145450 52178 145498
rect 42578 144914 42842 145450
rect 45696 145432 52178 145450
rect 45696 144914 51246 145432
rect 42578 144912 51246 144914
rect 52108 144912 52178 145432
rect 42578 144858 52178 144912
rect 598496 136498 601174 136596
rect 598496 135828 598684 136498
rect 601038 136256 601174 136498
rect 601038 136230 606976 136256
rect 601038 135964 605972 136230
rect 606926 135964 606976 136230
rect 601038 135936 606976 135964
rect 601038 135828 601174 135936
rect 598496 135712 601174 135828
rect 594072 132440 605388 132502
rect 594072 131900 594124 132440
rect 596856 132414 605388 132440
rect 596856 131914 602456 132414
rect 605326 131914 605388 132414
rect 596856 131900 605388 131914
rect 594072 131862 605388 131900
rect 42578 119446 52178 119498
rect 42578 118910 42832 119446
rect 45686 119438 52178 119446
rect 45686 118918 51242 119438
rect 52104 118918 52178 119438
rect 45686 118910 52178 118918
rect 42578 118858 52178 118910
rect 594072 106446 605388 106502
rect 594072 105906 594126 106446
rect 596858 106426 605388 106446
rect 596858 105926 602460 106426
rect 605330 105926 605388 106426
rect 596858 105906 605388 105926
rect 594072 105862 605388 105906
rect 598496 105620 601174 105676
rect 598496 105594 606976 105620
rect 598496 105578 605980 105594
rect 598496 104908 598684 105578
rect 601038 105326 605980 105578
rect 606942 105326 606976 105594
rect 601038 105300 606976 105326
rect 601038 104908 601174 105300
rect 598496 104792 601174 104908
rect 626002 98760 626322 102316
rect 656722 98804 657042 102238
rect 625442 98656 626852 98760
rect 625442 96074 625556 98656
rect 626744 96074 626852 98656
rect 636080 98622 636994 98758
rect 636080 96584 636216 98622
rect 636858 96584 636994 98622
rect 636080 96434 636994 96584
rect 656284 98712 657602 98804
rect 625442 95956 626852 96074
rect 636354 94448 636674 96434
rect 656284 96142 656422 98712
rect 657500 96142 657602 98712
rect 656284 96050 657602 96142
rect 42578 93444 52178 93498
rect 42578 92908 42828 93444
rect 45682 93434 52178 93444
rect 45682 92914 51246 93434
rect 52108 92914 52178 93434
rect 45682 92908 52178 92914
rect 42578 92858 52178 92908
rect 41864 82706 45778 82794
rect 41864 78242 41946 82706
rect 45672 78242 45778 82706
rect 632354 80924 632674 82062
rect 640354 81016 640674 82000
rect 632072 80776 633010 80924
rect 594072 80456 605388 80502
rect 594072 79916 594120 80456
rect 596852 80438 605388 80456
rect 596852 79938 602454 80438
rect 605324 79938 605388 80438
rect 596852 79916 605388 79938
rect 594072 79862 605388 79916
rect 41864 78154 45778 78242
rect 632072 78326 632200 80776
rect 632864 78326 633010 80776
rect 632072 78198 633010 78326
rect 640098 80900 640922 81016
rect 640098 78256 640210 80900
rect 640810 78256 640922 80900
rect 640098 78134 640922 78256
rect 41858 72802 45772 72890
rect 41858 68338 41922 72802
rect 45648 68338 45772 72802
rect 41858 68250 45772 68338
rect 41862 67438 52362 67498
rect 41862 66902 41936 67438
rect 45690 67436 52362 67438
rect 45690 66916 51444 67436
rect 52306 66916 52362 67436
rect 45690 66902 52362 66916
rect 41862 66858 52362 66902
rect 41874 51988 58536 52122
rect 41874 48404 42006 51988
rect 45590 51954 58536 51988
rect 45590 48404 54526 51954
rect 41874 48370 54526 48404
rect 58210 48370 58536 51954
rect 143324 50624 144738 50688
rect 143324 50004 143390 50624
rect 144652 50004 144738 50624
rect 143324 49936 144738 50004
rect 143860 49638 144040 49936
rect 41874 48222 58536 48370
rect 641936 47627 650202 48027
rect 142560 45396 142740 47256
rect 141776 45394 142866 45396
rect 141376 45306 142866 45394
rect 141376 44206 141442 45306
rect 142810 44206 142866 45306
rect 141376 44130 142866 44206
rect 143440 40762 143620 47296
rect 144740 41158 144920 47340
rect 241680 46616 246056 46692
rect 241680 42842 241740 46616
rect 245986 42842 246056 46616
rect 241680 42784 246056 42842
rect 251302 46630 255700 46684
rect 251302 42856 251392 46630
rect 255638 42856 255700 46630
rect 251302 42788 255700 42856
rect 641936 43988 643718 47627
rect 661270 47282 669426 47320
rect 648104 47124 649670 47188
rect 648104 46660 648166 47124
rect 649608 46660 649670 47124
rect 648104 46590 649670 46660
rect 641936 42198 641994 43988
rect 643660 42198 643718 43988
rect 653432 45026 656912 47054
rect 661270 47030 666460 47282
rect 669380 47030 669426 47282
rect 661270 46991 669426 47030
rect 653432 42634 653578 45026
rect 656772 42634 656912 45026
rect 653432 42488 656912 42634
rect 641936 42164 643718 42198
rect 144740 41148 150516 41158
rect 144740 40988 149618 41148
rect 150440 40988 150516 41148
rect 144740 40978 150516 40988
rect 143440 40752 148940 40762
rect 143440 40592 148086 40752
rect 148908 40592 148940 40752
rect 143440 40582 148940 40592
rect 208850 19412 209170 19578
rect 208850 18506 208868 19412
rect 209130 18506 209170 19412
rect 204960 18004 207956 18076
rect 204960 17128 205020 18004
rect 207872 17128 207956 18004
rect 204960 17072 207956 17128
rect 208850 16308 209170 18506
rect 210400 18010 210720 19578
rect 210400 17104 210420 18010
rect 210682 17104 210720 18010
rect 210400 16308 210720 17104
rect 211950 19426 212270 19578
rect 211950 18520 211980 19426
rect 212242 18520 212270 19426
rect 211950 16308 212270 18520
rect 213500 18014 213820 19578
rect 213500 17108 213514 18014
rect 213776 17108 213820 18014
rect 213500 16308 213820 17108
rect 215050 19422 215370 19578
rect 215050 18516 215070 19422
rect 215332 18516 215370 19422
rect 215050 16308 215370 18516
rect 216600 18018 216920 19578
rect 216600 17112 216622 18018
rect 216884 17112 216920 18018
rect 216600 16308 216920 17112
rect 218150 19422 218470 19578
rect 218150 18516 218164 19422
rect 218426 18516 218470 19422
rect 218150 16308 218470 18516
rect 219700 18010 220020 19578
rect 219700 17104 219726 18010
rect 219988 17104 220020 18010
rect 219700 16308 220020 17104
rect 221250 19434 221570 19578
rect 221250 18528 221272 19434
rect 221534 18528 221570 19434
rect 221250 16308 221570 18528
rect 222800 18036 223120 19578
rect 234818 19380 237824 19480
rect 234818 18544 234884 19380
rect 237754 18544 237824 19380
rect 234818 18470 237824 18544
rect 222800 17130 222828 18036
rect 223090 17130 223120 18036
rect 222800 16308 223120 17130
<< via4 >>
rect 575762 990884 580384 993314
rect 670928 995628 676500 996584
rect 585758 990898 590380 993328
rect 670976 990354 673264 992530
rect 47836 989738 49748 990276
rect 55820 989738 56394 990278
rect 50242 988774 52154 989312
rect 55824 988778 56398 989318
rect 658430 986872 663120 987376
rect 667268 986872 669770 987386
rect 41034 985878 43574 986448
rect 55804 985886 56378 986436
rect 44242 984918 46772 985498
rect 55804 984916 56408 985478
rect 52628 983968 53766 984510
rect 55802 983958 56376 984520
rect 658380 983984 663118 984492
rect 670858 983950 673384 984536
rect 658362 983028 663100 983536
rect 674056 982988 676582 983574
rect 44278 951976 46734 953030
rect 41068 950394 43524 951448
rect 674734 900074 675740 901112
rect 671566 898466 672596 899504
rect 674116 855052 675180 856116
rect 671570 853442 672638 854522
rect 47908 837800 49694 842324
rect 47908 827868 49694 832392
rect 667284 828630 669732 833206
rect 44278 826176 46734 827230
rect 41068 824594 43524 825648
rect 667270 818636 669718 823212
rect 44278 784576 46734 785630
rect 41068 782994 43524 784048
rect 44278 739776 46734 740830
rect 41068 738194 43524 739248
rect 44278 696576 46734 697630
rect 41068 694994 43524 696048
rect 44278 653376 46734 654430
rect 41068 651794 43524 652848
rect 44278 611236 46734 612290
rect 41068 609654 43524 610708
rect 44278 566976 46734 568030
rect 41068 565394 43524 566448
rect 667336 514056 669706 518582
rect 667350 504066 669720 508592
rect 50364 493250 52092 497732
rect 50352 483260 52080 487742
rect 44278 439376 46734 440430
rect 41068 437794 43524 438848
rect 664134 425684 666540 430390
rect 664112 415856 666528 420462
rect 44278 396176 46734 397230
rect 41068 394594 43524 395648
rect 44278 353976 46734 355030
rect 41068 352394 43524 353448
rect 44278 309776 46734 310830
rect 41068 308194 43524 309248
rect 44228 275888 46762 277262
rect 52652 276882 53730 278014
rect 658950 277842 663094 278344
rect 55790 276854 56378 277420
rect 55782 275898 56406 276442
rect 42830 269378 43528 275458
rect 55790 274944 56414 275488
rect 50248 272078 52134 273390
rect 55782 272052 56378 272618
rect 47848 270310 49746 271652
rect 55782 271088 56486 271656
rect 58532 266504 59082 269428
rect 48050 258676 49608 261338
rect 56554 258660 59352 261232
rect 62740 262500 63290 265424
rect 50450 254676 52008 257338
rect 56554 254660 60330 257232
rect 60826 254504 61370 257424
rect 52654 250538 53746 253402
rect 56204 250548 63216 253396
rect 41066 238362 43530 245388
rect 56394 242590 63344 245296
rect 63706 242510 64256 245434
rect 65618 250498 66168 253422
rect 393536 266556 394142 269370
rect 408538 262926 409192 265334
rect 394590 258566 395320 261336
rect 409786 254558 410720 257378
rect 211800 250572 212518 253384
rect 241900 250572 242618 253384
rect 272232 250572 272620 253384
rect 302162 250572 302714 253384
rect 332200 250572 332918 253384
rect 362300 250572 363018 253384
rect 392572 250572 393018 253384
rect 66582 246510 67132 249434
rect 196766 246554 197520 249384
rect 226866 246554 227620 249384
rect 256966 246554 257720 249384
rect 287156 246790 287658 249384
rect 317354 246554 317802 249324
rect 347266 246554 348020 249384
rect 377266 246554 378020 249384
rect 407266 246554 408020 249384
rect 658916 276900 663090 277396
rect 670884 276074 673364 277410
rect 674084 276820 676564 278356
rect 651612 250496 652172 253422
rect 650646 246514 651206 249440
rect 212622 242526 213464 245420
rect 242722 242526 243564 245420
rect 272982 242526 273314 245420
rect 303168 242526 303460 245420
rect 333022 242526 333864 245420
rect 363122 242526 363964 245420
rect 393210 242526 393800 245420
rect 44254 234532 46718 241358
rect 56424 238624 63344 241330
rect 64656 238506 65206 241430
rect 197632 238534 198322 241402
rect 227732 238534 228422 241402
rect 257832 238534 258522 241402
rect 288068 238534 288566 241402
rect 318226 238534 318574 241402
rect 348132 238534 348822 241402
rect 378132 238534 378822 241402
rect 408410 238534 408734 241402
rect 659050 274000 663076 274494
rect 667296 273206 669756 274502
rect 655458 266502 655992 269424
rect 654500 262500 655034 265422
rect 657374 258514 657908 261436
rect 656412 254496 656946 257418
rect 667058 246662 669642 249288
rect 674156 246616 676452 249296
rect 653536 242520 654058 245430
rect 652578 238518 653100 241428
rect 47980 234588 50678 237366
rect 56424 234594 63122 237372
rect 210958 234540 211722 237386
rect 241058 234540 241822 237386
rect 271344 234540 271922 237386
rect 301514 234540 302022 237290
rect 331414 234540 332122 237386
rect 361458 234540 362222 237386
rect 391834 234540 392222 237386
rect 56406 230606 63018 233340
rect 196058 230538 196556 233390
rect 226158 230538 226656 233390
rect 256258 230538 256756 233390
rect 286358 230538 286856 233390
rect 316458 230538 316956 233390
rect 346558 230538 347056 233390
rect 376558 230538 377056 233390
rect 406660 230538 407056 233390
rect 598598 209740 601098 212326
rect 607452 209740 609952 212326
rect 641152 209640 642010 212352
rect 596332 207926 597664 208442
rect 602456 207934 605326 208434
rect 51420 196934 52282 197454
rect 598684 197108 601038 197778
rect 606016 197238 606936 197492
rect 596116 183902 596848 184442
rect 602456 183918 605326 184418
rect 42002 173284 45608 176610
rect 42828 170908 45682 171444
rect 51312 170920 52174 171440
rect 598684 166468 601038 167138
rect 605986 166608 606932 166866
rect 594114 157906 596846 158446
rect 602430 157930 605300 158430
rect 42842 144914 45696 145450
rect 51246 144912 52108 145432
rect 598684 135828 601038 136498
rect 605972 135964 606926 136230
rect 594124 131900 596856 132440
rect 602456 131914 605326 132414
rect 42832 118910 45686 119446
rect 51242 118918 52104 119438
rect 594126 105906 596858 106446
rect 602460 105926 605330 106426
rect 598684 104908 601038 105578
rect 605980 105326 606942 105594
rect 625556 96074 626744 98656
rect 636216 96584 636858 98622
rect 656422 96142 657500 98712
rect 42828 92908 45682 93444
rect 51246 92914 52108 93434
rect 41946 78242 45672 82706
rect 594120 79916 596852 80456
rect 602454 79938 605324 80438
rect 632200 78326 632864 80776
rect 640210 78256 640810 80900
rect 41922 68338 45648 72802
rect 41936 66902 45690 67438
rect 51444 66916 52306 67436
rect 42006 48404 45590 51988
rect 54526 48370 58210 51954
rect 143390 50004 144652 50624
rect 141442 44206 142810 45306
rect 241740 42842 245986 46616
rect 251392 42856 255638 46630
rect 648166 46660 649608 47124
rect 666460 47030 669380 47282
rect 208868 18506 209130 19412
rect 205020 17128 207872 18004
rect 210420 17104 210682 18010
rect 211980 18520 212242 19426
rect 213514 17108 213776 18014
rect 215070 18516 215332 19422
rect 216622 17112 216884 18018
rect 218164 18516 218426 19422
rect 219726 17104 219988 18010
rect 221272 18528 221534 19434
rect 234884 18544 237754 19380
rect 222828 17130 223090 18036
<< metal5 >>
rect 52598 996584 676660 996702
rect 52598 995628 670928 996584
rect 676500 995628 676660 996584
rect 52598 995502 676660 995628
rect 47798 990276 49798 990466
rect 47798 989738 47836 990276
rect 49748 989738 49798 990276
rect 47798 842324 49798 989738
rect 47798 837800 47908 842324
rect 49694 837800 49798 842324
rect 47798 832392 49798 837800
rect 47798 827868 47908 832392
rect 49694 827868 49798 832392
rect 47798 271652 49798 827868
rect 47798 270310 47848 271652
rect 49746 270310 49798 271652
rect 47798 261338 49798 270310
rect 47798 258676 48050 261338
rect 49608 258676 49798 261338
rect 47798 258484 49798 258676
rect 50198 989312 52198 990466
rect 50198 988774 50242 989312
rect 52154 988774 52198 989312
rect 50198 497732 52198 988774
rect 50198 493250 50364 497732
rect 52092 493250 52198 497732
rect 50198 487742 52198 493250
rect 50198 483260 50352 487742
rect 52080 483260 52198 487742
rect 50198 273390 52198 483260
rect 50198 272078 50248 273390
rect 52134 272078 52198 273390
rect 50198 257338 52198 272078
rect 50198 254676 50450 257338
rect 52008 254676 52198 257338
rect 50198 254498 52198 254676
rect 52598 984510 53798 995502
rect 52598 983968 52628 984510
rect 53766 983968 53798 984510
rect 52598 278014 53798 983968
rect 52598 276882 52652 278014
rect 53730 276882 53798 278014
rect 52598 253402 53798 276882
rect 52598 250538 52654 253402
rect 53746 250538 53798 253402
rect 47836 237366 50836 237612
rect 47836 234588 47980 237366
rect 50678 234588 50836 237366
rect 47836 210498 50836 234588
rect 52598 217742 53798 250538
rect 54198 993902 676620 995102
rect 54198 983588 55398 993902
rect 575640 993328 666620 993396
rect 575640 993314 585758 993328
rect 575640 990884 575762 993314
rect 580384 990898 585758 993314
rect 590380 990898 666620 993328
rect 674020 992696 676620 993902
rect 580384 990884 666620 990898
rect 575640 990796 666620 990884
rect 55776 990278 56596 990308
rect 55776 989738 55820 990278
rect 56394 989738 56596 990278
rect 55776 989688 56596 989738
rect 55776 989318 57552 989348
rect 55776 988778 55824 989318
rect 56398 988778 57552 989318
rect 55776 988728 57552 988778
rect 664020 988388 666620 990796
rect 656038 987768 666620 988388
rect 655078 987376 663178 987428
rect 655078 986872 658430 987376
rect 663120 986872 663178 987376
rect 655078 986808 663178 986872
rect 55776 986436 60436 986468
rect 55776 985886 55804 986436
rect 56378 985886 60436 986436
rect 55776 985848 60436 985886
rect 55776 985478 61398 985508
rect 55776 984916 55804 985478
rect 56408 984916 61398 985478
rect 55776 984888 61398 984916
rect 55776 984520 62358 984548
rect 55776 983958 55802 984520
rect 56376 983958 62358 984520
rect 55776 983928 62358 983958
rect 652180 984492 663178 984548
rect 652180 983984 658380 984492
rect 663118 983984 663178 984492
rect 652180 983928 663178 983984
rect 54198 982968 63316 983588
rect 651228 983536 663178 983588
rect 651228 983028 658362 983536
rect 663100 983028 663178 983536
rect 651228 982968 663178 983028
rect 54198 278404 55398 982968
rect 664020 430390 666620 987768
rect 664020 425684 664134 430390
rect 666540 425684 666620 430390
rect 664020 420462 666620 425684
rect 664020 415856 664112 420462
rect 666528 415856 666620 420462
rect 54198 277784 63312 278404
rect 651226 278344 663158 278404
rect 651226 277842 658950 278344
rect 663094 277842 663158 278344
rect 651226 277784 663158 277842
rect 54198 249466 55398 277784
rect 55754 277420 62352 277444
rect 55754 276854 55790 277420
rect 56378 276854 62352 277420
rect 55754 276824 62352 276854
rect 652188 277396 663158 277444
rect 652188 276900 658916 277396
rect 663090 276900 663158 277396
rect 652188 276824 663158 276900
rect 55754 276442 61388 276484
rect 55754 275898 55782 276442
rect 56406 275898 61388 276442
rect 55754 275864 61388 275898
rect 55754 275488 60428 275524
rect 55754 274944 55790 275488
rect 56414 274944 60428 275488
rect 55754 274904 60428 274944
rect 655060 274494 663158 274564
rect 655060 274000 659050 274494
rect 663076 274000 663158 274494
rect 655060 273944 663158 274000
rect 664020 273604 666620 415856
rect 656026 272984 666620 273604
rect 55754 272618 57546 272644
rect 55754 272052 55782 272618
rect 56378 272052 57546 272618
rect 55754 272024 57546 272052
rect 55754 271656 56590 271684
rect 55754 271088 55782 271656
rect 56486 271088 56590 271656
rect 55754 271064 56590 271088
rect 664020 269466 666620 272984
rect 58388 269428 666620 269466
rect 58388 266504 58532 269428
rect 59082 269424 666620 269428
rect 59082 269370 655458 269424
rect 59082 266556 393536 269370
rect 394142 266556 655458 269370
rect 59082 266504 655458 266556
rect 58388 266502 655458 266504
rect 655992 266502 666620 269424
rect 58388 266466 666620 266502
rect 667220 987386 669820 987566
rect 667220 986872 667268 987386
rect 669770 986872 669820 987386
rect 667220 833206 669820 986872
rect 667220 828630 667284 833206
rect 669732 828630 669820 833206
rect 667220 823212 669820 828630
rect 667220 818636 667270 823212
rect 669718 818636 669820 823212
rect 667220 518582 669820 818636
rect 667220 514056 667336 518582
rect 669706 514056 669820 518582
rect 667220 508592 669820 514056
rect 667220 504066 667350 508592
rect 669720 504066 669820 508592
rect 667220 274502 669820 504066
rect 667220 273206 667296 274502
rect 669756 273206 669820 274502
rect 667220 265466 669820 273206
rect 62534 265424 669820 265466
rect 62534 262500 62740 265424
rect 63290 265422 669820 265424
rect 63290 265334 654500 265422
rect 63290 262926 408538 265334
rect 409192 262926 654500 265334
rect 63290 262500 654500 262926
rect 655034 262500 669820 265422
rect 62534 262466 669820 262500
rect 56370 261436 658090 261466
rect 56370 261336 657374 261436
rect 56370 261232 394590 261336
rect 56370 258660 56554 261232
rect 59352 258660 394590 261232
rect 56370 258566 394590 258660
rect 395320 258566 657374 261336
rect 56370 258514 657374 258566
rect 657908 258514 658090 261436
rect 56370 258466 658090 258514
rect 56370 257424 657076 257466
rect 56370 257232 60826 257424
rect 56370 254660 56554 257232
rect 60330 254660 60826 257232
rect 56370 254504 60826 254660
rect 61370 257418 657076 257424
rect 61370 257378 656412 257418
rect 61370 254558 409786 257378
rect 410720 254558 656412 257378
rect 61370 254504 656412 254558
rect 56370 254496 656412 254504
rect 656946 254496 657076 257418
rect 56370 254466 657076 254496
rect 56126 253422 670986 253466
rect 56126 253396 65618 253422
rect 56126 250548 56204 253396
rect 63216 250548 65618 253396
rect 56126 250498 65618 250548
rect 66168 253384 651612 253422
rect 66168 250572 211800 253384
rect 212518 250572 241900 253384
rect 242618 250572 272232 253384
rect 272620 250572 302162 253384
rect 302714 250572 332200 253384
rect 332918 250572 362300 253384
rect 363018 250572 392572 253384
rect 393018 250572 651612 253384
rect 66168 250498 651612 250572
rect 56126 250496 651612 250498
rect 652172 250496 670986 253422
rect 56126 250466 670986 250496
rect 54198 249440 669890 249466
rect 54198 249434 650646 249440
rect 54198 246510 66582 249434
rect 67132 249384 650646 249434
rect 67132 246554 196766 249384
rect 197520 246554 226866 249384
rect 227620 246554 256966 249384
rect 257720 246790 287156 249384
rect 287658 249324 347266 249384
rect 287658 246790 317354 249324
rect 257720 246554 317354 246790
rect 317802 246554 347266 249324
rect 348020 246554 377266 249384
rect 378020 246554 407266 249384
rect 408020 246554 650646 249384
rect 67132 246514 650646 246554
rect 651206 249288 669890 249440
rect 651206 246662 667058 249288
rect 669642 246662 669890 249288
rect 651206 246514 669890 246662
rect 67132 246510 669890 246514
rect 54198 246466 669890 246510
rect 54198 219342 55398 246466
rect 56278 245434 654222 245466
rect 56278 245296 63706 245434
rect 56278 242590 56394 245296
rect 63344 242590 63706 245296
rect 56278 242510 63706 242590
rect 64256 245430 654222 245434
rect 64256 245420 653536 245430
rect 64256 242526 212622 245420
rect 213464 242526 242722 245420
rect 243564 242526 272982 245420
rect 273314 242526 303168 245420
rect 303460 242526 333022 245420
rect 333864 242526 363122 245420
rect 363964 242526 393210 245420
rect 393800 242526 653536 245420
rect 64256 242520 653536 242526
rect 654058 242520 654222 245430
rect 64256 242510 654222 242520
rect 56278 242466 654222 242510
rect 56278 241430 653306 241466
rect 56278 241330 64656 241430
rect 56278 238624 56424 241330
rect 63344 238624 64656 241330
rect 56278 238506 64656 238624
rect 65206 241428 653306 241430
rect 65206 241402 652578 241428
rect 65206 238534 197632 241402
rect 198322 238534 227732 241402
rect 228422 238534 257832 241402
rect 258522 238534 288068 241402
rect 288566 238534 318226 241402
rect 318574 238534 348132 241402
rect 348822 238534 378132 241402
rect 378822 238534 408410 241402
rect 408734 238534 652578 241402
rect 65206 238518 652578 238534
rect 653100 238518 653306 241428
rect 65206 238506 653306 238518
rect 56278 238466 653306 238506
rect 56288 237386 605390 237466
rect 56288 237372 210958 237386
rect 56288 234594 56424 237372
rect 63122 234594 210958 237372
rect 56288 234540 210958 234594
rect 211722 234540 241058 237386
rect 241822 234540 271344 237386
rect 271922 237290 331414 237386
rect 271922 234540 301514 237290
rect 302022 234540 331414 237290
rect 332122 234540 361458 237386
rect 362222 234540 391834 237386
rect 392222 234540 605390 237386
rect 56288 234466 605390 234540
rect 56296 233390 601374 233466
rect 56296 233340 196058 233390
rect 56296 230606 56406 233340
rect 63018 230606 196058 233340
rect 56296 230538 196058 230606
rect 196556 230538 226158 233390
rect 226656 230538 256258 233390
rect 256756 230538 286358 233390
rect 286856 230538 316458 233390
rect 316956 230538 346558 233390
rect 347056 230538 376558 233390
rect 377056 230538 406660 233390
rect 407056 230538 601374 233390
rect 56296 230466 601374 230538
rect 598374 212326 601374 230466
rect 47836 209858 53232 210498
rect 574646 209858 596910 210498
rect 47836 184498 50836 209858
rect 596270 208502 596910 209858
rect 598374 209740 598598 212326
rect 601098 209740 601374 212326
rect 596270 208442 597742 208502
rect 596270 207926 596332 208442
rect 597664 207926 597742 208442
rect 596270 207862 597742 207926
rect 598374 197778 601374 209740
rect 598374 197498 598684 197778
rect 51344 197454 53216 197498
rect 51344 196934 51420 197454
rect 52282 196934 53216 197454
rect 51344 196858 53216 196934
rect 574646 197108 598684 197498
rect 601038 197108 601374 197778
rect 574646 196858 601374 197108
rect 47836 183858 53212 184498
rect 574646 184442 596910 184498
rect 574646 183902 596116 184442
rect 596848 183902 596910 184442
rect 574646 183858 596910 183902
rect 41768 176610 45768 176874
rect 41768 173284 42002 176610
rect 45608 173284 45768 176610
rect 41768 171444 45768 173284
rect 41768 170908 42828 171444
rect 45682 170908 45768 171444
rect 41768 145450 45768 170908
rect 47836 166788 50836 183858
rect 598374 171498 601374 196858
rect 51246 171440 53240 171498
rect 51246 170920 51312 171440
rect 52174 170920 53240 171440
rect 51246 170858 53240 170920
rect 574646 170858 601374 171498
rect 41768 144914 42842 145450
rect 45696 144914 45768 145450
rect 41768 119446 45768 144914
rect 41768 118910 42832 119446
rect 45686 118910 45768 119446
rect 41768 93444 45768 118910
rect 41768 92908 42828 93444
rect 45682 92908 45768 93444
rect 41768 82706 45768 92908
rect 41768 78242 41946 82706
rect 45672 78242 45768 82706
rect 41768 72802 45768 78242
rect 41768 68338 41922 72802
rect 45648 68338 45768 72802
rect 41768 67438 45768 68338
rect 41768 66902 41936 67438
rect 45690 66902 45768 67438
rect 41768 51988 45768 66902
rect 41768 48404 42006 51988
rect 45590 48404 45768 51988
rect 41768 48074 45768 48404
rect 46836 158498 50836 166788
rect 598374 167138 601374 170858
rect 598374 166468 598684 167138
rect 601038 166468 601374 167138
rect 46836 157858 53220 158498
rect 574646 158446 596910 158498
rect 574646 157906 594114 158446
rect 596846 157906 596910 158446
rect 574646 157858 596910 157906
rect 46836 132498 50836 157858
rect 598374 145498 601374 166468
rect 51178 145432 53266 145498
rect 51178 144912 51246 145432
rect 52108 144912 53266 145432
rect 51178 144858 53266 144912
rect 574646 144858 601374 145498
rect 598374 136498 601374 144858
rect 598374 135828 598684 136498
rect 601038 135828 601374 136498
rect 46836 131858 53206 132498
rect 574646 132440 596910 132498
rect 574646 131900 594124 132440
rect 596856 131900 596910 132440
rect 574646 131858 596910 131900
rect 46836 106498 50836 131858
rect 598374 119498 601374 135828
rect 51178 119438 53266 119498
rect 51178 118918 51242 119438
rect 52104 118918 53266 119438
rect 51178 118858 53266 118918
rect 574646 118858 601374 119498
rect 46836 105858 53222 106498
rect 574646 106446 596910 106498
rect 574646 105906 594126 106446
rect 596858 105906 596910 106446
rect 574646 105858 596910 105906
rect 46836 80498 50836 105858
rect 598374 105578 601374 118858
rect 598374 104908 598684 105578
rect 601038 104908 601374 105578
rect 598374 93498 601374 104908
rect 51178 93434 53266 93498
rect 51178 92914 51246 93434
rect 52108 92914 53266 93434
rect 51178 92858 53266 92914
rect 574646 92858 601374 93498
rect 46836 79858 53168 80498
rect 574646 80456 596910 80498
rect 574646 79916 594120 80456
rect 596852 79916 596910 80456
rect 574646 79858 596910 79916
rect 46836 46788 50836 79858
rect 598374 67498 601374 92858
rect 51362 67436 53172 67498
rect 51362 66916 51444 67436
rect 52306 66916 53172 67436
rect 51362 66858 53172 66916
rect 574754 66858 601374 67498
rect 598374 52222 601374 66858
rect 54374 51954 601374 52222
rect 54374 48370 54526 51954
rect 58210 50624 601374 51954
rect 58210 50004 143390 50624
rect 144652 50004 601374 50624
rect 58210 48370 601374 50004
rect 54374 48222 601374 48370
rect 602390 208434 605390 234466
rect 607252 212352 669426 212504
rect 607252 212326 641152 212352
rect 607252 209740 607452 212326
rect 609952 209740 641152 212326
rect 607252 209640 641152 209740
rect 642010 209640 669426 212352
rect 607252 209504 669426 209640
rect 602390 207934 602456 208434
rect 605326 207934 605390 208434
rect 602390 184418 605390 207934
rect 666426 197528 669426 209504
rect 605976 197492 607594 197528
rect 605976 197238 606016 197492
rect 606936 197238 607594 197492
rect 605976 197208 607594 197238
rect 665238 197208 669426 197528
rect 602390 183918 602456 184418
rect 605326 183918 605390 184418
rect 602390 182210 605390 183918
rect 602390 181890 607594 182210
rect 602390 158430 605390 181890
rect 666426 166892 669426 197208
rect 605952 166866 607594 166892
rect 605952 166608 605986 166866
rect 606932 166608 607594 166866
rect 605952 166572 607594 166608
rect 665206 166572 669426 166892
rect 602390 157930 602430 158430
rect 605300 157930 605390 158430
rect 602390 151574 605390 157930
rect 602390 151254 607594 151574
rect 602390 132414 605390 151254
rect 666426 136256 669426 166572
rect 605940 136230 607594 136256
rect 605940 135964 605972 136230
rect 606926 135964 607594 136230
rect 605940 135936 607594 135964
rect 665164 135936 669426 136256
rect 602390 131914 602456 132414
rect 605326 131914 605390 132414
rect 602390 120938 605390 131914
rect 602390 120618 607610 120938
rect 602390 106426 605390 120618
rect 602390 105926 602460 106426
rect 605330 105926 605390 106426
rect 602390 98956 605390 105926
rect 666426 105620 669426 135936
rect 605940 105594 607594 105620
rect 605940 105326 605980 105594
rect 606942 105326 607594 105594
rect 605940 105300 607594 105326
rect 665176 105300 669426 105620
rect 602390 98712 657728 98956
rect 602390 98656 656422 98712
rect 602390 96074 625556 98656
rect 626744 98622 656422 98656
rect 626744 96584 636216 98622
rect 636858 96584 656422 98622
rect 626744 96142 656422 96584
rect 657500 96142 657728 98712
rect 626744 96074 657728 96142
rect 602390 95956 657728 96074
rect 602390 80438 605390 95956
rect 624824 89474 627824 95956
rect 643544 93474 646544 93588
rect 641906 93154 646544 93474
rect 624824 89154 629362 89474
rect 624824 89012 627824 89154
rect 643544 85474 646544 93154
rect 650994 92590 653994 95956
rect 666426 93406 669426 105300
rect 662522 93086 669426 93406
rect 650994 92270 657754 92590
rect 650994 90958 653994 92270
rect 666426 91774 669426 93086
rect 662484 91454 669426 91774
rect 650994 90638 657784 90958
rect 650994 90522 653994 90638
rect 666426 90142 669426 91454
rect 662504 89822 669426 90142
rect 641968 85154 646544 85474
rect 643544 81082 646544 85154
rect 666426 81082 669426 89822
rect 602390 79938 602454 80438
rect 605324 79938 605390 80438
rect 602390 47188 605390 79938
rect 632002 80900 669426 81082
rect 632002 80776 640210 80900
rect 632002 78326 632200 80776
rect 632864 78326 640210 80776
rect 632002 78256 640210 78326
rect 640810 78256 669426 80900
rect 632002 78082 669426 78256
rect 666426 47282 669426 78082
rect 602390 47124 649668 47188
rect 602390 46788 648166 47124
rect 46836 46660 648166 46788
rect 649608 46660 649668 47124
rect 666426 47030 666460 47282
rect 669380 47030 669426 47282
rect 666426 46978 669426 47030
rect 46836 46630 649668 46660
rect 46836 46616 251392 46630
rect 46836 45306 241740 46616
rect 46836 44206 141442 45306
rect 142810 44206 241740 45306
rect 46836 42842 241740 44206
rect 245986 42856 251392 46616
rect 255638 46588 649668 46630
rect 255638 45788 605390 46588
rect 255638 42856 605396 45788
rect 245986 42842 605396 42856
rect 46836 42788 605396 42842
rect 205820 19434 237824 19472
rect 205820 19426 221272 19434
rect 205820 19412 211980 19426
rect 205820 18506 208868 19412
rect 209130 18520 211980 19412
rect 212242 19422 221272 19426
rect 212242 18520 215070 19422
rect 209130 18516 215070 18520
rect 215332 18516 218164 19422
rect 218426 18528 221272 19422
rect 221534 19380 237824 19434
rect 221534 18544 234884 19380
rect 237754 18544 237824 19380
rect 221534 18528 237824 18544
rect 218426 18516 237824 18528
rect 209130 18506 237824 18516
rect 205820 18472 237824 18506
rect 204580 18036 224806 18072
rect 204580 18018 222828 18036
rect 204580 18014 216622 18018
rect 204580 18010 213514 18014
rect 204580 18004 210420 18010
rect 204580 17128 205020 18004
rect 207872 17128 210420 18004
rect 204580 17104 210420 17128
rect 210682 17108 213514 18010
rect 213776 17112 216622 18014
rect 216884 18010 222828 18018
rect 216884 17112 219726 18010
rect 213776 17108 219726 17112
rect 210682 17104 219726 17108
rect 219988 17130 222828 18010
rect 223090 17130 224806 18036
rect 219988 17104 224806 17130
rect 204580 17072 224806 17104
rect 204580 14000 205380 17072
rect 225246 15690 226046 18472
rect 224498 15370 226046 15690
rect 204580 13680 205930 14000
rect 204580 10620 205380 13680
rect 225246 12310 226046 15370
rect 224464 11990 226046 12310
rect 204580 10300 205808 10620
rect 204580 8096 205380 10300
rect 225246 8930 226046 11990
rect 224586 8610 226046 8930
rect 225246 7838 226046 8610
<< comment >>
rect 0 1037400 717600 1037600
rect 0 200 200 1037400
rect 717400 200 717600 1037400
rect 0 0 717600 200
use gpio_control_power_routing  gpio_control_power_routing_0
timestamp 1637447660
transform 1 0 -10 0 1 0
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_1
timestamp 1637447660
transform 1 0 -10 0 1 43200
box 6032 203748 55470 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_14
timestamp 1637595202
transform -1 0 717846 0 1 -81600
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_13
timestamp 1637595202
transform -1 0 717846 0 1 -36400
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_12
timestamp 1637595202
transform -1 0 717846 0 1 8600
box 6032 203748 46226 221470
use gpio_control_power_routing  gpio_control_power_routing_2
timestamp 1637447660
transform 1 0 -10 0 1 86400
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_3
timestamp 1637447660
transform 1 0 -10 0 1 129600
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_4
timestamp 1637447660
transform 1 0 -10 0 1 172800
box 6032 203748 55470 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_11
timestamp 1637595202
transform -1 0 717846 0 1 53800
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_10
timestamp 1637595202
transform -1 0 717846 0 1 98800
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_9
timestamp 1637595202
transform -1 0 717846 0 1 143800
box 6032 203748 46226 221470
use gpio_control_power_routing  gpio_control_power_routing_5
timestamp 1637447660
transform 1 0 -10 0 1 216000
box 6032 203748 55470 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_8
timestamp 1637595202
transform -1 0 717846 0 1 189000
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_7
timestamp 1637595202
transform -1 0 717846 0 1 277200
box 6032 203748 46226 221470
use gpio_control_power_routing  gpio_control_power_routing_6
timestamp 1637447660
transform 1 0 -10 0 1 343600
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_7
timestamp 1637447660
transform 1 0 -10 0 1 386800
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_8
timestamp 1637447660
transform 1 0 -10 0 1 430000
box 6032 203748 55470 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_6
timestamp 1637595202
transform -1 0 717846 0 1 321200
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_5
timestamp 1637595202
transform -1 0 717846 0 1 366200
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_4
timestamp 1637595202
transform -1 0 717846 0 1 411400
box 6032 203748 46226 221470
use gpio_control_power_routing  gpio_control_power_routing_9
timestamp 1637447660
transform 1 0 -10 0 1 473200
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_11
timestamp 1637447660
transform 1 0 -10 0 1 559600
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_10
timestamp 1637447660
transform 1 0 -10 0 1 516400
box 6032 203748 55470 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_3
timestamp 1637595202
transform -1 0 717846 0 1 456400
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_2
timestamp 1637595202
transform -1 0 717846 0 1 501600
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_1
timestamp 1637595202
transform -1 0 717846 0 1 546600
box 6032 203748 46226 221470
use gpio_control_power_routing  gpio_control_power_routing_12
timestamp 1637447660
transform 1 0 -10 0 1 602800
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_13
timestamp 1637447660
transform 1 0 -10 0 1 728600
box 6032 203748 55470 221470
use gpio_control_power_routing_top  gpio_control_power_routing_top_0
timestamp 1637524495
transform 0 1 -105400 -1 0 1037728
box 6032 203748 43870 221470
use gpio_control_power_routing_top  gpio_control_power_routing_top_1
timestamp 1637524495
transform 0 1 -54000 -1 0 1037728
box 6032 203748 43870 221470
use gpio_control_power_routing_top  gpio_control_power_routing_top_3
timestamp 1637524495
transform 0 1 48800 -1 0 1037728
box 6032 203748 43870 221470
use gpio_control_power_routing_top  gpio_control_power_routing_top_2
timestamp 1637524495
transform 0 1 -2600 -1 0 1037728
box 6032 203748 43870 221470
use gpio_control_power_routing_top  gpio_control_power_routing_top_4
timestamp 1637524495
transform 0 1 100400 -1 0 1037728
box 6032 203748 43870 221470
use gpio_control_power_routing_top  gpio_control_power_routing_top_5
timestamp 1637524495
transform 0 1 150800 -1 0 1037728
box 6032 203748 43870 221470
use gpio_control_power_routing_top  gpio_control_power_routing_top_6
timestamp 1637524495
transform 0 1 218200 -1 0 1037728
box 6032 203748 43870 221470
use gpio_control_power_routing_top  gpio_control_power_routing_top_7
timestamp 1637524495
transform 0 1 295200 -1 0 1037728
box 6032 203748 43870 221470
use gpio_control_power_routing_top  gpio_control_power_routing_top_8
timestamp 1637524495
transform 0 1 346600 -1 0 1037728
box 6032 203748 43870 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_0
timestamp 1637595202
transform -1 0 717836 0 1 725000
box 6032 203748 46226 221470
<< labels >>
flabel metal5 54316 219436 55324 219998 0 FreeSans 1600 0 0 0 vccd1_core
flabel metal5 52692 217826 53700 218388 0 FreeSans 1600 0 0 0 vssd1_core
flabel metal5 184480 230750 189228 233134 0 FreeSans 16000 0 0 0 vccd_core
flabel metal5 184522 234770 189540 236910 0 FreeSans 16000 0 0 0 vssd_core
flabel metal5 182216 238830 190118 240864 0 FreeSans 16000 0 0 0 vccd2_core
flabel metal5 182126 242838 190088 244986 0 FreeSans 16000 0 0 0 vssd2_core
flabel metal5 181918 254572 189876 257076 0 FreeSans 16000 0 0 0 vdda2_core
flabel metal5 181918 258660 189876 261164 0 FreeSans 16000 0 0 0 vssa2_core
flabel metal5 621960 246802 629984 249230 0 FreeSans 16000 0 0 0 vccd1_core
flabel metal5 621948 250708 629990 253036 0 FreeSans 16000 0 0 0 vssd1_core
flabel metal5 621550 262640 629508 265144 0 FreeSans 16000 0 0 0 vdda1_core
flabel metal5 621514 266692 629472 269196 0 FreeSans 16000 0 0 0 vssa1_core
flabel metal5 590480 230750 595228 233134 0 FreeSans 16000 0 0 0 vccd_core
flabel metal5 590522 234770 595540 236910 0 FreeSans 16000 0 0 0 vssd_core
flabel metal5 42966 171382 45564 172780 0 FreeSans 3200 0 0 0 vccd_core
flabel metal5 664092 267180 666518 267904 0 FreeSans 3200 0 0 0 vssa1_core
flabel metal5 667280 263142 669706 263866 0 FreeSans 3200 0 0 0 vdda1_core
flabel metal5 634330 96284 638114 98514 0 FreeSans 16000 0 0 0 vssd_core
flabel metal5 633452 78554 637236 80784 0 FreeSans 16000 0 0 0 vccd_core
flabel metal5 206106 18628 207168 19326 0 FreeSans 4800 0 0 0 vccd_core
flabel metal5 206018 17180 207080 17878 0 FreeSans 4800 0 0 0 vssd_core
flabel metal5 182024 250550 190042 253308 0 FreeSans 16000 0 0 0 vssd1_core
flabel metal5 182160 246638 190178 249396 0 FreeSans 16000 0 0 0 vccd1_core
flabel metal5 181852 266620 189870 269378 0 FreeSans 16000 0 0 0 vssa1_core
flabel metal5 181950 262574 189968 265332 0 FreeSans 16000 0 0 0 vdda1_core
flabel metal5 47904 265444 49660 265998 0 FreeSans 3200 0 0 0 vssa2_core
flabel metal5 50338 265444 52094 265998 0 FreeSans 3200 0 0 0 vdda2_core
flabel metal5 621512 258708 630212 261250 0 FreeSans 16000 0 0 0 vssa2_core
flabel metal5 621598 254668 630298 257210 0 FreeSans 16000 0 0 0 vdda2_core
flabel metal5 621936 242776 630636 245318 0 FreeSans 16000 0 0 0 vssd2_core
flabel metal5 621794 238736 630494 241278 0 FreeSans 16000 0 0 0 vccd2_core
<< end >>
