magic
tech sky130A
magscale 1 2
timestamp 1666101175
<< obsli1 >>
rect 1104 1071 18860 13617
<< obsm1 >>
rect 1104 892 18860 13728
<< metal2 >>
rect 1122 14200 1178 15000
rect 2594 14200 2650 15000
rect 4066 14200 4122 15000
rect 5538 14200 5594 15000
rect 7010 14200 7066 15000
rect 8482 14200 8538 15000
rect 9954 14200 10010 15000
rect 11426 14200 11482 15000
rect 12898 14200 12954 15000
rect 14370 14200 14426 15000
rect 15842 14200 15898 15000
rect 17314 14200 17370 15000
rect 18786 14200 18842 15000
rect 4986 0 5042 800
rect 14922 0 14978 800
<< obsm2 >>
rect 1234 14144 2538 14362
rect 2706 14144 4010 14362
rect 4178 14144 5482 14362
rect 5650 14144 6954 14362
rect 7122 14144 8426 14362
rect 8594 14144 9898 14362
rect 10066 14144 11370 14362
rect 11538 14144 12842 14362
rect 13010 14144 14314 14362
rect 14482 14144 15786 14362
rect 15954 14144 17258 14362
rect 17426 14144 18730 14362
rect 1178 856 18842 14144
rect 1178 734 4930 856
rect 5098 734 14866 856
rect 15034 734 18842 856
<< metal3 >>
rect 0 13472 800 13592
rect 19200 13472 20000 13592
rect 0 12656 800 12776
rect 0 11840 800 11960
rect 0 11024 800 11144
rect 19200 11024 20000 11144
rect 0 10208 800 10328
rect 0 9392 800 9512
rect 0 8576 800 8696
rect 19200 8576 20000 8696
rect 0 7760 800 7880
rect 0 6944 800 7064
rect 0 6128 800 6248
rect 19200 6128 20000 6248
rect 0 5312 800 5432
rect 0 4496 800 4616
rect 0 3680 800 3800
rect 19200 3680 20000 3800
rect 0 2864 800 2984
rect 0 2048 800 2168
rect 0 1232 800 1352
rect 19200 1232 20000 1352
<< obsm3 >>
rect 880 13392 19120 13633
rect 800 12856 19200 13392
rect 880 12576 19200 12856
rect 800 12040 19200 12576
rect 880 11760 19200 12040
rect 800 11224 19200 11760
rect 880 10944 19120 11224
rect 800 10408 19200 10944
rect 880 10128 19200 10408
rect 800 9592 19200 10128
rect 880 9312 19200 9592
rect 800 8776 19200 9312
rect 880 8496 19120 8776
rect 800 7960 19200 8496
rect 880 7680 19200 7960
rect 800 7144 19200 7680
rect 880 6864 19200 7144
rect 800 6328 19200 6864
rect 880 6048 19120 6328
rect 800 5512 19200 6048
rect 880 5232 19200 5512
rect 800 4696 19200 5232
rect 880 4416 19200 4696
rect 800 3880 19200 4416
rect 880 3600 19120 3880
rect 800 3064 19200 3600
rect 880 2784 19200 3064
rect 800 2248 19200 2784
rect 880 1968 19200 2248
rect 800 1432 19200 1968
rect 880 1152 19120 1432
rect 800 1055 19200 1152
<< metal4 >>
rect 4208 1040 4528 13648
rect 8208 1040 8528 13648
rect 12208 1040 12528 13648
rect 16208 1040 16528 13648
<< metal5 >>
rect 1056 12210 18908 12530
rect 1056 8210 18908 8530
rect 1056 4210 18908 4530
<< labels >>
rlabel metal4 s 8208 1040 8528 13648 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 16208 1040 16528 13648 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 8210 18908 8530 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 1040 4528 13648 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12208 1040 12528 13648 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 4210 18908 4530 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 12210 18908 12530 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 1232 800 1352 6 clockp[0]
port 3 nsew signal output
rlabel metal3 s 0 2048 800 2168 6 clockp[1]
port 4 nsew signal output
rlabel metal3 s 0 7760 800 7880 6 dco
port 5 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 div[0]
port 6 nsew signal input
rlabel metal3 s 0 3680 800 3800 6 div[1]
port 7 nsew signal input
rlabel metal3 s 0 4496 800 4616 6 div[2]
port 8 nsew signal input
rlabel metal3 s 0 5312 800 5432 6 div[3]
port 9 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 div[4]
port 10 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 enable
port 11 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 ext_trim[0]
port 12 nsew signal input
rlabel metal2 s 5538 14200 5594 15000 6 ext_trim[10]
port 13 nsew signal input
rlabel metal2 s 7010 14200 7066 15000 6 ext_trim[11]
port 14 nsew signal input
rlabel metal2 s 8482 14200 8538 15000 6 ext_trim[12]
port 15 nsew signal input
rlabel metal2 s 9954 14200 10010 15000 6 ext_trim[13]
port 16 nsew signal input
rlabel metal2 s 11426 14200 11482 15000 6 ext_trim[14]
port 17 nsew signal input
rlabel metal2 s 12898 14200 12954 15000 6 ext_trim[15]
port 18 nsew signal input
rlabel metal2 s 14370 14200 14426 15000 6 ext_trim[16]
port 19 nsew signal input
rlabel metal2 s 15842 14200 15898 15000 6 ext_trim[17]
port 20 nsew signal input
rlabel metal2 s 17314 14200 17370 15000 6 ext_trim[18]
port 21 nsew signal input
rlabel metal2 s 18786 14200 18842 15000 6 ext_trim[19]
port 22 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 ext_trim[1]
port 23 nsew signal input
rlabel metal3 s 19200 13472 20000 13592 6 ext_trim[20]
port 24 nsew signal input
rlabel metal3 s 19200 11024 20000 11144 6 ext_trim[21]
port 25 nsew signal input
rlabel metal3 s 19200 8576 20000 8696 6 ext_trim[22]
port 26 nsew signal input
rlabel metal3 s 19200 6128 20000 6248 6 ext_trim[23]
port 27 nsew signal input
rlabel metal3 s 19200 3680 20000 3800 6 ext_trim[24]
port 28 nsew signal input
rlabel metal3 s 19200 1232 20000 1352 6 ext_trim[25]
port 29 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 ext_trim[2]
port 30 nsew signal input
rlabel metal3 s 0 11024 800 11144 6 ext_trim[3]
port 31 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 ext_trim[4]
port 32 nsew signal input
rlabel metal3 s 0 12656 800 12776 6 ext_trim[5]
port 33 nsew signal input
rlabel metal3 s 0 13472 800 13592 6 ext_trim[6]
port 34 nsew signal input
rlabel metal2 s 1122 14200 1178 15000 6 ext_trim[7]
port 35 nsew signal input
rlabel metal2 s 2594 14200 2650 15000 6 ext_trim[8]
port 36 nsew signal input
rlabel metal2 s 4066 14200 4122 15000 6 ext_trim[9]
port 37 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 osc
port 38 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 resetb
port 39 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 20000 15000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1263518
string GDS_FILE ../gds/digital_pll.gds
string GDS_START 348134
<< end >>

