VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO digital_pll
  CLASS BLOCK ;
  FOREIGN digital_pll ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 75.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 41.040 5.200 42.640 68.240 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 41.050 69.700 42.650 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 5.200 22.640 68.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 61.040 5.200 62.640 68.240 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 21.050 69.700 22.650 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 61.050 69.700 62.650 ;
    END
  END VPWR
  PIN clockp[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 4.000 2.680 ;
    END
  END clockp[0]
  PIN clockp[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 4.000 6.760 ;
    END
  END clockp[1]
  PIN dco
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END dco
  PIN div[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END div[0]
  PIN div[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 4.000 16.280 ;
    END
  END div[1]
  PIN div[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END div[2]
  PIN div[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END div[3]
  PIN div[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END div[4]
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END enable
  PIN ext_trim[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END ext_trim[0]
  PIN ext_trim[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 71.000 20.150 75.000 ;
    END
  END ext_trim[10]
  PIN ext_trim[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 71.000 26.130 75.000 ;
    END
  END ext_trim[11]
  PIN ext_trim[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 71.000 31.650 75.000 ;
    END
  END ext_trim[12]
  PIN ext_trim[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 71.000 37.630 75.000 ;
    END
  END ext_trim[13]
  PIN ext_trim[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 71.000 43.150 75.000 ;
    END
  END ext_trim[14]
  PIN ext_trim[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 71.000 49.130 75.000 ;
    END
  END ext_trim[15]
  PIN ext_trim[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 71.000 54.650 75.000 ;
    END
  END ext_trim[16]
  PIN ext_trim[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 71.000 60.630 75.000 ;
    END
  END ext_trim[17]
  PIN ext_trim[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 71.000 66.150 75.000 ;
    END
  END ext_trim[18]
  PIN ext_trim[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 71.000 72.130 75.000 ;
    END
  END ext_trim[19]
  PIN ext_trim[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END ext_trim[1]
  PIN ext_trim[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 68.040 75.000 68.640 ;
    END
  END ext_trim[20]
  PIN ext_trim[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 55.800 75.000 56.400 ;
    END
  END ext_trim[21]
  PIN ext_trim[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 43.560 75.000 44.160 ;
    END
  END ext_trim[22]
  PIN ext_trim[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 30.640 75.000 31.240 ;
    END
  END ext_trim[23]
  PIN ext_trim[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 18.400 75.000 19.000 ;
    END
  END ext_trim[24]
  PIN ext_trim[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 6.160 75.000 6.760 ;
    END
  END ext_trim[25]
  PIN ext_trim[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END ext_trim[2]
  PIN ext_trim[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END ext_trim[3]
  PIN ext_trim[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END ext_trim[4]
  PIN ext_trim[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END ext_trim[5]
  PIN ext_trim[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END ext_trim[6]
  PIN ext_trim[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 71.000 3.130 75.000 ;
    END
  END ext_trim[7]
  PIN ext_trim[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 71.000 8.650 75.000 ;
    END
  END ext_trim[8]
  PIN ext_trim[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 71.000 14.630 75.000 ;
    END
  END ext_trim[9]
  PIN osc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END osc
  PIN resetb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END resetb
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 69.460 68.085 ;
      LAYER met1 ;
        RECT 4.210 4.120 72.150 71.700 ;
      LAYER met2 ;
        RECT 3.410 70.720 8.090 72.605 ;
        RECT 8.930 70.720 14.070 72.605 ;
        RECT 14.910 70.720 19.590 72.605 ;
        RECT 20.430 70.720 25.570 72.605 ;
        RECT 26.410 70.720 31.090 72.605 ;
        RECT 31.930 70.720 37.070 72.605 ;
        RECT 37.910 70.720 42.590 72.605 ;
        RECT 43.430 70.720 48.570 72.605 ;
        RECT 49.410 70.720 54.090 72.605 ;
        RECT 54.930 70.720 60.070 72.605 ;
        RECT 60.910 70.720 65.590 72.605 ;
        RECT 66.430 70.720 71.570 72.605 ;
        RECT 3.130 4.280 72.120 70.720 ;
        RECT 3.130 2.195 18.210 4.280 ;
        RECT 19.050 2.195 55.470 4.280 ;
        RECT 56.310 2.195 72.120 4.280 ;
      LAYER met3 ;
        RECT 4.400 71.720 71.000 72.585 ;
        RECT 4.000 69.040 71.000 71.720 ;
        RECT 4.000 68.360 70.600 69.040 ;
        RECT 4.400 67.640 70.600 68.360 ;
        RECT 4.400 66.960 71.000 67.640 ;
        RECT 4.000 63.600 71.000 66.960 ;
        RECT 4.400 62.200 71.000 63.600 ;
        RECT 4.000 58.840 71.000 62.200 ;
        RECT 4.400 57.440 71.000 58.840 ;
        RECT 4.000 56.800 71.000 57.440 ;
        RECT 4.000 55.400 70.600 56.800 ;
        RECT 4.000 54.080 71.000 55.400 ;
        RECT 4.400 52.680 71.000 54.080 ;
        RECT 4.000 49.320 71.000 52.680 ;
        RECT 4.400 47.920 71.000 49.320 ;
        RECT 4.000 44.560 71.000 47.920 ;
        RECT 4.400 43.160 70.600 44.560 ;
        RECT 4.000 40.480 71.000 43.160 ;
        RECT 4.400 39.080 71.000 40.480 ;
        RECT 4.000 35.720 71.000 39.080 ;
        RECT 4.400 34.320 71.000 35.720 ;
        RECT 4.000 31.640 71.000 34.320 ;
        RECT 4.000 30.960 70.600 31.640 ;
        RECT 4.400 30.240 70.600 30.960 ;
        RECT 4.400 29.560 71.000 30.240 ;
        RECT 4.000 26.200 71.000 29.560 ;
        RECT 4.400 24.800 71.000 26.200 ;
        RECT 4.000 21.440 71.000 24.800 ;
        RECT 4.400 20.040 71.000 21.440 ;
        RECT 4.000 19.400 71.000 20.040 ;
        RECT 4.000 18.000 70.600 19.400 ;
        RECT 4.000 16.680 71.000 18.000 ;
        RECT 4.400 15.280 71.000 16.680 ;
        RECT 4.000 11.920 71.000 15.280 ;
        RECT 4.400 10.520 71.000 11.920 ;
        RECT 4.000 7.160 71.000 10.520 ;
        RECT 4.400 5.760 70.600 7.160 ;
        RECT 4.000 3.080 71.000 5.760 ;
        RECT 4.400 2.215 71.000 3.080 ;
      LAYER met4 ;
        RECT 31.575 38.935 40.640 67.825 ;
        RECT 43.040 38.935 51.225 67.825 ;
  END
END digital_pll
END LIBRARY

