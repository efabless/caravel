* NGSPICE file created from gpio_control_block.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfbbn_1 abstract view
.subckt sky130_fd_sc_hd__dfbbn_1 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_8 abstract view
.subckt sky130_fd_sc_hd__einvp_8 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for gpio_logic_high abstract view
.subckt gpio_logic_high gpio_logic1 vccd1 vssd1
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

.subckt gpio_control_block gpio_defaults[0] gpio_defaults[10] gpio_defaults[11] gpio_defaults[12]
+ gpio_defaults[1] gpio_defaults[2] gpio_defaults[3] gpio_defaults[4] gpio_defaults[5]
+ gpio_defaults[6] gpio_defaults[7] gpio_defaults[8] gpio_defaults[9] mgmt_gpio_in
+ mgmt_gpio_oeb mgmt_gpio_out one pad_gpio_ana_en pad_gpio_ana_pol pad_gpio_ana_sel
+ pad_gpio_dm[0] pad_gpio_dm[1] pad_gpio_dm[2] pad_gpio_holdover pad_gpio_ib_mode_sel
+ pad_gpio_in pad_gpio_inenb pad_gpio_out pad_gpio_outenb pad_gpio_slow_sel pad_gpio_vtrip_sel
+ resetn resetn_out serial_clock serial_clock_out serial_data_in serial_data_out serial_load
+ serial_load_out user_gpio_in user_gpio_oeb user_gpio_out vccd vccd1 vssd vssd1 zero
X_200_ _200_/A vssd vssd vccd vccd _201_/A sky130_fd_sc_hd__buf_1
X_131_ _131_/A vssd vssd vccd vccd _131_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_114_ _114_/A vssd vssd vccd vccd _114_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_5 user_gpio_oeb vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput31 _205_/X vssd vssd vccd vccd pad_gpio_outenb sky130_fd_sc_hd__buf_2
X_130_ _136_/A _132_/B vssd vssd vccd vccd _131_/A sky130_fd_sc_hd__or2b_1
X_113_ _187_/A _113_/B vssd vssd vccd vccd _114_/A sky130_fd_sc_hd__or2_1
XFILLER_9_45 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_69 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput32 _212_/Q vssd vssd vccd vccd pad_gpio_slow_sel sky130_fd_sc_hd__buf_2
XANTENNA_6 user_gpio_out vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput21 _220_/Q vssd vssd vccd vccd pad_gpio_ana_en sky130_fd_sc_hd__buf_2
X_189_ _189_/A _189_/B vssd vssd vccd vccd _190_/A sky130_fd_sc_hd__or2_1
Xhold10 _226_/D vssd vssd vccd vccd _211_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_112_ _202_/A vssd vssd vccd vccd _187_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_7 serial_data_in vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_80 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput33 _213_/Q vssd vssd vccd vccd pad_gpio_vtrip_sel sky130_fd_sc_hd__buf_2
Xoutput22 _222_/Q vssd vssd vccd vccd pad_gpio_ana_pol sky130_fd_sc_hd__buf_2
XFILLER_18_67 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_188_ _188_/A vssd vssd vccd vccd _188_/X sky130_fd_sc_hd__clkbuf_1
X_111_ _111_/A vssd vssd vccd vccd _111_/X sky130_fd_sc_hd__clkbuf_1
Xhold11 _224_/D vssd vssd vccd vccd _210_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xoutput34 _202_/X vssd vssd vccd vccd resetn_out sky130_fd_sc_hd__buf_2
Xoutput23 _221_/Q vssd vssd vccd vccd pad_gpio_ana_sel sky130_fd_sc_hd__buf_2
X_187_ _187_/A _189_/A vssd vssd vccd vccd _188_/A sky130_fd_sc_hd__or2b_1
XFILLER_4_92 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_57 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_110_ _136_/A _113_/B vssd vssd vccd vccd _111_/A sky130_fd_sc_hd__or2b_1
Xhold12 _230_/D vssd vssd vccd vccd _221_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xoutput24 _217_/Q vssd vssd vccd vccd pad_gpio_dm[0] sky130_fd_sc_hd__buf_2
Xoutput35 _203_/X vssd vssd vccd vccd serial_clock_out sky130_fd_sc_hd__clkbuf_1
X_186_ _186_/A vssd vssd vccd vccd _186_/X sky130_fd_sc_hd__buf_1
X_169_ _169_/A _171_/B vssd vssd vccd vccd _170_/A sky130_fd_sc_hd__or2b_1
Xhold13 _233_/D vssd vssd vccd vccd hold1/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xoutput36 _199_/X vssd vssd vccd vccd serial_data_out sky130_fd_sc_hd__buf_2
Xoutput25 _218_/Q vssd vssd vccd vccd pad_gpio_dm[1] sky130_fd_sc_hd__buf_2
XPHY_0 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_185_ _185_/A vssd vssd vccd vccd _186_/A sky130_fd_sc_hd__buf_1
X_168_ _168_/A vssd vssd vccd vccd _168_/X sky130_fd_sc_hd__buf_1
Xhold14 _231_/D vssd vssd vccd vccd _222_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_1_62 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_73 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_49 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_1 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput37 _204_/X vssd vssd vccd vccd serial_load_out sky130_fd_sc_hd__clkbuf_1
Xoutput26 _219_/Q vssd vssd vccd vccd pad_gpio_dm[2] sky130_fd_sc_hd__buf_2
XFILLER_18_49 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_184_ _184_/A vssd vssd vccd vccd _184_/X sky130_fd_sc_hd__clkbuf_1
Xconst_source vssd vssd vccd vccd one zero sky130_fd_sc_hd__conb_1
X_167_ _173_/A vssd vssd vccd vccd _168_/A sky130_fd_sc_hd__buf_1
Xhold15 _232_/D vssd vssd vccd vccd hold4/A sky130_fd_sc_hd__clkdlybuf4s25_1
X_219_ _129_/X hold8/X _133_/X _131_/X vssd vssd vccd vccd _219_/Q _219_/Q_N sky130_fd_sc_hd__dfbbn_1
XFILLER_1_30 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput27 _211_/Q vssd vssd vccd vccd pad_gpio_holdover sky130_fd_sc_hd__buf_2
XPHY_2 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_29 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_39 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_183_ _183_/A _183_/B vssd vssd vccd vccd _184_/A sky130_fd_sc_hd__or2_1
X_166_ _166_/A vssd vssd vccd vccd _166_/X sky130_fd_sc_hd__clkbuf_1
X_235_ _203_/A _235_/D _202_/A vssd vssd vccd vccd hold8/A sky130_fd_sc_hd__dfrtp_1
XFILLER_1_53 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput28 _215_/Q vssd vssd vccd vccd pad_gpio_ib_mode_sel sky130_fd_sc_hd__buf_2
Xhold16 _228_/D vssd vssd vccd vccd hold2/A sky130_fd_sc_hd__clkdlybuf4s25_1
X_149_ _149_/A vssd vssd vccd vccd _149_/X sky130_fd_sc_hd__buf_1
X_218_ _135_/X hold5/X _139_/X _137_/X vssd vssd vccd vccd _218_/Q _218_/Q_N sky130_fd_sc_hd__dfbbn_1
XPHY_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_29 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_182_ _182_/A vssd vssd vccd vccd _182_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_62 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_148_ _173_/A vssd vssd vccd vccd _149_/A sky130_fd_sc_hd__buf_1
X_165_ _183_/A _165_/B vssd vssd vccd vccd _166_/A sky130_fd_sc_hd__or2_1
X_217_ _141_/X hold6/X _146_/X _144_/X vssd vssd vccd vccd _217_/Q _206_/A0 sky130_fd_sc_hd__dfbbn_1
X_234_ _203_/A _234_/D _202_/A vssd vssd vccd vccd _235_/D sky130_fd_sc_hd__dfrtp_1
Xhold17 _234_/D vssd vssd vccd vccd hold6/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xoutput29 _214_/Q vssd vssd vccd vccd pad_gpio_inenb sky130_fd_sc_hd__buf_2
XPHY_4 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_181_ _187_/A _183_/B vssd vssd vccd vccd _182_/A sky130_fd_sc_hd__or2b_1
X_164_ _164_/A vssd vssd vccd vccd _164_/X sky130_fd_sc_hd__clkbuf_1
X_233_ _203_/A _233_/D _202_/A vssd vssd vccd vccd _234_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_18_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xhold18 _225_/D vssd vssd vccd vccd hold3/A sky130_fd_sc_hd__clkdlybuf4s25_1
X_216_ _149_/X hold3/X _153_/X _151_/X vssd vssd vccd vccd _216_/Q _216_/Q_N sky130_fd_sc_hd__dfbbn_1
X_147_ _147_/A vssd vssd vccd vccd _173_/A sky130_fd_sc_hd__buf_1
XFILLER_16_85 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_5 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_180_ _180_/A vssd vssd vccd vccd _180_/X sky130_fd_sc_hd__buf_1
X_232_ _203_/A _232_/D _202_/A vssd vssd vccd vccd _233_/D sky130_fd_sc_hd__dfrtp_1
X_163_ _169_/A _165_/B vssd vssd vccd vccd _164_/A sky130_fd_sc_hd__or2b_1
Xhold19 _235_/D vssd vssd vccd vccd hold5/A sky130_fd_sc_hd__clkdlybuf4s25_1
X_146_ _146_/A vssd vssd vccd vccd _146_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_88 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_215_ _155_/X hold2/X _160_/X _157_/X vssd vssd vccd vccd _215_/Q _215_/Q_N sky130_fd_sc_hd__dfbbn_1
XPHY_6 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_129_ _129_/A vssd vssd vccd vccd _129_/X sky130_fd_sc_hd__buf_1
XFILLER_16_75 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_231_ _231_/CLK _231_/D _202_/A vssd vssd vccd vccd _232_/D sky130_fd_sc_hd__dfrtp_1
X_162_ _162_/A vssd vssd vccd vccd _162_/X sky130_fd_sc_hd__buf_1
XFILLER_8_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_145_ _152_/A _145_/B vssd vssd vccd vccd _146_/A sky130_fd_sc_hd__or2_1
X_214_ _162_/X hold7/X _166_/X _164_/X vssd vssd vccd vccd _214_/Q _214_/Q_N sky130_fd_sc_hd__dfbbn_1
Xinput1 gpio_defaults[0] vssd vssd vccd vccd _189_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_1_35 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_7 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_128_ _140_/A vssd vssd vccd vccd _129_/A sky130_fd_sc_hd__buf_1
XFILLER_4_46 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_161_ _173_/A vssd vssd vccd vccd _162_/A sky130_fd_sc_hd__buf_1
X_230_ _231_/CLK _230_/D _202_/A vssd vssd vccd vccd _231_/D sky130_fd_sc_hd__dfrtp_1
Xinput2 gpio_defaults[10] vssd vssd vccd vccd _145_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_1_58 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xgpio_in_buf _197_/Y gpio_in_buf/TE vssd vssd vccd vccd user_gpio_in sky130_fd_sc_hd__einvp_8
X_144_ _144_/A vssd vssd vccd vccd _144_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_213_ _168_/X hold1/X _172_/X _170_/X vssd vssd vccd vccd _213_/Q _213_/Q_N sky130_fd_sc_hd__dfbbn_1
XPHY_8 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_127_ _127_/A vssd vssd vccd vccd _127_/X sky130_fd_sc_hd__clkbuf_1
X_212_ _174_/X hold4/X _178_/X _176_/X vssd vssd vccd vccd _212_/Q _212_/Q_N sky130_fd_sc_hd__dfbbn_1
X_143_ _169_/A _145_/B vssd vssd vccd vccd _144_/A sky130_fd_sc_hd__or2b_1
X_160_ _160_/A vssd vssd vccd vccd _160_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_26 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput3 gpio_defaults[11] vssd vssd vccd vccd _138_/B sky130_fd_sc_hd__clkbuf_1
XPHY_9 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_126_ _152_/A _126_/B vssd vssd vccd vccd _127_/A sky130_fd_sc_hd__or2_1
X_109_ _189_/B vssd vssd vccd vccd _136_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_60 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput4 gpio_defaults[12] vssd vssd vccd vccd _132_/B sky130_fd_sc_hd__clkbuf_1
X_211_ _180_/X _211_/D _184_/X _182_/X vssd vssd vccd vccd _211_/Q _211_/Q_N sky130_fd_sc_hd__dfbbn_1
X_125_ _189_/B vssd vssd vccd vccd _152_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_142_ _189_/B vssd vssd vccd vccd _169_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_26 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_70 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_108_ _202_/A vssd vssd vccd vccd _189_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_13_36 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_61 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_210_ _186_/X _210_/D _190_/X _188_/X vssd vssd vccd vccd _210_/Q _210_/Q_N sky130_fd_sc_hd__dfbbn_1
X_141_ _141_/A vssd vssd vccd vccd _141_/X sky130_fd_sc_hd__buf_1
XTAP_50 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_37 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput5 gpio_defaults[1] vssd vssd vccd vccd _152_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_1_39 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0_serial_clock clkbuf_0_serial_clock/X vssd vssd vccd vccd _203_/A sky130_fd_sc_hd__clkbuf_2
X_124_ _124_/A vssd vssd vccd vccd _124_/X sky130_fd_sc_hd__clkbuf_1
X_115__1 serial_load vssd vssd vccd vccd _200_/A sky130_fd_sc_hd__inv_2
XTAP_62 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_51 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_140_ _140_/A vssd vssd vccd vccd _141_/A sky130_fd_sc_hd__buf_1
Xinput6 gpio_defaults[2] vssd vssd vccd vccd _183_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_2_50 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_40 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_37 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_82 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput20 user_gpio_out vssd vssd vccd vccd _208_/A0 sky130_fd_sc_hd__clkbuf_1
X_123_ _136_/A _126_/B vssd vssd vccd vccd _124_/A sky130_fd_sc_hd__or2b_1
XTAP_63 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_115__2 serial_load vssd vssd vccd vccd _185_/A sky130_fd_sc_hd__inv_2
XTAP_52 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 gpio_defaults[3] vssd vssd vccd vccd _165_/B sky130_fd_sc_hd__clkbuf_1
XTAP_41 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_93 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_199_ _199_/A vssd vssd vccd vccd _199_/X sky130_fd_sc_hd__clkbuf_1
Xinput10 gpio_defaults[6] vssd vssd vccd vccd _119_/B sky130_fd_sc_hd__clkbuf_1
X_122_ _122_/A vssd vssd vccd vccd _122_/X sky130_fd_sc_hd__buf_1
X_115__3 serial_load vssd vssd vccd vccd _179_/A sky130_fd_sc_hd__inv_2
XTAP_64 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_53 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_198_ one hold8/A vssd vssd vccd vccd _199_/A sky130_fd_sc_hd__and2_1
XTAP_42 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 gpio_defaults[4] vssd vssd vccd vccd _159_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_2_41 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput11 gpio_defaults[7] vssd vssd vccd vccd _113_/B sky130_fd_sc_hd__clkbuf_1
X_121_ _140_/A vssd vssd vccd vccd _122_/A sky130_fd_sc_hd__buf_1
XFILLER_12_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_65 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_54 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_115__4 serial_load vssd vssd vccd vccd _147_/A sky130_fd_sc_hd__inv_2
Xinput9 gpio_defaults[5] vssd vssd vccd vccd _126_/B sky130_fd_sc_hd__clkbuf_1
XTAP_43 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput12 gpio_defaults[8] vssd vssd vccd vccd _177_/B sky130_fd_sc_hd__clkbuf_1
X_120_ _120_/A vssd vssd vccd vccd _120_/X sky130_fd_sc_hd__clkbuf_1
X_197_ _209_/A vssd vssd vccd vccd _197_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_75 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xhold1 hold1/A vssd vssd vccd vccd hold1/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_115__5 serial_load vssd vssd vccd vccd _116_/A sky130_fd_sc_hd__inv_2
XTAP_55 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_196_ _196_/A vssd vssd vccd vccd _206_/S sky130_fd_sc_hd__clkbuf_1
XTAP_44 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_32 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_179_ _179_/A vssd vssd vccd vccd _180_/A sky130_fd_sc_hd__buf_1
Xinput13 gpio_defaults[9] vssd vssd vccd vccd _171_/B sky130_fd_sc_hd__clkbuf_1
Xhold2 hold2/A vssd vssd vccd vccd hold2/X sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_56 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_45 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xgpio_logic_high gpio_in_buf/TE vccd1 vssd1 gpio_logic_high
X_195_ _219_/Q _218_/Q vssd vssd vccd vccd _196_/A sky130_fd_sc_hd__or2b_1
Xinput14 mgmt_gpio_oeb vssd vssd vccd vccd _207_/S sky130_fd_sc_hd__clkbuf_1
XFILLER_2_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_178_ _178_/A vssd vssd vccd vccd _178_/X sky130_fd_sc_hd__clkbuf_1
Xhold3 hold3/A vssd vssd vccd vccd hold3/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_10_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_57 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_46 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_194_ _194_/A vssd vssd vccd vccd _194_/X sky130_fd_sc_hd__clkbuf_1
X_177_ _183_/A _177_/B vssd vssd vccd vccd _178_/A sky130_fd_sc_hd__or2_1
Xinput15 mgmt_gpio_out vssd vssd vccd vccd _207_/A0 sky130_fd_sc_hd__clkbuf_1
Xhold4 hold4/A vssd vssd vccd vccd hold4/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_8_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_229_ _231_/CLK hold9/A _202_/A vssd vssd vccd vccd _230_/D sky130_fd_sc_hd__dfrtp_1
XTAP_58 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_43 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_47 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_193_ _216_/Q _207_/S vssd vssd vccd vccd _194_/A sky130_fd_sc_hd__and2_1
XPHY_20 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_46 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_176_ _176_/A vssd vssd vccd vccd _176_/X sky130_fd_sc_hd__clkbuf_1
X_159_ _183_/A _159_/B vssd vssd vccd vccd _160_/A sky130_fd_sc_hd__or2_1
X_228_ _231_/CLK _228_/D _202_/A vssd vssd vccd vccd hold9/A sky130_fd_sc_hd__dfrtp_1
Xinput16 pad_gpio_in vssd vssd vccd vccd _209_/A sky130_fd_sc_hd__clkbuf_1
Xhold5 hold5/A vssd vssd vccd vccd hold5/X sky130_fd_sc_hd__clkdlybuf4s25_1
XPHY_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_59 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_48 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_192_ _192_/A vssd vssd vccd vccd _192_/X sky130_fd_sc_hd__clkbuf_1
XPHY_10 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput17 resetn vssd vssd vccd vccd _202_/A sky130_fd_sc_hd__buf_6
X_175_ _187_/A _177_/B vssd vssd vccd vccd _176_/A sky130_fd_sc_hd__or2b_1
XFILLER_3_90 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_36 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_158_ _189_/B vssd vssd vccd vccd _183_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_17_11 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xhold6 hold6/A vssd vssd vccd vccd hold6/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_227_ _231_/CLK hold7/A _202_/A vssd vssd vccd vccd _228_/D sky130_fd_sc_hd__dfrtp_1
Xclkbuf_1_0_0_serial_clock clkbuf_0_serial_clock/X vssd vssd vccd vccd _231_/CLK sky130_fd_sc_hd__clkbuf_2
XTAP_49 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_38 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_33 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_57 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xclkbuf_0_serial_clock serial_clock vssd vssd vccd vccd clkbuf_0_serial_clock/X sky130_fd_sc_hd__clkbuf_16
XPHY_22 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_191_ _214_/Q _216_/Q vssd vssd vccd vccd _192_/A sky130_fd_sc_hd__or2b_1
XPHY_11 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_174_ _174_/A vssd vssd vccd vccd _174_/X sky130_fd_sc_hd__buf_1
X_226_ _231_/CLK _226_/D _202_/A vssd vssd vccd vccd hold7/A sky130_fd_sc_hd__dfrtp_1
X_157_ _157_/A vssd vssd vccd vccd _157_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_80 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput18 serial_data_in vssd vssd vccd vccd _223_/D sky130_fd_sc_hd__clkbuf_1
Xhold7 hold7/A vssd vssd vccd vccd hold7/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_209_ _209_/A _192_/X vssd vssd vccd vccd mgmt_gpio_in sky130_fd_sc_hd__ebufn_8
XFILLER_5_26 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_24 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_12 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_39 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_173_ _173_/A vssd vssd vccd vccd _174_/A sky130_fd_sc_hd__buf_1
XPHY_34 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_23 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_190_ _190_/A vssd vssd vccd vccd _190_/X sky130_fd_sc_hd__clkbuf_1
Xinput19 user_gpio_oeb vssd vssd vccd vccd _205_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_17_57 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_225_ _231_/CLK _225_/D _202_/A vssd vssd vccd vccd _226_/D sky130_fd_sc_hd__dfrtp_1
X_156_ _169_/A _159_/B vssd vssd vccd vccd _157_/A sky130_fd_sc_hd__or2b_1
Xhold8 hold8/A vssd vssd vccd vccd hold8/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_3_70 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_208_ _208_/A0 _207_/X _210_/Q vssd vssd vccd vccd _208_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_93 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_139_ _139_/A vssd vssd vccd vccd _139_/X sky130_fd_sc_hd__clkbuf_1
XPHY_35 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_24 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_13 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_172_ _172_/A vssd vssd vccd vccd _172_/X sky130_fd_sc_hd__clkbuf_1
X_224_ _231_/CLK _224_/D _202_/A vssd vssd vccd vccd _225_/D sky130_fd_sc_hd__dfrtp_1
X_155_ _155_/A vssd vssd vccd vccd _155_/X sky130_fd_sc_hd__buf_1
X_207_ _207_/A0 _206_/X _207_/S vssd vssd vccd vccd _207_/X sky130_fd_sc_hd__mux2_1
X_138_ _152_/A _138_/B vssd vssd vccd vccd _139_/A sky130_fd_sc_hd__or2_1
XFILLER_0_50 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xhold9 hold9/A vssd vssd vccd vccd hold9/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_171_ _183_/A _171_/B vssd vssd vccd vccd _172_/A sky130_fd_sc_hd__or2_1
XPHY_36 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_25 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_14 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_223_ _203_/A _223_/D _202_/A vssd vssd vccd vccd _224_/D sky130_fd_sc_hd__dfrtp_1
X_154_ _173_/A vssd vssd vccd vccd _155_/A sky130_fd_sc_hd__buf_1
X_206_ _206_/A0 _207_/A0 _206_/S vssd vssd vccd vccd _206_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_73 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_137_ _137_/A vssd vssd vccd vccd _137_/X sky130_fd_sc_hd__clkbuf_1
XPHY_37 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_26 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_170_ _170_/A vssd vssd vccd vccd _170_/X sky130_fd_sc_hd__clkbuf_1
X_153_ _153_/A vssd vssd vccd vccd _153_/X sky130_fd_sc_hd__clkbuf_1
X_205_ _205_/A0 _194_/X _210_/Q vssd vssd vccd vccd _205_/X sky130_fd_sc_hd__mux2_1
X_222_ _201_/X _222_/D _114_/X _111_/X vssd vssd vccd vccd _222_/Q _222_/Q_N sky130_fd_sc_hd__dfbbn_1
X_136_ _136_/A _138_/B vssd vssd vccd vccd _137_/A sky130_fd_sc_hd__or2b_1
X_119_ _187_/A _119_/B vssd vssd vccd vccd _120_/A sky130_fd_sc_hd__or2_1
XPHY_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_16 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_0 mgmt_gpio_oeb vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_152_ _152_/A _152_/B vssd vssd vccd vccd _153_/A sky130_fd_sc_hd__or2_1
X_221_ _140_/A _221_/D _120_/X _118_/X vssd vssd vccd vccd _221_/Q _221_/Q_N sky130_fd_sc_hd__dfbbn_1
X_204_ serial_load vssd vssd vccd vccd _204_/X sky130_fd_sc_hd__buf_2
X_118_ _118_/A vssd vssd vccd vccd _118_/X sky130_fd_sc_hd__clkbuf_1
X_135_ _135_/A vssd vssd vccd vccd _135_/X sky130_fd_sc_hd__buf_1
XPHY_28 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_17 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_52 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_1 mgmt_gpio_out vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_86 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_203_ _203_/A vssd vssd vccd vccd _203_/X sky130_fd_sc_hd__buf_2
X_151_ _151_/A vssd vssd vccd vccd _151_/X sky130_fd_sc_hd__clkbuf_1
X_134_ _140_/A vssd vssd vccd vccd _135_/A sky130_fd_sc_hd__buf_1
X_220_ _122_/X hold9/X _127_/X _124_/X vssd vssd vccd vccd _220_/Q _220_/Q_N sky130_fd_sc_hd__dfbbn_1
XFILLER_0_65 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_117_ _136_/A _119_/B vssd vssd vccd vccd _118_/A sky130_fd_sc_hd__or2b_1
XPHY_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_73 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_18 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_2 one vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_150_ _169_/A _152_/B vssd vssd vccd vccd _151_/A sky130_fd_sc_hd__or2b_1
X_133_ _133_/A vssd vssd vccd vccd _133_/X sky130_fd_sc_hd__clkbuf_1
X_202_ _202_/A vssd vssd vccd vccd _202_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_19 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_116_ _116_/A vssd vssd vccd vccd _140_/A sky130_fd_sc_hd__buf_1
XANTENNA_3 one vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_132_ _152_/A _132_/B vssd vssd vccd vccd _133_/A sky130_fd_sc_hd__or2_1
X_201_ _201_/A vssd vssd vccd vccd _201_/X sky130_fd_sc_hd__buf_1
XFILLER_18_85 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput30 _208_/X vssd vssd vccd vccd pad_gpio_out sky130_fd_sc_hd__buf_2
XANTENNA_4 pad_gpio_in vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
.ends

