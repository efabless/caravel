magic
tech sky130A
magscale 1 2
timestamp 1636250566
<< metal1 >>
rect 25840 629233 25846 629285
rect 25898 629273 25904 629285
rect 25898 629245 30798 629273
rect 25898 629233 25904 629245
rect 679888 302563 679894 302575
rect 679474 302535 679894 302563
rect 679888 302523 679894 302535
rect 679946 302523 679952 302575
rect 679696 256387 679702 256399
rect 679474 256359 679702 256387
rect 679696 256347 679702 256359
rect 679754 256347 679760 256399
rect 679792 210285 679798 210297
rect 679474 210257 679798 210285
rect 679792 210245 679798 210257
rect 679850 210245 679856 210297
<< via1 >>
rect 25846 629233 25898 629285
rect 679894 302523 679946 302575
rect 679702 256347 679754 256399
rect 679798 210245 679850 210297
<< metal2 >>
rect 148532 1016270 148588 1016279
rect 148532 1016205 148588 1016214
rect 250484 1016270 250540 1016279
rect 250484 1016205 250540 1016214
rect 353396 1016270 353452 1016279
rect 353396 1016205 353452 1016214
rect 148546 1013032 148574 1016205
rect 250498 1013032 250526 1016205
rect 353410 1013032 353438 1016205
rect 28820 932650 28876 932659
rect 28820 932585 28876 932594
rect 28834 932215 28862 932585
rect 28820 932206 28876 932215
rect 28820 932141 28876 932150
rect 685460 928950 685516 928959
rect 685460 928885 685516 928894
rect 685474 928515 685502 928885
rect 685460 928506 685516 928515
rect 685460 928441 685516 928450
rect 23060 806850 23116 806859
rect 23060 806785 23116 806794
rect 23074 806415 23102 806785
rect 23060 806406 23116 806415
rect 23060 806341 23116 806350
rect 23060 763634 23116 763643
rect 23060 763569 23116 763578
rect 23074 763199 23102 763569
rect 23060 763190 23116 763199
rect 23060 763125 23116 763134
rect 685460 750610 685516 750619
rect 685460 750545 685516 750554
rect 685474 750175 685502 750545
rect 685460 750166 685516 750175
rect 685460 750101 685516 750110
rect 23060 720418 23116 720427
rect 23060 720353 23116 720362
rect 23074 719835 23102 720353
rect 23060 719826 23116 719835
rect 23060 719761 23116 719770
rect 23060 677202 23116 677211
rect 23060 677137 23116 677146
rect 23074 676767 23102 677137
rect 23060 676758 23116 676767
rect 23060 676693 23116 676702
rect 685556 660478 685612 660487
rect 685556 660413 685612 660422
rect 685570 659895 685598 660413
rect 685556 659886 685612 659895
rect 685556 659821 685612 659830
rect 25844 642422 25900 642431
rect 25844 642357 25900 642366
rect 23156 633986 23212 633995
rect 23156 633921 23212 633930
rect 23170 633551 23198 633921
rect 23156 633542 23212 633551
rect 23156 633477 23212 633486
rect 25858 629291 25886 642357
rect 25846 629285 25898 629291
rect 25846 629227 25898 629233
rect 685460 615338 685516 615347
rect 685460 615273 685516 615282
rect 685474 614903 685502 615273
rect 685460 614894 685516 614903
rect 685460 614829 685516 614838
rect 23060 590770 23116 590779
rect 23060 590705 23116 590714
rect 23074 590335 23102 590705
rect 23060 590326 23116 590335
rect 23060 590261 23116 590270
rect 23060 547554 23116 547563
rect 23060 547489 23116 547498
rect 23074 547119 23102 547489
rect 23060 547110 23116 547119
rect 23060 547045 23116 547054
rect 685460 525206 685516 525215
rect 685460 525141 685516 525150
rect 685474 524771 685502 525141
rect 685460 524762 685516 524771
rect 685460 524697 685516 524706
rect 28820 419978 28876 419987
rect 28820 419913 28876 419922
rect 28834 419543 28862 419913
rect 28820 419534 28876 419543
rect 28820 419469 28876 419478
rect 685556 393042 685612 393051
rect 685556 392977 685612 392986
rect 685570 392607 685598 392977
rect 685556 392598 685612 392607
rect 685556 392533 685612 392542
rect 28820 376762 28876 376771
rect 28820 376697 28876 376706
rect 28834 376327 28862 376697
rect 28820 376318 28876 376327
rect 28820 376253 28876 376262
rect 685460 347754 685516 347763
rect 685460 347689 685516 347698
rect 685474 347319 685502 347689
rect 685460 347310 685516 347319
rect 685460 347245 685516 347254
rect 28820 333546 28876 333555
rect 28820 333481 28876 333490
rect 28834 333111 28862 333481
rect 28820 333102 28876 333111
rect 28820 333037 28876 333046
rect 679892 303354 679948 303363
rect 679892 303289 679948 303298
rect 679906 302919 679934 303289
rect 679892 302910 679948 302919
rect 679892 302845 679948 302854
rect 679796 302762 679852 302771
rect 679796 302697 679852 302706
rect 679810 302327 679838 302697
rect 679906 302581 679934 302845
rect 679894 302575 679946 302581
rect 679894 302517 679946 302523
rect 679796 302318 679852 302327
rect 679796 302253 679852 302262
rect 28820 290478 28876 290487
rect 28820 290413 28876 290422
rect 28834 289895 28862 290413
rect 28820 289886 28876 289895
rect 28820 289821 28876 289830
rect 679700 258362 679756 258371
rect 679700 258297 679756 258306
rect 679714 257779 679742 258297
rect 679700 257770 679756 257779
rect 679700 257705 679756 257714
rect 685460 257770 685516 257779
rect 685460 257705 685516 257714
rect 679714 256405 679742 257705
rect 685474 257335 685502 257705
rect 685460 257326 685516 257335
rect 685460 257261 685516 257270
rect 679702 256399 679754 256405
rect 679702 256341 679754 256347
rect 679796 213518 679852 213527
rect 679796 213453 679852 213462
rect 679810 212639 679838 213453
rect 679796 212630 679852 212639
rect 679796 212565 679852 212574
rect 685460 212630 685516 212639
rect 685460 212565 685516 212574
rect 679810 210303 679838 212565
rect 685474 212195 685502 212565
rect 685460 212186 685516 212195
rect 685460 212121 685516 212130
rect 679798 210297 679850 210303
rect 679798 210239 679850 210245
<< via2 >>
rect 148532 1016214 148588 1016270
rect 250484 1016214 250540 1016270
rect 353396 1016214 353452 1016270
rect 28820 932594 28876 932650
rect 28820 932150 28876 932206
rect 685460 928894 685516 928950
rect 685460 928450 685516 928506
rect 23060 806794 23116 806850
rect 23060 806350 23116 806406
rect 23060 763578 23116 763634
rect 23060 763134 23116 763190
rect 685460 750554 685516 750610
rect 685460 750110 685516 750166
rect 23060 720362 23116 720418
rect 23060 719770 23116 719826
rect 23060 677146 23116 677202
rect 23060 676702 23116 676758
rect 685556 660422 685612 660478
rect 685556 659830 685612 659886
rect 25844 642366 25900 642422
rect 23156 633930 23212 633986
rect 23156 633486 23212 633542
rect 685460 615282 685516 615338
rect 685460 614838 685516 614894
rect 23060 590714 23116 590770
rect 23060 590270 23116 590326
rect 23060 547498 23116 547554
rect 23060 547054 23116 547110
rect 685460 525150 685516 525206
rect 685460 524706 685516 524762
rect 28820 419922 28876 419978
rect 28820 419478 28876 419534
rect 685556 392986 685612 393042
rect 685556 392542 685612 392598
rect 28820 376706 28876 376762
rect 28820 376262 28876 376318
rect 685460 347698 685516 347754
rect 685460 347254 685516 347310
rect 28820 333490 28876 333546
rect 28820 333046 28876 333102
rect 679892 303298 679948 303354
rect 679892 302854 679948 302910
rect 679796 302706 679852 302762
rect 679796 302262 679852 302318
rect 28820 290422 28876 290478
rect 28820 289830 28876 289886
rect 679700 258306 679756 258362
rect 679700 257714 679756 257770
rect 685460 257714 685516 257770
rect 685460 257270 685516 257326
rect 679796 213462 679852 213518
rect 679796 212574 679852 212630
rect 685460 212574 685516 212630
rect 685460 212130 685516 212186
<< metal3 >>
rect 148527 1016272 148593 1016275
rect 250479 1016272 250545 1016275
rect 353391 1016272 353457 1016275
rect 98370 1016212 99390 1016272
rect 98370 1013032 98430 1016212
rect 99330 1015946 99390 1016212
rect 148527 1016270 150750 1016272
rect 148527 1016214 148532 1016270
rect 148588 1016214 150750 1016270
rect 148527 1016212 150750 1016214
rect 148527 1016209 148593 1016212
rect 149730 1015946 149790 1016212
rect 150690 1015946 150750 1016212
rect 200610 1016212 201726 1016272
rect 200610 1015946 200670 1016212
rect 201666 1015946 201726 1016212
rect 250479 1016270 253566 1016272
rect 250479 1016214 250484 1016270
rect 250540 1016214 253566 1016270
rect 250479 1016212 253566 1016214
rect 250479 1016209 250545 1016212
rect 252546 1015946 252606 1016212
rect 253506 1015946 253566 1016212
rect 353391 1016270 355518 1016272
rect 353391 1016214 353396 1016270
rect 353452 1016214 355518 1016270
rect 353391 1016212 355518 1016214
rect 353391 1016209 353457 1016212
rect 354498 1015946 354558 1016212
rect 355458 1015946 355518 1016212
rect 421890 1016212 422910 1016272
rect 421890 1013032 421950 1016212
rect 422850 1015946 422910 1016212
rect 550338 1016212 551358 1016272
rect 550338 1015946 550398 1016212
rect 551298 1006534 551358 1016212
rect 28866 932655 28926 932918
rect 28815 932650 28926 932655
rect 28815 932594 28820 932650
rect 28876 932594 28926 932650
rect 28815 932592 28926 932594
rect 28815 932589 28881 932592
rect 28815 932208 28881 932211
rect 28815 932206 28926 932208
rect 28815 932150 28820 932206
rect 28876 932150 28926 932206
rect 28815 932145 28926 932150
rect 28866 931882 28926 932145
rect 685506 928955 685566 929292
rect 685455 928950 685566 928955
rect 685455 928894 685460 928950
rect 685516 928894 685566 928950
rect 685455 928892 685566 928894
rect 685455 928889 685521 928892
rect 685455 928508 685521 928511
rect 685455 928506 685566 928508
rect 685455 928450 685460 928506
rect 685516 928450 685566 928506
rect 685455 928445 685566 928450
rect 685506 928182 685566 928445
rect 23106 806855 23166 807118
rect 23055 806850 23166 806855
rect 23055 806794 23060 806850
rect 23116 806794 23166 806850
rect 23055 806792 23166 806794
rect 23055 806789 23121 806792
rect 23055 806408 23121 806411
rect 23055 806406 23166 806408
rect 23055 806350 23060 806406
rect 23116 806350 23166 806406
rect 23055 806345 23166 806350
rect 23106 806008 23166 806345
rect 23106 763639 23166 763902
rect 23055 763634 23166 763639
rect 23055 763578 23060 763634
rect 23116 763578 23166 763634
rect 23055 763576 23166 763578
rect 23055 763573 23121 763576
rect 23055 763192 23121 763195
rect 23055 763190 23166 763192
rect 23055 763134 23060 763190
rect 23116 763134 23166 763190
rect 23055 763129 23166 763134
rect 23106 762866 23166 763129
rect 685506 750615 685566 750878
rect 685455 750610 685566 750615
rect 685455 750554 685460 750610
rect 685516 750554 685566 750610
rect 685455 750552 685566 750554
rect 685455 750549 685521 750552
rect 685455 750168 685521 750171
rect 685455 750166 685566 750168
rect 685455 750110 685460 750166
rect 685516 750110 685566 750166
rect 685455 750105 685566 750110
rect 685506 749842 685566 750105
rect 23106 720423 23166 720686
rect 23055 720418 23166 720423
rect 23055 720362 23060 720418
rect 23116 720362 23166 720418
rect 23055 720360 23166 720362
rect 23055 720357 23121 720360
rect 23055 719828 23121 719831
rect 23055 719826 23166 719828
rect 23055 719770 23060 719826
rect 23116 719770 23166 719826
rect 23055 719765 23166 719770
rect 23106 719650 23166 719765
rect 23106 677207 23166 677470
rect 23055 677202 23166 677207
rect 23055 677146 23060 677202
rect 23116 677146 23166 677202
rect 23055 677144 23166 677146
rect 23055 677141 23121 677144
rect 23055 676760 23121 676763
rect 23055 676758 23166 676760
rect 23055 676702 23060 676758
rect 23116 676702 23166 676758
rect 23055 676697 23166 676702
rect 23106 676434 23166 676697
rect 685506 660483 685566 660746
rect 685506 660478 685617 660483
rect 685506 660422 685556 660478
rect 685612 660422 685617 660478
rect 685506 660420 685617 660422
rect 685551 660417 685617 660420
rect 685551 659888 685617 659891
rect 685506 659886 685617 659888
rect 685506 659830 685556 659886
rect 685612 659830 685617 659886
rect 685506 659825 685617 659830
rect 685506 659562 685566 659825
rect 25794 642427 25854 642690
rect 25794 642422 25905 642427
rect 25794 642366 25844 642422
rect 25900 642366 25905 642422
rect 25794 642364 25905 642366
rect 25839 642361 25905 642364
rect 23106 633991 23166 634254
rect 23106 633986 23217 633991
rect 23106 633930 23156 633986
rect 23212 633930 23217 633986
rect 23106 633928 23217 633930
rect 23151 633925 23217 633928
rect 23151 633544 23217 633547
rect 23106 633542 23217 633544
rect 23106 633486 23156 633542
rect 23212 633486 23217 633542
rect 23106 633481 23217 633486
rect 23106 633218 23166 633481
rect 685506 615343 685566 615754
rect 685455 615338 685566 615343
rect 685455 615282 685460 615338
rect 685516 615282 685566 615338
rect 685455 615280 685566 615282
rect 685455 615277 685521 615280
rect 685455 614896 685521 614899
rect 685455 614894 685566 614896
rect 685455 614838 685460 614894
rect 685516 614838 685566 614894
rect 685455 614833 685566 614838
rect 685506 614570 685566 614833
rect 23106 590775 23166 591112
rect 23055 590770 23166 590775
rect 23055 590714 23060 590770
rect 23116 590714 23166 590770
rect 23055 590712 23166 590714
rect 23055 590709 23121 590712
rect 23055 590328 23121 590331
rect 23055 590326 23166 590328
rect 23055 590270 23060 590326
rect 23116 590270 23166 590326
rect 23055 590265 23166 590270
rect 23106 590002 23166 590265
rect 23106 547559 23166 547896
rect 23055 547554 23166 547559
rect 23055 547498 23060 547554
rect 23116 547498 23166 547554
rect 23055 547496 23166 547498
rect 23055 547493 23121 547496
rect 23055 547112 23121 547115
rect 23055 547110 23166 547112
rect 23055 547054 23060 547110
rect 23116 547054 23166 547110
rect 23055 547049 23166 547054
rect 23106 546786 23166 547049
rect 685506 525211 685566 525474
rect 685455 525206 685566 525211
rect 685455 525150 685460 525206
rect 685516 525150 685566 525206
rect 685455 525148 685566 525150
rect 685455 525145 685521 525148
rect 685455 524764 685521 524767
rect 685455 524762 685566 524764
rect 685455 524706 685460 524762
rect 685516 524706 685566 524762
rect 685455 524701 685566 524706
rect 685506 524438 685566 524701
rect 28866 419983 28926 420246
rect 28815 419978 28926 419983
rect 28815 419922 28820 419978
rect 28876 419922 28926 419978
rect 28815 419920 28926 419922
rect 28815 419917 28881 419920
rect 28815 419536 28881 419539
rect 28815 419534 28926 419536
rect 28815 419478 28820 419534
rect 28876 419478 28926 419534
rect 28815 419473 28926 419478
rect 28866 419210 28926 419473
rect 685506 393047 685566 393310
rect 685506 393042 685617 393047
rect 685506 392986 685556 393042
rect 685612 392986 685617 393042
rect 685506 392984 685617 392986
rect 685551 392981 685617 392984
rect 685551 392600 685617 392603
rect 685506 392598 685617 392600
rect 685506 392542 685556 392598
rect 685612 392542 685617 392598
rect 685506 392537 685617 392542
rect 685506 392200 685566 392537
rect 28866 376767 28926 377104
rect 28815 376762 28926 376767
rect 28815 376706 28820 376762
rect 28876 376706 28926 376762
rect 28815 376704 28926 376706
rect 28815 376701 28881 376704
rect 28815 376320 28881 376323
rect 28815 376318 28926 376320
rect 28815 376262 28820 376318
rect 28876 376262 28926 376318
rect 28815 376257 28926 376262
rect 28866 375994 28926 376257
rect 685506 347759 685566 348096
rect 685455 347754 685566 347759
rect 685455 347698 685460 347754
rect 685516 347698 685566 347754
rect 685455 347696 685566 347698
rect 685455 347693 685521 347696
rect 685455 347312 685521 347315
rect 685455 347310 685566 347312
rect 685455 347254 685460 347310
rect 685516 347254 685566 347310
rect 685455 347249 685566 347254
rect 685506 346986 685566 347249
rect 28866 333551 28926 333888
rect 28815 333546 28926 333551
rect 28815 333490 28820 333546
rect 28876 333490 28926 333546
rect 28815 333488 28926 333490
rect 28815 333485 28881 333488
rect 28815 333104 28881 333107
rect 28815 333102 28926 333104
rect 28815 333046 28820 333102
rect 28876 333046 28926 333102
rect 28815 333041 28926 333046
rect 28866 332778 28926 333041
rect 679938 303359 679998 303474
rect 679887 303354 679998 303359
rect 679887 303298 679892 303354
rect 679948 303298 679998 303354
rect 679887 303296 679998 303298
rect 679887 303293 679953 303296
rect 679746 302767 679806 303104
rect 679887 302912 679953 302915
rect 679887 302910 679998 302912
rect 679887 302854 679892 302910
rect 679948 302854 679998 302910
rect 679887 302849 679998 302854
rect 679746 302762 679857 302767
rect 679746 302706 679796 302762
rect 679852 302706 679857 302762
rect 679746 302704 679857 302706
rect 679791 302701 679857 302704
rect 679938 302586 679998 302849
rect 679791 302320 679857 302323
rect 679746 302318 679857 302320
rect 679746 302262 679796 302318
rect 679852 302262 679857 302318
rect 679746 302257 679857 302262
rect 679746 301994 679806 302257
rect 28866 290483 28926 290746
rect 28815 290478 28926 290483
rect 28815 290422 28820 290478
rect 28876 290422 28926 290478
rect 28815 290420 28926 290422
rect 28815 290417 28881 290420
rect 28815 289888 28881 289891
rect 28815 289886 28926 289888
rect 28815 289830 28820 289886
rect 28876 289830 28926 289886
rect 28815 289825 28926 289830
rect 28866 289562 28926 289825
rect 679746 258367 679806 258482
rect 679695 258362 679806 258367
rect 679695 258306 679700 258362
rect 679756 258306 679806 258362
rect 679695 258304 679806 258306
rect 679695 258301 679761 258304
rect 685506 257775 685566 258112
rect 679695 257772 679761 257775
rect 679695 257770 679806 257772
rect 679695 257714 679700 257770
rect 679756 257714 679806 257770
rect 679695 257709 679806 257714
rect 685455 257770 685566 257775
rect 685455 257714 685460 257770
rect 685516 257714 685566 257770
rect 685455 257712 685566 257714
rect 685455 257709 685521 257712
rect 679746 257594 679806 257709
rect 685455 257328 685521 257331
rect 685455 257326 685566 257328
rect 685455 257270 685460 257326
rect 685516 257270 685566 257326
rect 685455 257265 685566 257270
rect 685506 257002 685566 257265
rect 679791 213520 679857 213523
rect 679746 213518 679857 213520
rect 679746 213462 679796 213518
rect 679852 213462 679857 213518
rect 679746 213457 679857 213462
rect 679746 213342 679806 213457
rect 685506 212635 685566 212898
rect 679791 212632 679857 212635
rect 679746 212630 679857 212632
rect 679746 212574 679796 212630
rect 679852 212574 679857 212630
rect 679746 212569 679857 212574
rect 685455 212630 685566 212635
rect 685455 212574 685460 212630
rect 685516 212574 685566 212630
rect 685455 212572 685566 212574
rect 685455 212569 685521 212572
rect 679746 212306 679806 212569
rect 685455 212188 685521 212191
rect 685455 212186 685566 212188
rect 685455 212130 685460 212186
rect 685516 212130 685566 212186
rect 685455 212125 685566 212130
rect 685506 211862 685566 212125
<< metal5 >>
rect 78440 1018512 90960 1031002
rect 129840 1018512 142360 1031002
rect 181240 1018512 193760 1031002
rect 232640 1018512 245160 1031002
rect 284240 1018512 296760 1031002
rect 334810 1018624 346978 1030788
rect 386040 1018512 398560 1031002
rect 475040 1018512 487560 1031002
rect 526440 1018512 538960 1031002
rect 577010 1018624 589178 1030788
rect 628240 1018512 640760 1031002
rect 6598 956440 19088 968960
rect 698512 952840 711002 965360
rect 6167 914054 19619 924934
rect 697980 909666 711432 920546
rect 6811 871210 18975 883378
rect 698512 863640 711002 876160
rect 6811 829010 18975 841178
rect 698624 819822 710788 831990
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 698624 505222 710788 517390
rect 6811 484410 18975 496578
rect 697980 461866 711432 472746
rect 6167 442854 19619 453734
rect 698624 417022 710788 429190
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 698512 326640 711002 339160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 6811 111610 18975 123778
rect 698512 101240 711002 113760
rect 6167 70054 19619 80934
rect 80222 6811 92390 18975
rect 136713 7143 144149 18309
rect 187640 6598 200160 19088
rect 243266 6167 254146 19619
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18975
rect 624222 6811 636390 18975
use user_id_textblock  user_id_textblock_0
timestamp 1608324878
transform 1 0 96272 0 1 6890
box -656 1508 33720 10344
use open_source  open_source_0 hexdigits
timestamp 1635801696
transform 1 0 205230 0 1 2174
box 752 5164 29030 16242
use copyright_block  copyright_block_0
timestamp 1636248654
transform 1 0 149582 0 1 16298
box -262 -9464 35048 2764
use caravel_logo  caravel_logo_0
timestamp 1636495793
transform 1 0 270386 0 1 5116
box -2520 0 15000 15560
use gpio_defaults_block_1803  gpio_defaults_block_0
timestamp 1636219436
transform -1 0 709467 0 1 133600
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_1\[0\]
timestamp 1636130125
transform -1 0 710203 0 1 121000
box 750 416 34000 13000
use gpio_defaults_block_0402  gpio_defaults_block_37
timestamp 1636217749
transform -1 0 14347 0 1 215200
box -38 0 6018 2224
use gpio_defaults_block_0402  gpio_defaults_block_36
timestamp 1636217749
transform -1 0 14347 0 1 258400
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_2\[1\]
timestamp 1636130125
transform 1 0 7631 0 1 202600
box 750 416 34000 13000
use gpio_control_block  gpio_control_bidir_2\[0\]
timestamp 1636130125
transform 1 0 7631 0 1 245800
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_2\[16\]
timestamp 1636130125
transform 1 0 7631 0 1 289000
box 750 416 34000 13000
use gpio_defaults_block_1403  gpio_defaults_block_3
timestamp 1636219293
transform -1 0 709467 0 1 269000
box -38 0 6018 2224
use gpio_defaults_block_1403  gpio_defaults_block_2
timestamp 1636219293
transform -1 0 709467 0 1 223800
box -38 0 6018 2224
use gpio_defaults_block_1803  gpio_defaults_block_1
timestamp 1636219436
transform -1 0 709467 0 1 178800
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_1\[1\]
timestamp 1636130125
transform -1 0 710203 0 1 166200
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_1\[1\]
timestamp 1636130125
transform -1 0 710203 0 1 256400
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_1\[0\]
timestamp 1636130125
transform -1 0 710203 0 1 211200
box 750 416 34000 13000
use gpio_defaults_block_0402  gpio_defaults_block_35
timestamp 1636217749
transform -1 0 14347 0 1 301600
box -38 0 6018 2224
use gpio_defaults_block_0402  gpio_defaults_block_34
timestamp 1636217749
transform -1 0 14347 0 1 344800
box -38 0 6018 2224
use gpio_defaults_block_0402  gpio_defaults_block_33
timestamp 1636217749
transform -1 0 14347 0 1 388000
box -38 0 6018 2224
use gpio_defaults_block_0402  gpio_defaults_block_32
timestamp 1636217749
transform -1 0 14347 0 1 431200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[15\]
timestamp 1636130125
transform 1 0 7631 0 1 332200
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_2\[14\]
timestamp 1636130125
transform 1 0 7631 0 1 375400
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_2\[13\]
timestamp 1636130125
transform 1 0 7631 0 1 418600
box 750 416 34000 13000
use gpio_defaults_block_0402  gpio_defaults_block_6
timestamp 1636217749
transform -1 0 709467 0 1 404200
box -38 0 6018 2224
use gpio_defaults_block_0402  gpio_defaults_block_5
timestamp 1636217749
transform -1 0 709467 0 1 359000
box -38 0 6018 2224
use gpio_defaults_block_1403  gpio_defaults_block_4
timestamp 1636219293
transform -1 0 709467 0 1 314000
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[3\]
timestamp 1636130125
transform -1 0 710203 0 1 346400
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_1\[2\]
timestamp 1636130125
transform -1 0 710203 0 1 301400
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_1\[4\]
timestamp 1636130125
transform -1 0 710203 0 1 391600
box 750 416 34000 13000
use gpio_defaults_block_0402  gpio_defaults_block_7
timestamp 1636217749
transform -1 0 709467 0 1 492400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[5\]
timestamp 1636130125
transform -1 0 710203 0 1 479800
box 750 416 34000 13000
use gpio_defaults_block_0402  gpio_defaults_block_31
timestamp 1636217749
transform -1 0 14347 0 1 558800
box -38 0 6018 2224
use gpio_defaults_block_0402  gpio_defaults_block_30
timestamp 1636217749
transform -1 0 14347 0 1 602000
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[10\]
timestamp 1636130125
transform 1 0 7631 0 1 632600
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_2\[11\]
timestamp 1636130125
transform 1 0 7631 0 1 589400
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_2\[12\]
timestamp 1636130125
transform 1 0 7631 0 1 546200
box 750 416 34000 13000
use gpio_defaults_block_0402  gpio_defaults_block_10
timestamp 1636217749
transform -1 0 709467 0 1 626600
box -38 0 6018 2224
use gpio_defaults_block_0402  gpio_defaults_block_9
timestamp 1636217749
transform -1 0 709467 0 1 581400
box -38 0 6018 2224
use gpio_defaults_block_0402  gpio_defaults_block_8
timestamp 1636217749
transform -1 0 709467 0 1 536400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[6\]
timestamp 1636130125
transform -1 0 710203 0 1 523800
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_1\[7\]
timestamp 1636130125
transform -1 0 710203 0 1 568800
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_1\[8\]
timestamp 1636130125
transform -1 0 710203 0 1 614000
box 750 416 34000 13000
use gpio_defaults_block_0402  gpio_defaults_block_29
timestamp 1636217749
transform -1 0 14347 0 1 645200
box -38 0 6018 2224
use gpio_defaults_block_0402  gpio_defaults_block_28
timestamp 1636217749
transform -1 0 14347 0 1 688400
box -38 0 6018 2224
use gpio_defaults_block_0402  gpio_defaults_block_27
timestamp 1636217749
transform -1 0 14347 0 1 731600
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[7\]
timestamp 1636130125
transform 1 0 7631 0 1 762200
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_2\[8\]
timestamp 1636130125
transform 1 0 7631 0 1 719000
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_2\[9\]
timestamp 1636130125
transform 1 0 7631 0 1 675800
box 750 416 34000 13000
use gpio_defaults_block_0402  gpio_defaults_block_13
timestamp 1636217749
transform -1 0 709467 0 1 761800
box -38 0 6018 2224
use gpio_defaults_block_0402  gpio_defaults_block_12
timestamp 1636217749
transform -1 0 709467 0 1 716800
box -38 0 6018 2224
use gpio_defaults_block_0402  gpio_defaults_block_11
timestamp 1636217749
transform -1 0 709467 0 1 671600
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[10\]
timestamp 1636130125
transform -1 0 710203 0 1 704200
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_1\[11\]
timestamp 1636130125
transform -1 0 710203 0 1 749200
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_1\[9\]
timestamp 1636130125
transform -1 0 710203 0 1 659000
box 750 416 34000 13000
use gpio_defaults_block_0402  gpio_defaults_block_26
timestamp 1636217749
transform -1 0 14347 0 1 774800
box -38 0 6018 2224
use gpio_defaults_block_0402  gpio_defaults_block_25
timestamp 1636217749
transform -1 0 14347 0 1 818000
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[6\]
timestamp 1636130125
transform 1 0 7631 0 1 805400
box 750 416 34000 13000
use gpio_defaults_block_0402  gpio_defaults_block_24
timestamp 1636217749
transform 1 0 8367 0 1 943824
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[4\]
timestamp 1636130125
transform 0 1 97200 -1 0 1030077
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_2\[5\]
timestamp 1636130125
transform 1 0 7631 0 1 931224
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_2\[2\]
timestamp 1636130125
transform 0 1 200000 -1 0 1030077
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_2\[3\]
timestamp 1636130125
transform 0 1 148600 -1 0 1030077
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_1\[16\]
timestamp 1636130125
transform 0 1 353400 -1 0 1030077
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_2\[0\]
timestamp 1636130125
transform 0 1 303000 -1 0 1030077
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_2\[1\]
timestamp 1636130125
transform 0 1 251400 -1 0 1030077
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_1\[15\]
timestamp 1636130125
transform 0 1 420800 -1 0 1030077
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_1\[14\]
timestamp 1636130125
transform 0 1 497800 -1 0 1030077
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_1\[13\]
timestamp 1636130125
transform 0 1 549200 -1 0 1030077
box 750 416 34000 13000
use gpio_defaults_block_0402  gpio_defaults_block_14
timestamp 1636217749
transform -1 0 709467 0 1 940200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[12\]
timestamp 1636130125
transform -1 0 710203 0 1 927600
box 750 416 34000 13000
use gpio_defaults_block_0402  gpio_defaults_block_23
timestamp 1636217749
transform 0 1 109800 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block_0402  gpio_defaults_block_22
timestamp 1636217749
transform 0 1 161200 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block_0402  gpio_defaults_block_21
timestamp 1636217749
transform 0 1 212600 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block_0402  gpio_defaults_block_20
timestamp 1636217749
transform 0 1 264000 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block_0402  gpio_defaults_block_19
timestamp 1636217749
transform 0 1 315600 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block_0402  gpio_defaults_block_18
timestamp 1636217749
transform 0 1 366000 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block_0402  gpio_defaults_block_17
timestamp 1636217749
transform 0 1 433400 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block_0402  gpio_defaults_block_16
timestamp 1636217749
transform 0 1 510400 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block_0402  gpio_defaults_block_15
timestamp 1636217749
transform 0 1 561800 -1 0 1029341
box -38 0 6018 2224
use chip_io  padframe
timestamp 1624978002
transform 1 0 0 0 1 0
box -7 0 717607 1037600
<< labels >>
flabel metal5 s 187640 6598 200180 19088 0 FreeSans 16000 0 0 0 clock
port 0 nsew signal input
flabel metal5 s 351040 6598 363580 19088 0 FreeSans 16000 0 0 0 flash_clk
port 1 nsew signal tristate
flabel metal5 s 296240 6598 308780 19088 0 FreeSans 16000 0 0 0 flash_csb
port 2 nsew signal tristate
flabel metal5 s 405840 6598 418380 19088 0 FreeSans 16000 0 0 0 flash_io0
port 3 nsew signal tristate
flabel metal5 s 460640 6598 473180 19088 0 FreeSans 16000 0 0 0 flash_io1
port 4 nsew signal tristate
flabel metal5 s 515440 6598 527980 19088 0 FreeSans 16000 0 0 0 gpio
port 5 nsew signal bidirectional
flabel metal5 s 698512 101240 711002 113780 0 FreeSans 16000 0 0 0 mprj_io[0]
port 6 nsew signal bidirectional
flabel metal5 s 698512 684440 711002 696980 0 FreeSans 16000 0 0 0 mprj_io[10]
port 7 nsew signal bidirectional
flabel metal5 s 698512 729440 711002 741980 0 FreeSans 16000 0 0 0 mprj_io[11]
port 8 nsew signal bidirectional
flabel metal5 s 698512 774440 711002 786980 0 FreeSans 16000 0 0 0 mprj_io[12]
port 9 nsew signal bidirectional
flabel metal5 s 698512 863640 711002 876180 0 FreeSans 16000 0 0 0 mprj_io[13]
port 10 nsew signal bidirectional
flabel metal5 s 698512 952840 711002 965380 0 FreeSans 16000 0 0 0 mprj_io[14]
port 11 nsew signal bidirectional
flabel metal5 s 628220 1018512 640760 1031002 0 FreeSans 16000 0 0 0 mprj_io[15]
port 12 nsew signal bidirectional
flabel metal5 s 526420 1018512 538960 1031002 0 FreeSans 16000 0 0 0 mprj_io[16]
port 13 nsew signal bidirectional
flabel metal5 s 475020 1018512 487560 1031002 0 FreeSans 16000 0 0 0 mprj_io[17]
port 14 nsew signal bidirectional
flabel metal5 s 386020 1018512 398560 1031002 0 FreeSans 16000 0 0 0 mprj_io[18]
port 15 nsew signal bidirectional
flabel metal5 s 284220 1018512 296760 1031002 0 FreeSans 16000 0 0 0 mprj_io[19]
port 16 nsew signal bidirectional
flabel metal5 s 698512 146440 711002 158980 0 FreeSans 16000 0 0 0 mprj_io[1]
port 17 nsew signal bidirectional
flabel metal5 s 232620 1018512 245160 1031002 0 FreeSans 16000 0 0 0 mprj_io[20]
port 18 nsew signal bidirectional
flabel metal5 s 181220 1018512 193760 1031002 0 FreeSans 16000 0 0 0 mprj_io[21]
port 19 nsew signal bidirectional
flabel metal5 s 129820 1018512 142360 1031002 0 FreeSans 16000 0 0 0 mprj_io[22]
port 20 nsew signal bidirectional
flabel metal5 s 78420 1018512 90960 1031002 0 FreeSans 16000 0 0 0 mprj_io[23]
port 21 nsew signal bidirectional
flabel metal5 s 6598 956420 19088 968960 0 FreeSans 16000 0 0 0 mprj_io[24]
port 22 nsew signal bidirectional
flabel metal5 s 6598 786620 19088 799160 0 FreeSans 16000 0 0 0 mprj_io[25]
port 23 nsew signal bidirectional
flabel metal5 s 6598 743420 19088 755960 0 FreeSans 16000 0 0 0 mprj_io[26]
port 24 nsew signal bidirectional
flabel metal5 s 6598 700220 19088 712760 0 FreeSans 16000 0 0 0 mprj_io[27]
port 25 nsew signal bidirectional
flabel metal5 s 6598 657020 19088 669560 0 FreeSans 16000 0 0 0 mprj_io[28]
port 26 nsew signal bidirectional
flabel metal5 s 6598 613820 19088 626360 0 FreeSans 16000 0 0 0 mprj_io[29]
port 27 nsew signal bidirectional
flabel metal5 s 698512 191440 711002 203980 0 FreeSans 16000 0 0 0 mprj_io[2]
port 28 nsew signal bidirectional
flabel metal5 s 6598 570620 19088 583160 0 FreeSans 16000 0 0 0 mprj_io[30]
port 29 nsew signal bidirectional
flabel metal5 s 6598 527420 19088 539960 0 FreeSans 16000 0 0 0 mprj_io[31]
port 30 nsew signal bidirectional
flabel metal5 s 6598 399820 19088 412360 0 FreeSans 16000 0 0 0 mprj_io[32]
port 31 nsew signal bidirectional
flabel metal5 s 6598 356620 19088 369160 0 FreeSans 16000 0 0 0 mprj_io[33]
port 32 nsew signal bidirectional
flabel metal5 s 6598 313420 19088 325960 0 FreeSans 16000 0 0 0 mprj_io[34]
port 33 nsew signal bidirectional
flabel metal5 s 6598 270220 19088 282760 0 FreeSans 16000 0 0 0 mprj_io[35]
port 34 nsew signal bidirectional
flabel metal5 s 6598 227020 19088 239560 0 FreeSans 16000 0 0 0 mprj_io[36]
port 35 nsew signal bidirectional
flabel metal5 s 6598 183820 19088 196360 0 FreeSans 16000 0 0 0 mprj_io[37]
port 36 nsew signal bidirectional
flabel metal5 s 698512 236640 711002 249180 0 FreeSans 16000 0 0 0 mprj_io[3]
port 37 nsew signal bidirectional
flabel metal5 s 698512 281640 711002 294180 0 FreeSans 16000 0 0 0 mprj_io[4]
port 38 nsew signal bidirectional
flabel metal5 s 698512 326640 711002 339180 0 FreeSans 16000 0 0 0 mprj_io[5]
port 39 nsew signal bidirectional
flabel metal5 s 698512 371840 711002 384380 0 FreeSans 16000 0 0 0 mprj_io[6]
port 40 nsew signal bidirectional
flabel metal5 s 698512 549040 711002 561580 0 FreeSans 16000 0 0 0 mprj_io[7]
port 41 nsew signal bidirectional
flabel metal5 s 698512 594240 711002 606780 0 FreeSans 16000 0 0 0 mprj_io[8]
port 42 nsew signal bidirectional
flabel metal5 s 698512 639240 711002 651780 0 FreeSans 16000 0 0 0 mprj_io[9]
port 43 nsew signal bidirectional
flabel metal5 s 136713 7143 144149 18309 0 FreeSans 16000 0 0 0 resetb
port 44 nsew signal input
flabel metal5 s 6167 70054 19619 80934 0 FreeSans 16000 0 0 0 vccd
port 45 nsew signal bidirectional
flabel metal5 s 697980 909666 711432 920546 0 FreeSans 16000 0 0 0 vccd1
port 46 nsew signal bidirectional
flabel metal5 s 6167 914054 19619 924934 0 FreeSans 16000 0 0 0 vccd2
port 47 nsew signal bidirectional
flabel metal5 s 624222 6811 636390 18975 0 FreeSans 16000 0 0 0 vdda
port 48 nsew signal bidirectional
flabel metal5 s 698624 819822 710788 831990 0 FreeSans 16000 0 0 0 vdda1
port 49 nsew signal bidirectional
flabel metal5 s 698624 505222 710788 517390 0 FreeSans 16000 0 0 0 vdda1_2
port 50 nsew signal bidirectional
flabel metal5 s 6811 484410 18975 496578 0 FreeSans 16000 0 0 0 vdda2
port 51 nsew signal bidirectional
flabel metal5 s 6811 111610 18975 123778 0 FreeSans 16000 0 0 0 vddio
port 52 nsew signal bidirectional
flabel metal5 s 6811 871210 18975 883378 0 FreeSans 16000 0 0 0 vddio_2
port 53 nsew signal bidirectional
flabel metal5 s 80222 6811 92390 18975 0 FreeSans 16000 0 0 0 vssa
port 54 nsew signal bidirectional
flabel metal5 s 577010 1018624 589178 1030788 0 FreeSans 16000 0 0 0 vssa1
port 55 nsew signal bidirectional
flabel metal5 s 698624 417022 710788 429190 0 FreeSans 16000 0 0 0 vssa1_2
port 56 nsew signal bidirectional
flabel metal5 s 6811 829010 18975 841178 0 FreeSans 16000 0 0 0 vssa2
port 57 nsew signal bidirectional
flabel metal5 s 243266 6167 254146 19619 0 FreeSans 16000 0 0 0 vssd
port 58 nsew signal bidirectional
flabel metal5 s 697980 461866 711432 472746 0 FreeSans 16000 0 0 0 vssd1
port 59 nsew signal bidirectional
flabel metal5 s 6167 442854 19619 453734 0 FreeSans 16000 0 0 0 vssd2
port 60 nsew signal bidirectional
flabel metal5 s 570422 6811 582590 18975 0 FreeSans 16000 0 0 0 vssio
port 61 nsew signal bidirectional
flabel metal5 s 334810 1018624 346978 1030788 0 FreeSans 16000 0 0 0 vssio_2
port 62 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
