* NGSPICE file created from housekeeping.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufbuf_16 abstract view
.subckt sky130_fd_sc_hd__bufbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtn_1 abstract view
.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_2 abstract view
.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_16 abstract view
.subckt sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

.subckt housekeeping VGND VPWR debug_in debug_mode debug_oeb debug_out irq[0] irq[1]
+ irq[2] mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13]
+ mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18]
+ mask_rev_in[19] mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23]
+ mask_rev_in[24] mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4]
+ mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14]
+ mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19]
+ mgmt_gpio_in[1] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23]
+ mgmt_gpio_in[24] mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28]
+ mgmt_gpio_in[29] mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32]
+ mgmt_gpio_in[33] mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37]
+ mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7]
+ mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16]
+ mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20]
+ mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2]
+ mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[35] mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4]
+ mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18]
+ mgmt_gpio_out[19] mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22]
+ mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27]
+ mgmt_gpio_out[28] mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31]
+ mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36]
+ mgmt_gpio_out[37] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oeb
+ pad_flash_csb pad_flash_csb_oeb pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ieb
+ pad_flash_io0_oeb pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ieb pad_flash_io1_oeb
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1]
+ pll_div[2] pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0]
+ pll_trim[10] pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16]
+ pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22]
+ pll_trim[23] pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5]
+ pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out[0] pwr_ctrl_out[1]
+ pwr_ctrl_out[2] pwr_ctrl_out[3] qspi_enabled reset ser_rx ser_tx serial_clock serial_data_1
+ serial_data_2 serial_load serial_resetn spi_csb spi_enabled spi_sck spi_sdi spi_sdo
+ spi_sdoenb spimemio_flash_clk spimemio_flash_csb spimemio_flash_io0_di spimemio_flash_io0_do
+ spimemio_flash_io0_oeb spimemio_flash_io1_di spimemio_flash_io1_do spimemio_flash_io1_oeb
+ spimemio_flash_io2_di spimemio_flash_io2_do spimemio_flash_io2_oeb spimemio_flash_io3_di
+ spimemio_flash_io3_do spimemio_flash_io3_oeb trap uart_enabled user_clock usr1_vcc_pwrgood
+ usr1_vdd_pwrgood usr2_vcc_pwrgood usr2_vdd_pwrgood wb_ack_o wb_adr_i[0] wb_adr_i[10]
+ wb_adr_i[11] wb_adr_i[12] wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17]
+ wb_adr_i[18] wb_adr_i[19] wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23]
+ wb_adr_i[24] wb_adr_i[25] wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2]
+ wb_adr_i[30] wb_adr_i[31] wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7]
+ wb_adr_i[8] wb_adr_i[9] wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11]
+ wb_dat_i[12] wb_dat_i[13] wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18]
+ wb_dat_i[19] wb_dat_i[1] wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24]
+ wb_dat_i[25] wb_dat_i[26] wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30]
+ wb_dat_i[31] wb_dat_i[3] wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8]
+ wb_dat_i[9] wb_dat_o[0] wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14]
+ wb_dat_o[15] wb_dat_o[16] wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20]
+ wb_dat_o[21] wb_dat_o[22] wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27]
+ wb_dat_o[28] wb_dat_o[29] wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4]
+ wb_dat_o[5] wb_dat_o[6] wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0]
+ wb_sel_i[1] wb_sel_i[2] wb_sel_i[3] wb_stb_i wb_we_i
XFILLER_79_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6914_ _7122_/CLK _6914_/D fanout887/X VGND VGND VPWR VPWR _6914_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6845_ _7223_/CLK _6845_/D _6455_/A VGND VGND VPWR VPWR _6845_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3988_ hold646/X _6411_/A0 _3994_/S VGND VGND VPWR VPWR _6492_/D sky130_fd_sc_hd__mux2_1
X_6776_ _7225_/CLK _6776_/D fanout851/X VGND VGND VPWR VPWR _6776_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5727_ _7038_/Q wire694/X wire660/X wire534/X _5724_/X VGND VGND VPWR VPWR _5734_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_182_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5658_ _5665_/A _7173_/Q _5658_/S VGND VGND VPWR VPWR _7173_/D sky130_fd_sc_hd__mux2_1
XFILLER_190_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4609_ _4987_/A _4992_/B _4586_/B VGND VGND VPWR VPWR _4619_/A sky130_fd_sc_hd__o21ai_1
X_5589_ _5598_/A0 hold574/X _5593_/S VGND VGND VPWR VPWR _7144_/D sky130_fd_sc_hd__mux2_1
XFILLER_124_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold351 _4012_/X VGND VGND VPWR VPWR _6507_/D sky130_fd_sc_hd__bufbuf_16
Xhold362 _6831_/Q VGND VGND VPWR VPWR hold362/X sky130_fd_sc_hd__bufbuf_16
Xhold340 _3505_/A VGND VGND VPWR VPWR _3467_/A sky130_fd_sc_hd__bufbuf_16
Xhold373 _6896_/Q VGND VGND VPWR VPWR hold373/X sky130_fd_sc_hd__bufbuf_16
XFILLER_104_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold384 _7079_/Q VGND VGND VPWR VPWR hold384/X sky130_fd_sc_hd__bufbuf_16
Xhold395 _7027_/Q VGND VGND VPWR VPWR hold395/X sky130_fd_sc_hd__bufbuf_16
XFILLER_132_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout875 fanout890/X VGND VGND VPWR VPWR fanout875/X sky130_fd_sc_hd__buf_8
XFILLER_133_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout853 fanout855/X VGND VGND VPWR VPWR fanout853/X sky130_fd_sc_hd__buf_8
Xfanout864 fanout871/A VGND VGND VPWR VPWR fanout864/X sky130_fd_sc_hd__buf_8
Xfanout886 fanout888/X VGND VGND VPWR VPWR fanout886/X sky130_fd_sc_hd__buf_8
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_213 _3233_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_224 wire599/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_202 wire495/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_246 _5498_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_268 hold214/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_235 _4965_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_257 _3875_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_279 hold475/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4960_ _4949_/A _4949_/C _4959_/X _4907_/A VGND VGND VPWR VPWR _4974_/A sky130_fd_sc_hd__a31o_2
XFILLER_64_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4891_ _4986_/A _4617_/A _5005_/C _4757_/B VGND VGND VPWR VPWR _5174_/C sky130_fd_sc_hd__o22ai_4
XFILLER_60_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3911_ _7157_/Q _7159_/Q _7160_/Q _7158_/Q VGND VGND VPWR VPWR _3918_/B sky130_fd_sc_hd__or4b_2
XFILLER_44_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6630_ _6724_/CLK _6630_/D fanout858/X VGND VGND VPWR VPWR _6630_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3842_ _6487_/Q _6485_/Q _6664_/Q VGND VGND VPWR VPWR _3876_/S sky130_fd_sc_hd__and3_1
X_6561_ _7210_/CLK _6561_/D VGND VGND VPWR VPWR _6561_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_164_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3773_ _7045_/Q _5477_/A _3995_/A _6496_/Q _3772_/X VGND VGND VPWR VPWR _3773_/X
+ sky130_fd_sc_hd__a221o_1
X_5512_ wire739/A hold472/X _5512_/S VGND VGND VPWR VPWR _7076_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6492_ _6815_/CLK _6492_/D fanout855/X VGND VGND VPWR VPWR _6492_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_172_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5443_ _5578_/A0 hold389/X _5449_/S VGND VGND VPWR VPWR _7014_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5374_ hold150/X hold271/X _5377_/S VGND VGND VPWR VPWR _6953_/D sky130_fd_sc_hd__mux2_1
X_7113_ _7143_/CLK _7113_/D fanout880/X VGND VGND VPWR VPWR _7113_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_141_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4325_ _6409_/A0 _6770_/Q _4327_/S VGND VGND VPWR VPWR _6770_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4256_ _4256_/A _5378_/B VGND VGND VPWR VPWR _4261_/S sky130_fd_sc_hd__and2_4
XFILLER_86_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7044_ _7095_/CLK _7044_/D fanout862/X VGND VGND VPWR VPWR _7044_/Q sky130_fd_sc_hd__dfrtp_2
X_3207_ _7120_/Q VGND VGND VPWR VPWR _3207_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4187_ _6651_/Q _5579_/A0 _4189_/S VGND VGND VPWR VPWR _6651_/D sky130_fd_sc_hd__mux2_1
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6828_ _7091_/CLK _6828_/D fanout866/X VGND VGND VPWR VPWR _6828_/Q sky130_fd_sc_hd__dfrtp_2
Xwire506 _7048_/Q VGND VGND VPWR VPWR _3216_/A sky130_fd_sc_hd__buf_8
XFILLER_50_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire528 _6967_/Q VGND VGND VPWR VPWR wire528/X sky130_fd_sc_hd__buf_6
Xwire539 _6905_/Q VGND VGND VPWR VPWR wire539/X sky130_fd_sc_hd__buf_8
XFILLER_109_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6759_ _6806_/CLK _6759_/D fanout848/X VGND VGND VPWR VPWR _6759_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_164_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold170 wire445/X VGND VGND VPWR VPWR _3539_/B sky130_fd_sc_hd__bufbuf_16
Xhold181 _6897_/Q VGND VGND VPWR VPWR hold181/X sky130_fd_sc_hd__bufbuf_16
XFILLER_144_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold192 _3551_/A VGND VGND VPWR VPWR _5234_/A sky130_fd_sc_hd__bufbuf_16
XFILLER_144_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length693 _5684_/X VGND VGND VPWR VPWR wire692/A sky130_fd_sc_hd__buf_6
XFILLER_115_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length682 _5856_/A2 VGND VGND VPWR VPWR _5980_/A2 sky130_fd_sc_hd__buf_6
XFILLER_6_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5090_ _5121_/C _5121_/D _5140_/C _5118_/D VGND VGND VPWR VPWR _5091_/C sky130_fd_sc_hd__or4_1
X_4110_ _6587_/Q wire352/X _4111_/S VGND VGND VPWR VPWR _6587_/D sky130_fd_sc_hd__mux2_1
X_4041_ _5601_/A0 hold344/X hold73/X VGND VGND VPWR VPWR _4041_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5992_ _6014_/A _6036_/B VGND VGND VPWR VPWR _6020_/A sky130_fd_sc_hd__nor2_8
XFILLER_25_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4943_ _4745_/A _4697_/A _4756_/B VGND VGND VPWR VPWR _4943_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_91_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6613_ _6747_/CLK _6613_/D fanout874/X VGND VGND VPWR VPWR _6613_/Q sky130_fd_sc_hd__dfrtp_2
X_4874_ _5003_/A _4874_/B VGND VGND VPWR VPWR _5060_/A sky130_fd_sc_hd__nand2_1
XFILLER_193_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3825_ _6482_/Q _3825_/B VGND VGND VPWR VPWR _3826_/B sky130_fd_sc_hd__nand2_1
X_3756_ _6589_/Q _4112_/A _3739_/X VGND VGND VPWR VPWR _3759_/B sky130_fd_sc_hd__a21o_1
X_6544_ _6650_/CLK _6544_/D fanout858/X VGND VGND VPWR VPWR _6544_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_5_0_csclk clkbuf_3_5_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_5_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
X_6475_ _3957_/A1 _6475_/D _6430_/X VGND VGND VPWR VPWR _6475_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_146_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5426_ wire780/X hold636/X _5429_/S VGND VGND VPWR VPWR _6999_/D sky130_fd_sc_hd__mux2_1
X_3687_ _3687_/A _3687_/B _3687_/C VGND VGND VPWR VPWR _3727_/A sky130_fd_sc_hd__or3_1
Xoutput231 _6516_/Q VGND VGND VPWR VPWR mgmt_gpio_out[26] sky130_fd_sc_hd__buf_8
Xoutput242 _3930_/X VGND VGND VPWR VPWR mgmt_gpio_out[36] sky130_fd_sc_hd__buf_8
Xoutput220 _6669_/Q VGND VGND VPWR VPWR mgmt_gpio_out[16] sky130_fd_sc_hd__buf_8
XFILLER_161_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput253 _3955_/X VGND VGND VPWR VPWR pad_flash_csb sky130_fd_sc_hd__buf_8
X_5357_ _5600_/A0 hold436/X _5359_/S VGND VGND VPWR VPWR _5357_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput286 _6497_/Q VGND VGND VPWR VPWR pll_trim[1] sky130_fd_sc_hd__buf_8
Xoutput275 _6496_/Q VGND VGND VPWR VPWR pll_trim[0] sky130_fd_sc_hd__buf_8
Xoutput264 _6819_/Q VGND VGND VPWR VPWR pll_bypass sky130_fd_sc_hd__buf_8
X_5288_ _5288_/A _5594_/B VGND VGND VPWR VPWR _5296_/S sky130_fd_sc_hd__nand2_8
XFILLER_141_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput297 _6502_/Q VGND VGND VPWR VPWR pll_trim[6] sky130_fd_sc_hd__buf_8
X_4308_ hold713/X _6410_/A0 _4309_/S VGND VGND VPWR VPWR _6756_/D sky130_fd_sc_hd__mux2_1
XFILLER_75_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4239_ _6703_/Q _6706_/Q _6705_/Q _6707_/Q VGND VGND VPWR VPWR _4239_/X sky130_fd_sc_hd__or4_4
X_7027_ _7091_/CLK _7027_/D fanout867/X VGND VGND VPWR VPWR _7027_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_68_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire369 _3426_/X VGND VGND VPWR VPWR wire369/X sky130_fd_sc_hd__buf_6
XFILLER_109_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire358 _5539_/S VGND VGND VPWR VPWR _5536_/S sky130_fd_sc_hd__buf_6
XFILLER_99_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4590_ _4590_/A _4590_/B VGND VGND VPWR VPWR _4591_/B sky130_fd_sc_hd__or2_4
X_3610_ wire899/X _5245_/A _4124_/A _6601_/Q VGND VGND VPWR VPWR _3610_/X sky130_fd_sc_hd__a22o_1
XFILLER_190_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3541_ _6712_/Q _4250_/A _4268_/A _6727_/Q VGND VGND VPWR VPWR _3541_/X sky130_fd_sc_hd__a22o_2
XFILLER_155_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3472_ _3472_/A _3472_/B _3472_/C _3472_/D VGND VGND VPWR VPWR _3548_/A sky130_fd_sc_hd__or4_1
X_6260_ _7197_/Q _6309_/S _6258_/X _6259_/X VGND VGND VPWR VPWR _7197_/D sky130_fd_sc_hd__o22a_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5211_ hold704/X _6410_/A0 _5215_/S VGND VGND VPWR VPWR _6814_/D sky130_fd_sc_hd__mux2_1
X_6191_ wire521/X _5987_/Y _6191_/B1 _6923_/Q _6190_/X VGND VGND VPWR VPWR _6194_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_97_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5142_ _5142_/A _5142_/B _5124_/C VGND VGND VPWR VPWR _5143_/C sky130_fd_sc_hd__or3b_2
XFILLER_111_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5073_ _5079_/B _5073_/B _5073_/C _5073_/D VGND VGND VPWR VPWR _5145_/C sky130_fd_sc_hd__or4_1
X_4024_ hold853/X hold265/X _4024_/S VGND VGND VPWR VPWR _4024_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5975_ _6717_/Q wire702/X _5702_/X _6554_/Q _5974_/X VGND VGND VPWR VPWR _5976_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_52_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4926_ _4988_/A _4398_/Y _4660_/X _4746_/X VGND VGND VPWR VPWR _4926_/X sky130_fd_sc_hd__o22a_2
XFILLER_178_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4857_ _4622_/B _4845_/B _5071_/A _4849_/A VGND VGND VPWR VPWR _4857_/X sky130_fd_sc_hd__a211o_1
XFILLER_176_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3808_ _6485_/Q _3841_/B VGND VGND VPWR VPWR _3898_/A sky130_fd_sc_hd__nand2_4
XFILLER_193_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6527_ _7156_/CLK _6527_/D fanout882/X VGND VGND VPWR VPWR _6527_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4788_ _4758_/B _4652_/B _4758_/C _5136_/A VGND VGND VPWR VPWR _4802_/C sky130_fd_sc_hd__a31o_1
XFILLER_20_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3739_ _6925_/Q wire436/X _3739_/B1 _6981_/Q VGND VGND VPWR VPWR _3739_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6458_ _6458_/CLK _6458_/D _3878_/X VGND VGND VPWR VPWR _6458_/Q sky130_fd_sc_hd__dfstp_4
X_6389_ _4236_/B _6389_/A2 _6389_/B1 _4238_/B VGND VGND VPWR VPWR _6389_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5409_ hold640/X wire773/X _5413_/S VGND VGND VPWR VPWR _6984_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5760_ wire519/X _5678_/X wire670/X _6927_/Q _5759_/X VGND VGND VPWR VPWR _5763_/C
+ sky130_fd_sc_hd__a221o_2
XFILLER_98_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4711_ _4711_/A _4758_/A _4711_/C VGND VGND VPWR VPWR _4936_/A sky130_fd_sc_hd__and3_4
X_5691_ _5864_/B _5704_/B _5701_/C VGND VGND VPWR VPWR _5691_/X sky130_fd_sc_hd__and3_4
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4642_ _4642_/A _5069_/A _4922_/A _4641_/X VGND VGND VPWR VPWR _4642_/X sky130_fd_sc_hd__or4b_1
XFILLER_147_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4573_ _4947_/B _4875_/A VGND VGND VPWR VPWR _5128_/A sky130_fd_sc_hd__nor2_2
Xhold703 _6774_/Q VGND VGND VPWR VPWR hold703/X sky130_fd_sc_hd__bufbuf_16
Xhold714 _6879_/Q VGND VGND VPWR VPWR hold714/X sky130_fd_sc_hd__bufbuf_16
XFILLER_116_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3524_ _5252_/A _3543_/B VGND VGND VPWR VPWR _4292_/A sky130_fd_sc_hd__nor2_8
Xhold725 _7029_/Q VGND VGND VPWR VPWR hold725/X sky130_fd_sc_hd__bufbuf_16
Xhold736 _7099_/Q VGND VGND VPWR VPWR hold736/X sky130_fd_sc_hd__bufbuf_16
X_6312_ _6736_/Q wire642/X wire630/X _6788_/Q VGND VGND VPWR VPWR _6312_/X sky130_fd_sc_hd__a22o_1
XFILLER_170_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6243_ _6604_/Q wire645/X wire636/X _6614_/Q VGND VGND VPWR VPWR _6243_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3455_ _3540_/A _3543_/B VGND VGND VPWR VPWR _4130_/A sky130_fd_sc_hd__nor2_8
Xhold769 _6828_/Q VGND VGND VPWR VPWR hold769/X sky130_fd_sc_hd__bufbuf_16
Xhold758 _6810_/Q VGND VGND VPWR VPWR hold758/X sky130_fd_sc_hd__bufbuf_16
Xhold747 _6773_/Q VGND VGND VPWR VPWR hold747/X sky130_fd_sc_hd__bufbuf_16
XFILLER_143_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6174_ _6954_/Q wire637/X wire635/X _6930_/Q VGND VGND VPWR VPWR _6174_/X sky130_fd_sc_hd__a22o_1
X_3386_ _5225_/A hold87/A VGND VGND VPWR VPWR _3726_/A sky130_fd_sc_hd__nor2_8
XFILLER_111_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5125_ _4748_/A _4719_/X _4907_/C _4974_/A _5114_/B VGND VGND VPWR VPWR _5126_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_69_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5056_ _5056_/A _5056_/B _5157_/A _5056_/D VGND VGND VPWR VPWR _5057_/B sky130_fd_sc_hd__or4_1
XFILLER_85_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4007_ _6421_/B _4025_/A VGND VGND VPWR VPWR _4007_/X sky130_fd_sc_hd__and2b_4
XFILLER_84_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_1_wb_clk_i clkbuf_1_0_1_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_52_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5958_ _6612_/Q wire657/X wire651/X _6761_/Q _5957_/X VGND VGND VPWR VPWR _5959_/D
+ sky130_fd_sc_hd__a221o_1
X_4909_ _5145_/A _4909_/B _5075_/A _4909_/D VGND VGND VPWR VPWR _4910_/C sky130_fd_sc_hd__or4_1
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5889_ _6708_/Q wire680/X wire665/X _6614_/Q VGND VGND VPWR VPWR _5889_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_2_0_csclk clkbuf_2_3_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_5_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_146_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold30 hold70/X VGND VGND VPWR VPWR hold71/A sky130_fd_sc_hd__bufbuf_16
Xhold41 hold41/A VGND VGND VPWR VPWR hold41/X sky130_fd_sc_hd__bufbuf_16
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold52 hold52/A VGND VGND VPWR VPWR hold52/X sky130_fd_sc_hd__bufbuf_16
Xhold74 hold74/A VGND VGND VPWR VPWR hold74/X sky130_fd_sc_hd__bufbuf_16
XFILLER_152_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold63 hold63/A VGND VGND VPWR VPWR hold63/X sky130_fd_sc_hd__bufbuf_16
XFILLER_91_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold96 hold96/A VGND VGND VPWR VPWR hold96/X sky130_fd_sc_hd__bufbuf_16
XFILLER_29_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold85 hold85/A VGND VGND VPWR VPWR hold85/X sky130_fd_sc_hd__bufbuf_16
XFILLER_29_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_5 _6431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6930_ _6930_/CLK _6930_/D fanout887/X VGND VGND VPWR VPWR _6930_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_66_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6861_ _7133_/CLK _6861_/D fanout881/X VGND VGND VPWR VPWR _6861_/Q sky130_fd_sc_hd__dfstp_4
Xclkbuf_leaf_6_csclk _6744_/CLK VGND VGND VPWR VPWR _6727_/CLK sky130_fd_sc_hd__clkbuf_8
X_5812_ _6898_/Q wire674/X _5812_/B1 _7058_/Q VGND VGND VPWR VPWR _5812_/X sky130_fd_sc_hd__a22o_1
XFILLER_35_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6792_ _3957_/A1 _6792_/D _6450_/X VGND VGND VPWR VPWR _6792_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_179_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR clkbuf_1_0_1_mgmt_gpio_in[4]/A
+ sky130_fd_sc_hd__clkbuf_8
X_5743_ _5611_/A _7176_/Q wire381/A VGND VGND VPWR VPWR _5743_/X sky130_fd_sc_hd__a21o_1
XFILLER_62_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5674_ _5864_/B _5705_/B _5703_/B VGND VGND VPWR VPWR _5674_/X sky130_fd_sc_hd__and3_4
XFILLER_30_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4625_ _4995_/A _4749_/C VGND VGND VPWR VPWR _5114_/B sky130_fd_sc_hd__nor2_4
Xhold511 _7211_/Q VGND VGND VPWR VPWR hold511/X sky130_fd_sc_hd__bufbuf_16
XFILLER_190_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4556_ _5118_/A _4840_/A _4805_/A _4556_/D VGND VGND VPWR VPWR _4557_/D sky130_fd_sc_hd__or4_1
Xhold500 _5510_/X VGND VGND VPWR VPWR _7074_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_190_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold533 _6983_/Q VGND VGND VPWR VPWR hold533/X sky130_fd_sc_hd__bufbuf_16
Xhold522 _5545_/X VGND VGND VPWR VPWR _7105_/D sky130_fd_sc_hd__bufbuf_16
X_3507_ _6643_/Q _4172_/A _4286_/A _6742_/Q VGND VGND VPWR VPWR _3507_/X sky130_fd_sc_hd__a22o_2
Xhold544 _5253_/X VGND VGND VPWR VPWR _6845_/D sky130_fd_sc_hd__bufbuf_16
X_4487_ _4655_/A _5050_/A VGND VGND VPWR VPWR _4746_/A sky130_fd_sc_hd__or2_4
Xhold577 _4143_/X VGND VGND VPWR VPWR _6614_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold588 _6837_/Q VGND VGND VPWR VPWR hold588/X sky130_fd_sc_hd__bufbuf_16
Xhold555 _6742_/Q VGND VGND VPWR VPWR hold555/X sky130_fd_sc_hd__bufbuf_16
Xhold566 _6741_/Q VGND VGND VPWR VPWR hold566/X sky130_fd_sc_hd__bufbuf_16
X_6226_ _6876_/Q wire593/X wire591/X wire541/X _6225_/X VGND VGND VPWR VPWR _6231_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_106_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold599 _7088_/Q VGND VGND VPWR VPWR hold599/X sky130_fd_sc_hd__bufbuf_16
X_3438_ _6994_/Q _5414_/A _5540_/A _7106_/Q _3437_/X VGND VGND VPWR VPWR _3452_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3369_ _3369_/A _3672_/A VGND VGND VPWR VPWR _3369_/Y sky130_fd_sc_hd__nor2_8
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6157_ _6356_/A _6157_/B _6157_/C VGND VGND VPWR VPWR _6157_/X sky130_fd_sc_hd__or3_1
X_5108_ _5108_/A _5108_/B _5108_/C VGND VGND VPWR VPWR _5155_/A sky130_fd_sc_hd__or3_4
XFILLER_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6088_ _7135_/Q wire642/X wire630/X wire486/X VGND VGND VPWR VPWR _6088_/X sky130_fd_sc_hd__a22o_1
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5039_ _4832_/C _5050_/C _4689_/Y _4453_/Y VGND VGND VPWR VPWR _5039_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_45_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput120 wb_adr_i[29] VGND VGND VPWR VPWR input120/X sky130_fd_sc_hd__clkbuf_4
XFILLER_163_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput153 wb_dat_i[29] VGND VGND VPWR VPWR _6393_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput131 wb_cyc_i VGND VGND VPWR VPWR input131/X sky130_fd_sc_hd__clkbuf_4
Xinput142 wb_dat_i[19] VGND VGND VPWR VPWR _6387_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_163_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput164 wb_rstn_i VGND VGND VPWR VPWR input164/X sky130_fd_sc_hd__buf_6
XFILLER_63_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4410_ _4707_/B _4478_/C _4410_/C _4410_/D VGND VGND VPWR VPWR _4997_/A sky130_fd_sc_hd__or4_4
X_5390_ _5498_/A0 hold719/X _5395_/S VGND VGND VPWR VPWR _5390_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4341_ _4654_/A _4696_/A _4413_/C _4654_/B VGND VGND VPWR VPWR _4341_/X sky130_fd_sc_hd__a31o_2
XFILLER_160_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7060_ _7152_/CLK _7060_/D fanout886/X VGND VGND VPWR VPWR _7060_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_98_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4272_ hold487/X _5249_/A0 _4273_/S VGND VGND VPWR VPWR _4272_/X sky130_fd_sc_hd__mux2_1
X_3223_ _3223_/A VGND VGND VPWR VPWR _3223_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6011_ _6012_/A _6035_/A _6037_/C VGND VGND VPWR VPWR _6011_/X sky130_fd_sc_hd__and3_1
XFILLER_101_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6913_ _7096_/CLK _6913_/D fanout882/X VGND VGND VPWR VPWR _6913_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_82_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6844_ _6844_/CLK hold28/X _6420_/A VGND VGND VPWR VPWR _6844_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3987_ hold161/X hold152/X _3993_/S VGND VGND VPWR VPWR _3987_/X sky130_fd_sc_hd__mux2_8
X_6775_ _7225_/CLK _6775_/D fanout851/X VGND VGND VPWR VPWR _6775_/Q sky130_fd_sc_hd__dfstp_4
X_5726_ wire492/X _5685_/X wire670/X _6926_/Q VGND VGND VPWR VPWR _5726_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5657_ _5612_/B _5620_/Y _5656_/X _6680_/Q VGND VGND VPWR VPWR _5658_/S sky130_fd_sc_hd__a22o_1
XFILLER_184_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5588_ _5597_/A0 hold377/X _5593_/S VGND VGND VPWR VPWR _5588_/X sky130_fd_sc_hd__mux2_1
X_4608_ _4986_/B _4694_/A _4874_/B VGND VGND VPWR VPWR _4712_/B sky130_fd_sc_hd__o21ai_1
XFILLER_190_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold352 _6905_/Q VGND VGND VPWR VPWR hold352/X sky130_fd_sc_hd__bufbuf_16
Xhold330 _5382_/X VGND VGND VPWR VPWR _6960_/D sky130_fd_sc_hd__bufbuf_16
X_4539_ _4818_/A _4672_/A _4740_/A _4539_/D VGND VGND VPWR VPWR _4542_/B sky130_fd_sc_hd__and4_1
XFILLER_89_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold341 _3301_/Y VGND VGND VPWR VPWR _5450_/A sky130_fd_sc_hd__bufbuf_16
Xhold374 _5310_/X VGND VGND VPWR VPWR _6896_/D sky130_fd_sc_hd__bufbuf_16
Xhold385 _6508_/Q VGND VGND VPWR VPWR hold385/X sky130_fd_sc_hd__bufbuf_16
Xhold363 _6940_/Q VGND VGND VPWR VPWR hold363/X sky130_fd_sc_hd__bufbuf_16
XFILLER_104_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold396 _7134_/Q VGND VGND VPWR VPWR hold396/X sky130_fd_sc_hd__bufbuf_16
XFILLER_104_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout810 _3197_/Y VGND VGND VPWR VPWR _3921_/A sky130_fd_sc_hd__buf_6
X_6209_ _5611_/A _7194_/Q _5664_/X _6208_/X VGND VGND VPWR VPWR _6209_/X sky130_fd_sc_hd__a211o_1
Xfanout876 _6420_/A VGND VGND VPWR VPWR _6421_/A sky130_fd_sc_hd__buf_8
X_7189_ _7190_/CLK _7189_/D fanout869/X VGND VGND VPWR VPWR _7189_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout865 fanout867/X VGND VGND VPWR VPWR fanout865/X sky130_fd_sc_hd__buf_8
Xfanout854 fanout855/X VGND VGND VPWR VPWR fanout854/X sky130_fd_sc_hd__buf_8
Xfanout887 fanout888/X VGND VGND VPWR VPWR fanout887/X sky130_fd_sc_hd__buf_8
XFILLER_133_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_203 wire498/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_225 wire610/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_214 _3581_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_236 _5378_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_247 _5408_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_258 _3875_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_269 _6692_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length820 _3975_/B VGND VGND VPWR VPWR _3953_/A sky130_fd_sc_hd__buf_8
XFILLER_166_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length831 _5252_/C VGND VGND VPWR VPWR _6425_/B sky130_fd_sc_hd__buf_8
XFILLER_181_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_71_csclk _6744_/CLK VGND VGND VPWR VPWR _6724_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_49_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4890_ _4443_/X _4537_/X _4956_/C _5136_/B VGND VGND VPWR VPWR _5075_/A sky130_fd_sc_hd__a31o_1
XFILLER_83_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3910_ _5611_/A _3905_/X _3921_/B _6832_/Q _6677_/Q VGND VGND VPWR VPWR _6679_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_44_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3841_ _6664_/Q _3841_/B VGND VGND VPWR VPWR _3847_/B sky130_fd_sc_hd__nand2_1
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6560_ _7208_/CLK _6560_/D VGND VGND VPWR VPWR _6560_/Q sky130_fd_sc_hd__dfxtp_4
X_3772_ _6773_/Q _4328_/A _4172_/A _6639_/Q VGND VGND VPWR VPWR _3772_/X sky130_fd_sc_hd__a22o_1
XFILLER_192_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5511_ wire746/X hold777/X _5512_/S VGND VGND VPWR VPWR _7075_/D sky130_fd_sc_hd__mux2_1
X_6491_ _6771_/CLK _6491_/D fanout855/X VGND VGND VPWR VPWR _6491_/Q sky130_fd_sc_hd__dfstp_4
X_5442_ wire802/X _7013_/Q _5449_/S VGND VGND VPWR VPWR _7013_/D sky130_fd_sc_hd__mux2_1
X_5373_ wire773/X hold629/X _5377_/S VGND VGND VPWR VPWR _6952_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7112_ _7155_/CLK _7112_/D fanout884/X VGND VGND VPWR VPWR _7112_/Q sky130_fd_sc_hd__dfrtp_2
Xclkbuf_leaf_24_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _6974_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_141_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4324_ wire790/X hold469/X _4327_/S VGND VGND VPWR VPWR _6769_/D sky130_fd_sc_hd__mux2_1
X_7043_ _7132_/CLK _7043_/D fanout868/X VGND VGND VPWR VPWR _7043_/Q sky130_fd_sc_hd__dfrtp_2
X_4255_ _5599_/A0 hold365/X _4255_/S VGND VGND VPWR VPWR _6712_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3206_ _3206_/A VGND VGND VPWR VPWR _3206_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_39_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7122_/CLK sky130_fd_sc_hd__clkbuf_8
X_4186_ hold532/X _5247_/A0 _4189_/S VGND VGND VPWR VPWR _6650_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_1_0_csclk clkbuf_3_1_0_csclk/A VGND VGND VPWR VPWR _6744_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_55_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6827_ _7091_/CLK _6827_/D fanout866/X VGND VGND VPWR VPWR _6827_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire529 _6966_/Q VGND VGND VPWR VPWR wire529/X sky130_fd_sc_hd__buf_6
XFILLER_149_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire518 _7008_/Q VGND VGND VPWR VPWR _3221_/A sky130_fd_sc_hd__buf_8
XFILLER_6_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6758_ _6787_/CLK _6758_/D fanout854/X VGND VGND VPWR VPWR _6758_/Q sky130_fd_sc_hd__dfrtp_2
Xwire507 wire507/A VGND VGND VPWR VPWR wire507/X sky130_fd_sc_hd__buf_6
XFILLER_148_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5709_ _7045_/Q _5687_/X wire664/X _6949_/Q _5708_/X VGND VGND VPWR VPWR _5709_/X
+ sky130_fd_sc_hd__a221o_1
X_6689_ _7220_/CLK _6689_/D _6362_/B VGND VGND VPWR VPWR _6689_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_164_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold160 _6463_/Q VGND VGND VPWR VPWR hold160/X sky130_fd_sc_hd__bufbuf_16
XFILLER_151_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold171 _4097_/Y VGND VGND VPWR VPWR _4102_/S sky130_fd_sc_hd__bufbuf_16
XFILLER_2_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold182 _5311_/X VGND VGND VPWR VPWR _6897_/D sky130_fd_sc_hd__bufbuf_16
Xhold193 _5240_/X VGND VGND VPWR VPWR _6835_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length661 _5794_/B1 VGND VGND VPWR VPWR _5931_/A2 sky130_fd_sc_hd__buf_6
Xmax_length683 _5690_/X VGND VGND VPWR VPWR _5856_/A2 sky130_fd_sc_hd__buf_6
XFILLER_5_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4040_ _5600_/A0 hold478/X hold73/X VGND VGND VPWR VPWR _4040_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5991_ _6037_/A _6035_/C VGND VGND VPWR VPWR _6036_/B sky130_fd_sc_hd__nand2_8
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4942_ _4395_/D _4469_/Y _4689_/Y _4798_/C _4847_/A VGND VGND VPWR VPWR _5180_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_52_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6612_ _6747_/CLK hold84/X fanout874/X VGND VGND VPWR VPWR _6612_/Q sky130_fd_sc_hd__dfrtp_2
X_4873_ _4947_/B _4898_/B _4591_/B VGND VGND VPWR VPWR _5128_/B sky130_fd_sc_hd__a21oi_1
XFILLER_177_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3824_ _3840_/S _3824_/B _6481_/Q VGND VGND VPWR VPWR _3826_/A sky130_fd_sc_hd__or3b_2
XFILLER_118_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3755_ _6594_/Q _4118_/A wire390/X _6718_/Q _3734_/X VGND VGND VPWR VPWR _3759_/A
+ sky130_fd_sc_hd__a221o_4
X_6543_ _6650_/CLK _6543_/D fanout858/X VGND VGND VPWR VPWR _6543_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3686_ _6564_/Q _4082_/A _4142_/A _6615_/Q _3685_/X VGND VGND VPWR VPWR _3687_/C
+ sky130_fd_sc_hd__a221o_4
X_6474_ _3957_/A1 _6474_/D _6429_/X VGND VGND VPWR VPWR _6474_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_145_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput210 _3233_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[7] sky130_fd_sc_hd__buf_8
X_5425_ _5578_/A0 _6998_/Q _5429_/S VGND VGND VPWR VPWR _6998_/D sky130_fd_sc_hd__mux2_1
Xoutput232 _6517_/Q VGND VGND VPWR VPWR mgmt_gpio_out[27] sky130_fd_sc_hd__buf_8
Xoutput243 _3929_/X VGND VGND VPWR VPWR mgmt_gpio_out[37] sky130_fd_sc_hd__buf_8
Xoutput221 _6670_/Q VGND VGND VPWR VPWR mgmt_gpio_out[17] sky130_fd_sc_hd__buf_8
XFILLER_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5356_ hold150/X hold183/X _5359_/S VGND VGND VPWR VPWR _6937_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput254 _3956_/Y VGND VGND VPWR VPWR pad_flash_csb_oeb sky130_fd_sc_hd__buf_8
Xoutput265 _6799_/Q VGND VGND VPWR VPWR pll_dco_ena sky130_fd_sc_hd__buf_8
Xoutput276 _6490_/Q VGND VGND VPWR VPWR pll_trim[10] sky130_fd_sc_hd__buf_8
X_5287_ _5602_/A0 hold277/X _5287_/S VGND VGND VPWR VPWR _6876_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput298 _6503_/Q VGND VGND VPWR VPWR pll_trim[7] sky130_fd_sc_hd__buf_8
Xoutput287 _6815_/Q VGND VGND VPWR VPWR pll_trim[20] sky130_fd_sc_hd__buf_8
X_4307_ hold839/X _6409_/A0 _4309_/S VGND VGND VPWR VPWR _6755_/D sky130_fd_sc_hd__mux2_1
X_4238_ wire817/X _4238_/B VGND VGND VPWR VPWR _6376_/A sky130_fd_sc_hd__and2b_2
XFILLER_102_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7026_ _7091_/CLK _7026_/D fanout867/X VGND VGND VPWR VPWR _7026_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_114_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4169_ _5579_/A0 _6636_/Q _4171_/S VGND VGND VPWR VPWR _6636_/D sky130_fd_sc_hd__mux2_1
XFILLER_15_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3540_ _3540_/A _3733_/B VGND VGND VPWR VPWR _4268_/A sky130_fd_sc_hd__nor2_8
Xwire860 wire860/A VGND VGND VPWR VPWR wire860/X sky130_fd_sc_hd__buf_8
XFILLER_128_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3471_ wire480/X _5540_/A _4310_/A _6762_/Q _3469_/X VGND VGND VPWR VPWR _3472_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_6_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5210_ _6813_/Q wire780/X _5215_/S VGND VGND VPWR VPWR _6813_/D sky130_fd_sc_hd__mux2_1
X_6190_ _7123_/Q _6017_/Y _6030_/Y _7035_/Q VGND VGND VPWR VPWR _6190_/X sky130_fd_sc_hd__a22o_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5141_ _5172_/B _5171_/C _5172_/A VGND VGND VPWR VPWR _5169_/A sky130_fd_sc_hd__o21ba_1
X_5072_ _4748_/A _4689_/Y _4905_/C _4973_/C _4850_/B VGND VGND VPWR VPWR _5175_/A
+ sky130_fd_sc_hd__a2111o_4
XFILLER_96_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4023_ _6529_/Q hold21/X _4023_/S VGND VGND VPWR VPWR _4023_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5974_ _6663_/Q _5974_/A2 wire671/X _5963_/X VGND VGND VPWR VPWR _5974_/X sky130_fd_sc_hd__a22o_1
XFILLER_52_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4925_ _4930_/D _4586_/B _4933_/B _4748_/B VGND VGND VPWR VPWR _5022_/D sky130_fd_sc_hd__a22o_1
XFILLER_100_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4856_ _4586_/B _4845_/B _4850_/X _4855_/X _5116_/B VGND VGND VPWR VPWR _4856_/X
+ sky130_fd_sc_hd__a2111o_4
X_3807_ _6487_/Q _6486_/Q _6485_/Q VGND VGND VPWR VPWR _3843_/B sky130_fd_sc_hd__and3_4
XFILLER_20_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6526_ _6930_/CLK _6526_/D fanout885/X VGND VGND VPWR VPWR _6526_/Q sky130_fd_sc_hd__dfrtp_1
X_4787_ _4808_/A _4787_/B VGND VGND VPWR VPWR _5132_/A sky130_fd_sc_hd__or2_4
XFILLER_146_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3738_ _6563_/Q _4082_/A _4124_/A _6599_/Q VGND VGND VPWR VPWR _3738_/X sky130_fd_sc_hd__a22o_2
XFILLER_118_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3669_ _6729_/Q _4274_/A _4004_/A _6505_/Q VGND VGND VPWR VPWR _3669_/X sky130_fd_sc_hd__a22o_2
X_6457_ _6668_/CLK _6457_/D _6413_/X VGND VGND VPWR VPWR _6457_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6388_ _6387_/X hold79/A _6400_/S VGND VGND VPWR VPWR _7214_/D sky130_fd_sc_hd__mux2_1
XFILLER_121_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5408_ hold533/X _5408_/A1 _5413_/S VGND VGND VPWR VPWR _6983_/D sky130_fd_sc_hd__mux2_1
X_5339_ hold268/X wire758/X _5341_/S VGND VGND VPWR VPWR _6922_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7009_ _7105_/CLK _7009_/D fanout862/X VGND VGND VPWR VPWR _7009_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_28_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4710_ _5023_/A _4671_/A _5031_/B VGND VGND VPWR VPWR _4713_/C sky130_fd_sc_hd__a21oi_1
X_5690_ _7165_/Q _5704_/B _5701_/C VGND VGND VPWR VPWR _5690_/X sky130_fd_sc_hd__and3_4
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4641_ _4965_/A _5005_/C _4639_/X _4640_/X VGND VGND VPWR VPWR _4641_/X sky130_fd_sc_hd__o211a_1
XFILLER_147_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4572_ _4572_/A _4572_/B _5147_/A VGND VGND VPWR VPWR _4875_/A sky130_fd_sc_hd__or3_4
XFILLER_116_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold715 _6911_/Q VGND VGND VPWR VPWR hold715/X sky130_fd_sc_hd__bufbuf_16
Xhold726 _7149_/Q VGND VGND VPWR VPWR hold726/X sky130_fd_sc_hd__bufbuf_16
XFILLER_155_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire690 wire691/X VGND VGND VPWR VPWR wire690/X sky130_fd_sc_hd__buf_6
XFILLER_116_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3523_ _6857_/Q _5261_/A _5468_/A _7041_/Q VGND VGND VPWR VPWR _3523_/X sky130_fd_sc_hd__a22o_1
Xhold704 _6814_/Q VGND VGND VPWR VPWR hold704/X sky130_fd_sc_hd__bufbuf_16
Xhold737 _7083_/Q VGND VGND VPWR VPWR hold737/X sky130_fd_sc_hd__bufbuf_16
X_6311_ _6657_/Q _6311_/B VGND VGND VPWR VPWR _6311_/X sky130_fd_sc_hd__and2_1
XFILLER_131_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6242_ _6576_/Q wire599/X wire631/X _6785_/Q _6241_/X VGND VGND VPWR VPWR _6247_/B
+ sky130_fd_sc_hd__a221o_1
Xhold759 _6763_/Q VGND VGND VPWR VPWR hold759/X sky130_fd_sc_hd__bufbuf_16
Xhold748 _6530_/Q VGND VGND VPWR VPWR hold748/X sky130_fd_sc_hd__bufbuf_16
X_3454_ _3453_/X _6795_/Q _3928_/A VGND VGND VPWR VPWR _6795_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6173_ _7130_/Q wire598/X wire610/X _6173_/B2 _6172_/X VGND VGND VPWR VPWR _6182_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_97_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3385_ _7201_/Q _6830_/Q _6831_/Q VGND VGND VPWR VPWR _3385_/X sky130_fd_sc_hd__mux2_8
XFILLER_97_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5124_ _5142_/A _5124_/B _5124_/C _5124_/D VGND VGND VPWR VPWR _5131_/A sky130_fd_sc_hd__nand4b_2
XFILLER_57_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5055_ _5156_/B _5105_/C VGND VGND VPWR VPWR _5056_/D sky130_fd_sc_hd__or2_1
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4006_ _6408_/A0 _6505_/Q _4006_/S VGND VGND VPWR VPWR _6505_/D sky130_fd_sc_hd__mux2_1
XFILLER_25_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5957_ _6741_/Q wire700/X wire679/X _7224_/Q VGND VGND VPWR VPWR _5957_/X sky130_fd_sc_hd__a22o_1
XFILLER_25_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4908_ _4956_/C _4719_/X _5073_/C _4907_/X _4628_/Y VGND VGND VPWR VPWR _4909_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_33_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5888_ _6599_/Q _5964_/B1 wire653/X _6649_/Q _5887_/X VGND VGND VPWR VPWR _5893_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4839_ _5087_/B _5087_/C _4719_/C VGND VGND VPWR VPWR _4839_/X sky130_fd_sc_hd__o21a_2
XFILLER_193_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6509_ _6931_/CLK _6509_/D fanout885/X VGND VGND VPWR VPWR _6509_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_134_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold20 hold20/A VGND VGND VPWR VPWR hold20/X sky130_fd_sc_hd__bufbuf_16
Xhold31 hold72/X VGND VGND VPWR VPWR hold31/X sky130_fd_sc_hd__bufbuf_16
XFILLER_102_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold64 hold64/A VGND VGND VPWR VPWR hold64/X sky130_fd_sc_hd__bufbuf_16
Xhold53 hold53/A VGND VGND VPWR VPWR hold53/X sky130_fd_sc_hd__bufbuf_16
Xhold42 hold42/A VGND VGND VPWR VPWR hold42/X sky130_fd_sc_hd__bufbuf_16
Xhold75 hold75/A VGND VGND VPWR VPWR hold75/X sky130_fd_sc_hd__bufbuf_16
XFILLER_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold97 hold97/A VGND VGND VPWR VPWR hold97/X sky130_fd_sc_hd__bufbuf_16
Xhold86 hold86/A VGND VGND VPWR VPWR hold86/X sky130_fd_sc_hd__bufbuf_16
XFILLER_90_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_6 _6432_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6860_ _7082_/CLK _6860_/D fanout870/X VGND VGND VPWR VPWR _6860_/Q sky130_fd_sc_hd__dfrtp_2
X_5811_ wire490/X _5685_/X _5699_/X _6930_/Q VGND VGND VPWR VPWR _5811_/X sky130_fd_sc_hd__a22o_1
X_6791_ _3545_/A1 _6791_/D _6449_/X VGND VGND VPWR VPWR _6791_/Q sky130_fd_sc_hd__dfrtn_1
X_5742_ _6854_/Q _5722_/B _5734_/X _5741_/X _3197_/Y VGND VGND VPWR VPWR _5742_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_34_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5673_ _5864_/B _5707_/B _5701_/C VGND VGND VPWR VPWR _5673_/X sky130_fd_sc_hd__and3_4
XFILLER_175_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4624_ _4987_/A _4624_/B VGND VGND VPWR VPWR _4624_/Y sky130_fd_sc_hd__nand2_1
XFILLER_116_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4555_ _4987_/B _4845_/A _4552_/X _4554_/X VGND VGND VPWR VPWR _4556_/D sky130_fd_sc_hd__a211o_1
Xhold501 _7073_/Q VGND VGND VPWR VPWR hold501/X sky130_fd_sc_hd__bufbuf_16
Xhold512 hold512/A VGND VGND VPWR VPWR hold512/X sky130_fd_sc_hd__bufbuf_16
Xhold545 _6626_/Q VGND VGND VPWR VPWR hold545/X sky130_fd_sc_hd__bufbuf_16
Xhold534 _6986_/Q VGND VGND VPWR VPWR hold534/X sky130_fd_sc_hd__bufbuf_16
X_3506_ _3514_/A _5234_/B VGND VGND VPWR VPWR _4286_/A sky130_fd_sc_hd__nor2_8
Xhold523 _7089_/Q VGND VGND VPWR VPWR hold523/X sky130_fd_sc_hd__bufbuf_16
Xhold578 _7120_/Q VGND VGND VPWR VPWR hold578/X sky130_fd_sc_hd__bufbuf_16
X_4486_ _4735_/B _4486_/B _4507_/A VGND VGND VPWR VPWR _5118_/A sky130_fd_sc_hd__and3_4
XFILLER_143_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold556 _4291_/X VGND VGND VPWR VPWR _6742_/D sky130_fd_sc_hd__bufbuf_16
Xhold567 _4290_/X VGND VGND VPWR VPWR _6741_/D sky130_fd_sc_hd__bufbuf_16
X_6225_ _6964_/Q wire624/X wire613/X wire499/X VGND VGND VPWR VPWR _6225_/X sky130_fd_sc_hd__a22o_1
Xhold589 _6634_/Q VGND VGND VPWR VPWR hold589/X sky130_fd_sc_hd__bufbuf_16
X_3437_ _7074_/Q _5504_/A _5227_/A _3423_/X VGND VGND VPWR VPWR _3437_/X sky130_fd_sc_hd__a22o_1
X_6156_ _6156_/A _6156_/B _6156_/C _6156_/D VGND VGND VPWR VPWR _6157_/C sky130_fd_sc_hd__or4_4
X_3368_ _5225_/A _3368_/B VGND VGND VPWR VPWR _3368_/Y sky130_fd_sc_hd__nor2_8
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5107_ _4756_/B _5050_/C _4823_/X VGND VGND VPWR VPWR _5108_/C sky130_fd_sc_hd__o21ai_1
XFILLER_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6087_ _7063_/Q wire648/X wire633/X _6911_/Q VGND VGND VPWR VPWR _6087_/X sky130_fd_sc_hd__a22o_1
XFILLER_57_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3299_ _3505_/A _3668_/A VGND VGND VPWR VPWR _5414_/A sky130_fd_sc_hd__nor2_8
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5038_ _5156_/A _5158_/A VGND VGND VPWR VPWR _5038_/Y sky130_fd_sc_hd__nor2_1
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6989_ _7135_/CLK _6989_/D fanout863/X VGND VGND VPWR VPWR _6989_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_41_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput110 wb_adr_i[1] VGND VGND VPWR VPWR _4735_/A sky130_fd_sc_hd__buf_8
XFILLER_103_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput121 wb_adr_i[2] VGND VGND VPWR VPWR _4395_/D sky130_fd_sc_hd__buf_8
Xinput143 wb_dat_i[1] VGND VGND VPWR VPWR _6381_/B1 sky130_fd_sc_hd__clkbuf_4
Xinput154 wb_dat_i[2] VGND VGND VPWR VPWR _6383_/B1 sky130_fd_sc_hd__clkbuf_4
Xinput132 wb_dat_i[0] VGND VGND VPWR VPWR _6378_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_76_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput165 wb_sel_i[0] VGND VGND VPWR VPWR _6374_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4340_ _4654_/A _4340_/B VGND VGND VPWR VPWR _4408_/A sky130_fd_sc_hd__xor2_4
XFILLER_98_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4271_ hold546/X _5336_/A1 _4273_/S VGND VGND VPWR VPWR _6725_/D sky130_fd_sc_hd__mux2_1
X_3222_ _7000_/Q VGND VGND VPWR VPWR _3222_/Y sky130_fd_sc_hd__clkinv_2
X_6010_ _6036_/A _6010_/B VGND VGND VPWR VPWR _6010_/Y sky130_fd_sc_hd__nor2_8
XFILLER_79_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6912_ _6930_/CLK _6912_/D fanout887/X VGND VGND VPWR VPWR _6912_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_82_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6843_ _6844_/CLK _6843_/D _6420_/A VGND VGND VPWR VPWR _6843_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_90_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3986_ _6491_/Q _6410_/A0 _3994_/S VGND VGND VPWR VPWR _6491_/D sky130_fd_sc_hd__mux2_1
XFILLER_22_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6774_ _7225_/CLK _6774_/D fanout851/X VGND VGND VPWR VPWR _6774_/Q sky130_fd_sc_hd__dfrtp_2
X_5725_ _6894_/Q wire674/X _5812_/B1 _7054_/Q VGND VGND VPWR VPWR _5725_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5656_ _7159_/Q _7160_/Q _5610_/Y VGND VGND VPWR VPWR _5656_/X sky130_fd_sc_hd__or3b_1
XFILLER_163_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4607_ _4917_/A VGND VGND VPWR VPWR _4980_/C sky130_fd_sc_hd__inv_2
X_5587_ wire794/A _7142_/Q _5593_/S VGND VGND VPWR VPWR _7142_/D sky130_fd_sc_hd__mux2_1
Xhold320 _4162_/X VGND VGND VPWR VPWR _6630_/D sky130_fd_sc_hd__bufbuf_16
X_4538_ _4538_/A _4949_/B VGND VGND VPWR VPWR _4970_/B sky130_fd_sc_hd__nand2_1
Xhold353 _5320_/X VGND VGND VPWR VPWR _6905_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_104_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold342 _6782_/Q VGND VGND VPWR VPWR hold342/X sky130_fd_sc_hd__bufbuf_16
Xhold331 _6482_/Q VGND VGND VPWR VPWR hold331/X sky130_fd_sc_hd__bufbuf_16
Xhold386 _4014_/X VGND VGND VPWR VPWR _6508_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_171_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold364 _5359_/X VGND VGND VPWR VPWR _6940_/D sky130_fd_sc_hd__bufbuf_16
Xhold375 _6932_/Q VGND VGND VPWR VPWR hold375/X sky130_fd_sc_hd__bufbuf_16
X_4469_ _4469_/A _4663_/B VGND VGND VPWR VPWR _4469_/Y sky130_fd_sc_hd__nor2_8
XFILLER_117_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout800 hold514/X VGND VGND VPWR VPWR hold515/A sky130_fd_sc_hd__buf_6
XFILLER_77_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout822 _5663_/A VGND VGND VPWR VPWR _5611_/A sky130_fd_sc_hd__buf_8
X_6208_ _6859_/Q _6060_/B _6207_/X _3921_/A VGND VGND VPWR VPWR _6208_/X sky130_fd_sc_hd__o211a_1
Xhold397 _6638_/Q VGND VGND VPWR VPWR hold397/X sky130_fd_sc_hd__bufbuf_16
XFILLER_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7188_ _7220_/CLK _7188_/D fanout853/X VGND VGND VPWR VPWR _7188_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout855 fanout856/X VGND VGND VPWR VPWR fanout855/X sky130_fd_sc_hd__buf_8
Xfanout866 fanout867/X VGND VGND VPWR VPWR fanout866/X sky130_fd_sc_hd__buf_8
Xfanout888 fanout889/X VGND VGND VPWR VPWR fanout888/X sky130_fd_sc_hd__buf_8
Xfanout877 fanout890/X VGND VGND VPWR VPWR _6420_/A sky130_fd_sc_hd__buf_8
X_6139_ _7017_/Q _6139_/A2 _6139_/B1 _7041_/Q _6136_/X VGND VGND VPWR VPWR _6144_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_58_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_204 wire498/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_215 wire551/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_248 _5248_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_226 wire636/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_237 _4986_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_259 wire905/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3840_ _3839_/X _6477_/Q _3840_/S VGND VGND VPWR VPWR _6477_/D sky130_fd_sc_hd__mux2_1
XFILLER_32_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3771_ _6763_/Q _4316_/A _4196_/A _6659_/Q VGND VGND VPWR VPWR _3771_/X sky130_fd_sc_hd__a22o_1
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5510_ wire757/X hold499/X _5512_/S VGND VGND VPWR VPWR _5510_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6490_ _6815_/CLK _6490_/D fanout855/X VGND VGND VPWR VPWR _6490_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5441_ _5441_/A _5576_/B VGND VGND VPWR VPWR _5449_/S sky130_fd_sc_hd__nand2_8
X_5372_ _5597_/A0 hold335/X _5377_/S VGND VGND VPWR VPWR _6951_/D sky130_fd_sc_hd__mux2_1
X_7111_ _7111_/CLK _7111_/D fanout880/X VGND VGND VPWR VPWR _7111_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_114_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4323_ _5234_/C hold741/X _4327_/S VGND VGND VPWR VPWR _6768_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7042_ _7042_/CLK _7042_/D fanout865/X VGND VGND VPWR VPWR _7042_/Q sky130_fd_sc_hd__dfrtp_2
X_4254_ hold83/X hold230/X _4255_/S VGND VGND VPWR VPWR _4254_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4185_ hold586/X wire799/A _4189_/S VGND VGND VPWR VPWR _6649_/D sky130_fd_sc_hd__mux2_1
X_3205_ _7136_/Q VGND VGND VPWR VPWR _3205_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6826_ _7091_/CLK _6826_/D fanout866/X VGND VGND VPWR VPWR _6826_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6757_ _6824_/CLK _6757_/D fanout848/X VGND VGND VPWR VPWR _6757_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_183_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5708_ wire511/X _5688_/X wire651/A _7021_/Q _5670_/X VGND VGND VPWR VPWR _5708_/X
+ sky130_fd_sc_hd__a221o_1
X_3969_ _3969_/A _3969_/B VGND VGND VPWR VPWR _3969_/X sky130_fd_sc_hd__and2_1
Xwire519 _7007_/Q VGND VGND VPWR VPWR wire519/X sky130_fd_sc_hd__buf_6
XFILLER_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire508 _7040_/Q VGND VGND VPWR VPWR _3217_/A sky130_fd_sc_hd__buf_8
XFILLER_50_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6688_ _6992_/CLK _6688_/D fanout868/X VGND VGND VPWR VPWR _6688_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_191_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5639_ _7167_/Q _7166_/Q _6679_/Q VGND VGND VPWR VPWR _5648_/B sky130_fd_sc_hd__and3_2
Xhold150 hold150/A VGND VGND VPWR VPWR hold150/X sky130_fd_sc_hd__bufbuf_16
Xhold161 hold161/A VGND VGND VPWR VPWR hold161/X sky130_fd_sc_hd__bufbuf_16
Xhold183 _6937_/Q VGND VGND VPWR VPWR hold183/X sky130_fd_sc_hd__bufbuf_16
XFILLER_132_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold172 _4101_/X VGND VGND VPWR VPWR _6579_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_104_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold194 _6622_/Q VGND VGND VPWR VPWR hold194/X sky130_fd_sc_hd__bufbuf_16
XFILLER_120_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length695 _5683_/X VGND VGND VPWR VPWR _5803_/B1 sky130_fd_sc_hd__buf_6
XFILLER_5_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5990_ _7167_/Q _7166_/Q VGND VGND VPWR VPWR _6035_/C sky130_fd_sc_hd__nor2_8
XFILLER_52_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4941_ _5163_/A _4941_/B _4941_/C _4941_/D VGND VGND VPWR VPWR _4946_/A sky130_fd_sc_hd__or4_1
XFILLER_17_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4872_ _4953_/A _4899_/B VGND VGND VPWR VPWR _5099_/C sky130_fd_sc_hd__nor2_2
X_6611_ _6747_/CLK _6611_/D fanout874/X VGND VGND VPWR VPWR _6611_/Q sky130_fd_sc_hd__dfstp_4
X_3823_ _3845_/A _3828_/S VGND VGND VPWR VPWR _3824_/B sky130_fd_sc_hd__nor2_1
XFILLER_33_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3754_ _3754_/A _3754_/B _3754_/C _3754_/D VGND VGND VPWR VPWR _3794_/A sky130_fd_sc_hd__or4_4
X_6542_ _6591_/CLK _6542_/D fanout873/X VGND VGND VPWR VPWR _6542_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_173_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3685_ _6918_/Q _5333_/A _4112_/A _6590_/Q VGND VGND VPWR VPWR _3685_/X sky130_fd_sc_hd__a22o_1
X_6473_ _3957_/A1 _6473_/D _6428_/X VGND VGND VPWR VPWR _6473_/Q sky130_fd_sc_hd__dfrtp_2
Xoutput200 _3208_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[32] sky130_fd_sc_hd__buf_8
XFILLER_161_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5424_ _5532_/A0 _6997_/Q _5429_/S VGND VGND VPWR VPWR _6997_/D sky130_fd_sc_hd__mux2_1
Xoutput233 _6518_/Q VGND VGND VPWR VPWR mgmt_gpio_out[28] sky130_fd_sc_hd__buf_8
Xoutput222 _6671_/Q VGND VGND VPWR VPWR mgmt_gpio_out[18] sky130_fd_sc_hd__buf_8
XFILLER_160_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput211 _3232_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[8] sky130_fd_sc_hd__buf_8
Xoutput244 _6684_/Q VGND VGND VPWR VPWR mgmt_gpio_out[3] sky130_fd_sc_hd__buf_8
X_5355_ _5598_/A0 hold637/X _5359_/S VGND VGND VPWR VPWR _6936_/D sky130_fd_sc_hd__mux2_1
Xoutput277 _6491_/Q VGND VGND VPWR VPWR pll_trim[11] sky130_fd_sc_hd__buf_8
Xoutput266 _6800_/Q VGND VGND VPWR VPWR pll_div[0] sky130_fd_sc_hd__buf_8
Xoutput255 _3963_/X VGND VGND VPWR VPWR pad_flash_io0_do sky130_fd_sc_hd__buf_8
X_5286_ _5601_/A0 hold202/X _5287_/S VGND VGND VPWR VPWR _6875_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput299 _6488_/Q VGND VGND VPWR VPWR pll_trim[8] sky130_fd_sc_hd__buf_8
Xoutput288 _6816_/Q VGND VGND VPWR VPWR pll_trim[21] sky130_fd_sc_hd__buf_8
X_4306_ hold711/X _6408_/A0 _4309_/S VGND VGND VPWR VPWR _6754_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4237_ _6700_/Q _6704_/D _6701_/Q _6702_/Q VGND VGND VPWR VPWR _4237_/X sky130_fd_sc_hd__or4_2
X_7025_ _7105_/CLK _7025_/D fanout862/X VGND VGND VPWR VPWR _7025_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_114_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4168_ _5247_/A0 hold497/X _4171_/S VGND VGND VPWR VPWR _6635_/D sky130_fd_sc_hd__mux2_1
X_4099_ _5247_/A0 hold525/X _4102_/S VGND VGND VPWR VPWR _6577_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6809_ _6810_/CLK _6809_/D fanout853/X VGND VGND VPWR VPWR _6809_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_51_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_70_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7119_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_164_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_23_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7143_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_159_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_38_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7147_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_127_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire894 wire894/A VGND VGND VPWR VPWR _3972_/B sky130_fd_sc_hd__buf_6
XFILLER_170_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3470_ _3505_/A _3534_/A VGND VGND VPWR VPWR _4310_/A sky130_fd_sc_hd__nor2_8
XFILLER_170_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5140_ _5140_/A _5140_/B _5140_/C _5139_/X VGND VGND VPWR VPWR _5171_/C sky130_fd_sc_hd__or4b_4
XFILLER_142_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5071_ _5071_/A _5071_/B _5071_/C _5071_/D VGND VGND VPWR VPWR _5126_/A sky130_fd_sc_hd__or4_4
XFILLER_96_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4022_ hold494/X _4021_/X _4024_/S VGND VGND VPWR VPWR _4022_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5973_ _6638_/Q _5973_/A2 wire692/X _6727_/Q _5972_/X VGND VGND VPWR VPWR _5976_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_65_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4924_ _4756_/B _4660_/X _4624_/B _4930_/D VGND VGND VPWR VPWR _5098_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_80_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4855_ _4539_/D _4845_/B _4853_/X _4854_/X VGND VGND VPWR VPWR _4855_/X sky130_fd_sc_hd__a211o_1
XFILLER_138_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4786_ _4772_/A _4399_/Y _4453_/Y _4689_/Y VGND VGND VPWR VPWR _4798_/C sky130_fd_sc_hd__a22o_1
X_3806_ _6487_/Q _6486_/Q VGND VGND VPWR VPWR _3841_/B sky130_fd_sc_hd__and2_2
X_6525_ _6930_/CLK _6525_/D fanout885/X VGND VGND VPWR VPWR _6525_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3737_ _6877_/Q wire406/X _4055_/A _6540_/Q VGND VGND VPWR VPWR _3737_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3668_ _3668_/A _5234_/A VGND VGND VPWR VPWR _4004_/A sky130_fd_sc_hd__nor2_2
X_6456_ _6668_/CLK _6456_/D _6412_/X VGND VGND VPWR VPWR _6456_/Q sky130_fd_sc_hd__dfrtn_1
X_6387_ _4236_/B _6387_/A2 _6387_/B1 _4238_/B _6386_/X VGND VGND VPWR VPWR _6387_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5407_ _6982_/Q hold38/A _5413_/S VGND VGND VPWR VPWR hold18/A sky130_fd_sc_hd__mux2_1
XFILLER_88_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3599_ _7072_/Q _5504_/A _4166_/A _6637_/Q _3563_/X VGND VGND VPWR VPWR _3605_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_121_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5338_ hold343/X hold150/X _5341_/S VGND VGND VPWR VPWR _6921_/D sky130_fd_sc_hd__mux2_1
XFILLER_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5269_ hold380/X wire742/X _5269_/S VGND VGND VPWR VPWR _5269_/X sky130_fd_sc_hd__mux2_1
X_7008_ _7107_/CLK _7008_/D fanout865/X VGND VGND VPWR VPWR _7008_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_56_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4640_ _4603_/B _5005_/C _5135_/A VGND VGND VPWR VPWR _4640_/X sky130_fd_sc_hd__o21ba_1
XFILLER_175_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4571_ _4572_/B _5147_/A VGND VGND VPWR VPWR _4571_/Y sky130_fd_sc_hd__nor2_8
XFILLER_128_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6310_ _6622_/Q wire623/X wire612/X _6652_/Q VGND VGND VPWR VPWR _6310_/X sky130_fd_sc_hd__a22o_1
Xwire680 _5691_/X VGND VGND VPWR VPWR wire680/X sky130_fd_sc_hd__buf_8
Xwire691 _5685_/X VGND VGND VPWR VPWR wire691/X sky130_fd_sc_hd__buf_8
XFILLER_116_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3522_ _3522_/A _3522_/B _3522_/C _3522_/D VGND VGND VPWR VPWR _3547_/B sky130_fd_sc_hd__or4_1
XFILLER_7_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold705 _6801_/Q VGND VGND VPWR VPWR hold705/X sky130_fd_sc_hd__bufbuf_16
Xhold727 _7002_/Q VGND VGND VPWR VPWR hold727/X sky130_fd_sc_hd__bufbuf_16
Xhold716 _7093_/Q VGND VGND VPWR VPWR hold716/X sky130_fd_sc_hd__bufbuf_16
Xhold749 _6514_/Q VGND VGND VPWR VPWR hold749/X sky130_fd_sc_hd__bufbuf_16
XFILLER_171_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6241_ _6634_/Q wire712/X _6311_/B _6654_/Q VGND VGND VPWR VPWR _6241_/X sky130_fd_sc_hd__a22o_4
Xhold738 _6682_/Q VGND VGND VPWR VPWR hold738/X sky130_fd_sc_hd__bufbuf_16
X_3453_ wire351/X _6794_/Q _3857_/C VGND VGND VPWR VPWR _3453_/X sky130_fd_sc_hd__mux2_1
X_6172_ _6890_/Q wire602/X wire581/X _7146_/Q _6171_/X VGND VGND VPWR VPWR _6172_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5123_ _5129_/B _5123_/B _5123_/C _5123_/D VGND VGND VPWR VPWR _5124_/D sky130_fd_sc_hd__and4b_4
XFILLER_130_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3384_ _5234_/A _3520_/B VGND VGND VPWR VPWR _3384_/Y sky130_fd_sc_hd__nor2_4
XFILLER_85_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5054_ _4505_/X _4812_/C _5144_/B _4812_/X _4836_/X VGND VGND VPWR VPWR _5105_/C
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_97_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4005_ _5234_/C _6504_/Q _4006_/S VGND VGND VPWR VPWR _6504_/D sky130_fd_sc_hd__mux2_1
XFILLER_38_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5956_ _6788_/Q _5980_/A2 wire675/X _6657_/Q _5955_/X VGND VGND VPWR VPWR _5959_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_178_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5887_ _6576_/Q wire684/X wire671/X _5886_/X VGND VGND VPWR VPWR _5887_/X sky130_fd_sc_hd__a22o_1
X_4907_ _4907_/A _5071_/C _4907_/C _4907_/D VGND VGND VPWR VPWR _4907_/X sky130_fd_sc_hd__or4_1
XFILLER_40_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4838_ _5037_/A _4838_/B VGND VGND VPWR VPWR _4838_/X sky130_fd_sc_hd__or2_1
XFILLER_119_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4769_ _5013_/A _5135_/A VGND VGND VPWR VPWR _5142_/A sky130_fd_sc_hd__or2_4
XFILLER_5_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6508_ _6930_/CLK _6508_/D fanout884/X VGND VGND VPWR VPWR _6508_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_134_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6439_ _6446_/A _6447_/B VGND VGND VPWR VPWR _6439_/X sky130_fd_sc_hd__and2_1
XFILLER_136_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold10 hold10/A VGND VGND VPWR VPWR hold6/A sky130_fd_sc_hd__bufbuf_16
Xhold32 hold32/A VGND VGND VPWR VPWR hold32/X sky130_fd_sc_hd__bufbuf_16
Xhold21 hold21/A VGND VGND VPWR VPWR hold21/X sky130_fd_sc_hd__bufbuf_16
XFILLER_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold54 hold54/A VGND VGND VPWR VPWR hold54/X sky130_fd_sc_hd__bufbuf_16
Xhold65 hold65/A VGND VGND VPWR VPWR hold65/X sky130_fd_sc_hd__bufbuf_16
XFILLER_76_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold43 hold43/A VGND VGND VPWR VPWR hold43/X sky130_fd_sc_hd__bufbuf_16
XFILLER_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold76 hold80/X VGND VGND VPWR VPWR hold81/A sky130_fd_sc_hd__bufbuf_16
Xhold98 hold98/A VGND VGND VPWR VPWR hold98/X sky130_fd_sc_hd__bufbuf_16
Xhold87 hold87/A VGND VGND VPWR VPWR hold87/X sky130_fd_sc_hd__bufbuf_16
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3240__1 _3545_/A1 VGND VGND VPWR VPWR _6458_/CLK sky130_fd_sc_hd__inv_2
XFILLER_43_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_7 _6440_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5810_ _7002_/Q wire710/X wire689/X _7050_/Q VGND VGND VPWR VPWR _5810_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6790_ _3545_/A1 _6790_/D _6448_/X VGND VGND VPWR VPWR _6790_/Q sky130_fd_sc_hd__dfrtn_1
X_5741_ _5741_/A _5741_/B _5741_/C VGND VGND VPWR VPWR _5741_/X sky130_fd_sc_hd__or3_1
XFILLER_50_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5672_ _7164_/Q _7163_/Q VGND VGND VPWR VPWR _5701_/C sky130_fd_sc_hd__and2_4
XFILLER_30_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4623_ _4623_/A _4623_/B _4623_/C _4623_/D VGND VGND VPWR VPWR _4623_/X sky130_fd_sc_hd__and4_2
Xhold502 _6676_/Q VGND VGND VPWR VPWR hold502/X sky130_fd_sc_hd__bufbuf_16
X_4554_ _4554_/A _4554_/B VGND VGND VPWR VPWR _4554_/X sky130_fd_sc_hd__and2_4
Xhold513 _3979_/X VGND VGND VPWR VPWR hold513/X sky130_fd_sc_hd__bufbuf_16
XFILLER_116_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold524 _6819_/Q VGND VGND VPWR VPWR hold524/X sky130_fd_sc_hd__bufbuf_16
X_3505_ _3505_/A _5252_/B VGND VGND VPWR VPWR _4172_/A sky130_fd_sc_hd__nor2_8
Xhold535 _6595_/Q VGND VGND VPWR VPWR hold535/X sky130_fd_sc_hd__bufbuf_16
Xhold568 _6912_/Q VGND VGND VPWR VPWR hold568/X sky130_fd_sc_hd__bufbuf_16
Xhold579 _6904_/Q VGND VGND VPWR VPWR hold579/X sky130_fd_sc_hd__bufbuf_16
X_4485_ _4485_/A VGND VGND VPWR VPWR _4554_/A sky130_fd_sc_hd__inv_4
XFILLER_171_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6224_ _6908_/Q wire600/X wire646/X wire531/X _6223_/X VGND VGND VPWR VPWR _6231_/A
+ sky130_fd_sc_hd__a221o_1
Xhold546 _6725_/Q VGND VGND VPWR VPWR hold546/X sky130_fd_sc_hd__bufbuf_16
XFILLER_116_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold557 _6739_/Q VGND VGND VPWR VPWR hold557/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3436_ _3436_/A _3436_/B _3436_/C _3436_/D VGND VGND VPWR VPWR _3452_/A sky130_fd_sc_hd__or4_4
XFILLER_103_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6155_ _6977_/Q wire641/X wire639/X _6881_/Q _6154_/X VGND VGND VPWR VPWR _6156_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3367_ _3367_/A _3421_/C VGND VGND VPWR VPWR _3368_/B sky130_fd_sc_hd__or2_4
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _4745_/A _4947_/B _5017_/A VGND VGND VPWR VPWR _5108_/B sky130_fd_sc_hd__a21oi_1
XFILLER_85_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6086_ _7190_/Q _6110_/S _6084_/X _6085_/X VGND VGND VPWR VPWR _7190_/D sky130_fd_sc_hd__o22a_1
XFILLER_57_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5037_ _5037_/A _5037_/B _5003_/X VGND VGND VPWR VPWR _5158_/A sky130_fd_sc_hd__or3b_4
X_3298_ _3508_/A _3668_/A VGND VGND VPWR VPWR _3298_/Y sky130_fd_sc_hd__nor2_8
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6988_ _7136_/CLK _6988_/D fanout871/X VGND VGND VPWR VPWR _6988_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_53_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5939_ wire824/X _7185_/Q wire381/X VGND VGND VPWR VPWR _5939_/X sky130_fd_sc_hd__a21o_1
XFILLER_139_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput111 wb_adr_i[20] VGND VGND VPWR VPWR _4722_/A sky130_fd_sc_hd__buf_8
Xinput100 wb_adr_i[10] VGND VGND VPWR VPWR _4351_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_76_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput144 wb_dat_i[20] VGND VGND VPWR VPWR _6389_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput133 wb_dat_i[10] VGND VGND VPWR VPWR _6384_/B1 sky130_fd_sc_hd__clkbuf_4
Xinput122 wb_adr_i[30] VGND VGND VPWR VPWR _3892_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_49_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput155 wb_dat_i[30] VGND VGND VPWR VPWR _6396_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput166 wb_sel_i[1] VGND VGND VPWR VPWR _6371_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_48_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4270_ hold325/X wire790/A _4273_/S VGND VGND VPWR VPWR _4270_/X sky130_fd_sc_hd__mux2_1
X_3221_ _3221_/A VGND VGND VPWR VPWR _3221_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6911_ _7145_/CLK _6911_/D fanout883/X VGND VGND VPWR VPWR _6911_/Q sky130_fd_sc_hd__dfrtp_2
X_6842_ _6842_/CLK _6842_/D fanout857/X VGND VGND VPWR VPWR _6842_/Q sky130_fd_sc_hd__dfrtp_1
X_3985_ hold417/X hold79/X _3993_/S VGND VGND VPWR VPWR _3985_/X sky130_fd_sc_hd__mux2_8
X_6773_ _7225_/CLK _6773_/D fanout850/X VGND VGND VPWR VPWR _6773_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5724_ _6998_/Q wire710/X wire689/X _7046_/Q VGND VGND VPWR VPWR _5724_/X sky130_fd_sc_hd__a22o_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5655_ _6679_/Q _5653_/X _5654_/Y _7171_/Q VGND VGND VPWR VPWR _7171_/D sky130_fd_sc_hd__a22o_1
XFILLER_190_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4606_ _4775_/A _4694_/A VGND VGND VPWR VPWR _4917_/A sky130_fd_sc_hd__or2_4
Xhold310 _6694_/Q VGND VGND VPWR VPWR hold310/X sky130_fd_sc_hd__bufbuf_16
XFILLER_190_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5586_ _5595_/A0 hold730/X _5593_/S VGND VGND VPWR VPWR _7141_/D sky130_fd_sc_hd__mux2_1
X_4537_ _4533_/A _4533_/B _4537_/C _4538_/A VGND VGND VPWR VPWR _4537_/X sky130_fd_sc_hd__and4bb_4
XFILLER_132_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold343 _6921_/Q VGND VGND VPWR VPWR hold343/X sky130_fd_sc_hd__bufbuf_16
XFILLER_117_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold332 _3253_/X VGND VGND VPWR VPWR hold332/X sky130_fd_sc_hd__bufbuf_16
Xhold321 _7041_/Q VGND VGND VPWR VPWR hold321/X sky130_fd_sc_hd__bufbuf_16
Xhold387 _6843_/Q VGND VGND VPWR VPWR hold387/X sky130_fd_sc_hd__bufbuf_16
Xhold354 _7156_/Q VGND VGND VPWR VPWR hold354/X sky130_fd_sc_hd__bufbuf_16
Xhold376 _5350_/X VGND VGND VPWR VPWR _6932_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_131_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4468_ _4758_/A _5004_/A VGND VGND VPWR VPWR _4818_/C sky130_fd_sc_hd__nand2_2
Xhold365 _6712_/Q VGND VGND VPWR VPWR hold365/X sky130_fd_sc_hd__bufbuf_16
XFILLER_89_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold398 _6653_/Q VGND VGND VPWR VPWR hold398/X sky130_fd_sc_hd__bufbuf_16
X_3419_ hold43/X _3421_/C VGND VGND VPWR VPWR _3419_/X sky130_fd_sc_hd__or2_4
X_7187_ _7220_/CLK _7187_/D fanout854/X VGND VGND VPWR VPWR _7187_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout823 _6678_/Q VGND VGND VPWR VPWR _5663_/A sky130_fd_sc_hd__buf_8
X_6207_ _6232_/A _6207_/B _6207_/C _6207_/D VGND VGND VPWR VPWR _6207_/X sky130_fd_sc_hd__or4_1
X_4399_ _4400_/A _4513_/A VGND VGND VPWR VPWR _4399_/Y sky130_fd_sc_hd__nor2_4
X_6138_ _7025_/Q _6010_/Y wire616/X _7089_/Q _6137_/X VGND VGND VPWR VPWR _6144_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_58_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout856 wire860/A VGND VGND VPWR VPWR fanout856/X sky130_fd_sc_hd__buf_8
Xfanout867 fanout868/A VGND VGND VPWR VPWR fanout867/X sky130_fd_sc_hd__buf_8
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout889 fanout890/X VGND VGND VPWR VPWR fanout889/X sky130_fd_sc_hd__buf_8
XFILLER_133_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout878 fanout890/X VGND VGND VPWR VPWR fanout878/X sky130_fd_sc_hd__buf_8
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6069_ _7070_/Q _6009_/X wire627/X wire529/X VGND VGND VPWR VPWR _6069_/X sky130_fd_sc_hd__a22o_1
XFILLER_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_216 wire560/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_205 wire498/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_227 wire650/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_249 wire796/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_238 wire739/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3770_ wire479/X hold97/A _5185_/A _6785_/Q _3745_/X VGND VGND VPWR VPWR _3793_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5440_ wire739/X hold657/X _5440_/S VGND VGND VPWR VPWR _7012_/D sky130_fd_sc_hd__mux2_1
XFILLER_8_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5371_ wire794/A _6950_/Q _5377_/S VGND VGND VPWR VPWR _6950_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7110_ _7151_/CLK hold98/X fanout880/X VGND VGND VPWR VPWR _7110_/Q sky130_fd_sc_hd__dfstp_4
X_4322_ _4322_/A _6406_/B VGND VGND VPWR VPWR _4327_/S sky130_fd_sc_hd__nand2_4
X_4253_ _5408_/A1 hold692/X _4255_/S VGND VGND VPWR VPWR _6710_/D sky130_fd_sc_hd__mux2_1
X_7041_ _7129_/CLK _7041_/D fanout863/X VGND VGND VPWR VPWR _7041_/Q sky130_fd_sc_hd__dfrtp_2
X_3204_ _3204_/A VGND VGND VPWR VPWR _3204_/Y sky130_fd_sc_hd__inv_2
X_4184_ _4184_/A _5242_/B VGND VGND VPWR VPWR _4189_/S sky130_fd_sc_hd__and2_4
XFILLER_95_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A VGND VGND VPWR VPWR _3949_/A1 sky130_fd_sc_hd__clkbuf_8
X_6825_ _7103_/CLK _6825_/D fanout861/X VGND VGND VPWR VPWR _6825_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6756_ _6824_/CLK _6756_/D fanout848/X VGND VGND VPWR VPWR _6756_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3968_ _6706_/Q _3974_/B VGND VGND VPWR VPWR _6700_/D sky130_fd_sc_hd__and2_1
XFILLER_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5707_ _7165_/Q _5707_/B _5707_/C VGND VGND VPWR VPWR _5707_/X sky130_fd_sc_hd__and3_4
Xwire509 _7037_/Q VGND VGND VPWR VPWR wire509/X sky130_fd_sc_hd__buf_6
XFILLER_12_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3899_ _6664_/Q _3898_/A _3898_/Y _6666_/Q VGND VGND VPWR VPWR _6664_/D sky130_fd_sc_hd__a22o_1
X_6687_ _6851_/CLK _6687_/D _6447_/A VGND VGND VPWR VPWR _6687_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_164_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5638_ _7167_/Q _7166_/Q VGND VGND VPWR VPWR _6037_/B sky130_fd_sc_hd__and2_4
XFILLER_163_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5569_ _5578_/A0 hold394/X _5575_/S VGND VGND VPWR VPWR _7126_/D sky130_fd_sc_hd__mux2_1
Xhold151 _5563_/X VGND VGND VPWR VPWR _7121_/D sky130_fd_sc_hd__bufbuf_16
Xhold162 _3987_/X VGND VGND VPWR VPWR hold162/X sky130_fd_sc_hd__bufbuf_16
Xhold140 hold29/X VGND VGND VPWR VPWR hold140/X sky130_fd_sc_hd__bufbuf_16
Xhold195 _6465_/Q VGND VGND VPWR VPWR hold54/A sky130_fd_sc_hd__bufbuf_16
XFILLER_105_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold173 _6781_/Q VGND VGND VPWR VPWR hold85/A sky130_fd_sc_hd__bufbuf_16
Xhold184 _6477_/Q VGND VGND VPWR VPWR hold184/X sky130_fd_sc_hd__bufbuf_16
XFILLER_77_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length652 _5707_/X VGND VGND VPWR VPWR wire651/A sky130_fd_sc_hd__buf_6
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length685 _5689_/X VGND VGND VPWR VPWR _5814_/A2 sky130_fd_sc_hd__buf_6
Xmax_length663 _5703_/X VGND VGND VPWR VPWR _5794_/B1 sky130_fd_sc_hd__buf_6
Xmax_length696 wire697/X VGND VGND VPWR VPWR _5979_/A2 sky130_fd_sc_hd__buf_6
XFILLER_142_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4940_ _5034_/A _4940_/B _4940_/C _4940_/D VGND VGND VPWR VPWR _4941_/D sky130_fd_sc_hd__or4_1
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4871_ _4871_/A _5164_/B VGND VGND VPWR VPWR _4899_/B sky130_fd_sc_hd__and2_4
XFILLER_177_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6610_ _6747_/CLK _6610_/D fanout874/X VGND VGND VPWR VPWR _6610_/Q sky130_fd_sc_hd__dfrtp_2
X_3822_ _3821_/X _6483_/Q _3840_/S VGND VGND VPWR VPWR _6483_/D sky130_fd_sc_hd__mux2_1
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6541_ _6650_/CLK _6541_/D fanout858/X VGND VGND VPWR VPWR _6541_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_193_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3753_ _6973_/Q _5396_/A _4130_/A _6604_/Q _3752_/X VGND VGND VPWR VPWR _3754_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_9_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6472_ _3545_/A1 _6472_/D _6427_/X VGND VGND VPWR VPWR _6472_/Q sky130_fd_sc_hd__dfrtp_2
X_3684_ _7086_/Q _5522_/A _5513_/A _7078_/Q _3683_/X VGND VGND VPWR VPWR _3687_/B
+ sky130_fd_sc_hd__a221o_1
Xoutput201 _3207_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[33] sky130_fd_sc_hd__buf_8
XFILLER_145_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5423_ _5423_/A _5459_/B VGND VGND VPWR VPWR _5429_/S sky130_fd_sc_hd__nand2_8
Xoutput234 _6519_/Q VGND VGND VPWR VPWR mgmt_gpio_out[29] sky130_fd_sc_hd__buf_8
Xoutput223 _6672_/Q VGND VGND VPWR VPWR mgmt_gpio_out[19] sky130_fd_sc_hd__buf_8
X_5354_ _5498_/A0 hold729/X _5359_/S VGND VGND VPWR VPWR _6935_/D sky130_fd_sc_hd__mux2_1
Xoutput212 _3231_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[9] sky130_fd_sc_hd__buf_8
Xoutput245 _6685_/Q VGND VGND VPWR VPWR mgmt_gpio_out[4] sky130_fd_sc_hd__buf_8
Xoutput267 _6801_/Q VGND VGND VPWR VPWR pll_div[1] sky130_fd_sc_hd__buf_8
Xoutput256 _3960_/A VGND VGND VPWR VPWR pad_flash_io0_ieb sky130_fd_sc_hd__buf_8
X_4305_ hold771/X _6407_/A0 _4309_/S VGND VGND VPWR VPWR _6753_/D sky130_fd_sc_hd__mux2_1
X_5285_ _5600_/A0 hold474/X _5287_/S VGND VGND VPWR VPWR _6874_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput289 _6817_/Q VGND VGND VPWR VPWR pll_trim[22] sky130_fd_sc_hd__buf_8
Xoutput278 _6492_/Q VGND VGND VPWR VPWR pll_trim[12] sky130_fd_sc_hd__buf_8
X_4236_ _4236_/A _4236_/B _4236_/C VGND VGND VPWR VPWR _4238_/B sky130_fd_sc_hd__nor3_4
XFILLER_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7024_ _7095_/CLK _7024_/D fanout862/X VGND VGND VPWR VPWR _7024_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_74_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4167_ wire799/A hold589/X _4171_/S VGND VGND VPWR VPWR _6634_/D sky130_fd_sc_hd__mux2_1
X_4098_ _5487_/A0 hold794/X _4102_/S VGND VGND VPWR VPWR _6576_/D sky130_fd_sc_hd__mux2_1
XFILLER_82_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_4_csclk _6744_/CLK VGND VGND VPWR VPWR _6608_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6808_ _6810_/CLK _6808_/D fanout853/X VGND VGND VPWR VPWR _6808_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_51_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6739_ _6806_/CLK _6739_/D _6435_/A VGND VGND VPWR VPWR _6739_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_137_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire840 wire840/A VGND VGND VPWR VPWR _7227_/A sky130_fd_sc_hd__buf_6
XFILLER_183_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire895 wire895/A VGND VGND VPWR VPWR _3969_/A sky130_fd_sc_hd__buf_4
XFILLER_127_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5070_ _4749_/C _5005_/C _4965_/A VGND VGND VPWR VPWR _5076_/C sky130_fd_sc_hd__a21oi_1
X_4021_ hold344/X _5601_/A0 _4021_/S VGND VGND VPWR VPWR _4021_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5972_ _6549_/Q wire706/X wire686/X _6772_/Q VGND VGND VPWR VPWR _5972_/X sky130_fd_sc_hd__a22o_1
X_4923_ _4672_/A _4672_/B _4711_/C _4936_/B _4936_/C VGND VGND VPWR VPWR _5024_/C
+ sky130_fd_sc_hd__a311o_1
XFILLER_80_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4854_ _4409_/Y _4845_/B _4846_/X VGND VGND VPWR VPWR _4854_/X sky130_fd_sc_hd__a21o_1
XFILLER_21_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4785_ _4500_/A _4622_/B _4758_/C _4689_/Y VGND VGND VPWR VPWR _5180_/A sky130_fd_sc_hd__a22o_1
XFILLER_21_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3805_ _6664_/Q _3845_/A VGND VGND VPWR VPWR _3825_/B sky130_fd_sc_hd__nand2b_2
X_6524_ _6930_/CLK hold74/X fanout887/X VGND VGND VPWR VPWR _6524_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3736_ input43/X _3736_/A2 wire388/X wire559/X VGND VGND VPWR VPWR _3736_/X sky130_fd_sc_hd__a22o_2
XFILLER_146_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6455_ _6455_/A _6455_/B VGND VGND VPWR VPWR _6455_/X sky130_fd_sc_hd__and2_1
X_3667_ _3666_/X _6792_/Q _3928_/A VGND VGND VPWR VPWR _6792_/D sky130_fd_sc_hd__mux2_1
X_6386_ _4236_/C _6386_/A2 _6386_/B1 _4236_/A VGND VGND VPWR VPWR _6386_/X sky130_fd_sc_hd__a22o_1
X_5406_ hold581/X hold465/X _5413_/S VGND VGND VPWR VPWR _6981_/D sky130_fd_sc_hd__mux2_1
X_3598_ _3598_/A _3598_/B _3598_/C _3598_/D VGND VGND VPWR VPWR _3606_/C sky130_fd_sc_hd__or4_1
XFILLER_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5337_ hold628/X wire773/X _5341_/S VGND VGND VPWR VPWR _6920_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5268_ hold821/X _5547_/A0 _5269_/S VGND VGND VPWR VPWR _6859_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4219_ _5252_/B _5252_/C _4007_/X _3361_/Y wire729/A VGND VGND VPWR VPWR _4235_/S
+ sky130_fd_sc_hd__o221a_4
X_7007_ _7103_/CLK _7007_/D fanout861/X VGND VGND VPWR VPWR _7007_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_75_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5199_ _6411_/A0 hold634/X _5199_/S VGND VGND VPWR VPWR _6804_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4570_ _5071_/A VGND VGND VPWR VPWR _4623_/B sky130_fd_sc_hd__inv_2
XFILLER_162_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3521_ _6937_/Q _5351_/A _4280_/A _6737_/Q _3519_/X VGND VGND VPWR VPWR _3522_/D
+ sky130_fd_sc_hd__a221o_4
Xwire670 _5699_/X VGND VGND VPWR VPWR wire670/X sky130_fd_sc_hd__buf_8
Xhold717 _7063_/Q VGND VGND VPWR VPWR hold717/X sky130_fd_sc_hd__bufbuf_16
XFILLER_116_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire692 wire692/A VGND VGND VPWR VPWR wire692/X sky130_fd_sc_hd__buf_8
Xhold706 _7091_/Q VGND VGND VPWR VPWR hold706/X sky130_fd_sc_hd__bufbuf_16
Xhold728 _6721_/Q VGND VGND VPWR VPWR hold728/X sky130_fd_sc_hd__bufbuf_16
XFILLER_115_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6240_ _6535_/Q wire585/X _6352_/B1 _6639_/Q _6239_/X VGND VGND VPWR VPWR _6247_/A
+ sky130_fd_sc_hd__a221o_2
Xhold739 _4223_/X VGND VGND VPWR VPWR _6682_/D sky130_fd_sc_hd__bufbuf_16
X_3452_ _3452_/A _3452_/B _3452_/C _3452_/D VGND VGND VPWR VPWR _3452_/X sky130_fd_sc_hd__or4_1
X_6171_ _7114_/Q wire650/X _6021_/B _7154_/Q VGND VGND VPWR VPWR _6171_/X sky130_fd_sc_hd__a22o_1
XFILLER_170_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3383_ _3421_/A _3421_/B _3383_/C VGND VGND VPWR VPWR _5234_/B sky130_fd_sc_hd__or3_4
XFILLER_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5122_ _4749_/C _5005_/C _4898_/B _4953_/A VGND VGND VPWR VPWR _5124_/C sky130_fd_sc_hd__a31o_1
XFILLER_85_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5053_ _4745_/A _4648_/B _5164_/B _4818_/C _5052_/X VGND VGND VPWR VPWR _5157_/A
+ sky130_fd_sc_hd__o221ai_2
XFILLER_38_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4004_ _4004_/A _5576_/B VGND VGND VPWR VPWR _4006_/S sky130_fd_sc_hd__nand2_1
XFILLER_65_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5955_ _6751_/Q _5979_/A2 wire662/X _6543_/Q VGND VGND VPWR VPWR _5955_/X sky130_fd_sc_hd__a22o_1
X_5886_ _6624_/Q _5963_/B VGND VGND VPWR VPWR _5886_/X sky130_fd_sc_hd__or2_1
X_4906_ _5174_/C _4906_/B _4906_/C _4906_/D VGND VGND VPWR VPWR _4907_/D sky130_fd_sc_hd__or4_2
XFILLER_139_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4837_ _4898_/B _4717_/B _4757_/B _5164_/B VGND VGND VPWR VPWR _4837_/X sky130_fd_sc_hd__o22a_1
XFILLER_193_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4768_ _4772_/A _4409_/Y _4453_/Y _4656_/X VGND VGND VPWR VPWR _4796_/B sky130_fd_sc_hd__a22o_2
XFILLER_146_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4699_ _4595_/B _4697_/Y _4698_/Y _5165_/A VGND VGND VPWR VPWR _4713_/A sky130_fd_sc_hd__o31a_2
X_6507_ _6930_/CLK _6507_/D fanout884/X VGND VGND VPWR VPWR _6507_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_107_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3719_ input72/X wire432/X _4178_/A _6645_/Q _3718_/X VGND VGND VPWR VPWR _3725_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6438_ _6446_/A _6447_/B VGND VGND VPWR VPWR _6438_/X sky130_fd_sc_hd__and2_1
XFILLER_161_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_22_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7111_/CLK sky130_fd_sc_hd__clkbuf_8
X_6369_ _7209_/Q wire352/X _6370_/S VGND VGND VPWR VPWR _7209_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold11 hold6/X VGND VGND VPWR VPWR hold11/X sky130_fd_sc_hd__bufbuf_16
Xhold22 hold22/A VGND VGND VPWR VPWR hold22/X sky130_fd_sc_hd__bufbuf_16
XFILLER_48_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold55 hold55/A VGND VGND VPWR VPWR hold55/X sky130_fd_sc_hd__bufbuf_16
Xhold33 hold33/A VGND VGND VPWR VPWR hold33/X sky130_fd_sc_hd__bufbuf_16
XFILLER_88_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold44 hold44/A VGND VGND VPWR VPWR hold44/X sky130_fd_sc_hd__bufbuf_16
Xhold77 hold82/X VGND VGND VPWR VPWR hold83/A sky130_fd_sc_hd__bufbuf_16
Xhold66 hold66/A VGND VGND VPWR VPWR hold66/X sky130_fd_sc_hd__bufbuf_16
Xhold99 hold99/A VGND VGND VPWR VPWR hold99/X sky130_fd_sc_hd__bufbuf_16
Xhold88 hold88/A VGND VGND VPWR VPWR hold88/X sky130_fd_sc_hd__bufbuf_16
Xclkbuf_leaf_37_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7154_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_28_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_mgmt_gpio_in[4] mgmt_gpio_in[4] VGND VGND VPWR VPWR clkbuf_0_mgmt_gpio_in[4]/X
+ sky130_fd_sc_hd__clkbuf_8
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_8 _6442_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5740_ _6942_/Q wire657/X wire651/X _7022_/Q _5739_/X VGND VGND VPWR VPWR _5741_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_188_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5671_ _7162_/Q _7161_/Q VGND VGND VPWR VPWR _5707_/B sky130_fd_sc_hd__and2b_4
XFILLER_30_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4622_ _4987_/A _4622_/B VGND VGND VPWR VPWR _4623_/D sky130_fd_sc_hd__nand2_1
XFILLER_190_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4553_ _4553_/A _4553_/B _4986_/C VGND VGND VPWR VPWR _4554_/B sky130_fd_sc_hd__nor3_2
X_4484_ _4533_/A _4484_/B _4484_/C VGND VGND VPWR VPWR _4485_/A sky130_fd_sc_hd__or3_4
XFILLER_144_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold514 hold514/A VGND VGND VPWR VPWR hold514/X sky130_fd_sc_hd__bufbuf_16
XFILLER_116_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold525 _6577_/Q VGND VGND VPWR VPWR hold525/X sky130_fd_sc_hd__bufbuf_16
Xhold503 _7129_/Q VGND VGND VPWR VPWR hold503/X sky130_fd_sc_hd__bufbuf_16
Xhold536 _6645_/Q VGND VGND VPWR VPWR hold536/X sky130_fd_sc_hd__bufbuf_16
X_3504_ _3504_/A _3504_/B _3504_/C _3504_/D VGND VGND VPWR VPWR _3547_/A sky130_fd_sc_hd__or4_2
X_3435_ input57/X _4025_/A hold65/A _7154_/Q _3424_/X VGND VGND VPWR VPWR _3436_/D
+ sky130_fd_sc_hd__a221o_4
XFILLER_143_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6223_ _6956_/Q wire637/X wire635/X _6932_/Q VGND VGND VPWR VPWR _6223_/X sky130_fd_sc_hd__a22o_1
XFILLER_116_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold569 _6605_/Q VGND VGND VPWR VPWR hold569/X sky130_fd_sc_hd__bufbuf_16
Xhold558 _4288_/X VGND VGND VPWR VPWR _6739_/D sky130_fd_sc_hd__bufbuf_16
Xhold547 _6734_/Q VGND VGND VPWR VPWR hold547/X sky130_fd_sc_hd__bufbuf_16
X_6154_ _7065_/Q wire648/X wire633/X _6913_/Q VGND VGND VPWR VPWR _6154_/X sky130_fd_sc_hd__a22o_1
XFILLER_97_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3366_ _7084_/Q _5513_/A _5576_/A _7140_/Q VGND VGND VPWR VPWR _3366_/X sky130_fd_sc_hd__a22o_1
X_5105_ _5105_/A _5105_/B _5105_/C VGND VGND VPWR VPWR _5157_/B sky130_fd_sc_hd__or3_4
XFILLER_112_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6085_ _5611_/A _7189_/Q wire381/A VGND VGND VPWR VPWR _6085_/X sky130_fd_sc_hd__a21o_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3297_ _7012_/Q _5432_/A _5504_/A _7076_/Q _3296_/X VGND VGND VPWR VPWR _3379_/A
+ sky130_fd_sc_hd__a221o_1
X_5036_ _5036_/A _5101_/A _5036_/C VGND VGND VPWR VPWR _5036_/X sky130_fd_sc_hd__or3_4
XFILLER_57_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6987_ _6987_/CLK _6987_/D fanout870/X VGND VGND VPWR VPWR _6987_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_81_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5938_ _6532_/Q _5722_/B _5927_/X _5937_/X _6308_/S VGND VGND VPWR VPWR _5938_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5869_ wire488/X wire691/X wire665/X _6956_/Q VGND VGND VPWR VPWR _5869_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput101 wb_adr_i[11] VGND VGND VPWR VPWR _4351_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_150_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput112 wb_adr_i[21] VGND VGND VPWR VPWR _4368_/A sky130_fd_sc_hd__clkbuf_8
Xinput123 wb_adr_i[31] VGND VGND VPWR VPWR _3892_/A sky130_fd_sc_hd__clkbuf_4
Xinput145 wb_dat_i[21] VGND VGND VPWR VPWR _6392_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput134 wb_dat_i[11] VGND VGND VPWR VPWR _6386_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_103_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput167 wb_sel_i[2] VGND VGND VPWR VPWR _6372_/B sky130_fd_sc_hd__clkbuf_4
Xinput156 wb_dat_i[31] VGND VGND VPWR VPWR _6398_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_102_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3220_ _3220_/A VGND VGND VPWR VPWR _3220_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6910_ _7145_/CLK _6910_/D fanout883/X VGND VGND VPWR VPWR _6910_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_63_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6841_ _7122_/CLK _6841_/D fanout887/X VGND VGND VPWR VPWR _6841_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6772_ _6810_/CLK _6772_/D fanout853/X VGND VGND VPWR VPWR _6772_/Q sky130_fd_sc_hd__dfrtp_2
X_3984_ _6490_/Q _6409_/A0 _3994_/S VGND VGND VPWR VPWR _6490_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5723_ _5663_/Y _5721_/X _5722_/X wire381/A _7176_/Q VGND VGND VPWR VPWR _7176_/D
+ sky130_fd_sc_hd__a32o_1
X_5654_ _5654_/A _5654_/B VGND VGND VPWR VPWR _5654_/Y sky130_fd_sc_hd__nor2_1
XFILLER_176_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4605_ _5023_/A _4694_/A VGND VGND VPWR VPWR _4787_/B sky130_fd_sc_hd__nor2_1
Xhold311 _4246_/X VGND VGND VPWR VPWR _6694_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_163_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold300 _6717_/Q VGND VGND VPWR VPWR hold300/X sky130_fd_sc_hd__bufbuf_16
X_5585_ _5585_/A _5585_/B VGND VGND VPWR VPWR _5593_/S sky130_fd_sc_hd__nand2_8
XFILLER_7_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4536_ _4949_/B _4536_/B VGND VGND VPWR VPWR _4536_/X sky130_fd_sc_hd__and2_4
Xhold344 _6528_/Q VGND VGND VPWR VPWR hold344/X sky130_fd_sc_hd__bufbuf_16
XFILLER_116_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold333 _3254_/X VGND VGND VPWR VPWR hold333/X sky130_fd_sc_hd__bufbuf_16
Xhold322 _5473_/X VGND VGND VPWR VPWR _7041_/D sky130_fd_sc_hd__bufbuf_16
X_4467_ _4722_/A _4467_/B VGND VGND VPWR VPWR _4819_/B sky130_fd_sc_hd__nand2_8
Xhold355 _5602_/X VGND VGND VPWR VPWR _7156_/D sky130_fd_sc_hd__bufbuf_16
Xhold366 _7116_/Q VGND VGND VPWR VPWR hold366/X sky130_fd_sc_hd__bufbuf_16
Xhold377 _7143_/Q VGND VGND VPWR VPWR hold377/X sky130_fd_sc_hd__bufbuf_16
XFILLER_144_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold388 _5250_/X VGND VGND VPWR VPWR _6843_/D sky130_fd_sc_hd__bufbuf_16
Xhold399 _7113_/Q VGND VGND VPWR VPWR hold399/X sky130_fd_sc_hd__bufbuf_16
X_4398_ _4930_/D VGND VGND VPWR VPWR _4398_/Y sky130_fd_sc_hd__inv_2
X_6206_ _6206_/A _6206_/B _6206_/C _6206_/D VGND VGND VPWR VPWR _6207_/D sky130_fd_sc_hd__or4_4
X_3418_ _7130_/Q hold89/A _5558_/A wire475/X VGND VGND VPWR VPWR _3418_/X sky130_fd_sc_hd__a22o_1
XFILLER_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7186_ _7220_/CLK _7186_/D wire860/X VGND VGND VPWR VPWR _7186_/Q sky130_fd_sc_hd__dfrtp_1
X_6137_ _7137_/Q wire643/X wire631/X wire484/X VGND VGND VPWR VPWR _6137_/X sky130_fd_sc_hd__a22o_1
Xfanout846 _6447_/A VGND VGND VPWR VPWR _6446_/A sky130_fd_sc_hd__buf_8
X_3349_ _3514_/A hold87/X VGND VGND VPWR VPWR _5423_/A sky130_fd_sc_hd__nor2_8
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout857 fanout858/X VGND VGND VPWR VPWR fanout857/X sky130_fd_sc_hd__buf_8
XFILLER_112_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout879 fanout890/X VGND VGND VPWR VPWR fanout879/X sky130_fd_sc_hd__buf_8
XFILLER_100_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout868 fanout868/A VGND VGND VPWR VPWR fanout868/X sky130_fd_sc_hd__buf_8
XFILLER_133_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6068_ _6998_/Q wire603/X _6140_/B1 _6918_/Q _6067_/X VGND VGND VPWR VPWR _6071_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_206 wire500/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5019_ _5003_/X _5018_/X _5156_/A VGND VGND VPWR VPWR _5019_/X sky130_fd_sc_hd__a21o_1
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_228 wire650/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_217 wire565/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_239 _5547_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length801 wire802/X VGND VGND VPWR VPWR _5532_/A0 sky130_fd_sc_hd__buf_6
XFILLER_158_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_732 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5370_ _5487_/A0 _6949_/Q _5377_/S VGND VGND VPWR VPWR _6949_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4321_ hold635/X _6411_/A0 _4321_/S VGND VGND VPWR VPWR _6767_/D sky130_fd_sc_hd__mux2_1
X_4252_ wire794/X hold674/X _4255_/S VGND VGND VPWR VPWR _6709_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7040_ _7129_/CLK _7040_/D fanout863/X VGND VGND VPWR VPWR _7040_/Q sky130_fd_sc_hd__dfrtp_2
X_3203_ _7152_/Q VGND VGND VPWR VPWR _3203_/Y sky130_fd_sc_hd__clkinv_2
X_4183_ hold414/X _4303_/A0 _4183_/S VGND VGND VPWR VPWR _6648_/D sky130_fd_sc_hd__mux2_1
XFILLER_94_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6824_ _6824_/CLK _6824_/D _6435_/A VGND VGND VPWR VPWR _6824_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6755_ _6824_/CLK _6755_/D fanout848/X VGND VGND VPWR VPWR _6755_/Q sky130_fd_sc_hd__dfstp_2
X_3967_ _6703_/Q _3974_/B VGND VGND VPWR VPWR _6701_/D sky130_fd_sc_hd__and2_1
X_5706_ _7165_/Q _5706_/B _5707_/B VGND VGND VPWR VPWR _5706_/X sky130_fd_sc_hd__and3_4
X_6686_ _6994_/CLK _6686_/D fanout870/X VGND VGND VPWR VPWR _6686_/Q sky130_fd_sc_hd__dfrtp_2
X_3898_ _3898_/A _3898_/B VGND VGND VPWR VPWR _3898_/Y sky130_fd_sc_hd__nor2_1
XFILLER_148_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5637_ _5621_/X _5663_/B _7166_/Q VGND VGND VPWR VPWR _7166_/D sky130_fd_sc_hd__mux2_1
X_5568_ hold465/X _7125_/Q hold91/X VGND VGND VPWR VPWR _7125_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold152 _7215_/Q VGND VGND VPWR VPWR hold152/X sky130_fd_sc_hd__bufbuf_16
XFILLER_163_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold130 _5387_/Y VGND VGND VPWR VPWR _5395_/S sky130_fd_sc_hd__bufbuf_16
XFILLER_117_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4519_ _4871_/A _4995_/A VGND VGND VPWR VPWR _4519_/Y sky130_fd_sc_hd__nor2_1
XFILLER_104_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold141 hold253/X VGND VGND VPWR VPWR hold141/X sky130_fd_sc_hd__bufbuf_16
X_5499_ hold83/A hold106/X _5501_/S VGND VGND VPWR VPWR _5499_/X sky130_fd_sc_hd__mux2_1
Xhold163 hold163/A VGND VGND VPWR VPWR hold163/X sky130_fd_sc_hd__bufbuf_16
Xhold185 _3270_/X VGND VGND VPWR VPWR hold185/X sky130_fd_sc_hd__bufbuf_16
Xhold174 hold85/X VGND VGND VPWR VPWR hold174/X sky130_fd_sc_hd__bufbuf_16
Xhold196 hold54/X VGND VGND VPWR VPWR hold196/X sky130_fd_sc_hd__bufbuf_16
XFILLER_144_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7169_ _3949_/A1 _7169_/D fanout870/X VGND VGND VPWR VPWR _7169_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_58_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length620 _6140_/B1 VGND VGND VPWR VPWR _6340_/B1 sky130_fd_sc_hd__buf_6
XFILLER_6_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4870_ _4870_/A VGND VGND VPWR VPWR _4903_/A sky130_fd_sc_hd__inv_2
XFILLER_91_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3821_ _6482_/Q _3845_/A _3820_/X VGND VGND VPWR VPWR _3821_/X sky130_fd_sc_hd__a21o_1
XFILLER_177_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6540_ _6591_/CLK _6540_/D fanout873/X VGND VGND VPWR VPWR _6540_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_186_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3752_ _7125_/Q hold89/A _4097_/A _6576_/Q VGND VGND VPWR VPWR _3752_/X sky130_fd_sc_hd__a22o_1
XFILLER_185_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3683_ _6854_/Q _5261_/A _3683_/B1 wire534/X VGND VGND VPWR VPWR _3683_/X sky130_fd_sc_hd__a22o_1
X_6471_ _6668_/CLK _6471_/D _6426_/X VGND VGND VPWR VPWR _6471_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_118_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5422_ wire739/A hold590/X _5422_/S VGND VGND VPWR VPWR _5422_/X sky130_fd_sc_hd__mux2_1
X_5353_ wire794/A _6934_/Q _5359_/S VGND VGND VPWR VPWR _6934_/D sky130_fd_sc_hd__mux2_1
Xoutput202 _3206_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[34] sky130_fd_sc_hd__buf_8
XFILLER_160_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput213 wire458/X VGND VGND VPWR VPWR mgmt_gpio_out[0] sky130_fd_sc_hd__buf_8
Xoutput224 wire387/X VGND VGND VPWR VPWR mgmt_gpio_out[1] sky130_fd_sc_hd__buf_8
Xoutput235 _6683_/Q VGND VGND VPWR VPWR mgmt_gpio_out[2] sky130_fd_sc_hd__buf_8
Xoutput246 _6686_/Q VGND VGND VPWR VPWR mgmt_gpio_out[5] sky130_fd_sc_hd__buf_8
Xoutput268 _6802_/Q VGND VGND VPWR VPWR pll_div[2] sky130_fd_sc_hd__buf_8
Xoutput257 _3960_/Y VGND VGND VPWR VPWR pad_flash_io0_oeb sky130_fd_sc_hd__buf_8
X_4304_ _4304_/A _6406_/B VGND VGND VPWR VPWR _4309_/S sky130_fd_sc_hd__and2_4
X_5284_ _5599_/A0 hold305/X _5287_/S VGND VGND VPWR VPWR _6873_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput279 _6493_/Q VGND VGND VPWR VPWR pll_trim[13] sky130_fd_sc_hd__buf_8
XFILLER_87_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7023_ _7103_/CLK _7023_/D fanout861/X VGND VGND VPWR VPWR _7023_/Q sky130_fd_sc_hd__dfrtp_2
X_4235_ hold677/X _4234_/X _4235_/S VGND VGND VPWR VPWR _6688_/D sky130_fd_sc_hd__mux2_1
X_4166_ _4166_/A _5242_/B VGND VGND VPWR VPWR _4171_/S sky130_fd_sc_hd__nand2_4
X_4097_ _4097_/A _5242_/B VGND VGND VPWR VPWR _4097_/Y sky130_fd_sc_hd__nand2_8
XFILLER_83_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6807_ _6810_/CLK _6807_/D _6435_/A VGND VGND VPWR VPWR _6807_/Q sky130_fd_sc_hd__dfrtp_2
X_4999_ _5121_/C _5118_/C _5078_/C _4985_/Y VGND VGND VPWR VPWR _5001_/C sky130_fd_sc_hd__or4b_1
XFILLER_11_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6738_ _6806_/CLK _6738_/D fanout853/X VGND VGND VPWR VPWR _6738_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6669_ _6930_/CLK _6669_/D fanout887/X VGND VGND VPWR VPWR _6669_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_164_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire841 wire841/A VGND VGND VPWR VPWR _3959_/B sky130_fd_sc_hd__buf_6
XFILLER_80_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire896 wire896/A VGND VGND VPWR VPWR _3877_/C sky130_fd_sc_hd__buf_8
XFILLER_142_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4020_ hold647/X _4019_/X _4024_/S VGND VGND VPWR VPWR _4020_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5971_ _6623_/Q wire707/X _5681_/X _6598_/Q _5970_/X VGND VGND VPWR VPWR _5976_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_80_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4922_ _4922_/A _5142_/A VGND VGND VPWR VPWR _5034_/A sky130_fd_sc_hd__or2_1
XFILLER_80_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4853_ _4581_/B _4634_/B _4839_/X _4842_/X _5140_/A VGND VGND VPWR VPWR _4853_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_100_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4784_ _4724_/B _4756_/B _4519_/Y VGND VGND VPWR VPWR _4800_/C sky130_fd_sc_hd__o21bai_1
XFILLER_60_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3804_ _3797_/X _3803_/X _3801_/B VGND VGND VPWR VPWR _6485_/D sky130_fd_sc_hd__o21ba_1
X_6523_ _6930_/CLK hold39/X fanout885/X VGND VGND VPWR VPWR _6523_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3735_ _5225_/A _5225_/B VGND VGND VPWR VPWR _3735_/Y sky130_fd_sc_hd__nor2_1
XFILLER_109_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6454_ _6455_/A _6455_/B VGND VGND VPWR VPWR _6454_/X sky130_fd_sc_hd__and2_1
XFILLER_161_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5405_ _5405_/A _5585_/B VGND VGND VPWR VPWR _5413_/S sky130_fd_sc_hd__and2_4
X_3666_ _3665_/X _6791_/Q _3857_/C VGND VGND VPWR VPWR _3666_/X sky130_fd_sc_hd__mux2_1
X_6385_ _6384_/X hold9/A _6400_/S VGND VGND VPWR VPWR _7213_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3597_ input29/X _3283_/Y _3320_/Y input6/X _3562_/X VGND VGND VPWR VPWR _3598_/D
+ sky130_fd_sc_hd__a221o_4
X_5336_ hold540/X _5336_/A1 _5341_/S VGND VGND VPWR VPWR _6919_/D sky130_fd_sc_hd__mux2_1
XFILLER_125_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5267_ hold825/X wire753/X _5269_/S VGND VGND VPWR VPWR _5267_/X sky130_fd_sc_hd__mux2_1
X_4218_ hold502/X _4217_/X _4218_/S VGND VGND VPWR VPWR _6676_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7006_ _7103_/CLK _7006_/D fanout862/X VGND VGND VPWR VPWR _7006_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_56_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5198_ _6410_/A0 hold671/X _5199_/S VGND VGND VPWR VPWR _6803_/D sky130_fd_sc_hd__mux2_1
X_4149_ hold796/X _5487_/A0 _4153_/S VGND VGND VPWR VPWR _6619_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire660 _5704_/X VGND VGND VPWR VPWR wire660/X sky130_fd_sc_hd__buf_8
X_3520_ _4241_/A _3520_/B VGND VGND VPWR VPWR _4280_/A sky130_fd_sc_hd__nor2_8
Xhold718 _6871_/Q VGND VGND VPWR VPWR hold718/X sky130_fd_sc_hd__bufbuf_16
Xwire671 _5698_/B VGND VGND VPWR VPWR wire671/X sky130_fd_sc_hd__buf_8
XFILLER_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold707 _5529_/X VGND VGND VPWR VPWR _7091_/D sky130_fd_sc_hd__bufbuf_16
Xhold729 _6935_/Q VGND VGND VPWR VPWR hold729/X sky130_fd_sc_hd__bufbuf_16
X_3451_ _3451_/A _3451_/B _3451_/C _3451_/D VGND VGND VPWR VPWR _3452_/D sky130_fd_sc_hd__or4_1
XFILLER_97_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3382_ _3381_/X _6797_/Q _3928_/A VGND VGND VPWR VPWR _6797_/D sky130_fd_sc_hd__mux2_1
X_6170_ _6170_/A _6170_/B _6170_/C _6170_/D VGND VGND VPWR VPWR _6170_/X sky130_fd_sc_hd__or4_1
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_3_csclk _6744_/CLK VGND VGND VPWR VPWR _6650_/CLK sky130_fd_sc_hd__clkbuf_8
X_5121_ _5121_/A _5121_/B _5121_/C _5121_/D VGND VGND VPWR VPWR _5135_/D sky130_fd_sc_hd__or4_1
X_5052_ _4660_/X _4724_/B _4819_/B _4724_/A VGND VGND VPWR VPWR _5052_/X sky130_fd_sc_hd__a211o_2
XFILLER_38_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4003_ _6503_/Q wire739/X _4003_/S VGND VGND VPWR VPWR _6503_/D sky130_fd_sc_hd__mux2_1
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5954_ _6579_/Q wire684/X _5941_/X _5944_/X VGND VGND VPWR VPWR _5959_/B sky130_fd_sc_hd__a211o_4
XFILLER_80_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4905_ _4950_/B _4905_/B _4905_/C _4905_/D VGND VGND VPWR VPWR _4906_/D sky130_fd_sc_hd__or4_2
X_5885_ _6563_/Q wire672/X _5931_/A2 _6540_/Q _5884_/X VGND VGND VPWR VPWR _5893_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_33_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4836_ _4697_/A _5005_/C _4832_/B VGND VGND VPWR VPWR _4836_/X sky130_fd_sc_hd__a21o_1
XFILLER_166_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4767_ _4871_/A _4997_/A _4724_/B _4886_/B VGND VGND VPWR VPWR _4767_/X sky130_fd_sc_hd__o22a_1
X_6506_ _6930_/CLK _6506_/D fanout884/X VGND VGND VPWR VPWR _6506_/Q sky130_fd_sc_hd__dfrtp_2
X_4698_ _4745_/A _5147_/B VGND VGND VPWR VPWR _4698_/Y sky130_fd_sc_hd__nor2_2
X_3718_ _7102_/Q _5540_/A _4328_/A _6774_/Q VGND VGND VPWR VPWR _3718_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3649_ wire507/X _5477_/A _5207_/A _6813_/Q _3648_/X VGND VGND VPWR VPWR _3654_/B
+ sky130_fd_sc_hd__a221o_1
X_6437_ _6446_/A _6447_/B VGND VGND VPWR VPWR _6437_/X sky130_fd_sc_hd__and2_1
XFILLER_121_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6368_ _7208_/Q wire351/X _6370_/S VGND VGND VPWR VPWR _7208_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5319_ _5598_/A0 hold579/X _5323_/S VGND VGND VPWR VPWR _6904_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold23 hold23/A VGND VGND VPWR VPWR hold23/X sky130_fd_sc_hd__bufbuf_16
Xhold12 hold12/A VGND VGND VPWR VPWR hold7/A sky130_fd_sc_hd__bufbuf_16
X_6299_ _6621_/Q wire623/X wire612/X _6651_/Q VGND VGND VPWR VPWR _6299_/X sky130_fd_sc_hd__a22o_1
Xhold34 hold34/A VGND VGND VPWR VPWR hold34/X sky130_fd_sc_hd__bufbuf_16
Xhold56 hold56/A VGND VGND VPWR VPWR hold56/X sky130_fd_sc_hd__bufbuf_16
Xhold45 hold45/A VGND VGND VPWR VPWR hold45/X sky130_fd_sc_hd__bufbuf_16
XFILLER_102_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold78 hold78/A VGND VGND VPWR VPWR hold78/X sky130_fd_sc_hd__bufbuf_16
Xhold67 hold67/A VGND VGND VPWR VPWR hold67/X sky130_fd_sc_hd__bufbuf_16
Xhold89 hold89/A VGND VGND VPWR VPWR hold89/X sky130_fd_sc_hd__bufbuf_16
XFILLER_75_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_9 _6457_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_606 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5670_ _6997_/Q _5667_/X _5974_/A2 _7061_/Q VGND VGND VPWR VPWR _5670_/X sky130_fd_sc_hd__a22o_1
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4621_ _4988_/A _4986_/C _4619_/X _4620_/X VGND VGND VPWR VPWR _4623_/C sky130_fd_sc_hd__o211a_1
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4552_ _4376_/Y _4987_/B _4920_/A _5136_/A _4551_/X VGND VGND VPWR VPWR _4552_/X
+ sky130_fd_sc_hd__a2111o_1
X_4483_ _4533_/A _4484_/C VGND VGND VPWR VPWR _4693_/B sky130_fd_sc_hd__nor2_2
XFILLER_183_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold515 hold515/A VGND VGND VPWR VPWR wire802/A sky130_fd_sc_hd__bufbuf_16
Xhold526 _6541_/Q VGND VGND VPWR VPWR hold526/X sky130_fd_sc_hd__bufbuf_16
Xwire490 _7090_/Q VGND VGND VPWR VPWR wire490/X sky130_fd_sc_hd__buf_6
Xhold504 _5572_/X VGND VGND VPWR VPWR _7129_/D sky130_fd_sc_hd__bufbuf_16
X_3503_ _7017_/Q _5441_/A _4166_/A _6638_/Q _3502_/X VGND VGND VPWR VPWR _3504_/D
+ sky130_fd_sc_hd__a221o_1
X_3434_ input40/X _4023_/S _5333_/A _6922_/Q _3418_/X VGND VGND VPWR VPWR _3436_/C
+ sky130_fd_sc_hd__a221o_2
XFILLER_131_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold537 _6840_/Q VGND VGND VPWR VPWR hold537/X sky130_fd_sc_hd__bufbuf_16
Xhold559 _7104_/Q VGND VGND VPWR VPWR hold559/X sky130_fd_sc_hd__bufbuf_16
Xhold548 _4282_/X VGND VGND VPWR VPWR _6734_/D sky130_fd_sc_hd__bufbuf_16
X_6222_ _7132_/Q wire597/X wire611/X _7012_/Q _6221_/X VGND VGND VPWR VPWR _6232_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6153_ _6865_/Q _6179_/A2 _6029_/X wire505/X _6152_/X VGND VGND VPWR VPWR _6156_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3365_ _3365_/A _3552_/B VGND VGND VPWR VPWR _3365_/Y sky130_fd_sc_hd__nor2_2
X_5104_ _4588_/X _5050_/C _4754_/B VGND VGND VPWR VPWR _5104_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_112_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6084_ _6854_/Q _6357_/A2 _6071_/X _6083_/X _3197_/Y VGND VGND VPWR VPWR _6084_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_57_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3296_ _7052_/Q _5477_/A _3395_/A2 wire552/X _3287_/X VGND VGND VPWR VPWR _3296_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5035_ _5035_/A _5035_/B _5035_/C _5035_/D VGND VGND VPWR VPWR _5166_/C sky130_fd_sc_hd__or4_1
XFILLER_85_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6986_ _6986_/CLK _6986_/D fanout879/X VGND VGND VPWR VPWR _6986_/Q sky130_fd_sc_hd__dfrtp_2
X_5937_ _5937_/A _5937_/B _5937_/C _5937_/D VGND VGND VPWR VPWR _5937_/X sky130_fd_sc_hd__or4_1
XFILLER_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5868_ _7084_/Q wire677/X _5694_/X wire541/X _5867_/X VGND VGND VPWR VPWR _5871_/C
+ sky130_fd_sc_hd__a221o_1
X_4819_ _4819_/A _4819_/B _5005_/A _4819_/D VGND VGND VPWR VPWR _4820_/B sky130_fd_sc_hd__or4_1
X_5799_ _6985_/Q _5963_/B VGND VGND VPWR VPWR _5799_/X sky130_fd_sc_hd__or2_1
XFILLER_193_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput102 wb_adr_i[12] VGND VGND VPWR VPWR _4350_/B sky130_fd_sc_hd__clkbuf_4
Xinput124 wb_adr_i[3] VGND VGND VPWR VPWR _4469_/A sky130_fd_sc_hd__buf_8
XFILLER_193_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput113 wb_adr_i[22] VGND VGND VPWR VPWR _4345_/B sky130_fd_sc_hd__clkbuf_4
Xinput135 wb_dat_i[12] VGND VGND VPWR VPWR _6390_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_103_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput168 wb_sel_i[3] VGND VGND VPWR VPWR _6402_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput157 wb_dat_i[3] VGND VGND VPWR VPWR _6387_/B1 sky130_fd_sc_hd__clkbuf_4
Xinput146 wb_dat_i[22] VGND VGND VPWR VPWR _6395_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_91_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6840_ _6842_/CLK _6840_/D fanout857/X VGND VGND VPWR VPWR _6840_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_63_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6771_ _6771_/CLK _6771_/D fanout855/X VGND VGND VPWR VPWR _6771_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3983_ hold5/X hold9/X _3993_/S VGND VGND VPWR VPWR hold10/A sky130_fd_sc_hd__mux2_4
X_5722_ _6853_/Q _5722_/B VGND VGND VPWR VPWR _5722_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_21_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7145_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_175_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5653_ _6037_/B _6035_/A _6037_/C VGND VGND VPWR VPWR _5653_/X sky130_fd_sc_hd__and3_4
XFILLER_191_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4604_ _4694_/A _4898_/B VGND VGND VPWR VPWR _4887_/B sky130_fd_sc_hd__nor2_1
X_5584_ wire739/X hold654/X _5584_/S VGND VGND VPWR VPWR _5584_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4535_ _4533_/A _4533_/B _4537_/C _4956_/B VGND VGND VPWR VPWR _4536_/B sky130_fd_sc_hd__and4bb_4
Xclkbuf_leaf_36_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7155_/CLK sky130_fd_sc_hd__clkbuf_8
Xhold301 _7115_/Q VGND VGND VPWR VPWR hold301/X sky130_fd_sc_hd__bufbuf_16
XFILLER_144_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold323 _6670_/Q VGND VGND VPWR VPWR hold323/X sky130_fd_sc_hd__bufbuf_16
Xhold312 _7057_/Q VGND VGND VPWR VPWR hold312/X sky130_fd_sc_hd__bufbuf_16
XFILLER_132_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold334 _3505_/A VGND VGND VPWR VPWR _3514_/A sky130_fd_sc_hd__bufbuf_16
X_4466_ _4722_/A _4467_/B VGND VGND VPWR VPWR _5004_/A sky130_fd_sc_hd__and2_4
Xhold356 _6884_/Q VGND VGND VPWR VPWR hold356/X sky130_fd_sc_hd__bufbuf_16
Xhold367 _5557_/X VGND VGND VPWR VPWR _7116_/D sky130_fd_sc_hd__bufbuf_16
Xhold345 _4041_/X VGND VGND VPWR VPWR _6528_/D sky130_fd_sc_hd__bufbuf_16
Xhold378 _5588_/X VGND VGND VPWR VPWR _7143_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_116_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4397_ _4775_/A _4671_/A VGND VGND VPWR VPWR _4930_/D sky130_fd_sc_hd__nand2_4
Xfanout803 hold465/X VGND VGND VPWR VPWR _5487_/A0 sky130_fd_sc_hd__buf_8
X_6205_ _6979_/Q wire641/X wire639/X _6883_/Q _6204_/X VGND VGND VPWR VPWR _6206_/D
+ sky130_fd_sc_hd__a221o_1
X_7185_ _7220_/CLK _7185_/D wire860/X VGND VGND VPWR VPWR _7185_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout825 _6667_/Q VGND VGND VPWR VPWR _3845_/A sky130_fd_sc_hd__buf_8
Xhold389 _7014_/Q VGND VGND VPWR VPWR hold389/X sky130_fd_sc_hd__bufbuf_16
X_3417_ _3416_/X _6796_/Q _3928_/A VGND VGND VPWR VPWR _6796_/D sky130_fd_sc_hd__mux2_1
X_3348_ _7148_/Q _5585_/A _5297_/A _6892_/Q VGND VGND VPWR VPWR _3348_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6136_ _7081_/Q _6211_/B VGND VGND VPWR VPWR _6136_/X sky130_fd_sc_hd__and2_1
Xfanout858 wire860/X VGND VGND VPWR VPWR fanout858/X sky130_fd_sc_hd__buf_8
Xfanout847 _6447_/A VGND VGND VPWR VPWR _6435_/A sky130_fd_sc_hd__buf_8
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout869 fanout871/X VGND VGND VPWR VPWR fanout869/X sky130_fd_sc_hd__buf_8
X_6067_ _7118_/Q _6339_/A2 _6339_/B1 _7030_/Q VGND VGND VPWR VPWR _6067_/X sky130_fd_sc_hd__a22o_1
X_3279_ _3309_/A _3314_/B VGND VGND VPWR VPWR _5225_/A sky130_fd_sc_hd__or2_4
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_207 _3218_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5018_ _5037_/A _5037_/B _5018_/C VGND VGND VPWR VPWR _5018_/X sky130_fd_sc_hd__or3_1
XFILLER_85_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_229 _5812_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_218 wire569/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6969_ _6969_/CLK _6969_/D fanout880/X VGND VGND VPWR VPWR _6969_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_41_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4320_ hold684/X _6410_/A0 _4321_/S VGND VGND VPWR VPWR _6766_/D sky130_fd_sc_hd__mux2_1
XFILLER_153_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4251_ _5487_/A0 hold831/X _4255_/S VGND VGND VPWR VPWR _6708_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3202_ _3202_/A VGND VGND VPWR VPWR _3202_/Y sky130_fd_sc_hd__inv_2
X_4182_ hold731/X _6410_/A0 _4183_/S VGND VGND VPWR VPWR _6647_/D sky130_fd_sc_hd__mux2_1
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xnet899_2 _3545_/A1 VGND VGND VPWR VPWR _3953_/B sky130_fd_sc_hd__inv_2
XFILLER_94_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7172__918 VGND VGND VPWR VPWR _7172_/D _7172__918/LO sky130_fd_sc_hd__conb_1
XFILLER_63_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6823_ _7091_/CLK _6823_/D fanout866/X VGND VGND VPWR VPWR _6823_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3966_ _6705_/Q _3974_/B VGND VGND VPWR VPWR _6702_/D sky130_fd_sc_hd__and2_1
X_6754_ _7223_/CLK _6754_/D fanout850/X VGND VGND VPWR VPWR _6754_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5705_ _5864_/B _5705_/B _5706_/B VGND VGND VPWR VPWR _5705_/X sky130_fd_sc_hd__and3_4
X_6685_ _6994_/CLK _6685_/D fanout870/X VGND VGND VPWR VPWR _6685_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_10_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5636_ _5635_/Y _3241_/Y _5636_/S VGND VGND VPWR VPWR _7165_/D sky130_fd_sc_hd__mux2_1
XFILLER_12_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3897_ _6703_/Q _3883_/X _3915_/B _6698_/Q VGND VGND VPWR VPWR _6703_/D sky130_fd_sc_hd__a22o_1
XFILLER_163_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5567_ hold89/X _5585_/B VGND VGND VPWR VPWR hold90/A sky130_fd_sc_hd__nand2_2
XFILLER_117_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5498_ _5498_/A0 hold717/X _5501_/S VGND VGND VPWR VPWR _7063_/D sky130_fd_sc_hd__mux2_1
Xhold153 hold162/X VGND VGND VPWR VPWR hold163/A sky130_fd_sc_hd__bufbuf_16
Xhold131 _5389_/X VGND VGND VPWR VPWR _6966_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_144_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4518_ _4871_/A _4990_/A VGND VGND VPWR VPWR _5081_/A sky130_fd_sc_hd__nor2_1
XFILLER_117_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold120 _3295_/Y VGND VGND VPWR VPWR wire439/A sky130_fd_sc_hd__bufbuf_16
Xhold142 hold142/A VGND VGND VPWR VPWR wire729/A sky130_fd_sc_hd__bufbuf_16
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4449_ _4534_/B _4449_/B VGND VGND VPWR VPWR _4572_/B sky130_fd_sc_hd__nand2_4
Xhold164 _4039_/X VGND VGND VPWR VPWR _6526_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_132_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold175 _3265_/X VGND VGND VPWR VPWR hold86/A sky130_fd_sc_hd__bufbuf_16
Xhold186 _3271_/X VGND VGND VPWR VPWR hold94/A sky130_fd_sc_hd__bufbuf_16
Xhold197 _3991_/X VGND VGND VPWR VPWR hold55/A sky130_fd_sc_hd__bufbuf_16
XFILLER_144_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7168_ _3949_/A1 _7168_/D fanout870/X VGND VGND VPWR VPWR _7168_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_86_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6119_ _3213_/A _6009_/X _6020_/D _6968_/Q VGND VGND VPWR VPWR _6119_/X sky130_fd_sc_hd__a22o_1
XFILLER_58_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7099_ _7139_/CLK _7099_/D fanout867/X VGND VGND VPWR VPWR _7099_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length621 _6191_/B1 VGND VGND VPWR VPWR _6140_/B1 sky130_fd_sc_hd__buf_6
XFILLER_185_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length654 _5706_/X VGND VGND VPWR VPWR wire653/A sky130_fd_sc_hd__buf_6
Xmax_length687 _5688_/X VGND VGND VPWR VPWR _5855_/B1 sky130_fd_sc_hd__buf_6
Xmax_length676 _5693_/X VGND VGND VPWR VPWR wire675/A sky130_fd_sc_hd__buf_6
XFILLER_135_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length698 _5680_/X VGND VGND VPWR VPWR _5977_/A2 sky130_fd_sc_hd__buf_6
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3820_ _3845_/A _3820_/B _3820_/C VGND VGND VPWR VPWR _3820_/X sky130_fd_sc_hd__and3b_1
X_3751_ _6949_/Q _5369_/A _3473_/Y _6550_/Q _3750_/X VGND VGND VPWR VPWR _3754_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6470_ _6668_/CLK _6470_/D _6425_/X VGND VGND VPWR VPWR _6470_/Q sky130_fd_sc_hd__dfrtp_2
X_3682_ input15/X _3283_/Y _4280_/A _6734_/Q _3681_/X VGND VGND VPWR VPWR _3687_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5421_ wire746/X hold788/X _5422_/S VGND VGND VPWR VPWR _6995_/D sky130_fd_sc_hd__mux2_1
Xoutput225 _6673_/Q VGND VGND VPWR VPWR mgmt_gpio_out[20] sky130_fd_sc_hd__buf_8
Xoutput203 wire443/X VGND VGND VPWR VPWR mgmt_gpio_oeb[35] sky130_fd_sc_hd__buf_8
XFILLER_173_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5352_ _5595_/A0 _6933_/Q _5359_/S VGND VGND VPWR VPWR _6933_/D sky130_fd_sc_hd__mux2_1
Xoutput214 _3937_/X VGND VGND VPWR VPWR mgmt_gpio_out[10] sky130_fd_sc_hd__buf_8
XFILLER_99_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput236 _6520_/Q VGND VGND VPWR VPWR mgmt_gpio_out[30] sky130_fd_sc_hd__buf_8
XFILLER_126_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput247 wire459/X VGND VGND VPWR VPWR mgmt_gpio_out[6] sky130_fd_sc_hd__buf_8
X_4303_ _4303_/A0 hold401/X _4303_/S VGND VGND VPWR VPWR _6752_/D sky130_fd_sc_hd__mux2_1
Xoutput258 _7227_/X VGND VGND VPWR VPWR pad_flash_io1_do sky130_fd_sc_hd__buf_8
X_5283_ _5598_/A0 hold564/X _5287_/S VGND VGND VPWR VPWR _6872_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7022_ _7103_/CLK _7022_/D fanout861/X VGND VGND VPWR VPWR _7022_/Q sky130_fd_sc_hd__dfstp_4
Xoutput269 _6803_/Q VGND VGND VPWR VPWR pll_div[3] sky130_fd_sc_hd__buf_8
XFILLER_141_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4234_ hold489/X wire739/A _4234_/S VGND VGND VPWR VPWR _4234_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4165_ _4303_/A0 hold429/X _4165_/S VGND VGND VPWR VPWR _6633_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4096_ _6575_/Q wire353/X _4096_/S VGND VGND VPWR VPWR _6575_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6806_ _6806_/CLK _6806_/D _6435_/A VGND VGND VPWR VPWR _6806_/Q sky130_fd_sc_hd__dfstp_4
X_4998_ _5114_/C _5116_/C VGND VGND VPWR VPWR _5001_/B sky130_fd_sc_hd__or2_1
X_6737_ _6950_/CLK _6737_/D fanout875/X VGND VGND VPWR VPWR _6737_/Q sky130_fd_sc_hd__dfrtp_2
X_3949_ _6512_/Q _3949_/A1 _6834_/Q VGND VGND VPWR VPWR _3949_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6668_ _6668_/CLK _6668_/D _6447_/X VGND VGND VPWR VPWR _6668_/Q sky130_fd_sc_hd__dfrtp_2
X_6599_ _6950_/CLK _6599_/D fanout874/X VGND VGND VPWR VPWR _6599_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_109_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5619_ _7160_/Q _5616_/A _5618_/Y VGND VGND VPWR VPWR _7160_/D sky130_fd_sc_hd__o21a_1
XFILLER_164_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire842 wire842/A VGND VGND VPWR VPWR wire842/X sky130_fd_sc_hd__buf_6
XFILLER_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length440 _3295_/Y VGND VGND VPWR VPWR _3395_/A2 sky130_fd_sc_hd__buf_6
XFILLER_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire897 wire897/A VGND VGND VPWR VPWR _7229_/A sky130_fd_sc_hd__buf_6
XFILLER_115_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5970_ _6712_/Q wire680/X wire664/X _6618_/Q VGND VGND VPWR VPWR _5970_/X sky130_fd_sc_hd__a22o_1
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4921_ _4930_/D _4575_/B _4933_/B _4684_/Y VGND VGND VPWR VPWR _4941_/B sky130_fd_sc_hd__a22o_2
XFILLER_80_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4852_ _4986_/C _4989_/B VGND VGND VPWR VPWR _5118_/B sky130_fd_sc_hd__nor2_1
XFILLER_60_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3803_ _6485_/Q _6664_/Q VGND VGND VPWR VPWR _3803_/X sky130_fd_sc_hd__or2_1
X_4783_ _4920_/B _5047_/A VGND VGND VPWR VPWR _4802_/B sky130_fd_sc_hd__or2_2
X_6522_ _6930_/CLK _6522_/D fanout885/X VGND VGND VPWR VPWR _6522_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3734_ input71/X wire432/X _4234_/S wire911/A VGND VGND VPWR VPWR _3734_/X sky130_fd_sc_hd__a22o_4
XFILLER_174_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3665_ _3665_/A _3665_/B _3665_/C VGND VGND VPWR VPWR _3665_/X sky130_fd_sc_hd__or3_4
X_6453_ _6455_/A _6455_/B VGND VGND VPWR VPWR _6453_/X sky130_fd_sc_hd__and2_1
X_5404_ hold371/X _5602_/A0 _5404_/S VGND VGND VPWR VPWR _5404_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6384_ _4236_/C _6384_/A2 _6384_/B1 _4236_/A _6383_/X VGND VGND VPWR VPWR _6384_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_114_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3596_ _6814_/Q _5207_/A _3995_/A _6499_/Q _3564_/X VGND VGND VPWR VPWR _3598_/C
+ sky130_fd_sc_hd__a221o_2
X_5335_ _6918_/Q hold38/X _5341_/S VGND VGND VPWR VPWR _6918_/D sky130_fd_sc_hd__mux2_1
XFILLER_125_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5266_ hold482/X _5572_/A0 _5269_/S VGND VGND VPWR VPWR _6857_/D sky130_fd_sc_hd__mux2_1
X_4217_ hold314/X _5602_/A0 hold46/X VGND VGND VPWR VPWR _4217_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7005_ _7103_/CLK _7005_/D fanout861/X VGND VGND VPWR VPWR _7005_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_56_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5197_ _6409_/A0 _6802_/Q _5199_/S VGND VGND VPWR VPWR _6802_/D sky130_fd_sc_hd__mux2_1
X_4148_ _4148_/A _4154_/B VGND VGND VPWR VPWR _4153_/S sky130_fd_sc_hd__and2_4
XFILLER_83_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4079_ _6560_/Q wire351/X _4081_/S VGND VGND VPWR VPWR _6560_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire650 _6027_/B VGND VGND VPWR VPWR wire650/X sky130_fd_sc_hd__buf_8
XFILLER_7_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold719 _6967_/Q VGND VGND VPWR VPWR hold719/X sky130_fd_sc_hd__bufbuf_16
XFILLER_171_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire672 _5694_/X VGND VGND VPWR VPWR wire672/X sky130_fd_sc_hd__buf_6
Xwire694 _5683_/X VGND VGND VPWR VPWR wire694/X sky130_fd_sc_hd__buf_8
Xhold708 _6808_/Q VGND VGND VPWR VPWR hold708/X sky130_fd_sc_hd__bufbuf_16
XFILLER_171_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3450_ _3450_/A _3450_/B _3450_/C _3450_/D VGND VGND VPWR VPWR _3451_/D sky130_fd_sc_hd__or4_1
X_3381_ wire353/X _6796_/Q _3857_/C VGND VGND VPWR VPWR _3381_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5120_ _5135_/A _5137_/B _5120_/C _5135_/C VGND VGND VPWR VPWR _5120_/X sky130_fd_sc_hd__or4_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5051_ _4692_/C _5049_/X _5050_/X VGND VGND VPWR VPWR _5056_/B sky130_fd_sc_hd__a21bo_4
XFILLER_69_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4002_ _6502_/Q _5547_/A0 _4003_/S VGND VGND VPWR VPWR _6502_/D sky130_fd_sc_hd__mux2_1
XFILLER_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5953_ _5953_/A _5953_/B _5953_/C _5953_/D VGND VGND VPWR VPWR _5953_/X sky130_fd_sc_hd__or4_2
X_4904_ _4950_/A _5129_/A _4904_/C _4904_/D VGND VGND VPWR VPWR _4905_/D sky130_fd_sc_hd__or4_1
X_5884_ _6589_/Q _5977_/A2 wire690/X _6644_/Q VGND VGND VPWR VPWR _5884_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4835_ _4898_/B _4832_/A _4832_/B _5164_/B VGND VGND VPWR VPWR _4835_/X sky130_fd_sc_hd__o22a_1
X_4766_ _4766_/A _5151_/A VGND VGND VPWR VPWR _4802_/A sky130_fd_sc_hd__or2_4
X_6505_ _6815_/CLK _6505_/D fanout861/X VGND VGND VPWR VPWR _6505_/Q sky130_fd_sc_hd__dfstp_4
X_3717_ _3717_/A _3717_/B _3717_/C _3717_/D VGND VGND VPWR VPWR _3726_/C sky130_fd_sc_hd__or4_2
X_4697_ _4697_/A _5062_/C VGND VGND VPWR VPWR _4697_/Y sky130_fd_sc_hd__nor2_1
XFILLER_162_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6436_ _6446_/A _6447_/B VGND VGND VPWR VPWR _6436_/X sky130_fd_sc_hd__and2_1
XFILLER_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3648_ _7039_/Q _3334_/Y _4196_/A _6661_/Q VGND VGND VPWR VPWR _3648_/X sky130_fd_sc_hd__a22o_1
X_3579_ _6617_/Q _4142_/A _4250_/A _6711_/Q VGND VGND VPWR VPWR _3579_/X sky130_fd_sc_hd__a22o_1
X_6367_ _7207_/Q _6367_/A1 _6370_/S VGND VGND VPWR VPWR _7207_/D sky130_fd_sc_hd__mux2_1
X_5318_ _5498_/A0 hold722/X _5323_/S VGND VGND VPWR VPWR _6903_/D sky130_fd_sc_hd__mux2_1
Xhold13 hold7/X VGND VGND VPWR VPWR hold13/X sky130_fd_sc_hd__bufbuf_16
X_6298_ _6578_/Q wire600/X wire645/X _6606_/Q _6286_/X VGND VGND VPWR VPWR _6305_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold24 hold24/A VGND VGND VPWR VPWR hold2/A sky130_fd_sc_hd__bufbuf_16
Xhold35 hold51/X VGND VGND VPWR VPWR hold52/A sky130_fd_sc_hd__bufbuf_16
Xhold46 hold46/A VGND VGND VPWR VPWR hold46/X sky130_fd_sc_hd__bufbuf_16
XFILLER_102_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5249_ _5249_/A0 hold460/X _5249_/S VGND VGND VPWR VPWR _5249_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold57 hold57/A VGND VGND VPWR VPWR hold57/X sky130_fd_sc_hd__bufbuf_16
Xhold79 hold79/A VGND VGND VPWR VPWR hold79/X sky130_fd_sc_hd__bufbuf_16
XFILLER_29_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold68 hold68/A VGND VGND VPWR VPWR hold68/X sky130_fd_sc_hd__bufbuf_16
XFILLER_84_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4620_ _4986_/A _4617_/A _4749_/C _4988_/A _4893_/A VGND VGND VPWR VPWR _4620_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_156_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4551_ _5079_/A _5078_/A _4551_/C VGND VGND VPWR VPWR _4551_/X sky130_fd_sc_hd__or3_1
Xhold505 _7114_/Q VGND VGND VPWR VPWR hold505/X sky130_fd_sc_hd__bufbuf_16
X_4482_ _4694_/A _4986_/C VGND VGND VPWR VPWR _4980_/A sky130_fd_sc_hd__nor2_2
Xhold527 _7119_/Q VGND VGND VPWR VPWR hold527/X sky130_fd_sc_hd__bufbuf_16
X_3502_ _7073_/Q _5504_/A _4178_/A _6648_/Q VGND VGND VPWR VPWR _3502_/X sky130_fd_sc_hd__a22o_1
Xhold516 _5433_/X VGND VGND VPWR VPWR _7005_/D sky130_fd_sc_hd__bufbuf_16
Xwire480 _7105_/Q VGND VGND VPWR VPWR wire480/X sky130_fd_sc_hd__buf_6
Xwire491 _7088_/Q VGND VGND VPWR VPWR _3211_/A sky130_fd_sc_hd__buf_8
X_6221_ _6892_/Q wire602/X wire581/X _7148_/Q _6220_/X VGND VGND VPWR VPWR _6221_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_143_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold549 _6565_/Q VGND VGND VPWR VPWR hold549/X sky130_fd_sc_hd__bufbuf_16
XFILLER_89_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3433_ wire490/X _5522_/A _3301_/Y _7026_/Q _3425_/X VGND VGND VPWR VPWR _3436_/B
+ sky130_fd_sc_hd__a221o_4
Xhold538 _5247_/X VGND VGND VPWR VPWR _6840_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_131_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6152_ wire480/X wire711/X _6022_/B _6945_/Q VGND VGND VPWR VPWR _6152_/X sky130_fd_sc_hd__a22o_2
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _5095_/X _5101_/X _5161_/C _4928_/Y VGND VGND VPWR VPWR _5103_/X sky130_fd_sc_hd__o211a_2
XFILLER_106_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ _3508_/A _3375_/B VGND VGND VPWR VPWR _5513_/A sky130_fd_sc_hd__nor2_8
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _6356_/A _6083_/B _6083_/C VGND VGND VPWR VPWR _6083_/X sky130_fd_sc_hd__or3_1
XFILLER_58_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3295_ _3668_/A _3353_/B VGND VGND VPWR VPWR _3295_/Y sky130_fd_sc_hd__nor2_8
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _5034_/A _5034_/B _5095_/C _5102_/B VGND VGND VPWR VPWR _5036_/C sky130_fd_sc_hd__or4b_1
XFILLER_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6985_ _6985_/CLK _6985_/D fanout878/X VGND VGND VPWR VPWR _6985_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_81_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5936_ _6730_/Q wire710/X wire679/X wire469/X _5935_/X VGND VGND VPWR VPWR _5937_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5867_ _6884_/Q wire706/X wire689/X _7052_/Q VGND VGND VPWR VPWR _5867_/X sky130_fd_sc_hd__a22o_1
XFILLER_193_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4818_ _4818_/A _4818_/B _4818_/C VGND VGND VPWR VPWR _5003_/C sky130_fd_sc_hd__or3_4
X_5798_ wire484/X _5926_/A2 wire678/X _7073_/Q _5797_/X VGND VGND VPWR VPWR _5806_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_193_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4749_ _4812_/A _4819_/B _4749_/C VGND VGND VPWR VPWR _4935_/D sky130_fd_sc_hd__or3_4
XFILLER_147_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6419_ _6420_/A _6421_/B VGND VGND VPWR VPWR _6419_/X sky130_fd_sc_hd__and2_1
XFILLER_134_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput125 wb_adr_i[4] VGND VGND VPWR VPWR _5050_/A sky130_fd_sc_hd__buf_8
Xinput114 wb_adr_i[23] VGND VGND VPWR VPWR _4345_/A sky130_fd_sc_hd__clkbuf_4
Xinput103 wb_adr_i[13] VGND VGND VPWR VPWR _4350_/A sky130_fd_sc_hd__clkbuf_4
Xinput136 wb_dat_i[13] VGND VGND VPWR VPWR _6392_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_163_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput158 wb_dat_i[4] VGND VGND VPWR VPWR _6389_/B1 sky130_fd_sc_hd__clkbuf_4
Xinput147 wb_dat_i[23] VGND VGND VPWR VPWR _6399_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_103_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput169 wb_stb_i VGND VGND VPWR VPWR wire912/A sky130_fd_sc_hd__buf_6
XFILLER_186_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_2_csclk _6744_/CLK VGND VGND VPWR VPWR _6842_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_12_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6770_ _6810_/CLK _6770_/D fanout853/X VGND VGND VPWR VPWR _6770_/Q sky130_fd_sc_hd__dfstp_4
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3982_ hold476/X wire790/X _3994_/S VGND VGND VPWR VPWR _6489_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5721_ _7069_/Q wire678/X _5709_/X _5713_/X _5720_/X VGND VGND VPWR VPWR _5721_/X
+ sky130_fd_sc_hd__a2111o_4
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5652_ _7171_/Q _7170_/Q VGND VGND VPWR VPWR _6036_/A sky130_fd_sc_hd__nand2b_4
XFILLER_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4603_ _4871_/A _4603_/B VGND VGND VPWR VPWR _4922_/A sky130_fd_sc_hd__nor2_4
X_5583_ wire749/X hold413/X _5584_/S VGND VGND VPWR VPWR _7139_/D sky130_fd_sc_hd__mux2_1
X_4534_ _4655_/A _4534_/B VGND VGND VPWR VPWR _4956_/B sky130_fd_sc_hd__nor2_2
Xhold302 _5556_/X VGND VGND VPWR VPWR _7115_/D sky130_fd_sc_hd__bufbuf_16
Xhold324 _4206_/X VGND VGND VPWR VPWR _6670_/D sky130_fd_sc_hd__bufbuf_16
Xhold313 _5491_/X VGND VGND VPWR VPWR _7057_/D sky130_fd_sc_hd__bufbuf_16
Xhold335 _6951_/Q VGND VGND VPWR VPWR hold335/X sky130_fd_sc_hd__bufbuf_16
XFILLER_117_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4465_ _4685_/A _4651_/B VGND VGND VPWR VPWR _4812_/A sky130_fd_sc_hd__or2_4
Xhold357 _7148_/Q VGND VGND VPWR VPWR hold357/X sky130_fd_sc_hd__bufbuf_16
Xhold346 _6931_/Q VGND VGND VPWR VPWR hold346/X sky130_fd_sc_hd__bufbuf_16
Xhold368 _6972_/Q VGND VGND VPWR VPWR hold368/X sky130_fd_sc_hd__bufbuf_16
XFILLER_144_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout804 hold465/X VGND VGND VPWR VPWR _5595_/A0 sky130_fd_sc_hd__buf_8
X_4396_ _4672_/A _4413_/C VGND VGND VPWR VPWR _4671_/A sky130_fd_sc_hd__nand2_8
X_6204_ wire495/X wire648/X wire633/X _6915_/Q VGND VGND VPWR VPWR _6204_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold379 _6628_/Q VGND VGND VPWR VPWR hold379/X sky130_fd_sc_hd__bufbuf_16
X_7184_ _7190_/CLK _7184_/D wire860/X VGND VGND VPWR VPWR _7184_/Q sky130_fd_sc_hd__dfrtp_4
X_3416_ wire352/X _6795_/Q _3857_/C VGND VGND VPWR VPWR _3416_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3347_ _3543_/A _3375_/B VGND VGND VPWR VPWR _5297_/A sky130_fd_sc_hd__nor2_8
X_6135_ _7192_/Q _6110_/S _6134_/X VGND VGND VPWR VPWR _7192_/D sky130_fd_sc_hd__o21a_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout848 _6447_/A VGND VGND VPWR VPWR fanout848/X sky130_fd_sc_hd__buf_8
XFILLER_100_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout859 fanout891/X VGND VGND VPWR VPWR wire860/A sky130_fd_sc_hd__buf_6
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6066_ _7014_/Q wire575/X _6335_/B _7038_/Q _6063_/X VGND VGND VPWR VPWR _6071_/B
+ sky130_fd_sc_hd__a221o_1
X_5017_ _5017_/A _5050_/C VGND VGND VPWR VPWR _5047_/D sky130_fd_sc_hd__nor2_1
X_3278_ _3293_/B _3278_/B VGND VGND VPWR VPWR _3278_/X sky130_fd_sc_hd__or2_1
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_208 _3218_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_219 wire570/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6968_ _6971_/CLK _6968_/D fanout879/X VGND VGND VPWR VPWR _6968_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_41_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6899_ _7147_/CLK _6899_/D fanout887/X VGND VGND VPWR VPWR _6899_/Q sky130_fd_sc_hd__dfrtp_2
X_5919_ _6552_/Q _5702_/X wire656/X _6611_/Q VGND VGND VPWR VPWR _5919_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4250_ _4250_/A _5236_/B VGND VGND VPWR VPWR _4255_/S sky130_fd_sc_hd__nand2_4
XFILLER_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3201_ _6668_/Q VGND VGND VPWR VPWR _3201_/Y sky130_fd_sc_hd__inv_2
X_4181_ _6646_/Q _6409_/A0 _4183_/S VGND VGND VPWR VPWR _6646_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6822_ _7091_/CLK _6822_/D fanout866/X VGND VGND VPWR VPWR _6822_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_51_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3965_ _6473_/Q _3965_/B VGND VGND VPWR VPWR _3965_/X sky130_fd_sc_hd__and2b_4
X_6753_ _7223_/CLK _6753_/D fanout850/X VGND VGND VPWR VPWR _6753_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5704_ _5864_/B _5704_/B _5706_/B VGND VGND VPWR VPWR _5704_/X sky130_fd_sc_hd__and3_4
X_3896_ _6698_/Q _3915_/B VGND VGND VPWR VPWR _3896_/Y sky130_fd_sc_hd__nand2_1
X_6684_ _6992_/CLK _6684_/D fanout868/X VGND VGND VPWR VPWR _6684_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_191_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5635_ _5864_/B _5635_/B VGND VGND VPWR VPWR _5635_/Y sky130_fd_sc_hd__nand2_1
XFILLER_191_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5566_ wire742/X hold392/X _5566_/S VGND VGND VPWR VPWR _5566_/X sky130_fd_sc_hd__mux2_1
Xhold110 _3264_/X VGND VGND VPWR VPWR hold110/X sky130_fd_sc_hd__bufbuf_16
X_5497_ hold38/X hold216/X _5501_/S VGND VGND VPWR VPWR _7062_/D sky130_fd_sc_hd__mux2_1
XFILLER_163_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4517_ _4711_/A _4586_/B VGND VGND VPWR VPWR _4850_/A sky130_fd_sc_hd__and2_2
Xhold121 wire439/X VGND VGND VPWR VPWR _5270_/A sky130_fd_sc_hd__bufbuf_16
XFILLER_132_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold143 wire729/X VGND VGND VPWR VPWR _5459_/B sky130_fd_sc_hd__bufbuf_16
Xhold132 _6784_/Q VGND VGND VPWR VPWR hold132/X sky130_fd_sc_hd__bufbuf_16
X_4448_ _4707_/B _4445_/X _4440_/B VGND VGND VPWR VPWR _4449_/B sky130_fd_sc_hd__o21ai_4
XFILLER_144_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold154 hold154/A VGND VGND VPWR VPWR hold154/X sky130_fd_sc_hd__bufbuf_16
XFILLER_105_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold176 hold86/X VGND VGND VPWR VPWR _3421_/B sky130_fd_sc_hd__bufbuf_16
Xhold165 _6779_/Q VGND VGND VPWR VPWR hold165/X sky130_fd_sc_hd__bufbuf_16
Xhold198 hold55/X VGND VGND VPWR VPWR hold198/X sky130_fd_sc_hd__bufbuf_16
XFILLER_132_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold187 hold94/X VGND VGND VPWR VPWR _3281_/B sky130_fd_sc_hd__bufbuf_16
X_4379_ _4469_/A _5031_/A VGND VGND VPWR VPWR _4986_/B sky130_fd_sc_hd__or2_4
X_7167_ _3949_/A1 _7167_/D fanout879/X VGND VGND VPWR VPWR _7167_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_86_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6118_ _7120_/Q _6023_/D wire579/X _3218_/A _6117_/X VGND VGND VPWR VPWR _6121_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_58_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7098_ _7107_/CLK _7098_/D fanout865/X VGND VGND VPWR VPWR _7098_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6049_ _7061_/Q wire647/X wire618/X _7045_/Q VGND VGND VPWR VPWR _6049_/X sky130_fd_sc_hd__a22o_2
XFILLER_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_82_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6851_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_139_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length622 _6022_/D VGND VGND VPWR VPWR _6191_/B1 sky130_fd_sc_hd__buf_6
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length655 _5706_/X VGND VGND VPWR VPWR _5812_/B1 sky130_fd_sc_hd__buf_6
XFILLER_10_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length688 _5687_/X VGND VGND VPWR VPWR _5923_/B1 sky130_fd_sc_hd__buf_6
XFILLER_108_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_20_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7128_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_49_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_35_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7156_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_33_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3750_ _6619_/Q _4148_/A _4250_/A _6708_/Q VGND VGND VPWR VPWR _3750_/X sky130_fd_sc_hd__a22o_1
XFILLER_20_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3681_ _7038_/Q _5468_/A _5238_/A _6835_/Q VGND VGND VPWR VPWR _3681_/X sky130_fd_sc_hd__a22o_2
XFILLER_145_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5420_ wire757/X hold531/X _5422_/S VGND VGND VPWR VPWR _6994_/D sky130_fd_sc_hd__mux2_1
Xoutput226 _6674_/Q VGND VGND VPWR VPWR mgmt_gpio_out[21] sky130_fd_sc_hd__buf_8
XFILLER_173_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput204 _3932_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[36] sky130_fd_sc_hd__buf_8
X_5351_ _5351_/A _5594_/B VGND VGND VPWR VPWR _5359_/S sky130_fd_sc_hd__nand2_8
XFILLER_154_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput215 _6509_/Q VGND VGND VPWR VPWR mgmt_gpio_out[11] sky130_fd_sc_hd__buf_8
XFILLER_114_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput237 _6521_/Q VGND VGND VPWR VPWR mgmt_gpio_out[31] sky130_fd_sc_hd__buf_8
X_5282_ _5498_/A0 hold718/X _5287_/S VGND VGND VPWR VPWR _6871_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput248 _6688_/Q VGND VGND VPWR VPWR mgmt_gpio_out[7] sky130_fd_sc_hd__buf_8
Xoutput259 _3962_/Y VGND VGND VPWR VPWR pad_flash_io1_ieb sky130_fd_sc_hd__buf_8
X_4302_ _6410_/A0 hold662/X _4303_/S VGND VGND VPWR VPWR _6751_/D sky130_fd_sc_hd__mux2_1
X_7021_ _7103_/CLK _7021_/D fanout861/X VGND VGND VPWR VPWR _7021_/Q sky130_fd_sc_hd__dfstp_4
X_4233_ hold781/X _4232_/X _4235_/S VGND VGND VPWR VPWR _4233_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4164_ hold83/X _6632_/Q _4165_/S VGND VGND VPWR VPWR _4164_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4095_ _6574_/Q wire352/X _4096_/S VGND VGND VPWR VPWR _6574_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_532 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6805_ _6806_/CLK _6805_/D _6435_/A VGND VGND VPWR VPWR _6805_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_24_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4997_ _4997_/A _4997_/B VGND VGND VPWR VPWR _5116_/C sky130_fd_sc_hd__nor2_4
XFILLER_11_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6736_ _6736_/CLK _6736_/D wire860/X VGND VGND VPWR VPWR _6736_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_176_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3948_ _6513_/Q user_clock _6835_/Q VGND VGND VPWR VPWR _3948_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6667_ _3957_/A1 _6667_/D _6446_/X VGND VGND VPWR VPWR _6667_/Q sky130_fd_sc_hd__dfrtp_2
X_3879_ _6485_/Q _6459_/Q _3847_/B VGND VGND VPWR VPWR _3879_/X sky130_fd_sc_hd__a21o_1
XFILLER_164_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6598_ _6642_/CLK _6598_/D fanout856/X VGND VGND VPWR VPWR _6598_/Q sky130_fd_sc_hd__dfrtp_2
X_5618_ _7160_/Q _5616_/A _5617_/A VGND VGND VPWR VPWR _5618_/Y sky130_fd_sc_hd__a21boi_1
X_5549_ _5549_/A _5594_/B VGND VGND VPWR VPWR _5557_/S sky130_fd_sc_hd__and2_4
XFILLER_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7219_ _7220_/CLK _7219_/D _6362_/B VGND VGND VPWR VPWR _7219_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_48_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire843 wire843/A VGND VGND VPWR VPWR wire843/X sky130_fd_sc_hd__buf_6
Xwire821 wire821/A VGND VGND VPWR VPWR _3993_/S sky130_fd_sc_hd__buf_8
Xwire832 _5252_/C VGND VGND VPWR VPWR _6421_/B sky130_fd_sc_hd__buf_8
XFILLER_183_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire898 wire899/X VGND VGND VPWR VPWR _3970_/A sky130_fd_sc_hd__buf_6
XFILLER_108_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A VGND VGND VPWR VPWR _7194_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_69_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4920_ _4920_/A _4920_/B _4920_/C _5047_/A VGND VGND VPWR VPWR _5163_/A sky130_fd_sc_hd__or4_1
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4851_ _4478_/B _4851_/B VGND VGND VPWR VPWR _4989_/B sky130_fd_sc_hd__nand2b_4
XFILLER_60_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3802_ _3802_/A _3802_/B VGND VGND VPWR VPWR _6486_/D sky130_fd_sc_hd__and2_1
XFILLER_159_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4782_ _4775_/A _4990_/A _4756_/B _4745_/A VGND VGND VPWR VPWR _4800_/B sky130_fd_sc_hd__o22ai_2
X_6521_ _7147_/CLK _6521_/D fanout886/X VGND VGND VPWR VPWR _6521_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_158_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3733_ _4241_/A _3733_/B VGND VGND VPWR VPWR _5236_/A sky130_fd_sc_hd__nor2_1
XFILLER_174_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3664_ _3664_/A _3664_/B _3664_/C _3664_/D VGND VGND VPWR VPWR _3665_/C sky130_fd_sc_hd__or4_1
X_6452_ _6455_/A _6455_/B VGND VGND VPWR VPWR _6452_/X sky130_fd_sc_hd__and2_1
XFILLER_161_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5403_ hold317/X _5601_/A0 _5404_/S VGND VGND VPWR VPWR _5403_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6383_ _4236_/B _6383_/A2 _6383_/B1 _4238_/B VGND VGND VPWR VPWR _6383_/X sky130_fd_sc_hd__a22o_1
X_3595_ wire496/X wire430/X _4178_/A _6647_/Q _3558_/X VGND VGND VPWR VPWR _3598_/B
+ sky130_fd_sc_hd__a221o_2
X_5334_ hold580/X hold465/X _5341_/S VGND VGND VPWR VPWR _6917_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5265_ _6856_/Q wire769/X _5269_/S VGND VGND VPWR VPWR _6856_/D sky130_fd_sc_hd__mux2_1
X_7004_ _7152_/CLK _7004_/D fanout882/X VGND VGND VPWR VPWR _7004_/Q sky130_fd_sc_hd__dfrtp_2
X_4216_ hold415/X _4215_/X _4218_/S VGND VGND VPWR VPWR _6675_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5196_ _6408_/A0 hold705/X _5199_/S VGND VGND VPWR VPWR _6801_/D sky130_fd_sc_hd__mux2_1
X_4147_ _5599_/A0 hold316/X _4147_/S VGND VGND VPWR VPWR _6618_/D sky130_fd_sc_hd__mux2_1
XFILLER_18_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4078_ _6559_/Q _6367_/A1 _4081_/S VGND VGND VPWR VPWR _6559_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6719_ _6851_/CLK _6719_/D fanout850/X VGND VGND VPWR VPWR _6719_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire640 wire641/X VGND VGND VPWR VPWR wire640/X sky130_fd_sc_hd__buf_8
XFILLER_128_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire651 wire651/A VGND VGND VPWR VPWR wire651/X sky130_fd_sc_hd__buf_8
XFILLER_183_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire684 _5689_/X VGND VGND VPWR VPWR wire684/X sky130_fd_sc_hd__buf_8
XFILLER_128_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire673 _5694_/X VGND VGND VPWR VPWR wire673/X sky130_fd_sc_hd__buf_6
Xwire662 _5703_/X VGND VGND VPWR VPWR wire662/X sky130_fd_sc_hd__buf_8
Xhold709 _6642_/Q VGND VGND VPWR VPWR hold709/X sky130_fd_sc_hd__bufbuf_16
XFILLER_170_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3380_ _6470_/Q _6666_/Q VGND VGND VPWR VPWR _3928_/A sky130_fd_sc_hd__nand2_8
XFILLER_151_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5050_ _5050_/A _5050_/B _5050_/C VGND VGND VPWR VPWR _5050_/X sky130_fd_sc_hd__or3_1
XFILLER_111_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4001_ _6501_/Q wire753/A _4003_/S VGND VGND VPWR VPWR _6501_/D sky130_fd_sc_hd__mux2_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5952_ _6716_/Q wire702/X _5702_/X _6553_/Q _5951_/X VGND VGND VPWR VPWR _5953_/D
+ sky130_fd_sc_hd__a221o_4
X_4903_ _4903_/A _4936_/C _4903_/C _4878_/A VGND VGND VPWR VPWR _4904_/D sky130_fd_sc_hd__or4b_1
X_5883_ _5883_/A _5883_/B _5883_/C _5883_/D VGND VGND VPWR VPWR _5883_/X sky130_fd_sc_hd__or4_1
XFILLER_61_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4834_ _4834_/A _4834_/B _4834_/C _4834_/D VGND VGND VPWR VPWR _4838_/B sky130_fd_sc_hd__or4_4
XFILLER_147_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4765_ _4563_/X _4645_/X _4764_/X _4239_/X hold93/A VGND VGND VPWR VPWR _6778_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_193_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6504_ _6815_/CLK _6504_/D fanout861/X VGND VGND VPWR VPWR _6504_/Q sky130_fd_sc_hd__dfstp_4
X_3716_ _7006_/Q _5432_/A _3301_/Y _7022_/Q _3715_/X VGND VGND VPWR VPWR _3717_/D
+ sky130_fd_sc_hd__a221o_1
X_4696_ _4696_/A _4696_/B VGND VGND VPWR VPWR _5062_/C sky130_fd_sc_hd__nand2_8
XFILLER_174_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6435_ _6435_/A _6447_/B VGND VGND VPWR VPWR _6435_/X sky130_fd_sc_hd__and2_1
X_3647_ _6807_/Q _5200_/A _5185_/A _6787_/Q _3646_/X VGND VGND VPWR VPWR _3654_/A
+ sky130_fd_sc_hd__a221o_2
X_3578_ _3578_/A _3578_/B _3578_/C _3578_/D VGND VGND VPWR VPWR _3588_/C sky130_fd_sc_hd__or4_1
X_6366_ _7206_/Q _3606_/X _6370_/S VGND VGND VPWR VPWR _7206_/D sky130_fd_sc_hd__mux2_1
X_5317_ wire794/A _6902_/Q _5323_/S VGND VGND VPWR VPWR _6902_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold14 hold14/A VGND VGND VPWR VPWR hold14/X sky130_fd_sc_hd__bufbuf_16
X_6297_ _6745_/Q wire598/X wire610/X wire566/X _6296_/X VGND VGND VPWR VPWR _6306_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold47 hold47/A VGND VGND VPWR VPWR hold47/X sky130_fd_sc_hd__bufbuf_16
Xhold25 hold2/X VGND VGND VPWR VPWR hold25/X sky130_fd_sc_hd__bufbuf_16
Xhold36 hold36/A VGND VGND VPWR VPWR hold36/X sky130_fd_sc_hd__bufbuf_16
XFILLER_152_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5248_ _5248_/A0 hold243/X _5248_/S VGND VGND VPWR VPWR _5248_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold58 hold58/A VGND VGND VPWR VPWR hold58/X sky130_fd_sc_hd__bufbuf_16
XFILLER_130_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5179_ _5023_/A _4988_/A _5164_/B _4757_/B VGND VGND VPWR VPWR _5179_/X sky130_fd_sc_hd__o22a_1
XFILLER_102_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold69 hold69/A VGND VGND VPWR VPWR hold69/X sky130_fd_sc_hd__bufbuf_16
XFILLER_56_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4550_ _4987_/B _4575_/B _4519_/Y _4549_/X VGND VGND VPWR VPWR _4551_/C sky130_fd_sc_hd__a211o_1
XFILLER_190_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold506 _5555_/X VGND VGND VPWR VPWR _7114_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_143_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire470 _7147_/Q VGND VGND VPWR VPWR wire470/X sky130_fd_sc_hd__buf_6
X_4481_ _4558_/B _4663_/A VGND VGND VPWR VPWR _4986_/C sky130_fd_sc_hd__or2_4
XFILLER_128_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire492 _7086_/Q VGND VGND VPWR VPWR wire492/X sky130_fd_sc_hd__buf_6
Xhold517 _7101_/Q VGND VGND VPWR VPWR hold517/X sky130_fd_sc_hd__bufbuf_16
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire481 _7104_/Q VGND VGND VPWR VPWR _3209_/A sky130_fd_sc_hd__buf_8
X_3501_ _3508_/A _3534_/A VGND VGND VPWR VPWR _4178_/A sky130_fd_sc_hd__nor2_4
X_6220_ _7116_/Q wire650/X _6021_/B _7156_/Q VGND VGND VPWR VPWR _6220_/X sky130_fd_sc_hd__a22o_1
XFILLER_144_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3432_ wire556/X _5261_/A _3657_/A2 _7066_/Q _3431_/X VGND VGND VPWR VPWR _3436_/A
+ sky130_fd_sc_hd__a221o_1
Xhold528 _5561_/X VGND VGND VPWR VPWR _7119_/D sky130_fd_sc_hd__bufbuf_16
Xhold539 _6855_/Q VGND VGND VPWR VPWR hold539/X sky130_fd_sc_hd__bufbuf_16
X_6151_ _6873_/Q wire593/X wire591/X _6897_/Q _6150_/X VGND VGND VPWR VPWR _6156_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3363_ _3972_/B _4234_/S _5360_/A _6948_/Q _3360_/X VGND VGND VPWR VPWR _3377_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5102_ _5037_/B _5102_/B _5102_/C _5102_/D VGND VGND VPWR VPWR _5161_/C sky130_fd_sc_hd__and4b_1
XFILLER_112_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _6082_/A _6082_/B _6082_/C _6082_/D VGND VGND VPWR VPWR _6082_/X sky130_fd_sc_hd__or4_1
XFILLER_85_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3294_ _3309_/A _3304_/B VGND VGND VPWR VPWR _3294_/X sky130_fd_sc_hd__or2_4
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _5033_/A _5033_/B _5033_/C _5032_/X VGND VGND VPWR VPWR _5095_/C sky130_fd_sc_hd__or4b_4
XFILLER_97_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6984_ _6986_/CLK _6984_/D fanout879/X VGND VGND VPWR VPWR _6984_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_80_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5935_ wire566/X wire700/X wire686/X _6770_/Q VGND VGND VPWR VPWR _5935_/X sky130_fd_sc_hd__a22o_1
X_5866_ _7012_/Q wire701/X wire694/X _7044_/Q _5865_/X VGND VGND VPWR VPWR _5871_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4817_ _4817_/A _4817_/B _4817_/C _4817_/D VGND VGND VPWR VPWR _4834_/A sky130_fd_sc_hd__or4_1
XFILLER_139_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5797_ _6961_/Q _5673_/X _5681_/X _6921_/Q VGND VGND VPWR VPWR _5797_/X sky130_fd_sc_hd__a22o_1
X_4748_ _4748_/A _4748_/B VGND VGND VPWR VPWR _5123_/B sky130_fd_sc_hd__nand2_2
XFILLER_135_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4679_ _4920_/C _5047_/A _4679_/C VGND VGND VPWR VPWR _4680_/C sky130_fd_sc_hd__or3_1
XFILLER_119_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6418_ _6420_/A _6421_/B VGND VGND VPWR VPWR _6418_/X sky130_fd_sc_hd__and2_1
XFILLER_134_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6349_ _6623_/Q wire623/X wire612/X _6653_/Q VGND VGND VPWR VPWR _6349_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput126 wb_adr_i[5] VGND VGND VPWR VPWR _4665_/A sky130_fd_sc_hd__buf_6
Xinput115 wb_adr_i[24] VGND VGND VPWR VPWR _3887_/C sky130_fd_sc_hd__clkbuf_4
Xinput104 wb_adr_i[14] VGND VGND VPWR VPWR _4350_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput159 wb_dat_i[5] VGND VGND VPWR VPWR _6393_/B1 sky130_fd_sc_hd__clkbuf_4
Xinput137 wb_dat_i[14] VGND VGND VPWR VPWR _6395_/B1 sky130_fd_sc_hd__clkbuf_4
Xinput148 wb_dat_i[24] VGND VGND VPWR VPWR _6378_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3981_ hold50/X hold34/X _3991_/S VGND VGND VPWR VPWR hold51/A sky130_fd_sc_hd__mux2_8
XFILLER_62_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5720_ _5720_/A _5720_/B _5720_/C _5720_/D VGND VGND VPWR VPWR _5720_/X sky130_fd_sc_hd__or4_4
XFILLER_16_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5651_ _7171_/Q _7170_/Q VGND VGND VPWR VPWR _6037_/C sky130_fd_sc_hd__and2b_4
XFILLER_175_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4602_ _4603_/B _4947_/B VGND VGND VPWR VPWR _5069_/A sky130_fd_sc_hd__nor2_1
X_5582_ wire753/X hold827/X _5584_/S VGND VGND VPWR VPWR _7138_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4533_ _4533_/A _4533_/B _4533_/C VGND VGND VPWR VPWR _5147_/A sky130_fd_sc_hd__or3_4
XFILLER_129_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold314 _6697_/Q VGND VGND VPWR VPWR hold314/X sky130_fd_sc_hd__bufbuf_16
Xhold303 _7145_/Q VGND VGND VPWR VPWR hold303/X sky130_fd_sc_hd__bufbuf_16
Xhold325 _6724_/Q VGND VGND VPWR VPWR hold325/X sky130_fd_sc_hd__bufbuf_16
Xhold347 _6888_/Q VGND VGND VPWR VPWR hold347/X sky130_fd_sc_hd__bufbuf_16
X_4464_ _4685_/A _4651_/B VGND VGND VPWR VPWR _4758_/A sky130_fd_sc_hd__nor2_8
Xhold358 _5593_/X VGND VGND VPWR VPWR _7148_/D sky130_fd_sc_hd__bufbuf_16
Xhold369 _6916_/Q VGND VGND VPWR VPWR hold369/X sky130_fd_sc_hd__bufbuf_16
XFILLER_132_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold336 _6549_/Q VGND VGND VPWR VPWR hold336/X sky130_fd_sc_hd__bufbuf_16
X_6203_ wire553/X _6025_/D wire618/A _7051_/Q _6202_/X VGND VGND VPWR VPWR _6206_/C
+ sky130_fd_sc_hd__a221o_4
X_4395_ _4818_/A _4672_/A _4469_/A _4395_/D VGND VGND VPWR VPWR _4711_/A sky130_fd_sc_hd__and4_4
Xfanout805 hold514/X VGND VGND VPWR VPWR hold465/A sky130_fd_sc_hd__buf_8
XFILLER_131_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3415_ _3415_/A _3415_/B _3415_/C _3415_/D VGND VGND VPWR VPWR _3415_/X sky130_fd_sc_hd__or4_2
X_7183_ _7196_/CLK _7183_/D fanout870/X VGND VGND VPWR VPWR _7183_/Q sky130_fd_sc_hd__dfrtp_2
X_6134_ _5611_/A _7191_/Q wire381/A _6133_/X VGND VGND VPWR VPWR _6134_/X sky130_fd_sc_hd__a211o_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout849 _6447_/A VGND VGND VPWR VPWR _6455_/A sky130_fd_sc_hd__buf_8
X_3346_ _3552_/B _3375_/B VGND VGND VPWR VPWR _3346_/Y sky130_fd_sc_hd__nor2_8
XFILLER_100_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065_ _7022_/Q wire589/X wire615/X _7086_/Q _6064_/X VGND VGND VPWR VPWR _6071_/A
+ sky130_fd_sc_hd__a221o_2
X_5016_ _5016_/A _5156_/B _5016_/C _5015_/X VGND VGND VPWR VPWR _5018_/C sky130_fd_sc_hd__or4b_4
XFILLER_100_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3277_ _3953_/A hold125/X hold133/X VGND VGND VPWR VPWR _3277_/Y sky130_fd_sc_hd__o21bai_4
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_209 wire515/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6967_ _7145_/CLK _6967_/D fanout881/X VGND VGND VPWR VPWR _6967_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5918_ _7185_/Q _6309_/S _5917_/X VGND VGND VPWR VPWR _7185_/D sky130_fd_sc_hd__o21a_1
X_6898_ _7147_/CLK _6898_/D fanout887/X VGND VGND VPWR VPWR _6898_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_139_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5849_ _5849_/A _5849_/B _5849_/C _5849_/D VGND VGND VPWR VPWR _5849_/X sky130_fd_sc_hd__or4_2
XFILLER_108_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3200_ _6679_/Q VGND VGND VPWR VPWR _5663_/B sky130_fd_sc_hd__inv_4
X_4180_ hold536/X wire790/X _4183_/S VGND VGND VPWR VPWR _6645_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6821_ _7091_/CLK _6821_/D fanout866/X VGND VGND VPWR VPWR _6821_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6752_ _6752_/CLK _6752_/D fanout857/X VGND VGND VPWR VPWR _6752_/Q sky130_fd_sc_hd__dfrtp_2
X_3964_ _6474_/Q _3964_/B VGND VGND VPWR VPWR _3964_/X sky130_fd_sc_hd__and2b_4
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3895_ _3895_/A _3895_/B _3895_/C _3895_/D VGND VGND VPWR VPWR _3895_/Y sky130_fd_sc_hd__nor4_4
XFILLER_176_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5703_ _5864_/B _5703_/B _5704_/B VGND VGND VPWR VPWR _5703_/X sky130_fd_sc_hd__and3_4
X_6683_ _6992_/CLK _6683_/D fanout868/X VGND VGND VPWR VPWR _6683_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_136_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5634_ _7164_/Q _5635_/B _5633_/B _5636_/S VGND VGND VPWR VPWR _7164_/D sky130_fd_sc_hd__a31o_1
XFILLER_31_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold100 _3262_/X VGND VGND VPWR VPWR hold42/A sky130_fd_sc_hd__bufbuf_16
X_5565_ wire749/X hold420/X _5565_/S VGND VGND VPWR VPWR _5565_/X sky130_fd_sc_hd__mux2_1
Xhold122 _5270_/Y VGND VGND VPWR VPWR _5278_/S sky130_fd_sc_hd__bufbuf_16
Xhold144 _5297_/Y VGND VGND VPWR VPWR _5305_/S sky130_fd_sc_hd__bufbuf_16
XFILLER_144_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4516_ _4871_/A _4636_/A VGND VGND VPWR VPWR _5136_/A sky130_fd_sc_hd__nor2_4
Xhold111 _3266_/Y VGND VGND VPWR VPWR _3284_/B sky130_fd_sc_hd__bufbuf_16
X_5496_ _5532_/A0 _7061_/Q _5502_/S VGND VGND VPWR VPWR _7061_/D sky130_fd_sc_hd__mux2_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold133 _3258_/X VGND VGND VPWR VPWR hold133/X sky130_fd_sc_hd__bufbuf_16
X_4447_ _4696_/A _4446_/B _4445_/X _4707_/B VGND VGND VPWR VPWR _4510_/B sky130_fd_sc_hd__o2bb2a_1
Xhold155 hold155/A VGND VGND VPWR VPWR wire763/A sky130_fd_sc_hd__bufbuf_16
Xhold166 _3269_/X VGND VGND VPWR VPWR hold61/A sky130_fd_sc_hd__bufbuf_16
Xhold177 _3543_/B VGND VGND VPWR VPWR _3493_/B sky130_fd_sc_hd__bufbuf_16
Xhold199 hold199/A VGND VGND VPWR VPWR hold56/A sky130_fd_sc_hd__bufbuf_16
X_7166_ _3949_/A1 _7166_/D fanout879/X VGND VGND VPWR VPWR _7166_/Q sky130_fd_sc_hd__dfstp_4
Xhold188 _4086_/X VGND VGND VPWR VPWR _6566_/D sky130_fd_sc_hd__bufbuf_16
X_4378_ _4469_/A _5031_/A VGND VGND VPWR VPWR _4987_/B sky130_fd_sc_hd__nor2_8
X_6117_ wire522/A wire604/X _6022_/D _6920_/Q VGND VGND VPWR VPWR _6117_/X sky130_fd_sc_hd__a22o_1
XFILLER_86_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_1_csclk _6744_/CLK VGND VGND VPWR VPWR _6752_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7097_ _7133_/CLK _7097_/D fanout883/X VGND VGND VPWR VPWR _7097_/Q sky130_fd_sc_hd__dfrtp_2
X_3329_ _4241_/A hold45/X VGND VGND VPWR VPWR hold46/A sky130_fd_sc_hd__nor2_8
XFILLER_100_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6048_ _6885_/Q wire602/X wire581/X _7141_/Q _6047_/X VGND VGND VPWR VPWR _6058_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_100_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_0_0_mgmt_gpio_in[4] clkbuf_2_1_0_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR _3957_/A1
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_134_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3680_ _6958_/Q _5378_/A _3739_/B1 _6982_/Q VGND VGND VPWR VPWR _3680_/X sky130_fd_sc_hd__a22o_4
XFILLER_118_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput205 _3931_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[37] sky130_fd_sc_hd__buf_8
XFILLER_160_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5350_ _5602_/A0 hold375/X _5350_/S VGND VGND VPWR VPWR _5350_/X sky130_fd_sc_hd__mux2_1
Xoutput216 _6510_/Q VGND VGND VPWR VPWR mgmt_gpio_out[12] sky130_fd_sc_hd__buf_8
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput227 _6675_/Q VGND VGND VPWR VPWR mgmt_gpio_out[22] sky130_fd_sc_hd__buf_8
Xoutput238 wire464/X VGND VGND VPWR VPWR mgmt_gpio_out[32] sky130_fd_sc_hd__buf_8
X_5281_ wire794/A _6870_/Q _5287_/S VGND VGND VPWR VPWR _6870_/D sky130_fd_sc_hd__mux2_1
XFILLER_153_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput249 _3939_/X VGND VGND VPWR VPWR mgmt_gpio_out[8] sky130_fd_sc_hd__buf_8
XFILLER_5_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4301_ _6409_/A0 hold830/X _4303_/S VGND VGND VPWR VPWR _6750_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7020_ _7132_/CLK _7020_/D fanout868/X VGND VGND VPWR VPWR _7020_/Q sky130_fd_sc_hd__dfrtp_2
X_4232_ hold631/X _5259_/A0 _4232_/S VGND VGND VPWR VPWR _4232_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4163_ _5408_/A1 hold699/X _4165_/S VGND VGND VPWR VPWR _6631_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4094_ _6573_/Q wire351/X _4096_/S VGND VGND VPWR VPWR _6573_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4996_ _4996_/A _4997_/B VGND VGND VPWR VPWR _5136_/D sky130_fd_sc_hd__nor2_1
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6804_ _6806_/CLK _6804_/D _6435_/A VGND VGND VPWR VPWR _6804_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6735_ _6950_/CLK _6735_/D fanout875/X VGND VGND VPWR VPWR _6735_/Q sky130_fd_sc_hd__dfstp_4
X_3947_ _3239_/Y input2/X input1/X VGND VGND VPWR VPWR _3947_/X sky130_fd_sc_hd__mux2_4
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6666_ _3957_/A1 _6666_/D _6445_/X VGND VGND VPWR VPWR _6666_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_31_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3878_ _6455_/A _6455_/B VGND VGND VPWR VPWR _3878_/X sky130_fd_sc_hd__and2_1
XFILLER_137_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6597_ _6642_/CLK _6597_/D fanout856/X VGND VGND VPWR VPWR _6597_/Q sky130_fd_sc_hd__dfrtp_2
X_5617_ _5617_/A _5617_/B _5617_/C VGND VGND VPWR VPWR _7159_/D sky130_fd_sc_hd__and3_1
XFILLER_155_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5548_ wire739/X hold658/X _5548_/S VGND VGND VPWR VPWR _7108_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7218_ _7218_/CLK _7218_/D wire915/X VGND VGND VPWR VPWR _7218_/Q sky130_fd_sc_hd__dfrtp_4
X_5479_ _7046_/Q _5578_/A0 _5485_/S VGND VGND VPWR VPWR _7046_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7149_ _7151_/CLK _7149_/D fanout880/X VGND VGND VPWR VPWR _7149_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_101_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire833 wire833/A VGND VGND VPWR VPWR wire833/X sky130_fd_sc_hd__buf_6
XFILLER_128_616 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire811 _6109_/S VGND VGND VPWR VPWR _6308_/S sky130_fd_sc_hd__buf_8
Xmax_length420 hold46/A VGND VGND VPWR VPWR _3736_/A2 sky130_fd_sc_hd__buf_8
XFILLER_127_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire844 wire844/A VGND VGND VPWR VPWR wire844/X sky130_fd_sc_hd__buf_6
XFILLER_182_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire899 wire899/A VGND VGND VPWR VPWR wire899/X sky130_fd_sc_hd__buf_8
XFILLER_129_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length497 _7064_/Q VGND VGND VPWR VPWR _3214_/A sky130_fd_sc_hd__buf_6
XFILLER_163_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4850_ _4850_/A _4850_/B VGND VGND VPWR VPWR _4850_/X sky130_fd_sc_hd__or2_4
XFILLER_33_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3801_ _6486_/Q _3801_/B VGND VGND VPWR VPWR _3802_/B sky130_fd_sc_hd__or2_1
XFILLER_60_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6520_ _7147_/CLK _6520_/D fanout886/X VGND VGND VPWR VPWR _6520_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_158_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4781_ _4622_/B _4772_/A _5178_/A VGND VGND VPWR VPWR _4800_/A sky130_fd_sc_hd__a21o_1
XFILLER_119_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3732_ _5225_/A _3732_/B VGND VGND VPWR VPWR _5216_/A sky130_fd_sc_hd__nor2_1
XFILLER_173_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6451_ _6455_/A _6455_/B VGND VGND VPWR VPWR _6451_/X sky130_fd_sc_hd__and2_1
X_3663_ _3726_/A _3663_/B _3663_/C _3663_/D VGND VGND VPWR VPWR _3664_/D sky130_fd_sc_hd__or4_1
X_6382_ _6381_/X hold34/A _6400_/S VGND VGND VPWR VPWR _7212_/D sky130_fd_sc_hd__mux2_1
X_5402_ hold457/X _5600_/A0 _5404_/S VGND VGND VPWR VPWR _5402_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5333_ _5333_/A _5594_/B VGND VGND VPWR VPWR _5341_/S sky130_fd_sc_hd__and2_4
X_3594_ _6491_/Q _3978_/A _4298_/A _6751_/Q _3557_/X VGND VGND VPWR VPWR _3598_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_126_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5264_ hold539/X wire780/A _5269_/S VGND VGND VPWR VPWR _6855_/D sky130_fd_sc_hd__mux2_1
X_7003_ _7154_/CLK _7003_/D fanout886/X VGND VGND VPWR VPWR _7003_/Q sky130_fd_sc_hd__dfrtp_2
X_4215_ hold232/X _5601_/A0 hold46/X VGND VGND VPWR VPWR _4215_/X sky130_fd_sc_hd__mux2_1
X_5195_ _6407_/A0 hold752/X _5199_/S VGND VGND VPWR VPWR _6800_/D sky130_fd_sc_hd__mux2_1
X_4146_ hold83/X hold219/X _4147_/S VGND VGND VPWR VPWR _4146_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_81_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7223_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_141_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4077_ _6558_/Q _3606_/X _4081_/S VGND VGND VPWR VPWR _6558_/D sky130_fd_sc_hd__mux2_1
XFILLER_43_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4979_ _4913_/B _4977_/X _5060_/B VGND VGND VPWR VPWR _4979_/X sky130_fd_sc_hd__o21ba_1
X_6718_ _6842_/CLK _6718_/D fanout857/X VGND VGND VPWR VPWR _6718_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6649_ _6650_/CLK _6649_/D fanout858/X VGND VGND VPWR VPWR _6649_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_137_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_34_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7152_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_164_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_49_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7136_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_74_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire641 _6023_/B VGND VGND VPWR VPWR wire641/X sky130_fd_sc_hd__buf_8
Xwire630 wire631/X VGND VGND VPWR VPWR wire630/X sky130_fd_sc_hd__buf_8
XFILLER_143_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire674 _5694_/X VGND VGND VPWR VPWR wire674/X sky130_fd_sc_hd__buf_6
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4000_ _6500_/Q _6411_/A0 _4003_/S VGND VGND VPWR VPWR _6500_/D sky130_fd_sc_hd__mux2_1
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5951_ _6662_/Q _5974_/A2 wire671/X _5942_/X VGND VGND VPWR VPWR _5951_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_1_0_1_mgmt_gpio_in[4] clkbuf_1_0_1_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR clkbuf_2_1_0_mgmt_gpio_in[4]/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_53_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4902_ _4581_/A _4536_/X _4962_/A _4886_/Y VGND VGND VPWR VPWR _4904_/C sky130_fd_sc_hd__a211o_1
XFILLER_80_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5882_ _6594_/Q _5681_/X _5923_/B1 _6639_/Q _5881_/X VGND VGND VPWR VPWR _5883_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_178_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4833_ _4697_/A _5005_/C _4832_/X VGND VGND VPWR VPWR _4834_/D sky130_fd_sc_hd__a21oi_1
XFILLER_61_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4764_ _5003_/B _4763_/X _5156_/A _4720_/X VGND VGND VPWR VPWR _4764_/X sky130_fd_sc_hd__a211o_2
XFILLER_60_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6503_ _6771_/CLK _6503_/D fanout853/X VGND VGND VPWR VPWR _6503_/Q sky130_fd_sc_hd__dfstp_4
X_3715_ wire502/X _3298_/Y _5218_/A _6821_/Q VGND VGND VPWR VPWR _3715_/X sky130_fd_sc_hd__a22o_1
X_4695_ _4696_/A _4696_/B VGND VGND VPWR VPWR _4695_/X sky130_fd_sc_hd__and2_4
X_6434_ _6446_/A _6455_/B VGND VGND VPWR VPWR _6434_/X sky130_fd_sc_hd__and2_1
XFILLER_161_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3646_ _7223_/Q _6406_/A _5194_/A _6802_/Q VGND VGND VPWR VPWR _3646_/X sky130_fd_sc_hd__a22o_1
X_3577_ wire550/X _3374_/Y _4061_/A _6548_/Q _3576_/X VGND VGND VPWR VPWR _3578_/D
+ sky130_fd_sc_hd__a221o_2
X_6365_ _7205_/Q _3665_/X _6370_/S VGND VGND VPWR VPWR _7205_/D sky130_fd_sc_hd__mux2_1
X_5316_ _5595_/A0 _6901_/Q _5323_/S VGND VGND VPWR VPWR _6901_/D sky130_fd_sc_hd__mux2_1
X_6296_ _6552_/Q wire602/X wire581/X _6631_/Q _6295_/X VGND VGND VPWR VPWR _6296_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5247_ _5247_/A0 hold537/X _5249_/S VGND VGND VPWR VPWR _5247_/X sky130_fd_sc_hd__mux2_1
Xhold26 hold26/A VGND VGND VPWR VPWR hold3/A sky130_fd_sc_hd__bufbuf_16
Xhold15 hold49/X VGND VGND VPWR VPWR hold50/A sky130_fd_sc_hd__bufbuf_16
Xhold37 hold37/A VGND VGND VPWR VPWR hold37/X sky130_fd_sc_hd__bufbuf_16
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold48 hold48/A VGND VGND VPWR VPWR hold48/X sky130_fd_sc_hd__bufbuf_16
X_5178_ _5178_/A _5178_/B _5178_/C _5178_/D VGND VGND VPWR VPWR _5178_/X sky130_fd_sc_hd__or4_4
XFILLER_68_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold59 hold59/A VGND VGND VPWR VPWR hold59/X sky130_fd_sc_hd__bufbuf_16
XFILLER_29_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4129_ hold306/X _5599_/A0 _4129_/S VGND VGND VPWR VPWR _6603_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire460 wire461/X VGND VGND VPWR VPWR wire460/X sky130_fd_sc_hd__buf_6
X_3500_ _3508_/A hold44/X VGND VGND VPWR VPWR _4166_/A sky130_fd_sc_hd__nor2_8
Xwire471 _7144_/Q VGND VGND VPWR VPWR _3204_/A sky130_fd_sc_hd__buf_8
XFILLER_183_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold507 _6882_/Q VGND VGND VPWR VPWR hold507/X sky130_fd_sc_hd__bufbuf_16
XFILLER_156_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4480_ _4558_/B _4663_/A VGND VGND VPWR VPWR _4992_/B sky130_fd_sc_hd__nor2_2
XFILLER_144_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire482 _7103_/Q VGND VGND VPWR VPWR wire482/X sky130_fd_sc_hd__buf_6
Xwire493 _7085_/Q VGND VGND VPWR VPWR wire493/X sky130_fd_sc_hd__buf_6
Xhold518 _7017_/Q VGND VGND VPWR VPWR hold518/X sky130_fd_sc_hd__bufbuf_16
X_3431_ _6866_/Q wire439/X _5245_/A wire897/A VGND VGND VPWR VPWR _3431_/X sky130_fd_sc_hd__a22o_4
XFILLER_183_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold529 _7049_/Q VGND VGND VPWR VPWR hold529/X sky130_fd_sc_hd__bufbuf_16
X_6150_ _6961_/Q wire624/X wire613/X wire500/X VGND VGND VPWR VPWR _6150_/X sky130_fd_sc_hd__a22o_1
X_3362_ _3365_/A _3369_/A VGND VGND VPWR VPWR _5360_/A sky130_fd_sc_hd__nor2_8
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _5101_/A _5101_/B _5101_/C _5101_/D VGND VGND VPWR VPWR _5101_/X sky130_fd_sc_hd__or4_1
XFILLER_111_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _7062_/Q wire648/X wire633/X _6910_/Q _6080_/X VGND VGND VPWR VPWR _6082_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_85_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3293_ _3278_/B _3293_/B VGND VGND VPWR VPWR _3293_/Y sky130_fd_sc_hd__nand2b_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _5023_/A _4997_/A _5164_/B _4754_/B _4767_/X VGND VGND VPWR VPWR _5032_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_66_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6983_ _7081_/CLK _6983_/D fanout878/X VGND VGND VPWR VPWR _6983_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_80_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5934_ _6621_/Q wire707/X _5934_/B1 _6547_/Q _5933_/X VGND VGND VPWR VPWR _5937_/C
+ sky130_fd_sc_hd__a221o_4
XFILLER_15_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5865_ _6948_/Q wire656/A _5864_/X _5698_/B VGND VGND VPWR VPWR _5865_/X sky130_fd_sc_hd__a22o_2
X_4816_ _4687_/A _4832_/B _4729_/X VGND VGND VPWR VPWR _4817_/D sky130_fd_sc_hd__o21bai_1
XFILLER_193_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5796_ _5796_/A _5796_/B _5796_/C _5796_/D VGND VGND VPWR VPWR _5796_/X sky130_fd_sc_hd__or4_2
XFILLER_31_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4747_ _4728_/X _4735_/X _4746_/X _4740_/B _4745_/X VGND VGND VPWR VPWR _4753_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_147_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4678_ _4832_/C _4746_/B _4663_/B VGND VGND VPWR VPWR _4679_/C sky130_fd_sc_hd__a21oi_1
XFILLER_119_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6417_ _6420_/A _6421_/B VGND VGND VPWR VPWR _6417_/X sky130_fd_sc_hd__and2_1
XFILLER_162_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3629_ _3629_/A _3629_/B _3629_/C _3629_/D VGND VGND VPWR VPWR _3636_/C sky130_fd_sc_hd__or4_1
XFILLER_135_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6348_ _6580_/Q wire599/X wire645/X _6608_/Q _6347_/X VGND VGND VPWR VPWR _6355_/A
+ sky130_fd_sc_hd__a221o_1
Xinput127 wb_adr_i[6] VGND VGND VPWR VPWR _4654_/A sky130_fd_sc_hd__buf_8
Xinput116 wb_adr_i[25] VGND VGND VPWR VPWR input116/X sky130_fd_sc_hd__clkbuf_4
Xinput105 wb_adr_i[15] VGND VGND VPWR VPWR _4350_/C sky130_fd_sc_hd__clkbuf_4
X_6279_ _6660_/Q wire647/X wire632/X _6590_/Q VGND VGND VPWR VPWR _6279_/X sky130_fd_sc_hd__a22o_1
Xinput149 wb_dat_i[25] VGND VGND VPWR VPWR _6380_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput138 wb_dat_i[15] VGND VGND VPWR VPWR _6398_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_56_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3980_ hold746/X _5234_/C _3994_/S VGND VGND VPWR VPWR _6488_/D sky130_fd_sc_hd__mux2_1
XFILLER_62_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5650_ _5645_/Y _5649_/Y _5654_/B VGND VGND VPWR VPWR _7170_/D sky130_fd_sc_hd__a21oi_1
XFILLER_31_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4601_ _4603_/B _4965_/B VGND VGND VPWR VPWR _4642_/A sky130_fd_sc_hd__nor2_1
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5581_ wire763/X hold427/X _5581_/S VGND VGND VPWR VPWR _5581_/X sky130_fd_sc_hd__mux2_1
X_4532_ _4533_/A _4533_/B _4533_/C VGND VGND VPWR VPWR _4949_/C sky130_fd_sc_hd__nor3_4
XFILLER_190_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold315 _4249_/X VGND VGND VPWR VPWR _6697_/D sky130_fd_sc_hd__bufbuf_16
Xhold304 _5590_/X VGND VGND VPWR VPWR _7145_/D sky130_fd_sc_hd__bufbuf_16
X_4463_ _4654_/A _4958_/A VGND VGND VPWR VPWR _4651_/B sky130_fd_sc_hd__or2_4
XFILLER_144_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold326 _4270_/X VGND VGND VPWR VPWR _6724_/D sky130_fd_sc_hd__bufbuf_16
Xhold348 _5301_/X VGND VGND VPWR VPWR _6888_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_116_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6202_ _7107_/Q _5653_/X _6022_/B _6947_/Q VGND VGND VPWR VPWR _6202_/X sky130_fd_sc_hd__a22o_1
X_3414_ _3414_/A _3414_/B _3414_/C _3414_/D VGND VGND VPWR VPWR _3415_/D sky130_fd_sc_hd__or4_1
Xhold359 _7031_/Q VGND VGND VPWR VPWR hold359/X sky130_fd_sc_hd__bufbuf_16
Xhold337 _6484_/Q VGND VGND VPWR VPWR _3255_/B sky130_fd_sc_hd__bufbuf_16
X_4394_ _5031_/A _4663_/A VGND VGND VPWR VPWR _4775_/A sky130_fd_sc_hd__or2_4
X_7182_ _7196_/CLK _7182_/D fanout870/X VGND VGND VPWR VPWR _7182_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_131_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6133_ _6856_/Q _6060_/B _6121_/X _6132_/X _3197_/Y VGND VGND VPWR VPWR _6133_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_97_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout828 _6455_/B VGND VGND VPWR VPWR _6447_/B sky130_fd_sc_hd__buf_8
X_3345_ _7100_/Q _5531_/A _3995_/A _6503_/Q _3340_/X VGND VGND VPWR VPWR _3378_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_100_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6064_ _7134_/Q wire642/X _6212_/B1 _7094_/Q VGND VGND VPWR VPWR _6064_/X sky130_fd_sc_hd__a22o_1
X_3276_ _3365_/A _3508_/A VGND VGND VPWR VPWR _5504_/A sky130_fd_sc_hd__nor2_8
X_5015_ _4754_/B _4832_/C _5050_/B _4746_/X _5050_/C VGND VGND VPWR VPWR _5015_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_100_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6966_ _7153_/CLK _6966_/D fanout881/X VGND VGND VPWR VPWR _6966_/Q sky130_fd_sc_hd__dfstp_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5917_ wire824/X _7184_/Q wire381/X _5916_/X VGND VGND VPWR VPWR _5917_/X sky130_fd_sc_hd__a211o_1
XFILLER_53_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6897_ _7133_/CLK _6897_/D fanout882/X VGND VGND VPWR VPWR _6897_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_167_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5848_ wire526/X _5676_/X wire692/A _6995_/Q _5847_/X VGND VGND VPWR VPWR _5849_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_182_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5779_ _6904_/Q _5814_/A2 _5767_/X _5778_/X VGND VGND VPWR VPWR _5784_/A sky130_fd_sc_hd__a211o_4
XFILLER_139_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6820_ _7091_/CLK _6820_/D fanout866/X VGND VGND VPWR VPWR _6820_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3963_ wire842/X _3875_/B _6474_/Q VGND VGND VPWR VPWR _3963_/X sky130_fd_sc_hd__mux2_8
X_6751_ _7225_/CLK _6751_/D fanout851/X VGND VGND VPWR VPWR _6751_/Q sky130_fd_sc_hd__dfrtp_2
X_3894_ _4346_/S _4722_/B _3894_/C _3894_/D VGND VGND VPWR VPWR _3895_/D sky130_fd_sc_hd__or4_4
X_5702_ _5864_/B _5702_/B _5707_/C VGND VGND VPWR VPWR _5702_/X sky130_fd_sc_hd__and3_4
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_1_1_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
X_6682_ _7223_/CLK _6682_/D _6455_/A VGND VGND VPWR VPWR _6682_/Q sky130_fd_sc_hd__dfrtp_1
X_5633_ _7164_/Q _5633_/B VGND VGND VPWR VPWR _5636_/S sky130_fd_sc_hd__nor2_1
XFILLER_176_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5564_ _5600_/A0 hold480/X _5564_/S VGND VGND VPWR VPWR _5564_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4515_ _4996_/A _4871_/A VGND VGND VPWR VPWR _5078_/A sky130_fd_sc_hd__nor2_4
Xhold101 hold42/X VGND VGND VPWR VPWR _3421_/A sky130_fd_sc_hd__bufbuf_16
XFILLER_8_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold123 _5276_/X VGND VGND VPWR VPWR _6866_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_144_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold112 _3267_/Y VGND VGND VPWR VPWR _3367_/A sky130_fd_sc_hd__bufbuf_16
X_5495_ _5495_/A _5576_/B VGND VGND VPWR VPWR _5502_/S sky130_fd_sc_hd__nand2_4
Xhold134 _3259_/Y VGND VGND VPWR VPWR _3309_/B sky130_fd_sc_hd__bufbuf_16
X_4446_ _5050_/A _4446_/B VGND VGND VPWR VPWR _4534_/B sky130_fd_sc_hd__xnor2_4
Xhold145 _5303_/X VGND VGND VPWR VPWR _6890_/D sky130_fd_sc_hd__bufbuf_16
Xhold156 wire763/X VGND VGND VPWR VPWR hold156/X sky130_fd_sc_hd__bufbuf_16
Xhold167 hold61/X VGND VGND VPWR VPWR _3281_/A sky130_fd_sc_hd__bufbuf_16
XFILLER_144_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4377_ _4818_/A _4672_/A VGND VGND VPWR VPWR _5031_/A sky130_fd_sc_hd__nand2_8
X_7165_ _3949_/A1 _7165_/D fanout879/X VGND VGND VPWR VPWR _7165_/Q sky130_fd_sc_hd__dfstp_4
Xhold178 _4134_/X VGND VGND VPWR VPWR _6607_/D sky130_fd_sc_hd__bufbuf_16
Xhold189 _6783_/Q VGND VGND VPWR VPWR hold189/X sky130_fd_sc_hd__bufbuf_16
X_6116_ _3220_/A _6139_/A2 _6139_/B1 _3217_/A _6111_/X VGND VGND VPWR VPWR _6121_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_86_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3328_ _3383_/C hold43/X VGND VGND VPWR VPWR hold44/A sky130_fd_sc_hd__or2_4
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7096_ _7096_/CLK _7096_/D fanout883/X VGND VGND VPWR VPWR _7096_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_112_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6047_ _7077_/Q _6111_/B _6139_/B1 wire509/X _6046_/X VGND VGND VPWR VPWR _6047_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_100_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3259_ _3953_/A hold125/X hold133/X VGND VGND VPWR VPWR _3259_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_27_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6949_ _6950_/CLK _6949_/D fanout875/X VGND VGND VPWR VPWR _6949_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length668 _5700_/X VGND VGND VPWR VPWR wire667/A sky130_fd_sc_hd__buf_6
XFILLER_108_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold690 _6759_/Q VGND VGND VPWR VPWR hold690/X sky130_fd_sc_hd__bufbuf_16
XFILLER_150_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput217 _3950_/X VGND VGND VPWR VPWR mgmt_gpio_out[13] sky130_fd_sc_hd__buf_8
XFILLER_126_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput206 _3194_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[3] sky130_fd_sc_hd__buf_8
Xoutput228 _6676_/Q VGND VGND VPWR VPWR mgmt_gpio_out[23] sky130_fd_sc_hd__buf_8
Xoutput239 wire462/X VGND VGND VPWR VPWR mgmt_gpio_out[33] sky130_fd_sc_hd__buf_8
X_5280_ _5595_/A0 _6869_/Q _5287_/S VGND VGND VPWR VPWR _6869_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4300_ _6408_/A0 hold694/X _4303_/S VGND VGND VPWR VPWR _6749_/D sky130_fd_sc_hd__mux2_1
XFILLER_153_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4231_ hold680/X _4230_/X _4235_/S VGND VGND VPWR VPWR _4231_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4162_ wire790/A hold319/X _4165_/S VGND VGND VPWR VPWR _4162_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4093_ _6572_/Q _6367_/A1 _4096_/S VGND VGND VPWR VPWR _6572_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4995_ _4995_/A _4997_/B VGND VGND VPWR VPWR _5078_/C sky130_fd_sc_hd__nor2_1
X_6803_ _6806_/CLK _6803_/D _6435_/A VGND VGND VPWR VPWR _6803_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3946_ _3238_/Y _6458_/Q _5252_/C VGND VGND VPWR VPWR _3946_/X sky130_fd_sc_hd__mux2_8
X_6734_ _6736_/CLK _6734_/D wire860/X VGND VGND VPWR VPWR _6734_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3877_ _6833_/Q _6880_/Q _3877_/C VGND VGND VPWR VPWR _3877_/Y sky130_fd_sc_hd__nor3_4
X_6665_ _3957_/A1 _6665_/D _6444_/X VGND VGND VPWR VPWR _6665_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5616_ _5616_/A VGND VGND VPWR VPWR _5617_/C sky130_fd_sc_hd__inv_2
X_6596_ _6642_/CLK _6596_/D fanout856/X VGND VGND VPWR VPWR _6596_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_145_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5547_ _5547_/A0 hold820/X _5548_/S VGND VGND VPWR VPWR _7107_/D sky130_fd_sc_hd__mux2_1
XFILLER_155_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5478_ _7045_/Q wire802/X _5485_/S VGND VGND VPWR VPWR _7045_/D sky130_fd_sc_hd__mux2_1
X_7217_ _7218_/CLK _7217_/D wire915/X VGND VGND VPWR VPWR _7217_/Q sky130_fd_sc_hd__dfrtp_4
X_4429_ _4507_/A _4851_/B _4499_/C VGND VGND VPWR VPWR _4581_/B sky130_fd_sc_hd__and3_4
XFILLER_160_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7148_ _7156_/CLK _7148_/D fanout889/X VGND VGND VPWR VPWR _7148_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_101_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7079_ _7119_/CLK _7079_/D fanout869/X VGND VGND VPWR VPWR _7079_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_104_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire834 wire834/A VGND VGND VPWR VPWR wire834/X sky130_fd_sc_hd__buf_6
XFILLER_128_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire812 _3921_/A VGND VGND VPWR VPWR _6109_/S sky130_fd_sc_hd__buf_8
Xwire845 wire845/A VGND VGND VPWR VPWR _3932_/S sky130_fd_sc_hd__buf_8
XFILLER_10_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length454 _3355_/B VGND VGND VPWR VPWR _3672_/A sky130_fd_sc_hd__buf_8
XFILLER_89_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4780_ _4772_/A _4586_/B _4748_/B _4453_/Y VGND VGND VPWR VPWR _4799_/B sky130_fd_sc_hd__a22o_1
X_3800_ _6487_/Q _3802_/A VGND VGND VPWR VPWR _6487_/D sky130_fd_sc_hd__xnor2_1
XFILLER_21_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3731_ _5225_/A hold44/X VGND VGND VPWR VPWR _5223_/A sky130_fd_sc_hd__nor2_2
XFILLER_186_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_0_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7225_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_173_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6450_ _6455_/A _6455_/B VGND VGND VPWR VPWR _6450_/X sky130_fd_sc_hd__and2_1
X_3662_ _6999_/Q _5423_/A _4322_/A _6770_/Q VGND VGND VPWR VPWR _3663_/D sky130_fd_sc_hd__a22o_1
X_6381_ _4236_/B _6381_/A2 _6381_/B1 _4238_/B _6380_/X VGND VGND VPWR VPWR _6381_/X
+ sky130_fd_sc_hd__a221o_1
X_5401_ hold267/X hold150/X _5404_/S VGND VGND VPWR VPWR _6977_/D sky130_fd_sc_hd__mux2_1
X_3593_ _3593_/A _3593_/B _3593_/C _3593_/D VGND VGND VPWR VPWR _3606_/B sky130_fd_sc_hd__or4_2
X_5332_ _5602_/A0 hold369/X _5332_/S VGND VGND VPWR VPWR _6916_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5263_ hold467/X _5578_/A0 _5269_/S VGND VGND VPWR VPWR _6854_/D sky130_fd_sc_hd__mux2_1
X_4214_ hold851/X hold47/X _4218_/S VGND VGND VPWR VPWR hold48/A sky130_fd_sc_hd__mux2_1
X_7002_ _7042_/CLK _7002_/D fanout865/X VGND VGND VPWR VPWR _7002_/Q sky130_fd_sc_hd__dfrtp_2
X_5194_ _5194_/A _6406_/B VGND VGND VPWR VPWR _5199_/S sky130_fd_sc_hd__nand2_4
X_4145_ _5498_/A0 hold753/X _4147_/S VGND VGND VPWR VPWR _6616_/D sky130_fd_sc_hd__mux2_1
XFILLER_18_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4076_ _6557_/Q _3665_/X _4081_/S VGND VGND VPWR VPWR _6557_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_670 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4978_ _4980_/C _4978_/B _4567_/X VGND VGND VPWR VPWR _5060_/B sky130_fd_sc_hd__or3b_1
XFILLER_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3929_ _6844_/Q input91/X _3932_/S VGND VGND VPWR VPWR _3929_/X sky130_fd_sc_hd__mux2_8
XFILLER_177_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6717_ _6747_/CLK _6717_/D fanout875/X VGND VGND VPWR VPWR _6717_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_109_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6648_ _6724_/CLK _6648_/D fanout858/X VGND VGND VPWR VPWR _6648_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6579_ _6623_/CLK _6579_/D fanout890/X VGND VGND VPWR VPWR _6579_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_59_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire631 _6011_/X VGND VGND VPWR VPWR wire631/X sky130_fd_sc_hd__buf_8
Xwire642 _5998_/X VGND VGND VPWR VPWR wire642/X sky130_fd_sc_hd__buf_8
XFILLER_183_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire653 wire653/A VGND VGND VPWR VPWR wire653/X sky130_fd_sc_hd__buf_8
Xwire664 wire665/X VGND VGND VPWR VPWR wire664/X sky130_fd_sc_hd__buf_6
Xwire675 wire675/A VGND VGND VPWR VPWR wire675/X sky130_fd_sc_hd__buf_6
XFILLER_171_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire697 _5682_/X VGND VGND VPWR VPWR wire697/X sky130_fd_sc_hd__buf_8
Xwire686 _5688_/X VGND VGND VPWR VPWR wire686/X sky130_fd_sc_hd__buf_8
XFILLER_124_675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5950_ _6637_/Q _5973_/A2 wire692/X _6726_/Q _5949_/X VGND VGND VPWR VPWR _5953_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_53_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4901_ _4987_/A _4624_/B _4736_/B _4719_/X VGND VGND VPWR VPWR _4907_/C sky130_fd_sc_hd__a22o_2
XFILLER_46_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5881_ _6723_/Q _5684_/X wire659/X _6604_/Q VGND VGND VPWR VPWR _5881_/X sky130_fd_sc_hd__a22o_2
XFILLER_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4832_ _4832_/A _4832_/B _4832_/C _4832_/D VGND VGND VPWR VPWR _4832_/X sky130_fd_sc_hd__and4_1
XFILLER_60_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_190 _4232_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4763_ _4808_/A _4763_/B _4980_/B _4763_/D VGND VGND VPWR VPWR _4763_/X sky130_fd_sc_hd__or4_1
X_4694_ _4694_/A _5005_/C VGND VGND VPWR VPWR _5069_/B sky130_fd_sc_hd__nor2_8
X_6502_ _6771_/CLK _6502_/D fanout853/X VGND VGND VPWR VPWR _6502_/Q sky130_fd_sc_hd__dfstp_4
X_3714_ wire472/X _3714_/A2 _4316_/A _6764_/Q _3713_/X VGND VGND VPWR VPWR _3717_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6433_ _6446_/A _6447_/B VGND VGND VPWR VPWR _6433_/X sky130_fd_sc_hd__and2_1
XFILLER_174_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3645_ _3645_/A _3645_/B _3645_/C _3645_/D VGND VGND VPWR VPWR _3665_/B sky130_fd_sc_hd__or4_2
XFILLER_161_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3576_ _6880_/Q wire406/X _4082_/A _6566_/Q VGND VGND VPWR VPWR _3576_/X sky130_fd_sc_hd__a22o_1
X_6364_ _7204_/Q _3727_/X _6370_/S VGND VGND VPWR VPWR _7204_/D sky130_fd_sc_hd__mux2_1
X_5315_ _5315_/A _5594_/B VGND VGND VPWR VPWR _5323_/S sky130_fd_sc_hd__nand2_8
X_6295_ wire562/X wire650/X _6295_/B1 _6720_/Q VGND VGND VPWR VPWR _6295_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5246_ wire799/A hold592/X _5249_/S VGND VGND VPWR VPWR _5246_/X sky130_fd_sc_hd__mux2_1
Xhold27 hold3/X VGND VGND VPWR VPWR hold27/X sky130_fd_sc_hd__bufbuf_16
Xhold16 hold52/X VGND VGND VPWR VPWR hold36/A sky130_fd_sc_hd__bufbuf_16
Xhold38 hold38/A VGND VGND VPWR VPWR hold38/X sky130_fd_sc_hd__bufbuf_16
XFILLER_130_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold49 hold49/A VGND VGND VPWR VPWR hold49/X sky130_fd_sc_hd__bufbuf_16
X_5177_ _5048_/A _5177_/B VGND VGND VPWR VPWR _5178_/D sky130_fd_sc_hd__nand2b_1
X_4128_ hold146/X hold83/X _4129_/S VGND VGND VPWR VPWR _4128_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4059_ _5249_/A0 hold456/X _4060_/S VGND VGND VPWR VPWR _6543_/D sky130_fd_sc_hd__mux2_1
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_80_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6824_/CLK sky130_fd_sc_hd__clkbuf_8
Xwire450 _5423_/A VGND VGND VPWR VPWR wire450/X sky130_fd_sc_hd__buf_8
XFILLER_167_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire472 _7142_/Q VGND VGND VPWR VPWR wire472/X sky130_fd_sc_hd__buf_6
Xwire461 _3936_/X VGND VGND VPWR VPWR wire461/X sky130_fd_sc_hd__buf_6
Xwire494 _7072_/Q VGND VGND VPWR VPWR _3213_/A sky130_fd_sc_hd__buf_8
Xwire483 _7101_/Q VGND VGND VPWR VPWR wire483/X sky130_fd_sc_hd__buf_6
Xhold508 _6993_/Q VGND VGND VPWR VPWR hold508/X sky130_fd_sc_hd__bufbuf_16
XFILLER_171_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3430_ _6501_/Q _3995_/A _3368_/Y input17/X VGND VGND VPWR VPWR _3430_/X sky130_fd_sc_hd__a22o_2
Xhold519 _7009_/Q VGND VGND VPWR VPWR hold519/X sky130_fd_sc_hd__bufbuf_16
XFILLER_171_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3361_ _5252_/A _5252_/B VGND VGND VPWR VPWR _3361_/Y sky130_fd_sc_hd__nor2_8
X_6080_ _6974_/Q wire641/X wire639/X wire546/X VGND VGND VPWR VPWR _6080_/X sky130_fd_sc_hd__a22o_1
X_5100_ _4414_/B _5165_/A _5119_/A _4932_/C VGND VGND VPWR VPWR _5101_/D sky130_fd_sc_hd__a211o_1
XFILLER_97_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _5031_/A _5031_/B _4584_/A VGND VGND VPWR VPWR _5102_/B sky130_fd_sc_hd__or3b_2
XFILLER_112_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3292_ _3421_/A _3421_/B hold62/X VGND VGND VPWR VPWR _3292_/X sky130_fd_sc_hd__or3_4
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6982_ _7081_/CLK hold18/X fanout878/X VGND VGND VPWR VPWR _6982_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_19_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_33_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7096_/CLK sky130_fd_sc_hd__clkbuf_8
X_5933_ _6710_/Q wire680/X wire659/X _6606_/Q VGND VGND VPWR VPWR _5933_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5864_ _6988_/Q _5864_/B VGND VGND VPWR VPWR _5864_/X sky130_fd_sc_hd__or2_1
XFILLER_179_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4815_ _4687_/A _4728_/X _4881_/B VGND VGND VPWR VPWR _4817_/C sky130_fd_sc_hd__o21ai_4
XFILLER_21_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5795_ _6929_/Q wire670/X wire651/A _7025_/Q _5794_/X VGND VGND VPWR VPWR _5796_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_193_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4746_ _4746_/A _4746_/B VGND VGND VPWR VPWR _4746_/X sky130_fd_sc_hd__or2_4
XFILLER_147_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_48_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7137_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_31_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4677_ _4690_/A _5062_/B VGND VGND VPWR VPWR _4746_/B sky130_fd_sc_hd__or2_4
XFILLER_147_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6416_ _6420_/A _6421_/B VGND VGND VPWR VPWR _6416_/X sky130_fd_sc_hd__and2_1
X_3628_ input54/X _4025_/A _4292_/A _6745_/Q _3617_/X VGND VGND VPWR VPWR _3629_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6347_ _6618_/Q wire636/X wire634/X _6603_/Q VGND VGND VPWR VPWR _6347_/X sky130_fd_sc_hd__a22o_1
XFILLER_163_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3559_ wire477/X hold97/A _5227_/A _6827_/Q VGND VGND VPWR VPWR _3559_/X sky130_fd_sc_hd__a22o_2
Xinput117 wb_adr_i[26] VGND VGND VPWR VPWR input117/X sky130_fd_sc_hd__clkbuf_4
Xinput106 wb_adr_i[16] VGND VGND VPWR VPWR _4349_/B sky130_fd_sc_hd__clkbuf_4
X_6278_ _6536_/Q wire585/X _6352_/B1 _6640_/Q _6277_/X VGND VGND VPWR VPWR _6281_/C
+ sky130_fd_sc_hd__a221o_2
Xinput128 wb_adr_i[7] VGND VGND VPWR VPWR _4958_/A sky130_fd_sc_hd__buf_8
Xinput139 wb_dat_i[16] VGND VGND VPWR VPWR _6377_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_69_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5229_ wire769/X hold595/X _5233_/S VGND VGND VPWR VPWR _6827_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_90 _5314_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_121_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4600_ _4617_/A _4749_/C VGND VGND VPWR VPWR _4850_/B sky130_fd_sc_hd__nor2_2
X_5580_ wire770/X hold485/X _5580_/S VGND VGND VPWR VPWR _7136_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4531_ _4529_/B _4529_/C _4650_/B VGND VGND VPWR VPWR _4537_/C sky130_fd_sc_hd__a21bo_1
XFILLER_175_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold305 _6873_/Q VGND VGND VPWR VPWR hold305/X sky130_fd_sc_hd__bufbuf_16
X_4462_ _4707_/B _5050_/A VGND VGND VPWR VPWR _4685_/A sky130_fd_sc_hd__or2_4
Xhold316 _6618_/Q VGND VGND VPWR VPWR hold316/X sky130_fd_sc_hd__bufbuf_16
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6201_ _6875_/Q wire593/X wire591/X wire542/X _6200_/X VGND VGND VPWR VPWR _6206_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_144_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold349 _6985_/Q VGND VGND VPWR VPWR hold349/X sky130_fd_sc_hd__bufbuf_16
Xhold327 _6623_/Q VGND VGND VPWR VPWR hold327/X sky130_fd_sc_hd__bufbuf_16
XFILLER_89_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold338 _3255_/X VGND VGND VPWR VPWR hold338/X sky130_fd_sc_hd__bufbuf_16
X_3413_ wire901/X _3322_/Y _3368_/Y input18/X _3412_/X VGND VGND VPWR VPWR _3414_/D
+ sky130_fd_sc_hd__a221o_4
X_4393_ _5031_/A _4663_/A VGND VGND VPWR VPWR _4772_/A sky130_fd_sc_hd__nor2_8
X_7181_ _7196_/CLK _7181_/D fanout870/X VGND VGND VPWR VPWR _7181_/Q sky130_fd_sc_hd__dfrtp_4
X_6132_ _6306_/A _6132_/B _6132_/C _6132_/D VGND VGND VPWR VPWR _6132_/X sky130_fd_sc_hd__or4_4
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3344_ _5225_/A _5252_/B VGND VGND VPWR VPWR _3995_/A sky130_fd_sc_hd__nor2_8
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout829 _6425_/B VGND VGND VPWR VPWR _6455_/B sky130_fd_sc_hd__buf_8
Xfanout818 wire821/A VGND VGND VPWR VPWR _3975_/B sky130_fd_sc_hd__buf_8
XFILLER_112_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3275_ _3314_/A _3293_/B _3309_/B VGND VGND VPWR VPWR _3508_/A sky130_fd_sc_hd__or3_4
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6063_ _7078_/Q _6211_/B VGND VGND VPWR VPWR _6063_/X sky130_fd_sc_hd__and2_1
X_5014_ _4561_/Y _4758_/B _4725_/A _4839_/X VGND VGND VPWR VPWR _5016_/C sky130_fd_sc_hd__a211o_1
XFILLER_100_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6965_ _7153_/CLK _6965_/D fanout881/X VGND VGND VPWR VPWR _6965_/Q sky130_fd_sc_hd__dfstp_4
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5916_ _6531_/Q _5722_/B _5915_/X _6308_/S VGND VGND VPWR VPWR _5916_/X sky130_fd_sc_hd__o211a_1
XFILLER_53_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6896_ _7122_/CLK _6896_/D fanout887/X VGND VGND VPWR VPWR _6896_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_166_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5847_ _7043_/Q _5683_/X _5702_/X _6891_/Q VGND VGND VPWR VPWR _5847_/X sky130_fd_sc_hd__a22o_1
X_5778_ _6912_/Q wire699/X wire666/X _6864_/Q _5768_/X VGND VGND VPWR VPWR _5778_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_166_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4729_ _4740_/A _4819_/A _4729_/C VGND VGND VPWR VPWR _4729_/X sky130_fd_sc_hd__and3_1
XFILLER_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold850 _6515_/Q VGND VGND VPWR VPWR hold850/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6750_ _7225_/CLK _6750_/D fanout851/X VGND VGND VPWR VPWR _6750_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_188_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5701_ _5864_/B _5702_/B _5701_/C VGND VGND VPWR VPWR _5701_/X sky130_fd_sc_hd__and3_4
X_3962_ _3962_/A VGND VGND VPWR VPWR _3962_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3893_ _3893_/A _3893_/B input120/X input117/X VGND VGND VPWR VPWR _3894_/D sky130_fd_sc_hd__or4bb_1
XFILLER_149_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6681_ _7223_/CLK _6681_/D _6455_/A VGND VGND VPWR VPWR _6681_/Q sky130_fd_sc_hd__dfrtp_2
X_5632_ _7164_/Q _7163_/Q VGND VGND VPWR VPWR _5703_/B sky130_fd_sc_hd__nor2_8
X_5563_ hold150/X hold848/X _5564_/S VGND VGND VPWR VPWR _5563_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4514_ _4671_/A _4995_/A VGND VGND VPWR VPWR _5079_/A sky130_fd_sc_hd__nor2_4
XFILLER_172_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5494_ _5602_/A0 hold294/X _5494_/S VGND VGND VPWR VPWR _5494_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold124 _6483_/Q VGND VGND VPWR VPWR hold124/X sky130_fd_sc_hd__bufbuf_16
Xhold102 _3292_/X VGND VGND VPWR VPWR _3668_/A sky130_fd_sc_hd__bufbuf_16
Xhold135 _3309_/X VGND VGND VPWR VPWR _3552_/B sky130_fd_sc_hd__bufbuf_16
Xhold113 _3368_/B VGND VGND VPWR VPWR _3528_/B sky130_fd_sc_hd__bufbuf_16
X_4445_ _4735_/A _4672_/A _4469_/A _4395_/D _5050_/A VGND VGND VPWR VPWR _4445_/X
+ sky130_fd_sc_hd__o2111a_2
Xhold146 _6602_/Q VGND VGND VPWR VPWR hold146/X sky130_fd_sc_hd__bufbuf_16
XFILLER_132_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold157 _5518_/X VGND VGND VPWR VPWR _7081_/D sky130_fd_sc_hd__bufbuf_16
Xhold168 _3342_/Y VGND VGND VPWR VPWR _3421_/C sky130_fd_sc_hd__bufbuf_16
Xhold179 _7097_/Q VGND VGND VPWR VPWR hold179/X sky130_fd_sc_hd__bufbuf_16
XFILLER_171_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7164_ _3949_/A1 _7164_/D fanout879/X VGND VGND VPWR VPWR _7164_/Q sky130_fd_sc_hd__dfrtp_2
X_4376_ _4996_/A VGND VGND VPWR VPWR _4376_/Y sky130_fd_sc_hd__clkinv_2
X_6115_ wire513/A _6010_/Y wire616/X _3211_/A _6112_/X VGND VGND VPWR VPWR _6121_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_100_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3327_ _3369_/A _5225_/B VGND VGND VPWR VPWR _3327_/Y sky130_fd_sc_hd__nor2_8
XFILLER_86_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7095_ _7095_/CLK _7095_/D fanout862/X VGND VGND VPWR VPWR _7095_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ _6941_/Q _6301_/B1 wire610/X wire520/X VGND VGND VPWR VPWR _6046_/X sky130_fd_sc_hd__a22o_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3258_ _3257_/X hold132/X _3953_/A VGND VGND VPWR VPWR _3258_/X sky130_fd_sc_hd__mux2_4
XFILLER_170_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6948_ _7036_/CLK _6948_/D fanout869/X VGND VGND VPWR VPWR _6948_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_41_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6879_ _7145_/CLK _6879_/D fanout881/X VGND VGND VPWR VPWR _6879_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_139_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length614 wire615/X VGND VGND VPWR VPWR _6337_/B1 sky130_fd_sc_hd__buf_6
XFILLER_154_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length669 wire670/X VGND VGND VPWR VPWR _5964_/B1 sky130_fd_sc_hd__buf_6
Xmax_length658 _5705_/X VGND VGND VPWR VPWR wire656/A sky130_fd_sc_hd__buf_6
XFILLER_118_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold680 _6686_/Q VGND VGND VPWR VPWR hold680/X sky130_fd_sc_hd__bufbuf_16
XFILLER_110_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold691 _6536_/Q VGND VGND VPWR VPWR hold691/X sky130_fd_sc_hd__bufbuf_16
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput207 _3236_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[4] sky130_fd_sc_hd__buf_8
Xoutput229 _6514_/Q VGND VGND VPWR VPWR mgmt_gpio_out[24] sky130_fd_sc_hd__buf_8
XFILLER_153_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput218 _3949_/X VGND VGND VPWR VPWR mgmt_gpio_out[14] sky130_fd_sc_hd__clkbuf_4
XFILLER_141_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4230_ hold644/X wire757/X _4234_/S VGND VGND VPWR VPWR _4230_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4161_ _5487_/A0 hold791/X _4165_/S VGND VGND VPWR VPWR _6629_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4092_ _6571_/Q _3606_/X _4096_/S VGND VGND VPWR VPWR _6571_/D sky130_fd_sc_hd__mux2_1
XFILLER_82_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6802_ _6806_/CLK _6802_/D _6435_/A VGND VGND VPWR VPWR _6802_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4994_ _4399_/Y _4539_/D _4586_/B _4987_/X VGND VGND VPWR VPWR _5000_/C sky130_fd_sc_hd__o31a_4
X_6733_ _6974_/CLK _6733_/D fanout875/X VGND VGND VPWR VPWR _6733_/Q sky130_fd_sc_hd__dfrtp_2
X_3945_ _6681_/Q input3/X input1/X VGND VGND VPWR VPWR _3945_/X sky130_fd_sc_hd__mux2_4
XFILLER_176_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6664_ _6668_/CLK _6664_/D _6443_/X VGND VGND VPWR VPWR _6664_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_176_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5615_ _7157_/Q _7158_/Q _7159_/Q _5615_/D VGND VGND VPWR VPWR _5616_/A sky130_fd_sc_hd__and4_2
X_3876_ _6459_/Q _3875_/X _3876_/S VGND VGND VPWR VPWR _6459_/D sky130_fd_sc_hd__mux2_1
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6595_ _6646_/CLK _6595_/D fanout856/X VGND VGND VPWR VPWR _6595_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_129_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5546_ wire753/X hold815/X _5548_/S VGND VGND VPWR VPWR _7106_/D sky130_fd_sc_hd__mux2_1
XFILLER_191_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5477_ _5477_/A _5576_/B VGND VGND VPWR VPWR _5485_/S sky130_fd_sc_hd__and2_4
X_7216_ _7218_/CLK _7216_/D wire915/X VGND VGND VPWR VPWR hold23/A sky130_fd_sc_hd__dfrtp_1
X_4428_ _4711_/A _5165_/A _4428_/C VGND VGND VPWR VPWR _5140_/A sky130_fd_sc_hd__and3_2
XFILLER_144_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4359_ _4672_/A _4735_/A VGND VGND VPWR VPWR _4558_/B sky130_fd_sc_hd__nand2b_4
X_7147_ _7147_/CLK hold58/X fanout888/X VGND VGND VPWR VPWR _7147_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_98_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7078_ _7135_/CLK _7078_/D fanout864/X VGND VGND VPWR VPWR _7078_/Q sky130_fd_sc_hd__dfstp_1
X_6029_ _6037_/C _6035_/C _6032_/C VGND VGND VPWR VPWR _6029_/X sky130_fd_sc_hd__and3_4
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire813 _3916_/A VGND VGND VPWR VPWR wire813/X sky130_fd_sc_hd__buf_6
Xwire802 wire802/A VGND VGND VPWR VPWR wire802/X sky130_fd_sc_hd__buf_8
Xwire824 _5663_/A VGND VGND VPWR VPWR wire824/X sky130_fd_sc_hd__buf_8
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length400 _5513_/A VGND VGND VPWR VPWR _3638_/B1 sky130_fd_sc_hd__buf_6
XFILLER_182_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length433 _4023_/S VGND VGND VPWR VPWR _4021_/S sky130_fd_sc_hd__buf_6
Xwire835 wire835/A VGND VGND VPWR VPWR wire835/X sky130_fd_sc_hd__buf_6
Xmax_length422 hold129/X VGND VGND VPWR VPWR wire421/A sky130_fd_sc_hd__buf_6
XFILLER_6_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_22 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_350 _5234_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3730_ _6474_/Q _6459_/Q _6824_/Q VGND VGND VPWR VPWR _3730_/X sky130_fd_sc_hd__or3_4
XFILLER_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3661_ _5225_/A _3543_/B _4049_/A _6537_/Q VGND VGND VPWR VPWR _3663_/C sky130_fd_sc_hd__a2bb2o_1
X_6380_ _4236_/C _6380_/A2 _6380_/B1 _4236_/A VGND VGND VPWR VPWR _6380_/X sky130_fd_sc_hd__a22o_1
X_5400_ hold602/X wire773/X _5404_/S VGND VGND VPWR VPWR _6976_/D sky130_fd_sc_hd__mux2_1
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3592_ _6788_/Q _5185_/A _5194_/A _6803_/Q _3556_/X VGND VGND VPWR VPWR _3593_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5331_ _5601_/A0 _6915_/Q _5332_/S VGND VGND VPWR VPWR _5331_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7001_ _7137_/CLK _7001_/D fanout871/X VGND VGND VPWR VPWR _7001_/Q sky130_fd_sc_hd__dfrtp_2
X_5262_ hold663/X wire802/X _5269_/S VGND VGND VPWR VPWR _6853_/D sky130_fd_sc_hd__mux2_1
X_4213_ _6695_/Q hold27/X hold46/X VGND VGND VPWR VPWR hold47/A sky130_fd_sc_hd__mux2_1
XFILLER_141_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5193_ _6408_/A0 _6799_/Q _5193_/S VGND VGND VPWR VPWR _6799_/D sky130_fd_sc_hd__mux2_1
X_4144_ wire794/X hold675/X _4147_/S VGND VGND VPWR VPWR _6615_/D sky130_fd_sc_hd__mux2_1
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4075_ _6556_/Q _3727_/X _4081_/S VGND VGND VPWR VPWR _6556_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_3_4_0_csclk clkbuf_3_5_0_csclk/A VGND VGND VPWR VPWR _6708_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_64_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6716_ _6747_/CLK hold78/X _6420_/A VGND VGND VPWR VPWR _6716_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4977_ _5132_/A _5142_/B _5069_/D _4977_/D VGND VGND VPWR VPWR _4977_/X sky130_fd_sc_hd__or4_1
X_3928_ _3928_/A _3928_/B VGND VGND VPWR VPWR _6458_/D sky130_fd_sc_hd__and2_1
X_3859_ _6666_/Q _3859_/B VGND VGND VPWR VPWR _3859_/Y sky130_fd_sc_hd__nand2_8
X_6647_ _6724_/CLK _6647_/D fanout858/X VGND VGND VPWR VPWR _6647_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6578_ _6720_/CLK _6578_/D fanout874/X VGND VGND VPWR VPWR _6578_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_118_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5529_ wire746/X hold706/X _5530_/S VGND VGND VPWR VPWR _5529_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire632 _6020_/C VGND VGND VPWR VPWR wire632/X sky130_fd_sc_hd__buf_8
Xwire610 _6033_/X VGND VGND VPWR VPWR wire610/X sky130_fd_sc_hd__buf_8
Xwire643 _5998_/X VGND VGND VPWR VPWR wire643/X sky130_fd_sc_hd__buf_6
XFILLER_7_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire665 _5701_/X VGND VGND VPWR VPWR wire665/X sky130_fd_sc_hd__buf_8
XFILLER_143_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4900_ _4947_/B _4898_/B _4591_/B VGND VGND VPWR VPWR _5075_/B sky130_fd_sc_hd__a21oi_1
XFILLER_80_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5880_ _6728_/Q wire710/X _5879_/X VGND VGND VPWR VPWR _5883_/C sky130_fd_sc_hd__a21o_1
XFILLER_61_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4831_ _4707_/B _4746_/B _4728_/X _4886_/B VGND VGND VPWR VPWR _4832_/D sky130_fd_sc_hd__o211a_1
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_180 _6817_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_191 _4232_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4762_ _4949_/B _4537_/X _4565_/Y _4759_/Y VGND VGND VPWR VPWR _4763_/D sky130_fd_sc_hd__a31o_4
XFILLER_159_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4693_ _4774_/C _4693_/B VGND VGND VPWR VPWR _4711_/C sky130_fd_sc_hd__and2_4
X_6501_ _6771_/CLK _6501_/D fanout853/X VGND VGND VPWR VPWR _6501_/Q sky130_fd_sc_hd__dfstp_4
X_3713_ _6759_/Q _4310_/A _5191_/A _6799_/Q VGND VGND VPWR VPWR _3713_/X sky130_fd_sc_hd__a22o_2
XFILLER_174_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3644_ _7023_/Q _3301_/Y _4274_/A _6730_/Q _3643_/X VGND VGND VPWR VPWR _3645_/D
+ sky130_fd_sc_hd__a221o_1
X_6432_ _6446_/A _6455_/B VGND VGND VPWR VPWR _6432_/X sky130_fd_sc_hd__and2_1
XFILLER_146_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3575_ _3236_/A _5297_/A _5405_/A _6984_/Q _3574_/X VGND VGND VPWR VPWR _3578_/C
+ sky130_fd_sc_hd__a221o_4
X_6363_ _7203_/Q wire350/X _6370_/S VGND VGND VPWR VPWR _7203_/D sky130_fd_sc_hd__mux2_1
X_5314_ _5602_/A0 hold290/X _5314_/S VGND VGND VPWR VPWR _5314_/X sky130_fd_sc_hd__mux2_1
X_6294_ _6656_/Q _6311_/B _6289_/X _6291_/X _6293_/X VGND VGND VPWR VPWR _6294_/X
+ sky130_fd_sc_hd__a2111o_1
X_5245_ _5245_/A _5594_/B VGND VGND VPWR VPWR _5248_/S sky130_fd_sc_hd__nand2_4
XFILLER_130_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold28 hold28/A VGND VGND VPWR VPWR hold28/X sky130_fd_sc_hd__bufbuf_16
Xhold17 hold37/X VGND VGND VPWR VPWR hold38/A sky130_fd_sc_hd__bufbuf_16
XFILLER_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold39 hold39/A VGND VGND VPWR VPWR hold39/X sky130_fd_sc_hd__bufbuf_16
XFILLER_152_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5176_ _4947_/B _4757_/B _5050_/C _4717_/B _4837_/X VGND VGND VPWR VPWR _5177_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_84_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4127_ _6601_/Q _5498_/A0 _4129_/S VGND VGND VPWR VPWR _6601_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4058_ _5336_/A1 _6542_/Q _4060_/S VGND VGND VPWR VPWR _6542_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_5_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A VGND VGND VPWR VPWR _7190_/CLK sky130_fd_sc_hd__clkbuf_8
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire451 _3510_/B VGND VGND VPWR VPWR _3733_/B sky130_fd_sc_hd__buf_8
XFILLER_171_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold509 _6954_/Q VGND VGND VPWR VPWR hold509/X sky130_fd_sc_hd__bufbuf_16
Xwire484 _7097_/Q VGND VGND VPWR VPWR wire484/X sky130_fd_sc_hd__buf_6
XFILLER_144_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire462 wire463/X VGND VGND VPWR VPWR wire462/X sky130_fd_sc_hd__buf_6
Xwire473 _7131_/Q VGND VGND VPWR VPWR wire473/X sky130_fd_sc_hd__buf_6
XFILLER_7_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire495 _7067_/Q VGND VGND VPWR VPWR wire495/X sky130_fd_sc_hd__buf_6
X_3360_ _7132_/Q hold88/A _5441_/A _7020_/Q VGND VGND VPWR VPWR _3360_/X sky130_fd_sc_hd__a22o_1
XFILLER_112_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5030_ _4500_/A _4758_/A _5004_/A _5099_/C _4932_/A VGND VGND VPWR VPWR _5034_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_112_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3291_ _3505_/A hold96/X VGND VGND VPWR VPWR _5477_/A sky130_fd_sc_hd__nor2_8
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6981_ _6981_/CLK _6981_/D fanout878/X VGND VGND VPWR VPWR _6981_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_38_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5932_ _6656_/Q wire675/X wire651/X _6760_/Q _5931_/X VGND VGND VPWR VPWR _5937_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_53_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5863_ _6996_/Q wire692/X _5703_/X _6876_/Q _5862_/X VGND VGND VPWR VPWR _5871_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4814_ _5095_/A _4950_/B _4814_/C _4812_/X VGND VGND VPWR VPWR _4817_/B sky130_fd_sc_hd__or4b_2
XFILLER_166_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5794_ _7081_/Q wire675/A _5794_/B1 wire548/X VGND VGND VPWR VPWR _5794_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4745_ _4745_/A _4745_/B VGND VGND VPWR VPWR _4745_/X sky130_fd_sc_hd__or2_1
XFILLER_159_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4676_ _4685_/A _5062_/B _4696_/B VGND VGND VPWR VPWR _4832_/C sky130_fd_sc_hd__or3b_4
XFILLER_147_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6415_ _6420_/A _6421_/B VGND VGND VPWR VPWR _6415_/X sky130_fd_sc_hd__and2_1
X_3627_ _6983_/Q _3739_/B1 _4256_/A _6715_/Q _3616_/X VGND VGND VPWR VPWR _3629_/C
+ sky130_fd_sc_hd__a221o_1
X_6346_ wire564/X wire597/X wire611/X _6742_/Q _6345_/X VGND VGND VPWR VPWR _6356_/C
+ sky130_fd_sc_hd__a221o_1
X_3558_ _7088_/Q _5522_/A _4043_/A _6533_/Q VGND VGND VPWR VPWR _3558_/X sky130_fd_sc_hd__a22o_1
XFILLER_163_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput107 wb_adr_i[17] VGND VGND VPWR VPWR _4349_/A sky130_fd_sc_hd__clkbuf_4
Xinput118 wb_adr_i[27] VGND VGND VPWR VPWR _3893_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_130_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3489_ _3540_/A _3520_/B VGND VGND VPWR VPWR _4136_/A sky130_fd_sc_hd__nor2_8
XFILLER_88_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6277_ _6635_/Q wire712/X wire625/X wire570/X VGND VGND VPWR VPWR _6277_/X sky130_fd_sc_hd__a22o_1
Xinput129 wb_adr_i[8] VGND VGND VPWR VPWR _4351_/B sky130_fd_sc_hd__clkbuf_4
X_5228_ _5572_/A0 hold491/X _5233_/S VGND VGND VPWR VPWR _6826_/D sky130_fd_sc_hd__mux2_1
XFILLER_186_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5159_ _4414_/B _5165_/A _4922_/A _4704_/X _5156_/B VGND VGND VPWR VPWR _5159_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_72_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_1_0_csclk clkbuf_2_1_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_3_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_91 _5681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_80 _4267_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4530_ _4529_/B _4529_/C _4650_/B VGND VGND VPWR VPWR _4533_/C sky130_fd_sc_hd__a21boi_4
XFILLER_156_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4461_ _4707_/B _5050_/A VGND VGND VPWR VPWR _4719_/B sky130_fd_sc_hd__nor2_1
Xhold306 _6603_/Q VGND VGND VPWR VPWR hold306/X sky130_fd_sc_hd__bufbuf_16
Xhold317 _6979_/Q VGND VGND VPWR VPWR hold317/X sky130_fd_sc_hd__bufbuf_16
XFILLER_144_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6200_ _6963_/Q wire624/X wire613/X _7059_/Q VGND VGND VPWR VPWR _6200_/X sky130_fd_sc_hd__a22o_1
Xhold328 _6567_/Q VGND VGND VPWR VPWR hold328/X sky130_fd_sc_hd__bufbuf_16
X_7180_ _7194_/CLK _7180_/D fanout870/X VGND VGND VPWR VPWR _7180_/Q sky130_fd_sc_hd__dfrtp_4
Xhold339 _3256_/Y VGND VGND VPWR VPWR hold339/X sky130_fd_sc_hd__bufbuf_16
X_3412_ input27/X _3302_/Y _3371_/Y _7123_/Q VGND VGND VPWR VPWR _3412_/X sky130_fd_sc_hd__a22o_1
X_6131_ _6131_/A _6131_/B _6131_/C _6131_/D VGND VGND VPWR VPWR _6132_/D sky130_fd_sc_hd__or4_1
X_4392_ _4469_/A _4395_/D VGND VGND VPWR VPWR _4663_/A sky130_fd_sc_hd__or2_4
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout808 _3241_/Y VGND VGND VPWR VPWR _5864_/B sky130_fd_sc_hd__buf_8
XFILLER_112_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3343_ _3343_/A _3421_/C VGND VGND VPWR VPWR _5252_/B sky130_fd_sc_hd__or2_4
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _7110_/Q wire650/X _6295_/B1 _7150_/Q VGND VGND VPWR VPWR _6062_/X sky130_fd_sc_hd__a22o_1
XFILLER_85_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3274_ _3505_/A _3365_/A VGND VGND VPWR VPWR _5432_/A sky130_fd_sc_hd__nor2_8
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5013_ _5013_/A _5013_/B VGND VGND VPWR VPWR _5156_/B sky130_fd_sc_hd__or2_4
XFILLER_85_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6964_ _7152_/CLK _6964_/D fanout886/X VGND VGND VPWR VPWR _6964_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6895_ _7128_/CLK _6895_/D _6421_/A VGND VGND VPWR VPWR _6895_/Q sky130_fd_sc_hd__dfrtp_2
X_5915_ _5915_/A _5915_/B _5915_/C _5915_/D VGND VGND VPWR VPWR _5915_/X sky130_fd_sc_hd__or4_1
XFILLER_34_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5846_ wire532/X wire660/X _5705_/X _6947_/Q _5845_/X VGND VGND VPWR VPWR _5849_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5777_ _5777_/A _5777_/B _5777_/C _5777_/D VGND VGND VPWR VPWR _5777_/X sky130_fd_sc_hd__or4_4
X_4728_ _4728_/A _4746_/B VGND VGND VPWR VPWR _4728_/X sky130_fd_sc_hd__or2_4
XFILLER_135_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4659_ _4659_/A _4758_/B VGND VGND VPWR VPWR _4832_/B sky130_fd_sc_hd__nand2_8
XFILLER_162_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold851 _6674_/Q VGND VGND VPWR VPWR hold851/X sky130_fd_sc_hd__bufbuf_16
XFILLER_107_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold840 _6946_/Q VGND VGND VPWR VPWR hold840/X sky130_fd_sc_hd__bufbuf_16
XFILLER_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6329_ _6538_/Q wire585/X _6352_/B1 _6642_/Q _6328_/X VGND VGND VPWR VPWR _6330_/D
+ sky130_fd_sc_hd__a221o_4
XFILLER_103_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_32_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7133_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_95_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_47_csclk clkbuf_opt_1_0_csclk/X VGND VGND VPWR VPWR _7081_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_75_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3961_ _6473_/Q _3961_/B VGND VGND VPWR VPWR _3962_/A sky130_fd_sc_hd__or2_4
X_5700_ _5864_/B _5703_/B _5707_/B VGND VGND VPWR VPWR _5700_/X sky130_fd_sc_hd__and3_4
X_3892_ _3892_/A _3892_/B input131/X wire912/X VGND VGND VPWR VPWR _3894_/C sky130_fd_sc_hd__or4bb_1
XFILLER_148_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6680_ _7194_/CLK _6680_/D fanout866/X VGND VGND VPWR VPWR _6680_/Q sky130_fd_sc_hd__dfrtp_2
X_5631_ _7163_/Q _5629_/B _5635_/B _5630_/Y VGND VGND VPWR VPWR _7163_/D sky130_fd_sc_hd__a31o_1
XFILLER_31_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5562_ _5598_/A0 hold578/X _5564_/S VGND VGND VPWR VPWR _7120_/D sky130_fd_sc_hd__mux2_1
XFILLER_148_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4513_ _4513_/A _4513_/B VGND VGND VPWR VPWR _4990_/A sky130_fd_sc_hd__or2_4
X_5493_ _5601_/A0 hold228/X _5494_/S VGND VGND VPWR VPWR _7059_/D sky130_fd_sc_hd__mux2_1
Xhold114 _3473_/Y VGND VGND VPWR VPWR _4067_/A sky130_fd_sc_hd__bufbuf_16
Xhold125 hold339/X VGND VGND VPWR VPWR hold125/X sky130_fd_sc_hd__bufbuf_16
Xhold103 _3298_/Y VGND VGND VPWR VPWR wire438/A sky130_fd_sc_hd__bufbuf_16
X_4444_ _4958_/B _4444_/B VGND VGND VPWR VPWR _4572_/A sky130_fd_sc_hd__nand2_8
Xhold147 _4128_/X VGND VGND VPWR VPWR _6602_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_144_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold158 _6592_/Q VGND VGND VPWR VPWR hold158/X sky130_fd_sc_hd__bufbuf_16
Xhold136 _3322_/Y VGND VGND VPWR VPWR hold136/X sky130_fd_sc_hd__bufbuf_16
X_4375_ _4553_/A _4400_/A VGND VGND VPWR VPWR _4996_/A sky130_fd_sc_hd__or2_4
X_7163_ _3949_/A1 _7163_/D fanout879/X VGND VGND VPWR VPWR _7163_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_98_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold169 _3419_/X VGND VGND VPWR VPWR _3732_/B sky130_fd_sc_hd__bufbuf_16
X_6114_ _6976_/Q wire641/X wire633/X _3233_/A VGND VGND VPWR VPWR _6131_/B sky130_fd_sc_hd__a22o_1
X_3326_ _6924_/Q _5333_/A _5324_/A _6916_/Q VGND VGND VPWR VPWR _3326_/X sky130_fd_sc_hd__a22o_1
XFILLER_112_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7094_ _7129_/CLK _7094_/D fanout863/X VGND VGND VPWR VPWR _7094_/Q sky130_fd_sc_hd__dfstp_4
X_6045_ _7117_/Q _6023_/D _6293_/B1 _6989_/Q _6044_/X VGND VGND VPWR VPWR _6059_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_100_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3257_ hold331/X _3845_/A hold124/X VGND VGND VPWR VPWR _3257_/X sky130_fd_sc_hd__a21o_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6947_ _7072_/CLK _6947_/D fanout870/X VGND VGND VPWR VPWR _6947_/Q sky130_fd_sc_hd__dfrtp_2
X_6878_ _7111_/CLK _6878_/D fanout881/X VGND VGND VPWR VPWR _6878_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_167_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5829_ _5611_/A _7180_/Q wire381/A VGND VGND VPWR VPWR _5829_/X sky130_fd_sc_hd__a21o_1
XFILLER_22_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length626 _6022_/B VGND VGND VPWR VPWR _6301_/B1 sky130_fd_sc_hd__buf_6
XFILLER_147_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold681 _4231_/X VGND VGND VPWR VPWR _6686_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_1_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold670 _6757_/Q VGND VGND VPWR VPWR hold670/X sky130_fd_sc_hd__bufbuf_16
Xhold692 _6710_/Q VGND VGND VPWR VPWR hold692/X sky130_fd_sc_hd__bufbuf_16
XFILLER_103_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput208 _3235_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[5] sky130_fd_sc_hd__buf_8
Xoutput219 _3948_/X VGND VGND VPWR VPWR mgmt_gpio_out[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_126_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4160_ _4160_/A _5236_/B VGND VGND VPWR VPWR _4165_/S sky130_fd_sc_hd__nand2_8
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4091_ _6570_/Q _3665_/X _4096_/S VGND VGND VPWR VPWR _6570_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6801_ _6806_/CLK _6801_/D _6435_/A VGND VGND VPWR VPWR _6801_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4993_ _4478_/B _4992_/Y _4991_/X VGND VGND VPWR VPWR _5118_/C sky130_fd_sc_hd__o21ai_4
XFILLER_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6732_ _6771_/CLK _6732_/D fanout854/X VGND VGND VPWR VPWR _6732_/Q sky130_fd_sc_hd__dfrtp_2
X_3944_ _6473_/Q _3965_/B _3942_/X _3943_/Y VGND VGND VPWR VPWR _3944_/X sky130_fd_sc_hd__a22o_1
XFILLER_149_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3875_ _6486_/Q _3875_/B VGND VGND VPWR VPWR _3875_/X sky130_fd_sc_hd__and2b_1
X_6663_ _6851_/CLK _6663_/D fanout850/X VGND VGND VPWR VPWR _6663_/Q sky130_fd_sc_hd__dfrtp_2
X_5614_ _7157_/Q _7158_/Q _5615_/D _7159_/Q VGND VGND VPWR VPWR _5617_/B sky130_fd_sc_hd__a31o_1
XFILLER_176_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6594_ _6727_/CLK _6594_/D fanout858/X VGND VGND VPWR VPWR _6594_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_129_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5545_ _5572_/A0 hold521/X _5548_/S VGND VGND VPWR VPWR _5545_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5476_ wire739/X hold687/X _5476_/S VGND VGND VPWR VPWR _7044_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_3_0_0_csclk clkbuf_3_1_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_0_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
X_7215_ _7218_/CLK _7215_/D wire915/X VGND VGND VPWR VPWR _7215_/Q sky130_fd_sc_hd__dfrtp_2
X_4427_ _5165_/A _4428_/C VGND VGND VPWR VPWR _5023_/B sky130_fd_sc_hd__nand2_2
X_7146_ _7147_/CLK _7146_/D fanout888/X VGND VGND VPWR VPWR _7146_/Q sky130_fd_sc_hd__dfrtp_2
X_4358_ _4553_/A _4774_/A _4484_/B VGND VGND VPWR VPWR _4478_/B sky130_fd_sc_hd__or3b_4
XFILLER_171_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4289_ _6409_/A0 _6740_/Q _4291_/S VGND VGND VPWR VPWR _6740_/D sky130_fd_sc_hd__mux2_1
X_3309_ _3309_/A _3309_/B _3293_/B VGND VGND VPWR VPWR _3309_/X sky130_fd_sc_hd__or3b_4
X_7077_ _7135_/CLK _7077_/D fanout863/X VGND VGND VPWR VPWR _7077_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_86_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6028_ _6037_/C _6033_/C _6035_/C VGND VGND VPWR VPWR _6028_/X sky130_fd_sc_hd__and3_4
XFILLER_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire814 _6707_/Q VGND VGND VPWR VPWR _4236_/C sky130_fd_sc_hd__buf_8
XFILLER_167_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length434 _3310_/Y VGND VGND VPWR VPWR _4023_/S sky130_fd_sc_hd__buf_8
XFILLER_129_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire836 wire836/A VGND VGND VPWR VPWR wire836/X sky130_fd_sc_hd__buf_6
Xmax_length423 wire424/X VGND VGND VPWR VPWR _5324_/A sky130_fd_sc_hd__buf_8
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length412 _3346_/Y VGND VGND VPWR VPWR _3714_/A2 sky130_fd_sc_hd__buf_6
XFILLER_155_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_340 hold633/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_351 _3972_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3660_ wire563/X _4298_/A _4184_/A _6651_/Q _3659_/X VGND VGND VPWR VPWR _3663_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3591_ _6657_/Q _4190_/A _6406_/A _7224_/Q _3565_/X VGND VGND VPWR VPWR _3593_/C
+ sky130_fd_sc_hd__a221o_1
X_5330_ _5600_/A0 hold475/X _5332_/S VGND VGND VPWR VPWR _6914_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5261_ _5261_/A _5459_/B VGND VGND VPWR VPWR _5269_/S sky130_fd_sc_hd__and2_4
XFILLER_5_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4212_ hold409/X _4211_/X _4218_/S VGND VGND VPWR VPWR _4212_/X sky130_fd_sc_hd__mux2_1
X_7000_ _7096_/CLK _7000_/D fanout882/X VGND VGND VPWR VPWR _7000_/Q sky130_fd_sc_hd__dfrtp_2
X_5192_ _6407_/A0 hold803/X _5193_/S VGND VGND VPWR VPWR _6798_/D sky130_fd_sc_hd__mux2_1
X_4143_ hold465/X hold576/X _4147_/S VGND VGND VPWR VPWR _4143_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4074_ _6555_/Q wire350/X _4081_/S VGND VGND VPWR VPWR _6555_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6715_ _6747_/CLK _6715_/D _6420_/A VGND VGND VPWR VPWR _6715_/Q sky130_fd_sc_hd__dfstp_4
X_4976_ _4976_/A _4976_/B _4976_/C _4638_/X VGND VGND VPWR VPWR _4977_/D sky130_fd_sc_hd__or4b_1
XFILLER_137_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3927_ _6665_/Q _6668_/Q _3196_/Y VGND VGND VPWR VPWR _3928_/B sky130_fd_sc_hd__o21ai_1
XFILLER_192_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3858_ _3864_/B VGND VGND VPWR VPWR _3858_/Y sky130_fd_sc_hd__inv_2
X_6646_ _6646_/CLK _6646_/D fanout856/X VGND VGND VPWR VPWR _6646_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_166_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6577_ _6650_/CLK _6577_/D fanout858/X VGND VGND VPWR VPWR _6577_/Q sky130_fd_sc_hd__dfrtp_2
X_3789_ wire838/X _3280_/Y _3308_/Y _4274_/A _6728_/Q VGND VGND VPWR VPWR _3789_/X
+ sky130_fd_sc_hd__a32o_1
X_5528_ wire753/X hold816/X _5530_/S VGND VGND VPWR VPWR _5528_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5459_ _5459_/A _5459_/B VGND VGND VPWR VPWR _5467_/S sky130_fd_sc_hd__nand2_8
XFILLER_133_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7129_ _7129_/CLK _7129_/D fanout864/X VGND VGND VPWR VPWR _7129_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_87_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire600 _6021_/A VGND VGND VPWR VPWR wire600/X sky130_fd_sc_hd__buf_8
XFILLER_128_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire633 _6020_/C VGND VGND VPWR VPWR wire633/X sky130_fd_sc_hd__buf_8
Xwire611 _6033_/X VGND VGND VPWR VPWR wire611/X sky130_fd_sc_hd__buf_8
Xwire666 _5700_/X VGND VGND VPWR VPWR wire666/X sky130_fd_sc_hd__buf_8
Xwire644 _5998_/X VGND VGND VPWR VPWR _6020_/B sky130_fd_sc_hd__buf_6
XFILLER_6_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire677 _5693_/X VGND VGND VPWR VPWR wire677/X sky130_fd_sc_hd__buf_8
Xwire699 _5680_/X VGND VGND VPWR VPWR wire699/X sky130_fd_sc_hd__buf_8
XFILLER_108_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4830_ _4672_/B _4737_/Y _4829_/X _4692_/C VGND VGND VPWR VPWR _4834_/C sky130_fd_sc_hd__o31a_2
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_170 input22/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_181 wire350/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_192 _4232_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4761_ _4965_/B _4832_/A VGND VGND VPWR VPWR _5073_/B sky130_fd_sc_hd__nor2_1
XFILLER_21_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4692_ _4711_/A _4758_/A _4692_/C VGND VGND VPWR VPWR _5035_/A sky130_fd_sc_hd__and3_1
XFILLER_119_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6500_ _6810_/CLK _6500_/D fanout853/X VGND VGND VPWR VPWR _6500_/Q sky130_fd_sc_hd__dfstp_4
X_3712_ wire478/X hold97/A _5200_/A _6806_/Q wire366/X VGND VGND VPWR VPWR _3717_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3643_ input26/X _3283_/Y _4190_/A _6656_/Q VGND VGND VPWR VPWR _3643_/X sky130_fd_sc_hd__a22o_1
X_6431_ _6446_/A _6447_/B VGND VGND VPWR VPWR _6431_/X sky130_fd_sc_hd__and2_1
XFILLER_161_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6362_ _6704_/D _6362_/B VGND VGND VPWR VPWR _6370_/S sky130_fd_sc_hd__and2_4
X_3574_ _7152_/Q hold65/A _5558_/A _7120_/Q VGND VGND VPWR VPWR _3574_/X sky130_fd_sc_hd__a22o_1
X_5313_ _5601_/A0 hold206/X _5314_/S VGND VGND VPWR VPWR _5313_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6293_ _6626_/Q _6028_/X _6293_/B1 _6725_/Q _6292_/X VGND VGND VPWR VPWR _6293_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_115_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5244_ _5247_/A0 hold541/X _5244_/S VGND VGND VPWR VPWR _5244_/X sky130_fd_sc_hd__mux2_1
X_5175_ _5175_/A _5175_/B _5175_/C _5175_/D VGND VGND VPWR VPWR _5175_/X sky130_fd_sc_hd__or4_4
Xhold18 hold18/A VGND VGND VPWR VPWR hold18/X sky130_fd_sc_hd__bufbuf_16
Xhold29 hold29/A VGND VGND VPWR VPWR hold29/X sky130_fd_sc_hd__bufbuf_16
X_4126_ hold446/X wire794/A _4129_/S VGND VGND VPWR VPWR _6600_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4057_ _5247_/A0 hold526/X _4060_/S VGND VGND VPWR VPWR _6541_/D sky130_fd_sc_hd__mux2_1
XFILLER_45_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4959_ _4959_/A _4959_/B VGND VGND VPWR VPWR _4959_/X sky130_fd_sc_hd__and2_2
XFILLER_177_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6629_ _6633_/CLK _6629_/D fanout872/X VGND VGND VPWR VPWR _6629_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_193_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire441 _6146_/X VGND VGND VPWR VPWR wire441/X sky130_fd_sc_hd__buf_4
XFILLER_129_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire430 _5495_/A VGND VGND VPWR VPWR wire430/X sky130_fd_sc_hd__buf_6
XFILLER_51_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire474 _7128_/Q VGND VGND VPWR VPWR _3206_/A sky130_fd_sc_hd__buf_6
Xwire485 _7096_/Q VGND VGND VPWR VPWR wire485/X sky130_fd_sc_hd__buf_6
XFILLER_116_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire463 _3935_/X VGND VGND VPWR VPWR wire463/X sky130_fd_sc_hd__buf_6
Xwire452 hold44/X VGND VGND VPWR VPWR hold45/A sky130_fd_sc_hd__buf_8
Xwire496 _7064_/Q VGND VGND VPWR VPWR wire496/X sky130_fd_sc_hd__buf_6
XFILLER_171_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3290_ hold95/X _3343_/A VGND VGND VPWR VPWR hold96/A sky130_fd_sc_hd__or2_4
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6980_ _6980_/CLK _6980_/D fanout884/X VGND VGND VPWR VPWR _6980_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_38_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5931_ _6542_/Q _5931_/A2 _5930_/X wire671/X VGND VGND VPWR VPWR _5931_/X sky130_fd_sc_hd__a22o_4
XFILLER_81_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5862_ _7068_/Q _5669_/X _5692_/X _7076_/Q VGND VGND VPWR VPWR _5862_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4813_ _4395_/D _4470_/B _4656_/X _4494_/Y VGND VGND VPWR VPWR _4814_/C sky130_fd_sc_hd__a31o_1
X_5793_ _7001_/Q _5667_/X _5792_/X VGND VGND VPWR VPWR _5796_/C sky130_fd_sc_hd__a21o_1
XFILLER_33_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4744_ _4672_/A _4566_/A _4745_/B _4742_/X _4743_/X VGND VGND VPWR VPWR _4753_/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_193_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4675_ _4719_/B _4692_/C _4696_/B VGND VGND VPWR VPWR _4748_/B sky130_fd_sc_hd__and3_4
X_3626_ _6919_/Q _5333_/A _4061_/A _6547_/Q _3615_/X VGND VGND VPWR VPWR _3629_/B
+ sky130_fd_sc_hd__a221o_1
X_6414_ _6446_/A _6447_/B VGND VGND VPWR VPWR _6414_/X sky130_fd_sc_hd__and2_1
X_6345_ _6554_/Q wire601/X wire580/X _6633_/Q _6344_/X VGND VGND VPWR VPWR _6345_/X
+ sky130_fd_sc_hd__a221o_2
X_3557_ _7048_/Q _5477_/A _4172_/A _6642_/Q VGND VGND VPWR VPWR _3557_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6276_ _6541_/Q wire592/X wire590/X _6564_/Q _6275_/X VGND VGND VPWR VPWR _6281_/B
+ sky130_fd_sc_hd__a221o_1
Xinput108 wb_adr_i[18] VGND VGND VPWR VPWR _4349_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_142_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3488_ _3488_/A _3488_/B _3488_/C _3488_/D VGND VGND VPWR VPWR _3548_/B sky130_fd_sc_hd__or4_2
XFILLER_88_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5227_ _5227_/A _5576_/B VGND VGND VPWR VPWR _5233_/S sky130_fd_sc_hd__nand2_8
Xinput119 wb_adr_i[28] VGND VGND VPWR VPWR _3893_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_130_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5158_ _5158_/A _5158_/B VGND VGND VPWR VPWR _5158_/Y sky130_fd_sc_hd__nor2_1
XFILLER_57_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5089_ _4871_/A _4749_/C _4953_/A VGND VGND VPWR VPWR _5118_/D sky130_fd_sc_hd__a21oi_1
X_4109_ _6586_/Q wire351/X _4111_/S VGND VGND VPWR VPWR _6586_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_81 _4267_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_92 _5734_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_70 _3792_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold307 _6737_/Q VGND VGND VPWR VPWR hold307/X sky130_fd_sc_hd__bufbuf_16
XFILLER_117_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4460_ _4694_/A _4989_/A VGND VGND VPWR VPWR _5003_/A sky130_fd_sc_hd__or2_4
Xhold329 _6960_/Q VGND VGND VPWR VPWR hold329/X sky130_fd_sc_hd__bufbuf_16
Xhold318 _5403_/X VGND VGND VPWR VPWR _6979_/D sky130_fd_sc_hd__bufbuf_16
X_4391_ _4513_/A _4405_/B VGND VGND VPWR VPWR _4988_/A sky130_fd_sc_hd__or2_4
XFILLER_125_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3411_ _6995_/Q _5414_/A _3544_/A2 _6494_/Q _3388_/X VGND VGND VPWR VPWR _3414_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_171_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6130_ _6864_/Q _6179_/A2 _6029_/X _3216_/A _6129_/X VGND VGND VPWR VPWR _6131_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_98_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3342_ _3281_/A hold94/X VGND VGND VPWR VPWR _3342_/Y sky130_fd_sc_hd__nand2b_4
XFILLER_112_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6061_ _5663_/Y _6059_/X _6060_/X wire381/A _7189_/Q VGND VGND VPWR VPWR _7189_/D
+ sky130_fd_sc_hd__a32o_1
X_3273_ _3367_/A hold62/X VGND VGND VPWR VPWR _3365_/A sky130_fd_sc_hd__or2_4
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _5012_/A _5105_/B _5011_/X VGND VGND VPWR VPWR _5016_/A sky130_fd_sc_hd__or3b_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6963_ _7147_/CLK _6963_/D fanout887/X VGND VGND VPWR VPWR _6963_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_53_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6894_ _7128_/CLK _6894_/D _6421_/A VGND VGND VPWR VPWR _6894_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_81_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5914_ _6786_/Q _5980_/A2 wire675/X _6655_/Q _5913_/X VGND VGND VPWR VPWR _5915_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5845_ _7011_/Q wire701/X wire697/X _7019_/Q VGND VGND VPWR VPWR _5845_/X sky130_fd_sc_hd__a22o_2
XFILLER_179_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5776_ _6976_/Q _5676_/X _5702_/X _3236_/A _5775_/X VGND VGND VPWR VPWR _5777_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4727_ _4663_/A _4729_/C _4725_/A VGND VGND VPWR VPWR _4727_/Y sky130_fd_sc_hd__a21oi_2
X_4658_ _4470_/B _4656_/X _4653_/Y _4957_/A _5135_/A VGND VGND VPWR VPWR _4708_/C
+ sky130_fd_sc_hd__a2111o_1
XFILLER_190_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput90 spimemio_flash_io2_oeb VGND VGND VPWR VPWR input90/X sky130_fd_sc_hd__clkbuf_4
XFILLER_162_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3609_ _5234_/A hold44/X VGND VGND VPWR VPWR _5238_/A sky130_fd_sc_hd__nor2_8
Xhold830 _6750_/Q VGND VGND VPWR VPWR hold830/X sky130_fd_sc_hd__bufbuf_16
XFILLER_190_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4589_ _4593_/A _4693_/B VGND VGND VPWR VPWR _4590_/B sky130_fd_sc_hd__nand2_1
Xhold841 _6691_/Q VGND VGND VPWR VPWR hold841/X sky130_fd_sc_hd__bufbuf_16
XFILLER_107_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold852 _7081_/Q VGND VGND VPWR VPWR hold852/X sky130_fd_sc_hd__bufbuf_16
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6328_ _6637_/Q wire712/X wire625/X _6612_/Q VGND VGND VPWR VPWR _6328_/X sky130_fd_sc_hd__a22o_1
XFILLER_107_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6259_ _5611_/A _7196_/Q wire381/A VGND VGND VPWR VPWR _6259_/X sky130_fd_sc_hd__a21o_2
XFILLER_190_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3960_ _3960_/A VGND VGND VPWR VPWR _3960_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3891_ _4345_/A _4345_/B VGND VGND VPWR VPWR _4722_/B sky130_fd_sc_hd__or2_4
XFILLER_189_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5630_ _5633_/B VGND VGND VPWR VPWR _5630_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5561_ wire780/A hold527/X _5566_/S VGND VGND VPWR VPWR _5561_/X sky130_fd_sc_hd__mux2_1
X_4512_ _4513_/A _4513_/B VGND VGND VPWR VPWR _4624_/B sky130_fd_sc_hd__nor2_8
X_5492_ _5600_/A0 hold433/X _5494_/S VGND VGND VPWR VPWR _7058_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold115 _4067_/Y VGND VGND VPWR VPWR _4072_/S sky130_fd_sc_hd__bufbuf_16
Xhold104 wire438/X VGND VGND VPWR VPWR _5486_/A sky130_fd_sc_hd__bufbuf_16
XFILLER_117_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold126 _3277_/Y VGND VGND VPWR VPWR _3278_/B sky130_fd_sc_hd__bufbuf_16
Xhold137 _4025_/Y VGND VGND VPWR VPWR _4033_/S sky130_fd_sc_hd__bufbuf_16
X_4443_ _4958_/B _4444_/B VGND VGND VPWR VPWR _4443_/X sky130_fd_sc_hd__and2_4
Xhold148 hold160/X VGND VGND VPWR VPWR hold161/A sky130_fd_sc_hd__bufbuf_16
Xhold159 _4116_/X VGND VGND VPWR VPWR _6592_/D sky130_fd_sc_hd__bufbuf_16
X_4374_ _4507_/A _4992_/A VGND VGND VPWR VPWR _4400_/A sky130_fd_sc_hd__nand2_4
X_7162_ _3949_/A1 _7162_/D fanout879/X VGND VGND VPWR VPWR _7162_/Q sky130_fd_sc_hd__dfstp_4
X_6113_ _3214_/A wire648/X wire639/X _6880_/Q VGND VGND VPWR VPWR _6131_/A sky130_fd_sc_hd__a22o_1
XFILLER_113_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7093_ _7105_/CLK _7093_/D fanout862/X VGND VGND VPWR VPWR _7093_/Q sky130_fd_sc_hd__dfstp_1
X_3325_ _3353_/B _3355_/B VGND VGND VPWR VPWR _3325_/Y sky130_fd_sc_hd__nor2_8
X_6044_ _6917_/Q _6022_/D wire612/X wire503/X VGND VGND VPWR VPWR _6044_/X sky130_fd_sc_hd__a22o_1
XFILLER_85_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3256_ hold124/X _3845_/A hold338/X VGND VGND VPWR VPWR _3256_/Y sky130_fd_sc_hd__a21oi_4
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6946_ _7082_/CLK _6946_/D fanout870/X VGND VGND VPWR VPWR _6946_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_54_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6877_ _7153_/CLK _6877_/D fanout881/X VGND VGND VPWR VPWR _6877_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_169_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5828_ wire556/X _5698_/Y _5826_/X _5827_/X _3921_/A VGND VGND VPWR VPWR _5828_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_155_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5759_ _6903_/Q wire684/X _5707_/X wire515/X VGND VGND VPWR VPWR _5759_/X sky130_fd_sc_hd__a22o_1
XFILLER_147_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold671 _6803_/Q VGND VGND VPWR VPWR hold671/X sky130_fd_sc_hd__bufbuf_16
Xhold660 _7047_/Q VGND VGND VPWR VPWR wire507/A sky130_fd_sc_hd__bufbuf_16
XFILLER_131_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold693 _6625_/Q VGND VGND VPWR VPWR hold693/X sky130_fd_sc_hd__bufbuf_16
XFILLER_104_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold682 _7028_/Q VGND VGND VPWR VPWR hold682/X sky130_fd_sc_hd__bufbuf_16
XFILLER_76_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput209 _3234_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[6] sky130_fd_sc_hd__buf_8
XFILLER_4_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4090_ _6569_/Q _3727_/X _4096_/S VGND VGND VPWR VPWR _6569_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6800_ _6806_/CLK _6800_/D _6435_/A VGND VGND VPWR VPWR _6800_/Q sky130_fd_sc_hd__dfrtp_2
X_4992_ _4992_/A _4992_/B VGND VGND VPWR VPWR _4992_/Y sky130_fd_sc_hd__nand2_2
XFILLER_90_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6731_ _6771_/CLK _6731_/D fanout855/X VGND VGND VPWR VPWR _6731_/Q sky130_fd_sc_hd__dfrtp_2
X_3943_ _6475_/Q _3202_/Y _6473_/Q VGND VGND VPWR VPWR _3943_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_177_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3874_ wire903/X hold49/A _3874_/S VGND VGND VPWR VPWR _6460_/D sky130_fd_sc_hd__mux2_1
X_6662_ _6752_/CLK _6662_/D fanout857/X VGND VGND VPWR VPWR _6662_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5613_ _3920_/Y _5610_/Y _5612_/Y _5605_/Y _7158_/Q VGND VGND VPWR VPWR _7158_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_191_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6593_ _6650_/CLK _6593_/D fanout858/X VGND VGND VPWR VPWR _6593_/Q sky130_fd_sc_hd__dfrtp_2
X_5544_ wire769/X hold559/X _5548_/S VGND VGND VPWR VPWR _7104_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5475_ wire746/X hold710/X _5476_/S VGND VGND VPWR VPWR _7043_/D sky130_fd_sc_hd__mux2_1
X_7214_ _7218_/CLK _7214_/D wire915/X VGND VGND VPWR VPWR hold79/A sky130_fd_sc_hd__dfrtp_2
X_4426_ _4426_/A _4776_/A VGND VGND VPWR VPWR _4428_/C sky130_fd_sc_hd__nor2_2
XFILLER_160_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7145_ _7145_/CLK _7145_/D fanout883/X VGND VGND VPWR VPWR _7145_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_160_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4357_ _4372_/B _4372_/C VGND VGND VPWR VPWR _4484_/B sky130_fd_sc_hd__nand2_1
XFILLER_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4288_ _6408_/A0 hold557/X _4291_/S VGND VGND VPWR VPWR _4288_/X sky130_fd_sc_hd__mux2_1
X_3308_ _3672_/A VGND VGND VPWR VPWR _3308_/Y sky130_fd_sc_hd__inv_2
X_7076_ _7132_/CLK _7076_/D fanout868/X VGND VGND VPWR VPWR _7076_/Q sky130_fd_sc_hd__dfrtp_2
X_6027_ _6037_/C _6027_/B _6027_/C _6027_/D VGND VGND VPWR VPWR _6027_/X sky130_fd_sc_hd__or4_2
XFILLER_86_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3239_ _6856_/Q VGND VGND VPWR VPWR _3239_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_31_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7153_/CLK sky130_fd_sc_hd__clkbuf_8
X_6929_ _7153_/CLK _6929_/D fanout882/X VGND VGND VPWR VPWR _6929_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_168_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire815 _6706_/Q VGND VGND VPWR VPWR _4236_/A sky130_fd_sc_hd__buf_8
XFILLER_22_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire837 wire838/X VGND VGND VPWR VPWR wire837/X sky130_fd_sc_hd__buf_6
Xwire826 _6476_/Q VGND VGND VPWR VPWR _3939_/S sky130_fd_sc_hd__buf_6
XFILLER_10_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_46_csclk _6987_/CLK VGND VGND VPWR VPWR _6985_/CLK sky130_fd_sc_hd__clkbuf_8
Xmax_length468 _3552_/B VGND VGND VPWR VPWR _5252_/A sky130_fd_sc_hd__buf_8
XFILLER_89_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold490 _5260_/X VGND VGND VPWR VPWR _6852_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_151_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_1_0_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_89_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_352 hold32/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_341 hold691/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_330 _3877_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3590_ _6808_/Q _5200_/A _3551_/Y wire836/X _3559_/X VGND VGND VPWR VPWR _3593_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_126_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5260_ wire739/A hold489/X _5260_/S VGND VGND VPWR VPWR _5260_/X sky130_fd_sc_hd__mux2_1
X_4211_ hold310/X _5599_/A0 hold46/X VGND VGND VPWR VPWR _4211_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5191_ _5191_/A _6406_/B VGND VGND VPWR VPWR _5193_/S sky130_fd_sc_hd__nand2_1
X_4142_ _4142_/A _4154_/B VGND VGND VPWR VPWR _4147_/S sky130_fd_sc_hd__nand2_8
XFILLER_96_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4073_ _6702_/Q _6362_/B VGND VGND VPWR VPWR _4081_/S sky130_fd_sc_hd__and2_4
XFILLER_56_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4975_ _5075_/A _5075_/C _4975_/C VGND VGND VPWR VPWR _4976_/B sky130_fd_sc_hd__or3_1
X_6714_ _6747_/CLK _6714_/D fanout874/X VGND VGND VPWR VPWR _6714_/Q sky130_fd_sc_hd__dfrtp_2
X_3926_ _3196_/Y _3898_/Y _3843_/B _6667_/Q VGND VGND VPWR VPWR _6666_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_51_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6645_ _6724_/CLK _6645_/D fanout858/X VGND VGND VPWR VPWR _6645_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3857_ _3841_/B _6664_/Q _3857_/C _3857_/D VGND VGND VPWR VPWR _3864_/B sky130_fd_sc_hd__and4b_4
XFILLER_50_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6576_ _6621_/CLK _6576_/D fanout872/X VGND VGND VPWR VPWR _6576_/Q sky130_fd_sc_hd__dfrtp_2
X_3788_ wire503/X _3298_/Y _4184_/A _6649_/Q _3787_/X VGND VGND VPWR VPWR _3792_/B
+ sky130_fd_sc_hd__a221o_4
XFILLER_192_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5527_ _5572_/A0 hold523/X _5530_/S VGND VGND VPWR VPWR _7089_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5458_ wire739/X hold682/X _5458_/S VGND VGND VPWR VPWR _7028_/D sky130_fd_sc_hd__mux2_1
X_5389_ hold38/X _6966_/Q _5395_/S VGND VGND VPWR VPWR _5389_/X sky130_fd_sc_hd__mux2_1
X_4409_ _4513_/B _4410_/D VGND VGND VPWR VPWR _4409_/Y sky130_fd_sc_hd__nor2_4
XFILLER_132_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7128_ _7128_/CLK hold92/X _6420_/A VGND VGND VPWR VPWR _7128_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7059_ _7154_/CLK _7059_/D fanout884/X VGND VGND VPWR VPWR _7059_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_86_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire623 _6022_/C VGND VGND VPWR VPWR wire623/X sky130_fd_sc_hd__buf_8
Xwire612 _6032_/X VGND VGND VPWR VPWR wire612/X sky130_fd_sc_hd__buf_8
Xwire634 _6025_/C VGND VGND VPWR VPWR wire634/X sky130_fd_sc_hd__buf_8
Xwire601 _6020_/A VGND VGND VPWR VPWR wire601/X sky130_fd_sc_hd__buf_8
XFILLER_11_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire645 wire646/X VGND VGND VPWR VPWR wire645/X sky130_fd_sc_hd__buf_8
Xwire667 wire667/A VGND VGND VPWR VPWR wire667/X sky130_fd_sc_hd__buf_6
Xwire656 wire656/A VGND VGND VPWR VPWR wire656/X sky130_fd_sc_hd__buf_6
XFILLER_7_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire689 _5687_/X VGND VGND VPWR VPWR wire689/X sky130_fd_sc_hd__buf_8
Xwire678 _5692_/X VGND VGND VPWR VPWR wire678/X sky130_fd_sc_hd__buf_8
XFILLER_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_160 wb_clk_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_193 wire438/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_171 input16/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_182 wire353/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4760_ _4947_/B _4832_/A VGND VGND VPWR VPWR _5047_/B sky130_fd_sc_hd__nor2_1
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3711_ input53/X _4025_/A _4209_/S input44/X VGND VGND VPWR VPWR _3711_/X sky130_fd_sc_hd__a22o_4
X_4691_ _4746_/B _4707_/B _5050_/A VGND VGND VPWR VPWR _4756_/B sky130_fd_sc_hd__or3b_4
XFILLER_159_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3642_ wire501/X _3298_/Y _3384_/Y _6828_/Q _3641_/X VGND VGND VPWR VPWR _3645_/C
+ sky130_fd_sc_hd__a221o_1
X_6430_ _6455_/A _6455_/B VGND VGND VPWR VPWR _6430_/X sky130_fd_sc_hd__and2_1
XFILLER_174_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6361_ _7202_/Q _3896_/Y _6360_/Y _3916_/B _6704_/D VGND VGND VPWR VPWR _7202_/D
+ sky130_fd_sc_hd__a32o_1
X_5312_ _5600_/A0 hold432/X _5314_/S VGND VGND VPWR VPWR _6898_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3573_ _6960_/Q _3305_/Y wire388/X wire557/X _3572_/X VGND VGND VPWR VPWR _3578_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_154_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6292_ wire469/X _6009_/X _6020_/D _6710_/Q VGND VGND VPWR VPWR _6292_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5243_ wire799/A hold588/X _5244_/S VGND VGND VPWR VPWR _6837_/D sky130_fd_sc_hd__mux2_1
Xhold19 hold19/A VGND VGND VPWR VPWR hold19/X sky130_fd_sc_hd__bufbuf_16
X_5174_ _5174_/A _5174_/B _5174_/C _5174_/D VGND VGND VPWR VPWR _5175_/D sky130_fd_sc_hd__or4_1
XFILLER_114_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4125_ hold774/X _5487_/A0 _4129_/S VGND VGND VPWR VPWR _6599_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4056_ _5487_/A0 hold785/X _4060_/S VGND VGND VPWR VPWR _6540_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4958_ _4958_/A _4958_/B VGND VGND VPWR VPWR _4959_/B sky130_fd_sc_hd__nor2_4
XFILLER_61_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4889_ _5005_/C _4832_/A _4575_/Y VGND VGND VPWR VPWR _5073_/C sky130_fd_sc_hd__o21ai_2
X_3909_ _5611_/A _3921_/B VGND VGND VPWR VPWR _3909_/Y sky130_fd_sc_hd__nand2_1
XFILLER_165_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6628_ _6632_/CLK _6628_/D fanout872/X VGND VGND VPWR VPWR _6628_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6559_ _7208_/CLK _6559_/D VGND VGND VPWR VPWR _6559_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_193_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire431 hold97/X VGND VGND VPWR VPWR _5549_/A sky130_fd_sc_hd__buf_8
Xwire442 _3947_/X VGND VGND VPWR VPWR wire442/X sky130_fd_sc_hd__buf_6
XFILLER_11_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire475 _7122_/Q VGND VGND VPWR VPWR wire475/X sky130_fd_sc_hd__buf_6
XFILLER_156_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire464 wire465/X VGND VGND VPWR VPWR wire464/X sky130_fd_sc_hd__buf_6
Xwire453 _3672_/A VGND VGND VPWR VPWR _4034_/A sky130_fd_sc_hd__buf_8
XFILLER_171_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire486 _7095_/Q VGND VGND VPWR VPWR wire486/X sky130_fd_sc_hd__buf_6
XFILLER_124_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5930_ _6626_/Q _5963_/B VGND VGND VPWR VPWR _5930_/X sky130_fd_sc_hd__or2_1
XFILLER_65_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5861_ _5861_/A _5861_/B _5861_/C _5861_/D VGND VGND VPWR VPWR _5861_/X sky130_fd_sc_hd__or4_2
XFILLER_33_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4812_ _4812_/A _5005_/A _4812_/C VGND VGND VPWR VPWR _4812_/X sky130_fd_sc_hd__or3_4
XFILLER_178_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5792_ wire539/X _5689_/X wire656/A _6945_/Q VGND VGND VPWR VPWR _5792_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4743_ _4488_/X _4724_/A _4724_/B _4819_/B VGND VGND VPWR VPWR _4743_/X sky130_fd_sc_hd__a211o_1
XFILLER_166_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4674_ _4745_/A _4832_/A VGND VGND VPWR VPWR _5047_/A sky130_fd_sc_hd__nor2_2
X_6413_ _6446_/A _6447_/B VGND VGND VPWR VPWR _6413_/X sky130_fd_sc_hd__and2_1
X_3625_ _6951_/Q _5369_/A wire390/X _6720_/Q _3610_/X VGND VGND VPWR VPWR _3629_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_135_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3556_ _7056_/Q wire438/X _3638_/B1 _7080_/Q VGND VGND VPWR VPWR _3556_/X sky130_fd_sc_hd__a22o_4
X_6344_ _6767_/Q wire649/X wire594/X _6722_/Q VGND VGND VPWR VPWR _6344_/X sky130_fd_sc_hd__a22o_4
XFILLER_103_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6275_ _6620_/Q wire623/X wire612/X _6650_/Q VGND VGND VPWR VPWR _6275_/X sky130_fd_sc_hd__a22o_1
Xinput109 wb_adr_i[19] VGND VGND VPWR VPWR _4349_/C sky130_fd_sc_hd__clkbuf_4
X_3487_ _7113_/Q _5549_/A _5369_/A _6953_/Q _3486_/X VGND VGND VPWR VPWR _3488_/D
+ sky130_fd_sc_hd__a221o_4
XFILLER_115_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5226_ hold800/X _3735_/Y _5576_/B _5225_/X VGND VGND VPWR VPWR _6825_/D sky130_fd_sc_hd__o211a_1
XFILLER_130_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5157_ _5157_/A _5157_/B _5157_/C VGND VGND VPWR VPWR _5158_/B sky130_fd_sc_hd__or3_4
XFILLER_84_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5088_ _4507_/A _5087_/X _4985_/Y VGND VGND VPWR VPWR _5140_/C sky130_fd_sc_hd__a21bo_4
X_4108_ _6585_/Q _4108_/A1 _4111_/S VGND VGND VPWR VPWR _6585_/D sky130_fd_sc_hd__mux2_1
X_4039_ hold150/X hold843/X hold73/X VGND VGND VPWR VPWR _4039_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_82 _4566_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_93 _5784_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_60 _3687_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_71 _3801_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_670 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold308 _6613_/Q VGND VGND VPWR VPWR hold308/X sky130_fd_sc_hd__bufbuf_16
XFILLER_117_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4390_ _4513_/A _4405_/B VGND VGND VPWR VPWR _4622_/B sky130_fd_sc_hd__nor2_8
X_3410_ _6931_/Q wire436/X _5387_/A _6971_/Q _3409_/X VGND VGND VPWR VPWR _3414_/B
+ sky130_fd_sc_hd__a221o_4
Xhold319 _6630_/Q VGND VGND VPWR VPWR hold319/X sky130_fd_sc_hd__bufbuf_16
XFILLER_98_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3341_ _3508_/A _5225_/B VGND VGND VPWR VPWR _5531_/A sky130_fd_sc_hd__nor2_8
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6060_ _6853_/Q _6060_/B VGND VGND VPWR VPWR _6060_/X sky130_fd_sc_hd__or2_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ hold61/X _3281_/B VGND VGND VPWR VPWR hold62/A sky130_fd_sc_hd__or2_4
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5011_ _5005_/C _4832_/B _5144_/B _5010_/X VGND VGND VPWR VPWR _5011_/X sky130_fd_sc_hd__o211a_1
XFILLER_97_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6962_ _7154_/CLK _6962_/D fanout887/X VGND VGND VPWR VPWR _6962_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_179_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6893_ _7133_/CLK _6893_/D fanout881/X VGND VGND VPWR VPWR _6893_/Q sky130_fd_sc_hd__dfstp_4
X_5913_ _6749_/Q _5979_/A2 wire662/X _6541_/Q VGND VGND VPWR VPWR _5913_/X sky130_fd_sc_hd__a22o_1
X_5844_ _7035_/Q _5855_/B1 _5856_/A2 _7099_/Q _5843_/X VGND VGND VPWR VPWR _5849_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_61_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5775_ _3214_/A _5921_/A2 _5698_/B _6984_/Q _5697_/X VGND VGND VPWR VPWR _5775_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_175_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4726_ _4740_/B _4832_/A VGND VGND VPWR VPWR _4729_/C sky130_fd_sc_hd__nor2_1
X_4657_ _4692_/C _4657_/B VGND VGND VPWR VPWR _4754_/B sky130_fd_sc_hd__nand2_8
XFILLER_175_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput91 spimemio_flash_io3_do VGND VGND VPWR VPWR input91/X sky130_fd_sc_hd__clkbuf_4
XFILLER_174_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold820 _7107_/Q VGND VGND VPWR VPWR hold820/X sky130_fd_sc_hd__bufbuf_16
Xinput80 spi_sck VGND VGND VPWR VPWR input80/X sky130_fd_sc_hd__clkbuf_4
X_3608_ _3607_/X _6793_/Q _3928_/A VGND VGND VPWR VPWR _6793_/D sky130_fd_sc_hd__mux2_1
XFILLER_190_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold842 _6690_/Q VGND VGND VPWR VPWR hold842/X sky130_fd_sc_hd__bufbuf_16
Xhold853 _6513_/Q VGND VGND VPWR VPWR hold853/X sky130_fd_sc_hd__bufbuf_16
XFILLER_150_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4588_ _4663_/A _4740_/B VGND VGND VPWR VPWR _4588_/X sky130_fd_sc_hd__or2_4
XFILLER_131_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold831 _6708_/Q VGND VGND VPWR VPWR hold831/X sky130_fd_sc_hd__bufbuf_16
XFILLER_122_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6327_ _6543_/Q wire592/X wire590/X _6566_/Q _6310_/X VGND VGND VPWR VPWR _6330_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3539_ _3540_/A _3539_/B VGND VGND VPWR VPWR _4250_/A sky130_fd_sc_hd__nor2_8
XFILLER_107_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6258_ _6530_/Q _6357_/A2 _6248_/X _6257_/X _6308_/S VGND VGND VPWR VPWR _6258_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_67_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5209_ _6812_/Q _5578_/A0 _5215_/S VGND VGND VPWR VPWR _6812_/D sky130_fd_sc_hd__mux2_1
X_6189_ _7083_/Q _6211_/B wire575/X _7019_/Q _6186_/X VGND VGND VPWR VPWR _6194_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_123_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3890_ _4368_/A _4722_/A VGND VGND VPWR VPWR _4529_/A sky130_fd_sc_hd__nand2_4
XFILLER_188_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5560_ wire796/X _7118_/Q _5566_/S VGND VGND VPWR VPWR hold53/A sky130_fd_sc_hd__mux2_1
X_4511_ _4956_/A _4538_/A VGND VGND VPWR VPWR _4953_/A sky130_fd_sc_hd__nand2_8
X_5491_ _5599_/A0 hold312/X _5494_/S VGND VGND VPWR VPWR _5491_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4442_ _4529_/C _4442_/B VGND VGND VPWR VPWR _4444_/B sky130_fd_sc_hd__nand2b_4
Xhold105 _5486_/Y VGND VGND VPWR VPWR _5494_/S sky130_fd_sc_hd__bufbuf_16
Xhold116 _4071_/X VGND VGND VPWR VPWR _6553_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_156_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold138 _4027_/X VGND VGND VPWR VPWR _6515_/D sky130_fd_sc_hd__bufbuf_16
Xhold149 hold163/X VGND VGND VPWR VPWR hold154/A sky130_fd_sc_hd__bufbuf_16
XFILLER_171_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold127 _3293_/Y VGND VGND VPWR VPWR _3304_/B sky130_fd_sc_hd__bufbuf_16
XFILLER_172_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4373_ _4655_/A _4478_/C VGND VGND VPWR VPWR _4992_/A sky130_fd_sc_hd__nor2_8
XFILLER_98_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7161_ _7194_/CLK _7161_/D fanout868/X VGND VGND VPWR VPWR _7161_/Q sky130_fd_sc_hd__dfrtp_2
X_6112_ _7136_/Q wire643/X wire631/X wire485/X VGND VGND VPWR VPWR _6112_/X sky130_fd_sc_hd__a22o_1
X_3324_ hold96/A _3543_/A VGND VGND VPWR VPWR _3324_/Y sky130_fd_sc_hd__nor2_4
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7092_ _7095_/CLK _7092_/D fanout862/X VGND VGND VPWR VPWR _7092_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_140_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6043_ _6997_/Q wire604/X _6139_/A2 _7013_/Q _6042_/X VGND VGND VPWR VPWR _6059_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ _3845_/A _3255_/B VGND VGND VPWR VPWR _3255_/X sky130_fd_sc_hd__and2b_2
XFILLER_85_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6945_ _7140_/CLK _6945_/D fanout862/X VGND VGND VPWR VPWR _6945_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_42_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
X_6876_ _7152_/CLK _6876_/D fanout886/X VGND VGND VPWR VPWR _6876_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5827_ _5827_/A _5827_/B _5827_/C VGND VGND VPWR VPWR _5827_/X sky130_fd_sc_hd__or3_1
XFILLER_50_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5758_ _6999_/Q _5667_/X _5803_/B1 _7039_/Q _5757_/X VGND VGND VPWR VPWR _5763_/B
+ sky130_fd_sc_hd__a221o_1
Xmax_length617 wire618/X VGND VGND VPWR VPWR _6352_/B1 sky130_fd_sc_hd__buf_6
XFILLER_185_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4709_ _4436_/B _5165_/A _4702_/A _4704_/X _4708_/X VGND VGND VPWR VPWR _4713_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_154_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5689_ _5864_/B _5704_/B _5707_/C VGND VGND VPWR VPWR _5689_/X sky130_fd_sc_hd__and3_4
XFILLER_162_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold650 _6772_/Q VGND VGND VPWR VPWR hold650/X sky130_fd_sc_hd__bufbuf_16
Xhold672 _7020_/Q VGND VGND VPWR VPWR hold672/X sky130_fd_sc_hd__bufbuf_16
Xhold661 _7015_/Q VGND VGND VPWR VPWR hold661/X sky130_fd_sc_hd__bufbuf_16
Xhold683 _6620_/Q VGND VGND VPWR VPWR hold683/X sky130_fd_sc_hd__bufbuf_16
XFILLER_104_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold694 _6749_/Q VGND VGND VPWR VPWR hold694/X sky130_fd_sc_hd__bufbuf_16
XFILLER_103_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4991_ _4818_/A _4672_/A _4566_/A _4648_/B VGND VGND VPWR VPWR _4991_/X sky130_fd_sc_hd__a211o_2
XFILLER_91_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6730_ _6771_/CLK _6730_/D fanout854/X VGND VGND VPWR VPWR _6730_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3942_ _6475_/Q _3942_/B VGND VGND VPWR VPWR _3942_/X sky130_fd_sc_hd__or2_1
X_3873_ hold49/A hold5/A _3874_/S VGND VGND VPWR VPWR _6461_/D sky130_fd_sc_hd__mux2_1
XFILLER_149_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6661_ _6752_/CLK _6661_/D fanout857/X VGND VGND VPWR VPWR _6661_/Q sky130_fd_sc_hd__dfstp_4
X_6592_ _6623_/CLK _6592_/D fanout890/X VGND VGND VPWR VPWR _6592_/Q sky130_fd_sc_hd__dfrtp_2
X_5612_ _5612_/A _5612_/B VGND VGND VPWR VPWR _5612_/Y sky130_fd_sc_hd__nor2_1
XFILLER_164_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5543_ wire780/X hold618/X _5548_/S VGND VGND VPWR VPWR _5543_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5474_ _5519_/A0 hold835/X _5476_/S VGND VGND VPWR VPWR _7042_/D sky130_fd_sc_hd__mux2_1
X_7213_ _7218_/CLK _7213_/D wire915/X VGND VGND VPWR VPWR hold9/A sky130_fd_sc_hd__dfrtp_4
XFILLER_172_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4425_ _4422_/Y _4423_/X _4424_/Y _4414_/B VGND VGND VPWR VPWR _4776_/A sky130_fd_sc_hd__a211o_4
XFILLER_144_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7144_ _7152_/CLK _7144_/D fanout888/X VGND VGND VPWR VPWR _7144_/Q sky130_fd_sc_hd__dfrtp_2
X_4356_ _4722_/A _4529_/B _4486_/B VGND VGND VPWR VPWR _4372_/C sky130_fd_sc_hd__nand3b_4
XFILLER_132_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3307_ hold62/X _3343_/A VGND VGND VPWR VPWR _3355_/B sky130_fd_sc_hd__or2_4
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7075_ _7082_/CLK _7075_/D fanout870/X VGND VGND VPWR VPWR _7075_/Q sky130_fd_sc_hd__dfrtp_2
X_4287_ _6407_/A0 _6738_/Q _4291_/S VGND VGND VPWR VPWR _4287_/X sky130_fd_sc_hd__mux2_1
X_6026_ _6037_/C _6027_/B _6027_/C _6027_/D VGND VGND VPWR VPWR _6232_/A sky130_fd_sc_hd__nor4_4
XFILLER_100_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3238_ _3238_/A VGND VGND VPWR VPWR _3238_/Y sky130_fd_sc_hd__inv_2
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6928_ _6930_/CLK _6928_/D fanout887/X VGND VGND VPWR VPWR _6928_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_167_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6859_ _7042_/CLK _6859_/D fanout865/X VGND VGND VPWR VPWR _6859_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_168_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire816 _6705_/Q VGND VGND VPWR VPWR _4236_/B sky130_fd_sc_hd__buf_8
XFILLER_167_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length425 _3582_/A2 VGND VGND VPWR VPWR _5333_/A sky130_fd_sc_hd__buf_6
Xwire827 _6475_/Q VGND VGND VPWR VPWR _3938_/S sky130_fd_sc_hd__buf_6
XFILLER_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire838 wire838/A VGND VGND VPWR VPWR wire838/X sky130_fd_sc_hd__buf_6
Xmax_length414 _3338_/Y VGND VGND VPWR VPWR _3443_/A2 sky130_fd_sc_hd__buf_6
XFILLER_136_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length447 _3371_/Y VGND VGND VPWR VPWR wire446/A sky130_fd_sc_hd__buf_6
XFILLER_163_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold480 _7122_/Q VGND VGND VPWR VPWR hold480/X sky130_fd_sc_hd__bufbuf_16
XFILLER_151_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold491 _6826_/Q VGND VGND VPWR VPWR hold491/X sky130_fd_sc_hd__bufbuf_16
XFILLER_77_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_342 hold847/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_331 _3973_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_320 wire739/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_353 hold465/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_3_0_mgmt_gpio_in[4] clkbuf_2_3_0_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR _3938_/A1
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_173_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4210_ hold750/X _4209_/X _4218_/S VGND VGND VPWR VPWR _4210_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5190_ _6411_/A0 hold625/X _5190_/S VGND VGND VPWR VPWR _6789_/D sky130_fd_sc_hd__mux2_1
X_4141_ _5599_/A0 hold308/X _4141_/S VGND VGND VPWR VPWR _6613_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4072_ _4303_/A0 hold439/X _4072_/S VGND VGND VPWR VPWR _6554_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4974_ _4974_/A _5145_/B _5073_/D _4974_/D VGND VGND VPWR VPWR _4975_/C sky130_fd_sc_hd__or4_1
X_6713_ _6747_/CLK _6713_/D fanout874/X VGND VGND VPWR VPWR _6713_/Q sky130_fd_sc_hd__dfrtp_2
X_3925_ _6667_/Q _3898_/A _3924_/X VGND VGND VPWR VPWR _6667_/D sky130_fd_sc_hd__a21bo_1
XFILLER_165_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6644_ _6646_/CLK _6644_/D fanout856/X VGND VGND VPWR VPWR _6644_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_177_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3856_ _3875_/B _6470_/Q _3856_/S VGND VGND VPWR VPWR _6470_/D sky130_fd_sc_hd__mux2_1
XFILLER_164_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3787_ _6853_/Q _5261_/A _5238_/A _6836_/Q VGND VGND VPWR VPWR _3787_/X sky130_fd_sc_hd__a22o_2
X_6575_ _7210_/CLK _6575_/D VGND VGND VPWR VPWR _6575_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_117_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5526_ wire769/X hold599/X _5530_/S VGND VGND VPWR VPWR _7088_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5457_ wire749/X hold395/X _5458_/S VGND VGND VPWR VPWR _7027_/D sky130_fd_sc_hd__mux2_1
X_4408_ _4408_/A _4408_/B VGND VGND VPWR VPWR _4410_/D sky130_fd_sc_hd__nand2_4
XFILLER_105_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5388_ _5595_/A0 _6965_/Q _5395_/S VGND VGND VPWR VPWR _6965_/D sky130_fd_sc_hd__mux2_1
XFILLER_182_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7127_ _7145_/CLK hold14/X fanout883/X VGND VGND VPWR VPWR _7127_/Q sky130_fd_sc_hd__dfrtp_2
X_4339_ _4696_/A _4413_/C VGND VGND VPWR VPWR _4340_/B sky130_fd_sc_hd__nand2_8
XFILLER_59_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7058_ _7147_/CLK _7058_/D fanout886/X VGND VGND VPWR VPWR _7058_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_59_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6009_ _6037_/B _6037_/C _6032_/C VGND VGND VPWR VPWR _6009_/X sky130_fd_sc_hd__and3_4
XFILLER_86_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire602 _6020_/A VGND VGND VPWR VPWR wire602/X sky130_fd_sc_hd__buf_8
Xwire624 _6022_/C VGND VGND VPWR VPWR wire624/X sky130_fd_sc_hd__buf_8
Xwire613 _6032_/X VGND VGND VPWR VPWR wire613/X sky130_fd_sc_hd__buf_8
XFILLER_183_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire646 _6025_/A VGND VGND VPWR VPWR wire646/X sky130_fd_sc_hd__buf_8
Xwire635 _6025_/C VGND VGND VPWR VPWR wire635/X sky130_fd_sc_hd__buf_8
Xwire657 _5705_/X VGND VGND VPWR VPWR wire657/X sky130_fd_sc_hd__buf_8
XFILLER_10_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire679 _5692_/X VGND VGND VPWR VPWR wire679/X sky130_fd_sc_hd__buf_8
XFILLER_156_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_161 wb_dat_i[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_150 _6828_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_172 input117/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_194 wire450/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_183 wire353/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3710_ _6635_/Q _4166_/A _3701_/X _3709_/X VGND VGND VPWR VPWR _3726_/B sky130_fd_sc_hd__a211o_1
XFILLER_186_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4690_ _4690_/A _4746_/A _5062_/B VGND VGND VPWR VPWR _4757_/B sky130_fd_sc_hd__or3_4
XFILLER_147_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3641_ _6765_/Q _4316_/A _4304_/A _6755_/Q VGND VGND VPWR VPWR _3641_/X sky130_fd_sc_hd__a22o_1
X_3572_ _6607_/Q _4130_/A _4148_/A _6622_/Q VGND VGND VPWR VPWR _3572_/X sky130_fd_sc_hd__a22o_2
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6360_ _6360_/A _6704_/Q VGND VGND VPWR VPWR _6360_/Y sky130_fd_sc_hd__nand2_1
X_5311_ hold150/X hold181/X _5314_/S VGND VGND VPWR VPWR _5311_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6291_ _6755_/Q _6339_/A2 _6339_/B1 _6770_/Q _6290_/X VGND VGND VPWR VPWR _6291_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_102_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5242_ _5242_/A _5242_/B VGND VGND VPWR VPWR _5244_/S sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_30_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7151_/CLK sky130_fd_sc_hd__clkbuf_8
X_5173_ _5120_/C _5171_/X _5172_/Y VGND VGND VPWR VPWR _5184_/A sky130_fd_sc_hd__o21a_1
X_4124_ _4124_/A _5378_/B VGND VGND VPWR VPWR _4129_/S sky130_fd_sc_hd__and2_4
XFILLER_56_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput1 debug_mode VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__clkbuf_4
X_4055_ _4055_/A _4154_/B VGND VGND VPWR VPWR _4060_/S sky130_fd_sc_hd__nand2_8
Xclkbuf_leaf_45_csclk _6987_/CLK VGND VGND VPWR VPWR _7068_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_37_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4957_ _4957_/A _5099_/C _4976_/C VGND VGND VPWR VPWR _5128_/D sky130_fd_sc_hd__or3_1
XFILLER_101_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4888_ _4956_/C _4758_/B _4652_/B _5078_/B VGND VGND VPWR VPWR _4909_/B sky130_fd_sc_hd__a31o_1
XFILLER_20_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3908_ _3921_/A _3920_/B VGND VGND VPWR VPWR _5665_/A sky130_fd_sc_hd__nor2_4
XFILLER_192_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6627_ _6632_/CLK _6627_/D fanout872/X VGND VGND VPWR VPWR _6627_/Q sky130_fd_sc_hd__dfrtp_2
X_3839_ _3191_/Y _3875_/B _3845_/A VGND VGND VPWR VPWR _3839_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6558_ _7208_/CLK _6558_/D VGND VGND VPWR VPWR _6558_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_152_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6489_ _6771_/CLK _6489_/D fanout855/X VGND VGND VPWR VPWR _6489_/Q sky130_fd_sc_hd__dfstp_2
X_5509_ _5572_/A0 hold501/X _5512_/S VGND VGND VPWR VPWR _7073_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire421 wire421/A VGND VGND VPWR VPWR _5387_/A sky130_fd_sc_hd__buf_8
Xwire410 hold64/X VGND VGND VPWR VPWR hold65/A sky130_fd_sc_hd__buf_8
Xwire432 _3310_/Y VGND VGND VPWR VPWR wire432/X sky130_fd_sc_hd__buf_6
Xwire476 _7121_/Q VGND VGND VPWR VPWR wire476/X sky130_fd_sc_hd__buf_6
XFILLER_171_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire443 wire444/X VGND VGND VPWR VPWR wire443/X sky130_fd_sc_hd__buf_6
XFILLER_128_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire465 _3934_/X VGND VGND VPWR VPWR wire465/X sky130_fd_sc_hd__buf_6
Xwire498 _7062_/Q VGND VGND VPWR VPWR wire498/X sky130_fd_sc_hd__buf_6
Xwire487 _7093_/Q VGND VGND VPWR VPWR wire487/X sky130_fd_sc_hd__buf_6
XFILLER_124_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5860_ _7004_/Q _5667_/X _5702_/X _6892_/Q _5859_/X VGND VGND VPWR VPWR _5861_/D
+ sky130_fd_sc_hd__a221o_4
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4811_ _4736_/B _4758_/B _4695_/X _5105_/A _4810_/Y VGND VGND VPWR VPWR _4817_/A
+ sky130_fd_sc_hd__a311o_1
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5791_ _7033_/Q _5688_/X _5702_/X _6889_/Q _5790_/X VGND VGND VPWR VPWR _5796_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4742_ _4740_/A _4740_/B _4832_/B _4740_/X _4881_/B VGND VGND VPWR VPWR _4742_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_147_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4673_ _4697_/A _4832_/A VGND VGND VPWR VPWR _4920_/C sky130_fd_sc_hd__nor2_1
XFILLER_119_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3624_ _6631_/Q _4160_/A _3613_/X _3622_/X _3623_/X VGND VGND VPWR VPWR _3636_/B
+ sky130_fd_sc_hd__a2111o_2
X_6412_ _6446_/A _6447_/B VGND VGND VPWR VPWR _6412_/X sky130_fd_sc_hd__and2_1
XFILLER_174_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3555_ _3202_/A _3310_/Y _4292_/A wire565/X VGND VGND VPWR VPWR _3555_/X sky130_fd_sc_hd__a22o_1
X_6343_ _6343_/A _6343_/B _6343_/C _6343_/D VGND VGND VPWR VPWR _6356_/B sky130_fd_sc_hd__or4_1
XFILLER_142_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6274_ _6577_/Q wire599/X wire645/X _6605_/Q _6273_/X VGND VGND VPWR VPWR _6281_/A
+ sky130_fd_sc_hd__a221o_1
X_3486_ _6549_/Q _4061_/A _4043_/A _6534_/Q VGND VGND VPWR VPWR _3486_/X sky130_fd_sc_hd__a22o_4
X_5225_ _5225_/A _5225_/B _5234_/C VGND VGND VPWR VPWR _5225_/X sky130_fd_sc_hd__or3_1
XFILLER_130_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5156_ _5156_/A _5156_/B _5156_/C VGND VGND VPWR VPWR _5157_/C sky130_fd_sc_hd__or3_1
XFILLER_111_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5087_ _5087_/A _5087_/B _5087_/C _5087_/D VGND VGND VPWR VPWR _5087_/X sky130_fd_sc_hd__or4_4
XFILLER_84_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4107_ _6584_/Q _3606_/X _4111_/S VGND VGND VPWR VPWR _6584_/D sky130_fd_sc_hd__mux2_1
X_4038_ _5598_/A0 hold562/X hold73/X VGND VGND VPWR VPWR _4038_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5989_ _7170_/Q _7171_/Q VGND VGND VPWR VPWR _6014_/A sky130_fd_sc_hd__or2_4
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_50 _3546_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_83 _4575_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_61 _3687_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 _3802_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_94 _5802_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput190 _3217_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[23] sky130_fd_sc_hd__buf_8
XFILLER_153_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold309 _6908_/Q VGND VGND VPWR VPWR hold309/X sky130_fd_sc_hd__bufbuf_16
XFILLER_109_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_4_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A VGND VGND VPWR VPWR _7196_/CLK sky130_fd_sc_hd__clkbuf_8
X_3340_ _6908_/Q _3443_/A2 _5459_/A _7036_/Q VGND VGND VPWR VPWR _3340_/X sky130_fd_sc_hd__a22o_1
XFILLER_152_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _4697_/A _4832_/B _4812_/C _4505_/X VGND VGND VPWR VPWR _5010_/X sky130_fd_sc_hd__o22a_1
X_3271_ hold185/X hold93/X _3953_/A VGND VGND VPWR VPWR _3271_/X sky130_fd_sc_hd__mux2_8
XFILLER_3_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6961_ _7151_/CLK _6961_/D fanout880/X VGND VGND VPWR VPWR _6961_/Q sky130_fd_sc_hd__dfrtp_2
X_6892_ _7152_/CLK _6892_/D fanout882/X VGND VGND VPWR VPWR _6892_/Q sky130_fd_sc_hd__dfrtp_2
X_5912_ _6577_/Q wire684/X _5901_/X _5911_/X VGND VGND VPWR VPWR _5915_/C sky130_fd_sc_hd__a211o_2
XFILLER_53_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5843_ _7059_/Q _5706_/X _5842_/X _5698_/B VGND VGND VPWR VPWR _5843_/X sky130_fd_sc_hd__a22o_4
XFILLER_34_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5774_ _6880_/Q _5674_/X _5688_/X _3218_/A _5773_/X VGND VGND VPWR VPWR _5777_/C
+ sky130_fd_sc_hd__a221o_1
X_4725_ _4725_/A VGND VGND VPWR VPWR _4725_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4656_ _4692_/C _4657_/B VGND VGND VPWR VPWR _4656_/X sky130_fd_sc_hd__and2_4
XFILLER_174_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold810 _6506_/Q VGND VGND VPWR VPWR hold810/X sky130_fd_sc_hd__bufbuf_16
X_4587_ _4663_/A _4740_/B VGND VGND VPWR VPWR _4956_/C sky130_fd_sc_hd__nor2_8
XFILLER_107_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput70 mgmt_gpio_in[7] VGND VGND VPWR VPWR wire894/A sky130_fd_sc_hd__buf_6
Xhold821 _6859_/Q VGND VGND VPWR VPWR hold821/X sky130_fd_sc_hd__bufbuf_16
Xinput81 spi_sdo VGND VGND VPWR VPWR input81/X sky130_fd_sc_hd__clkbuf_4
X_3607_ _3606_/X _6792_/Q _3857_/C VGND VGND VPWR VPWR _3607_/X sky130_fd_sc_hd__mux2_1
Xinput92 spimemio_flash_io3_oeb VGND VGND VPWR VPWR input92/X sky130_fd_sc_hd__clkbuf_4
Xhold843 _6526_/Q VGND VGND VPWR VPWR hold843/X sky130_fd_sc_hd__bufbuf_16
X_3538_ _6865_/Q wire439/X _5387_/A _6969_/Q _3537_/X VGND VGND VPWR VPWR _3546_/B
+ sky130_fd_sc_hd__a221o_4
X_6326_ _6579_/Q wire599/X wire645/X _6607_/Q _6325_/X VGND VGND VPWR VPWR _6331_/C
+ sky130_fd_sc_hd__a221o_4
Xhold832 _6537_/Q VGND VGND VPWR VPWR hold832/X sky130_fd_sc_hd__bufbuf_16
XFILLER_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6257_ _6356_/A _6257_/B _6257_/C _6257_/D VGND VGND VPWR VPWR _6257_/X sky130_fd_sc_hd__or4_1
X_3469_ _6752_/Q _4298_/A _4184_/A _6653_/Q VGND VGND VPWR VPWR _3469_/X sky130_fd_sc_hd__a22o_2
XFILLER_190_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5208_ hold787/X _6407_/A0 _5215_/S VGND VGND VPWR VPWR _6811_/D sky130_fd_sc_hd__mux2_1
X_6188_ _7027_/Q wire589/X wire615/X wire489/X _6187_/X VGND VGND VPWR VPWR _6194_/A
+ sky130_fd_sc_hd__a221o_1
X_5139_ _4400_/A _4410_/D _4997_/B _5138_/Y VGND VGND VPWR VPWR _5139_/X sky130_fd_sc_hd__o31a_1
XFILLER_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4510_ _4534_/B _4510_/B VGND VGND VPWR VPWR _4538_/A sky130_fd_sc_hd__and2_4
XFILLER_184_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5490_ _5598_/A0 hold622/X _5494_/S VGND VGND VPWR VPWR _7056_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold106 _7064_/Q VGND VGND VPWR VPWR hold106/X sky130_fd_sc_hd__bufbuf_16
X_4441_ _4654_/A _4696_/A _4446_/B _4958_/A VGND VGND VPWR VPWR _4442_/B sky130_fd_sc_hd__a31o_2
XFILLER_144_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold117 hold342/X VGND VGND VPWR VPWR hold117/X sky130_fd_sc_hd__bufbuf_16
X_7160_ _7194_/CLK _7160_/D fanout866/X VGND VGND VPWR VPWR _7160_/Q sky130_fd_sc_hd__dfrtp_2
Xhold139 _6456_/Q VGND VGND VPWR VPWR hold29/A sky130_fd_sc_hd__bufbuf_16
Xhold128 _3304_/X VGND VGND VPWR VPWR _3369_/A sky130_fd_sc_hd__bufbuf_16
X_4372_ _4533_/A _4372_/B _4372_/C _4484_/C VGND VGND VPWR VPWR _4410_/C sky130_fd_sc_hd__nand4b_4
XFILLER_171_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6111_ _7080_/Q _6111_/B VGND VGND VPWR VPWR _6111_/X sky130_fd_sc_hd__and2_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7091_ _7091_/CLK _7091_/D fanout867/X VGND VGND VPWR VPWR _7091_/Q sky130_fd_sc_hd__dfrtp_2
X_3323_ input10/X _3320_/Y _3322_/Y wire900/X _3318_/X VGND VGND VPWR VPWR _3331_/C
+ sky130_fd_sc_hd__a221o_1
X_6042_ wire483/X wire711/X _6028_/X _6981_/Q VGND VGND VPWR VPWR _6042_/X sky130_fd_sc_hd__a22o_1
XFILLER_112_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3254_ hold332/X hold189/X _3953_/A VGND VGND VPWR VPWR _3254_/X sky130_fd_sc_hd__mux2_8
XFILLER_85_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6944_ _7068_/CLK _6944_/D fanout878/X VGND VGND VPWR VPWR _6944_/Q sky130_fd_sc_hd__dfrtp_2
X_6875_ _6930_/CLK _6875_/D fanout885/X VGND VGND VPWR VPWR _6875_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5826_ _5826_/A _5826_/B _5826_/C _5826_/D VGND VGND VPWR VPWR _5826_/X sky130_fd_sc_hd__or4_1
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5757_ _6887_/Q _5702_/X _5756_/X wire671/X VGND VGND VPWR VPWR _5757_/X sky130_fd_sc_hd__a22o_2
Xmax_length607 _6037_/X VGND VGND VPWR VPWR _6139_/B1 sky130_fd_sc_hd__buf_6
X_4708_ _4708_/A _4708_/B _4708_/C _4708_/D VGND VGND VPWR VPWR _4708_/X sky130_fd_sc_hd__or4_2
Xmax_length629 wire630/X VGND VGND VPWR VPWR _6212_/B1 sky130_fd_sc_hd__buf_6
X_5688_ _7165_/Q _5704_/B _5707_/C VGND VGND VPWR VPWR _5688_/X sky130_fd_sc_hd__and3_4
XFILLER_162_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4639_ _4871_/A _4965_/A _4574_/Y _4637_/X _4638_/X VGND VGND VPWR VPWR _4639_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_190_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold640 _6984_/Q VGND VGND VPWR VPWR hold640/X sky130_fd_sc_hd__bufbuf_16
Xhold651 _6762_/Q VGND VGND VPWR VPWR hold651/X sky130_fd_sc_hd__bufbuf_16
Xhold662 _6751_/Q VGND VGND VPWR VPWR hold662/X sky130_fd_sc_hd__bufbuf_16
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6309_ _7199_/Q _6308_/X _6309_/S VGND VGND VPWR VPWR _7199_/D sky130_fd_sc_hd__mux2_1
Xhold673 _7084_/Q VGND VGND VPWR VPWR hold673/X sky130_fd_sc_hd__bufbuf_16
Xhold684 _6766_/Q VGND VGND VPWR VPWR hold684/X sky130_fd_sc_hd__bufbuf_16
Xhold695 _6786_/Q VGND VGND VPWR VPWR hold695/X sky130_fd_sc_hd__bufbuf_16
XFILLER_77_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4990_ _4990_/A _4997_/B VGND VGND VPWR VPWR _5114_/C sky130_fd_sc_hd__nor2_1
X_3941_ _6682_/Q _6797_/Q _6455_/B VGND VGND VPWR VPWR _3942_/B sky130_fd_sc_hd__mux2_1
X_3872_ hold5/A _6462_/Q _3874_/S VGND VGND VPWR VPWR _6462_/D sky130_fd_sc_hd__mux2_1
XFILLER_149_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6660_ _6752_/CLK _6660_/D fanout857/X VGND VGND VPWR VPWR _6660_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_32_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6591_ _6591_/CLK _6591_/D fanout873/X VGND VGND VPWR VPWR _6591_/Q sky130_fd_sc_hd__dfstp_4
X_5611_ _5611_/A _6680_/Q VGND VGND VPWR VPWR _5612_/B sky130_fd_sc_hd__nor2_1
XFILLER_176_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5542_ _5578_/A0 _7102_/Q _5548_/S VGND VGND VPWR VPWR _7102_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5473_ hold156/X hold321/X _5476_/S VGND VGND VPWR VPWR _5473_/X sky130_fd_sc_hd__mux2_1
X_7212_ _7218_/CLK _7212_/D wire915/X VGND VGND VPWR VPWR hold34/A sky130_fd_sc_hd__dfrtp_2
X_4424_ _4711_/A _4422_/B _4958_/A VGND VGND VPWR VPWR _4424_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_172_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4355_ _4529_/B _4486_/B _4722_/A VGND VGND VPWR VPWR _4372_/B sky130_fd_sc_hd__a21bo_2
X_7143_ _7143_/CLK _7143_/D fanout880/X VGND VGND VPWR VPWR _7143_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_132_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3306_ _3668_/A _3369_/A VGND VGND VPWR VPWR _3306_/Y sky130_fd_sc_hd__nor2_4
X_7074_ _7082_/CLK _7074_/D fanout870/X VGND VGND VPWR VPWR _7074_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_58_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4286_ _4286_/A _6406_/B VGND VGND VPWR VPWR _4291_/S sky130_fd_sc_hd__nand2_4
X_6025_ _6025_/A _6025_/B _6025_/C _6025_/D VGND VGND VPWR VPWR _6027_/D sky130_fd_sc_hd__or4_4
X_3237_ _3237_/A VGND VGND VPWR VPWR _3237_/Y sky130_fd_sc_hd__inv_2
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6927_ _6951_/CLK _6927_/D _6421_/A VGND VGND VPWR VPWR _6927_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_167_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6858_ _7042_/CLK _6858_/D fanout865/X VGND VGND VPWR VPWR _6858_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire806 _3965_/X VGND VGND VPWR VPWR wire806/X sky130_fd_sc_hd__buf_6
X_5809_ _7180_/Q _6110_/S _5808_/X VGND VGND VPWR VPWR _7180_/D sky130_fd_sc_hd__o21a_1
XFILLER_155_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire817 _6703_/Q VGND VGND VPWR VPWR wire817/X sky130_fd_sc_hd__buf_6
Xwire839 wire839/A VGND VGND VPWR VPWR _3961_/B sky130_fd_sc_hd__buf_6
Xmax_length415 _3978_/A VGND VGND VPWR VPWR _3544_/A2 sky130_fd_sc_hd__buf_6
X_6789_ _7225_/CLK _6789_/D fanout851/X VGND VGND VPWR VPWR _6789_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_136_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length426 _3324_/Y VGND VGND VPWR VPWR _3582_/A2 sky130_fd_sc_hd__buf_6
XFILLER_6_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold481 _5564_/X VGND VGND VPWR VPWR _7122_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_145_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold470 _7132_/Q VGND VGND VPWR VPWR hold470/X sky130_fd_sc_hd__bufbuf_16
Xhold492 _6947_/Q VGND VGND VPWR VPWR hold492/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_310 _6498_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_343 hold851/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_332 _7190_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_321 _5547_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_354 hold557/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4140_ hold83/X _6612_/Q _4141_/S VGND VGND VPWR VPWR hold84/A sky130_fd_sc_hd__mux2_1
XFILLER_96_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4071_ hold83/X _6553_/Q _4072_/S VGND VGND VPWR VPWR _4071_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4973_ _5174_/D _5071_/D _4973_/C _4973_/D VGND VGND VPWR VPWR _4974_/D sky130_fd_sc_hd__or4_4
X_6712_ _6712_/CLK _6712_/D fanout873/X VGND VGND VPWR VPWR _6712_/Q sky130_fd_sc_hd__dfrtp_2
X_3924_ _6457_/Q _6459_/Q _3924_/C VGND VGND VPWR VPWR _3924_/X sky130_fd_sc_hd__or3_1
XFILLER_189_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6643_ _6787_/CLK _6643_/D fanout856/X VGND VGND VPWR VPWR _6643_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_177_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3855_ _3857_/D _6487_/Q _6664_/Q VGND VGND VPWR VPWR _3856_/S sky130_fd_sc_hd__or3b_1
XFILLER_164_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6574_ _7210_/CLK _6574_/D VGND VGND VPWR VPWR _6574_/Q sky130_fd_sc_hd__dfxtp_2
X_3786_ _6811_/Q _5207_/A _5191_/A _6798_/Q _3744_/X VGND VGND VPWR VPWR _3792_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_145_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5525_ wire786/X hold257/X _5530_/S VGND VGND VPWR VPWR _5525_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5456_ wire753/X hold818/X _5458_/S VGND VGND VPWR VPWR _7026_/D sky130_fd_sc_hd__mux2_1
X_4407_ _4408_/A _4408_/B VGND VGND VPWR VPWR _4499_/C sky130_fd_sc_hd__and2_2
XFILLER_132_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5387_ _5387_/A _5594_/B VGND VGND VPWR VPWR _5387_/Y sky130_fd_sc_hd__nand2_8
XFILLER_99_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4338_ _4564_/A _4566_/A VGND VGND VPWR VPWR _4501_/A sky130_fd_sc_hd__or2_4
XFILLER_115_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7126_ _7135_/CLK _7126_/D fanout864/X VGND VGND VPWR VPWR _7126_/Q sky130_fd_sc_hd__dfstp_1
X_7057_ _7111_/CLK _7057_/D _6421_/A VGND VGND VPWR VPWR _7057_/Q sky130_fd_sc_hd__dfrtp_2
X_4269_ hold799/X _5487_/A0 _4273_/S VGND VGND VPWR VPWR _6723_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6008_ _6037_/A _6037_/B _6018_/A VGND VGND VPWR VPWR _6020_/C sky130_fd_sc_hd__and3_4
XFILLER_46_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire625 _6022_/B VGND VGND VPWR VPWR wire625/X sky130_fd_sc_hd__buf_8
Xwire603 _5987_/Y VGND VGND VPWR VPWR wire603/X sky130_fd_sc_hd__buf_8
XFILLER_10_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire647 _5996_/X VGND VGND VPWR VPWR wire647/X sky130_fd_sc_hd__buf_8
Xwire636 _6022_/A VGND VGND VPWR VPWR wire636/X sky130_fd_sc_hd__buf_8
XFILLER_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_140 mgmt_gpio_in[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_151 _7174_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_173 _6392_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_162 wb_dat_i[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_184 wire353/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_195 wire459/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3640_ input5/X _3320_/Y _3995_/A _6498_/Q _3639_/X VGND VGND VPWR VPWR _3645_/B
+ sky130_fd_sc_hd__a221o_1
X_3571_ wire908/X _3571_/A2 _5576_/A _7136_/Q _3570_/X VGND VGND VPWR VPWR _3578_/A
+ sky130_fd_sc_hd__a221o_1
X_5310_ wire773/A hold373/X _5314_/S VGND VGND VPWR VPWR _5310_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6290_ _6730_/Q wire603/X _6340_/B1 _6596_/Q VGND VGND VPWR VPWR _6290_/X sky130_fd_sc_hd__a22o_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5241_ hold465/X hold530/X _5241_/S VGND VGND VPWR VPWR _6836_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5172_ _5172_/A _5172_/B VGND VGND VPWR VPWR _5172_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4123_ hold406/X _4303_/A0 _4123_/S VGND VGND VPWR VPWR _6598_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput2 debug_oeb VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_4
X_4054_ _6539_/Q _6411_/A0 _4054_/S VGND VGND VPWR VPWR _6539_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_opt_1_0_csclk _6987_/CLK VGND VGND VPWR VPWR clkbuf_opt_1_0_csclk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_83_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4956_ _4956_/A _4956_/B _4956_/C VGND VGND VPWR VPWR _4976_/C sky130_fd_sc_hd__and3_4
XFILLER_51_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4887_ _4980_/A _4887_/B VGND VGND VPWR VPWR _4978_/B sky130_fd_sc_hd__or2_1
XFILLER_20_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3907_ _3920_/B _5612_/A _7159_/Q _7160_/Q VGND VGND VPWR VPWR _3921_/B sky130_fd_sc_hd__and4b_2
XFILLER_137_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6626_ _6626_/CLK _6626_/D fanout873/X VGND VGND VPWR VPWR _6626_/Q sky130_fd_sc_hd__dfstp_2
X_3838_ _6477_/Q _3837_/Y _3836_/X VGND VGND VPWR VPWR _6478_/D sky130_fd_sc_hd__a21o_1
XFILLER_165_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6557_ _7208_/CLK _6557_/D VGND VGND VPWR VPWR _6557_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_20_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3769_ _6545_/Q _4061_/A _3764_/X _3768_/X _3476_/Y VGND VGND VPWR VPWR _3794_/C
+ sky130_fd_sc_hd__a2111o_1
X_5508_ wire770/X hold496/X _5512_/S VGND VGND VPWR VPWR _7072_/D sky130_fd_sc_hd__mux2_1
XFILLER_193_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6488_ _6771_/CLK _6488_/D fanout855/X VGND VGND VPWR VPWR _6488_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_161_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5439_ _5547_/A0 hold819/X _5440_/S VGND VGND VPWR VPWR _7011_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7109_ _7151_/CLK _7109_/D fanout889/X VGND VGND VPWR VPWR _7109_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_101_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_718 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire411 _3346_/Y VGND VGND VPWR VPWR _5585_/A sky130_fd_sc_hd__buf_8
XFILLER_7_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire444 _3933_/X VGND VGND VPWR VPWR wire444/X sky130_fd_sc_hd__buf_6
Xwire466 _5234_/B VGND VGND VPWR VPWR _3520_/B sky130_fd_sc_hd__buf_8
Xwire455 _3369_/A VGND VGND VPWR VPWR _3540_/A sky130_fd_sc_hd__buf_8
Xwire499 _7060_/Q VGND VGND VPWR VPWR wire499/X sky130_fd_sc_hd__buf_6
Xwire477 _7112_/Q VGND VGND VPWR VPWR wire477/X sky130_fd_sc_hd__buf_4
XFILLER_124_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire488 _7092_/Q VGND VGND VPWR VPWR wire488/X sky130_fd_sc_hd__buf_4
XFILLER_124_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4810_ _4745_/B _4660_/X _4809_/X VGND VGND VPWR VPWR _4810_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5790_ _6969_/Q wire680/X wire665/X _6953_/Q VGND VGND VPWR VPWR _5790_/X sky130_fd_sc_hd__a22o_2
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4741_ _4956_/C _4748_/B VGND VGND VPWR VPWR _4881_/B sky130_fd_sc_hd__nand2_4
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4672_ _4672_/A _4672_/B _4758_/B VGND VGND VPWR VPWR _5024_/A sky130_fd_sc_hd__and3_2
XFILLER_174_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3623_ _6621_/Q _4148_/A _4268_/A _6725_/Q _3619_/X VGND VGND VPWR VPWR _3623_/X
+ sky130_fd_sc_hd__a221o_1
X_6411_ _6411_/A0 hold616/X _6411_/S VGND VGND VPWR VPWR _7225_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3554_ _6944_/Q wire401/X _5369_/A _6952_/Q VGND VGND VPWR VPWR _3554_/X sky130_fd_sc_hd__a22o_1
X_6342_ _6628_/Q _6028_/X _6342_/B1 _6727_/Q _6341_/X VGND VGND VPWR VPWR _6343_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_170_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6273_ _6615_/Q wire636/X wire634/X _6600_/Q VGND VGND VPWR VPWR _6273_/X sky130_fd_sc_hd__a22o_1
X_3485_ _5234_/A _5252_/B VGND VGND VPWR VPWR _4043_/A sky130_fd_sc_hd__nor2_8
XFILLER_103_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5224_ _6407_/A0 hold804/X _5224_/S VGND VGND VPWR VPWR _5224_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5155_ _5155_/A _5155_/B _5178_/C VGND VGND VPWR VPWR _5155_/X sky130_fd_sc_hd__or3_4
XFILLER_96_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5086_ _5086_/A _5086_/B VGND VGND VPWR VPWR _5121_/D sky130_fd_sc_hd__or2_1
X_4106_ _6583_/Q _3665_/X _4111_/S VGND VGND VPWR VPWR _6583_/D sky130_fd_sc_hd__mux2_1
X_4037_ _5248_/A0 hold844/X hold73/X VGND VGND VPWR VPWR hold74/A sky130_fd_sc_hd__mux2_1
XFILLER_84_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5988_ _7170_/Q _7171_/Q VGND VGND VPWR VPWR _6018_/A sky130_fd_sc_hd__nor2_8
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4939_ _4622_/B _4772_/A _4849_/A _4938_/Y VGND VGND VPWR VPWR _4940_/D sky130_fd_sc_hd__a211o_1
XFILLER_52_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_40 _3451_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6609_ _6747_/CLK _6609_/D fanout874/X VGND VGND VPWR VPWR _6609_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_84 _5118_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_51 _3546_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 _3830_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_62 _3687_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_95 _5826_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput191 _3216_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[24] sky130_fd_sc_hd__buf_8
Xoutput180 _3226_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[14] sky130_fd_sc_hd__buf_8
XFILLER_153_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_44_csclk _6987_/CLK VGND VGND VPWR VPWR _6986_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_140_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3270_ hold184/X _3875_/B _3845_/A VGND VGND VPWR VPWR _3270_/X sky130_fd_sc_hd__mux2_2
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_59_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7139_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_112_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6960_ _7154_/CLK _6960_/D fanout885/X VGND VGND VPWR VPWR _6960_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_66_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5911_ _6590_/Q _5977_/A2 wire667/X _6536_/Q _5897_/X VGND VGND VPWR VPWR _5911_/X
+ sky130_fd_sc_hd__a221o_1
X_6891_ _7154_/CLK _6891_/D fanout884/X VGND VGND VPWR VPWR _6891_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_179_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5842_ _6987_/Q _5864_/B VGND VGND VPWR VPWR _5842_/X sky130_fd_sc_hd__or2_1
XFILLER_62_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5773_ _3209_/A _5675_/X _5684_/X _3223_/A VGND VGND VPWR VPWR _5773_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4724_ _4724_/A _4724_/B _4812_/C VGND VGND VPWR VPWR _4725_/A sky130_fd_sc_hd__nor3_4
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4655_ _4655_/A _5050_/A _4696_/B VGND VGND VPWR VPWR _4657_/B sky130_fd_sc_hd__and3_4
XFILLER_174_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4586_ _4868_/A _4586_/B VGND VGND VPWR VPWR _4881_/A sky130_fd_sc_hd__nand2_2
Xinput60 mgmt_gpio_in[31] VGND VGND VPWR VPWR wire900/A sky130_fd_sc_hd__buf_6
XFILLER_116_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput71 mgmt_gpio_in[8] VGND VGND VPWR VPWR input71/X sky130_fd_sc_hd__clkbuf_4
Xhold811 _7067_/Q VGND VGND VPWR VPWR hold811/X sky130_fd_sc_hd__bufbuf_16
Xhold800 _6825_/Q VGND VGND VPWR VPWR hold800/X sky130_fd_sc_hd__bufbuf_16
Xinput82 spi_sdoenb VGND VGND VPWR VPWR input82/X sky130_fd_sc_hd__clkbuf_4
X_3606_ _3606_/A _3606_/B _3606_/C _3606_/D VGND VGND VPWR VPWR _3606_/X sky130_fd_sc_hd__or4_4
XFILLER_190_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold844 _6524_/Q VGND VGND VPWR VPWR hold844/X sky130_fd_sc_hd__bufbuf_16
X_3537_ _6929_/Q _5342_/A _5396_/A _6977_/Q VGND VGND VPWR VPWR _3537_/X sky130_fd_sc_hd__a22o_1
XFILLER_116_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6325_ _6617_/Q wire636/X wire634/X _6602_/Q VGND VGND VPWR VPWR _6325_/X sky130_fd_sc_hd__a22o_1
Xhold822 _7098_/Q VGND VGND VPWR VPWR hold822/X sky130_fd_sc_hd__bufbuf_16
Xhold833 _7018_/Q VGND VGND VPWR VPWR hold833/X sky130_fd_sc_hd__bufbuf_16
Xinput93 trap VGND VGND VPWR VPWR wire838/A sky130_fd_sc_hd__buf_6
XFILLER_143_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6256_ _7221_/Q _6009_/X _6253_/X _6255_/X VGND VGND VPWR VPWR _6257_/D sky130_fd_sc_hd__a211o_1
X_3468_ _3505_/A _3733_/B VGND VGND VPWR VPWR _4184_/A sky130_fd_sc_hd__nor2_8
XFILLER_97_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5207_ _5207_/A _6406_/B VGND VGND VPWR VPWR _5215_/S sky130_fd_sc_hd__and2_4
X_3399_ _7099_/Q _5531_/A _5513_/A _7083_/Q _3391_/X VGND VGND VPWR VPWR _3399_/X
+ sky130_fd_sc_hd__a221o_2
X_6187_ _7139_/Q wire642/X _6212_/B1 _7099_/Q VGND VGND VPWR VPWR _6187_/X sky130_fd_sc_hd__a22o_1
X_5138_ _4868_/A _4634_/B _4581_/B VGND VGND VPWR VPWR _5138_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_123_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5069_ _5069_/A _5069_/B _5069_/C _5069_/D VGND VGND VPWR VPWR _5076_/B sky130_fd_sc_hd__or4_1
XFILLER_38_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold107 _5499_/X VGND VGND VPWR VPWR _7064_/D sky130_fd_sc_hd__bufbuf_16
X_4440_ _4654_/A _4440_/B VGND VGND VPWR VPWR _4958_/B sky130_fd_sc_hd__xor2_4
XFILLER_172_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold129 _3327_/Y VGND VGND VPWR VPWR hold129/X sky130_fd_sc_hd__bufbuf_16
Xhold118 hold237/X VGND VGND VPWR VPWR _3260_/A sky130_fd_sc_hd__bufbuf_16
XFILLER_171_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4371_ _4533_/A _4372_/B _4372_/C _4484_/C VGND VGND VPWR VPWR _4507_/A sky130_fd_sc_hd__and4b_4
XFILLER_125_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6110_ _7191_/Q _6109_/X _6110_/S VGND VGND VPWR VPWR _7191_/D sky130_fd_sc_hd__mux2_1
XFILLER_3_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3322_ _3552_/B _5225_/B VGND VGND VPWR VPWR _3322_/Y sky130_fd_sc_hd__nor2_8
X_7090_ _7091_/CLK _7090_/D fanout868/X VGND VGND VPWR VPWR _7090_/Q sky130_fd_sc_hd__dfrtp_2
X_6041_ _7109_/Q wire650/X _6039_/X _6040_/X VGND VGND VPWR VPWR _6059_/A sky130_fd_sc_hd__a211o_2
XFILLER_98_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ hold331/X _3249_/B _3845_/A VGND VGND VPWR VPWR _3253_/X sky130_fd_sc_hd__mux2_2
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6943_ _7140_/CLK _6943_/D fanout862/X VGND VGND VPWR VPWR _6943_/Q sky130_fd_sc_hd__dfrtp_2
X_6874_ _7122_/CLK _6874_/D fanout887/X VGND VGND VPWR VPWR _6874_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_179_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5825_ wire527/X _5676_/X _5702_/X _6890_/Q _5824_/X VGND VGND VPWR VPWR _5826_/D
+ sky130_fd_sc_hd__a221o_4
XFILLER_50_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5756_ _6983_/Q _5963_/B VGND VGND VPWR VPWR _5756_/X sky130_fd_sc_hd__or2_1
Xmax_length608 _6211_/B VGND VGND VPWR VPWR _6311_/B sky130_fd_sc_hd__buf_6
X_4707_ _4707_/A _4707_/B _4773_/A _4930_/C VGND VGND VPWR VPWR _5031_/B sky130_fd_sc_hd__or4bb_4
X_5687_ _7165_/Q _5702_/B _5706_/B VGND VGND VPWR VPWR _5687_/X sky130_fd_sc_hd__and3_4
Xmax_length619 _6029_/X VGND VGND VPWR VPWR wire618/A sky130_fd_sc_hd__buf_6
XFILLER_163_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4638_ _4819_/B _4819_/D _4947_/B VGND VGND VPWR VPWR _4638_/X sky130_fd_sc_hd__or3_4
Xhold630 _6968_/Q VGND VGND VPWR VPWR hold630/X sky130_fd_sc_hd__bufbuf_16
XFILLER_118_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4569_ _4749_/C _4990_/A VGND VGND VPWR VPWR _5071_/A sky130_fd_sc_hd__nor2_2
XFILLER_104_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold641 _6594_/Q VGND VGND VPWR VPWR hold641/X sky130_fd_sc_hd__bufbuf_16
XFILLER_78_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold663 _6853_/Q VGND VGND VPWR VPWR hold663/X sky130_fd_sc_hd__bufbuf_16
Xhold652 _6643_/Q VGND VGND VPWR VPWR hold652/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold685 _6547_/Q VGND VGND VPWR VPWR hold685/X sky130_fd_sc_hd__bufbuf_16
Xhold674 _6709_/Q VGND VGND VPWR VPWR hold674/X sky130_fd_sc_hd__bufbuf_16
XFILLER_89_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6308_ _7198_/Q _6307_/X _6308_/S VGND VGND VPWR VPWR _6308_/X sky130_fd_sc_hd__mux2_1
Xhold696 _5187_/X VGND VGND VPWR VPWR _6786_/D sky130_fd_sc_hd__bufbuf_16
X_6239_ _6659_/Q wire647/X wire640/X _6713_/Q VGND VGND VPWR VPWR _6239_/X sky130_fd_sc_hd__a22o_1
XFILLER_77_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3940_ _6687_/Q input77/X _3969_/B VGND VGND VPWR VPWR _3940_/X sky130_fd_sc_hd__mux2_8
XFILLER_189_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3871_ _6462_/Q _6463_/Q _3874_/S VGND VGND VPWR VPWR _6463_/D sky130_fd_sc_hd__mux2_1
XFILLER_177_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6590_ _6650_/CLK _6590_/D fanout858/X VGND VGND VPWR VPWR _6590_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5610_ _7157_/Q _7158_/Q VGND VGND VPWR VPWR _5610_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5541_ wire802/X hold517/X _5548_/S VGND VGND VPWR VPWR _7101_/D sky130_fd_sc_hd__mux2_1
X_7211_ _7218_/CLK _7211_/D wire915/X VGND VGND VPWR VPWR _7211_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_145_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5472_ wire769/X hold603/X _5476_/S VGND VGND VPWR VPWR _5472_/X sky130_fd_sc_hd__mux2_1
X_4423_ _4696_/A _4711_/A _4654_/A VGND VGND VPWR VPWR _4423_/X sky130_fd_sc_hd__a21o_1
X_4354_ _4696_/A _4413_/C _4436_/B VGND VGND VPWR VPWR _4486_/B sky130_fd_sc_hd__and3_4
X_7142_ _7145_/CLK _7142_/D fanout883/X VGND VGND VPWR VPWR _7142_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_125_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3305_ hold63/X _3540_/A VGND VGND VPWR VPWR _3305_/Y sky130_fd_sc_hd__nor2_8
XFILLER_59_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7073_ _7129_/CLK _7073_/D fanout863/X VGND VGND VPWR VPWR _7073_/Q sky130_fd_sc_hd__dfrtp_2
X_4285_ _5599_/A0 hold307/X _4285_/S VGND VGND VPWR VPWR _6737_/D sky130_fd_sc_hd__mux2_1
X_6024_ _6024_/A _6024_/B _6024_/C _6024_/D VGND VGND VPWR VPWR _6027_/C sky130_fd_sc_hd__or4_4
XFILLER_101_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3236_ _3236_/A VGND VGND VPWR VPWR _3236_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6926_ _6951_/CLK _6926_/D _6421_/A VGND VGND VPWR VPWR _6926_/Q sky130_fd_sc_hd__dfstp_2
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6857_ _7140_/CLK _6857_/D fanout862/X VGND VGND VPWR VPWR _6857_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5808_ _5611_/A _7179_/Q wire381/A _5807_/X VGND VGND VPWR VPWR _5808_/X sky130_fd_sc_hd__a211o_2
Xwire807 _3964_/X VGND VGND VPWR VPWR wire807/X sky130_fd_sc_hd__buf_6
XFILLER_13_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6788_ _7223_/CLK _6788_/D fanout850/X VGND VGND VPWR VPWR _6788_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length405 _3356_/Y VGND VGND VPWR VPWR _3683_/B1 sky130_fd_sc_hd__buf_6
Xmax_length416 _3335_/Y VGND VGND VPWR VPWR _3978_/A sky130_fd_sc_hd__buf_6
X_5739_ _7006_/Q wire700/X wire679/X _7070_/Q VGND VGND VPWR VPWR _5739_/X sky130_fd_sc_hd__a22o_1
XFILLER_163_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length449 hold88/A VGND VGND VPWR VPWR _3583_/A2 sky130_fd_sc_hd__buf_6
XFILLER_136_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold460 _6842_/Q VGND VGND VPWR VPWR hold460/X sky130_fd_sc_hd__bufbuf_16
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold471 _5575_/X VGND VGND VPWR VPWR _7132_/D sky130_fd_sc_hd__bufbuf_16
Xhold493 _5367_/X VGND VGND VPWR VPWR _6947_/D sky130_fd_sc_hd__bufbuf_16
Xhold482 _6857_/Q VGND VGND VPWR VPWR hold482/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_300 _5685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_333 hold212/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_322 wire753/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_311 _6500_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_344 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_355 hold566/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4070_ _5498_/A0 hold723/X _4072_/S VGND VGND VPWR VPWR _6552_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4972_ _4536_/X _4959_/A _5129_/B _4971_/X _4903_/A VGND VGND VPWR VPWR _4973_/D
+ sky130_fd_sc_hd__a2111o_4
XFILLER_24_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6711_ _6712_/CLK _6711_/D fanout872/X VGND VGND VPWR VPWR _6711_/Q sky130_fd_sc_hd__dfrtp_2
X_3923_ _6459_/Q _6664_/Q _3843_/B _6668_/Q VGND VGND VPWR VPWR _6668_/D sky130_fd_sc_hd__a31o_1
XFILLER_149_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3854_ _6486_/Q _6485_/Q VGND VGND VPWR VPWR _3857_/D sky130_fd_sc_hd__nand2b_1
X_6642_ _6642_/CLK _6642_/D fanout856/X VGND VGND VPWR VPWR _6642_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_32_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6573_ _7208_/CLK _6573_/D VGND VGND VPWR VPWR _6573_/Q sky130_fd_sc_hd__dfxtp_4
X_3785_ _3785_/A _3785_/B _3785_/C _3785_/D VGND VGND VPWR VPWR _3793_/C sky130_fd_sc_hd__or4_1
XFILLER_145_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR clkbuf_1_1_1_mgmt_gpio_in[4]/A
+ sky130_fd_sc_hd__clkbuf_8
X_5524_ _5578_/A0 _7086_/Q _5530_/S VGND VGND VPWR VPWR _7086_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5455_ _5572_/A0 hold520/X _5458_/S VGND VGND VPWR VPWR _7025_/D sky130_fd_sc_hd__mux2_1
X_4406_ _4707_/B _4478_/C _4410_/C VGND VGND VPWR VPWR _4513_/B sky130_fd_sc_hd__or3_4
X_7125_ _7128_/CLK _7125_/D _6420_/A VGND VGND VPWR VPWR _7125_/Q sky130_fd_sc_hd__dfstp_4
X_5386_ _5602_/A0 hold288/X _5386_/S VGND VGND VPWR VPWR _6964_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4337_ _4818_/A _4469_/A _4395_/D VGND VGND VPWR VPWR _4413_/C sky130_fd_sc_hd__and3_4
X_7056_ _7096_/CLK _7056_/D fanout883/X VGND VGND VPWR VPWR _7056_/Q sky130_fd_sc_hd__dfrtp_2
X_4268_ _4268_/A _5236_/B VGND VGND VPWR VPWR _4273_/S sky130_fd_sc_hd__and2_4
XFILLER_115_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3219_ _3219_/A VGND VGND VPWR VPWR _3219_/Y sky130_fd_sc_hd__inv_2
X_6007_ _6032_/A _6018_/A _6032_/C VGND VGND VPWR VPWR _6025_/C sky130_fd_sc_hd__and3_4
XFILLER_75_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4199_ _5579_/A0 _6661_/Q _4201_/S VGND VGND VPWR VPWR _6661_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6909_ _7151_/CLK _6909_/D fanout880/X VGND VGND VPWR VPWR _6909_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_70_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire615 wire616/X VGND VGND VPWR VPWR wire615/X sky130_fd_sc_hd__buf_8
Xwire604 _5987_/Y VGND VGND VPWR VPWR wire604/X sky130_fd_sc_hd__buf_8
XFILLER_11_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire637 _6022_/A VGND VGND VPWR VPWR wire637/X sky130_fd_sc_hd__buf_8
Xwire648 _5996_/X VGND VGND VPWR VPWR wire648/X sky130_fd_sc_hd__buf_8
Xwire659 _5704_/X VGND VGND VPWR VPWR wire659/X sky130_fd_sc_hd__buf_8
XFILLER_6_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold290 _6900_/Q VGND VGND VPWR VPWR hold290/X sky130_fd_sc_hd__bufbuf_16
XFILLER_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout781 _5336_/A1 VGND VGND VPWR VPWR _5498_/A0 sky130_fd_sc_hd__buf_8
XFILLER_65_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout792 wire796/X VGND VGND VPWR VPWR _5578_/A0 sky130_fd_sc_hd__buf_8
XFILLER_92_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_141 mgmt_gpio_in[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_152 spi_csb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_130 mask_rev_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_174 _6395_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_163 wb_dat_i[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_185 _3331_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_196 wire470/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3570_ _6736_/Q _4280_/A _4268_/A _6726_/Q VGND VGND VPWR VPWR _3570_/X sky130_fd_sc_hd__a22o_4
XFILLER_154_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5240_ hold38/X _6835_/Q _5241_/S VGND VGND VPWR VPWR _5240_/X sky130_fd_sc_hd__mux2_1
Xmax_length791 wire790/A VGND VGND VPWR VPWR _5247_/A0 sky130_fd_sc_hd__buf_6
XFILLER_114_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5171_ _5171_/A _5171_/B _5171_/C _5170_/X VGND VGND VPWR VPWR _5171_/X sky130_fd_sc_hd__or4b_4
XFILLER_69_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4122_ hold459/X _5249_/A0 _4123_/S VGND VGND VPWR VPWR _6597_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4053_ _6538_/Q _6410_/A0 _4054_/S VGND VGND VPWR VPWR _6538_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput3 debug_out VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_4
XFILLER_91_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4955_ _4443_/X _4537_/X _4956_/C _5136_/B _5075_/C VGND VGND VPWR VPWR _5128_/C
+ sky130_fd_sc_hd__a311o_1
XFILLER_101_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3906_ _7157_/Q _7158_/Q VGND VGND VPWR VPWR _5612_/A sky130_fd_sc_hd__nor2_1
X_4886_ _5005_/C _4886_/B VGND VGND VPWR VPWR _4886_/Y sky130_fd_sc_hd__nor2_1
XFILLER_137_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6625_ _6632_/CLK _6625_/D fanout872/X VGND VGND VPWR VPWR _6625_/Q sky130_fd_sc_hd__dfrtp_2
X_3837_ hold59/A _3825_/B _3840_/S VGND VGND VPWR VPWR _3837_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_20_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6556_ _7208_/CLK _6556_/D VGND VGND VPWR VPWR _6556_/Q sky130_fd_sc_hd__dfxtp_4
X_3768_ _6748_/Q _4298_/A _5242_/A _6837_/Q _3767_/X VGND VGND VPWR VPWR _3768_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_106_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5507_ wire786/X hold360/X _5512_/S VGND VGND VPWR VPWR _7071_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6487_ _6668_/CLK _6487_/D _6442_/X VGND VGND VPWR VPWR _6487_/Q sky130_fd_sc_hd__dfrtp_2
X_3699_ _3699_/A _3699_/B _3699_/C _3699_/D VGND VGND VPWR VPWR _3727_/C sky130_fd_sc_hd__or4_2
XFILLER_160_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput340 _6583_/Q VGND VGND VPWR VPWR wb_dat_o[2] sky130_fd_sc_hd__buf_8
X_5438_ wire753/X hold823/X _5440_/S VGND VGND VPWR VPWR _7010_/D sky130_fd_sc_hd__mux2_1
X_5369_ _5369_/A _5594_/B VGND VGND VPWR VPWR _5377_/S sky130_fd_sc_hd__nand2_8
XFILLER_120_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7108_ _7140_/CLK _7108_/D fanout865/X VGND VGND VPWR VPWR _7108_/Q sky130_fd_sc_hd__dfrtp_2
X_7039_ _7135_/CLK _7039_/D fanout864/X VGND VGND VPWR VPWR _7039_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_74_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire401 _5360_/A VGND VGND VPWR VPWR wire401/X sky130_fd_sc_hd__buf_8
XFILLER_183_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire467 _5252_/A VGND VGND VPWR VPWR _4241_/A sky130_fd_sc_hd__buf_8
Xwire445 _3419_/X VGND VGND VPWR VPWR wire445/X sky130_fd_sc_hd__buf_8
Xwire456 _3353_/B VGND VGND VPWR VPWR _3543_/A sky130_fd_sc_hd__buf_8
XFILLER_164_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire478 _7110_/Q VGND VGND VPWR VPWR wire478/X sky130_fd_sc_hd__buf_6
XFILLER_109_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire489 _7091_/Q VGND VGND VPWR VPWR wire489/X sky130_fd_sc_hd__buf_6
XFILLER_3_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4740_ _4740_/A _4740_/B _4832_/C VGND VGND VPWR VPWR _4740_/X sky130_fd_sc_hd__or3_4
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4671_ _4671_/A _4745_/B VGND VGND VPWR VPWR _5099_/A sky130_fd_sc_hd__nor2_2
XFILLER_186_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3622_ _6591_/Q _4112_/A _4250_/A _6710_/Q _3614_/X VGND VGND VPWR VPWR _3622_/X
+ sky130_fd_sc_hd__a221o_1
X_6410_ _6410_/A0 hold664/X _6411_/S VGND VGND VPWR VPWR _7224_/D sky130_fd_sc_hd__mux2_1
XFILLER_162_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6341_ _7225_/Q _6009_/X wire627/X _6712_/Q VGND VGND VPWR VPWR _6341_/X sky130_fd_sc_hd__a22o_1
X_3553_ _7104_/Q _5540_/A _4316_/A _6766_/Q VGND VGND VPWR VPWR _3553_/X sky130_fd_sc_hd__a22o_1
XFILLER_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3484_ _3543_/A _3520_/B VGND VGND VPWR VPWR _4061_/A sky130_fd_sc_hd__nor2_8
XFILLER_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6272_ _6744_/Q wire597/X wire611/X _6739_/Q _6271_/X VGND VGND VPWR VPWR _6282_/B
+ sky130_fd_sc_hd__a221o_1
X_5223_ _5223_/A _6406_/B VGND VGND VPWR VPWR _5224_/S sky130_fd_sc_hd__nand2_1
X_5154_ _5154_/A _5154_/B VGND VGND VPWR VPWR _5178_/C sky130_fd_sc_hd__or2_2
XFILLER_111_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4105_ _6582_/Q _3727_/X _4111_/S VGND VGND VPWR VPWR _6582_/D sky130_fd_sc_hd__mux2_1
X_5085_ _4986_/A _4844_/B _4935_/D VGND VGND VPWR VPWR _5086_/B sky130_fd_sc_hd__o21ai_1
X_4036_ hold38/X hold845/X hold73/X VGND VGND VPWR VPWR hold39/A sky130_fd_sc_hd__mux2_1
XFILLER_112_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5987_ _6036_/A _6004_/A VGND VGND VPWR VPWR _5987_/Y sky130_fd_sc_hd__nor2_8
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4938_ _4745_/A _4697_/A _4757_/B VGND VGND VPWR VPWR _4938_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_30 _5563_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4869_ _4737_/Y _5087_/D _4949_/C VGND VGND VPWR VPWR _4870_/A sky130_fd_sc_hd__o21ai_2
XFILLER_177_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_41 _3461_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6608_ _6608_/CLK _6608_/D fanout858/X VGND VGND VPWR VPWR _6608_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_74 _3830_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_52 _3560_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_63 _3687_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_85 _4558_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_96 _5861_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6539_ _6824_/CLK _6539_/D _6435_/A VGND VGND VPWR VPWR _6539_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_137_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput192 _3215_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[25] sky130_fd_sc_hd__buf_8
Xoutput181 _3225_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[15] sky130_fd_sc_hd__buf_8
XFILLER_102_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5910_ _5910_/A _5910_/B _5910_/C _5910_/D VGND VGND VPWR VPWR _5915_/B sky130_fd_sc_hd__or4_2
X_6890_ _7154_/CLK _6890_/D fanout886/X VGND VGND VPWR VPWR _6890_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_34_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5841_ wire495/X _5669_/X _5703_/X _6875_/Q _5840_/X VGND VGND VPWR VPWR _5849_/A
+ sky130_fd_sc_hd__a221o_1
X_5772_ _6960_/Q _5673_/X _5681_/X _6920_/Q _5771_/X VGND VGND VPWR VPWR _5777_/B
+ sky130_fd_sc_hd__a221o_1
X_4723_ _4592_/B _4898_/B _4886_/B VGND VGND VPWR VPWR _4723_/X sky130_fd_sc_hd__a21o_1
XFILLER_166_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4654_ _4654_/A _4654_/B VGND VGND VPWR VPWR _4696_/B sky130_fd_sc_hd__nor2_8
XFILLER_174_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4585_ _4634_/B _4586_/B VGND VGND VPWR VPWR _5123_/C sky130_fd_sc_hd__nand2_4
Xinput50 mgmt_gpio_in[22] VGND VGND VPWR VPWR wire906/A sky130_fd_sc_hd__buf_6
Xinput61 mgmt_gpio_in[32] VGND VGND VPWR VPWR input61/X sky130_fd_sc_hd__clkbuf_4
XFILLER_135_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold801 _6624_/Q VGND VGND VPWR VPWR hold801/X sky130_fd_sc_hd__bufbuf_16
Xinput72 mgmt_gpio_in[9] VGND VGND VPWR VPWR input72/X sky130_fd_sc_hd__buf_4
Xhold812 _7223_/Q VGND VGND VPWR VPWR hold812/X sky130_fd_sc_hd__bufbuf_16
X_3605_ _3605_/A _3605_/B _3605_/C _3605_/D VGND VGND VPWR VPWR _3606_/D sky130_fd_sc_hd__or4_1
Xhold845 _6523_/Q VGND VGND VPWR VPWR hold845/X sky130_fd_sc_hd__bufbuf_16
Xinput83 spimemio_flash_clk VGND VGND VPWR VPWR wire844/A sky130_fd_sc_hd__buf_6
Xinput94 uart_enabled VGND VGND VPWR VPWR _3969_/B sky130_fd_sc_hd__clkbuf_4
X_6324_ wire565/X wire597/X wire611/X _6741_/Q _6323_/X VGND VGND VPWR VPWR _6331_/B
+ sky130_fd_sc_hd__a221o_1
Xhold823 _7010_/Q VGND VGND VPWR VPWR hold823/X sky130_fd_sc_hd__bufbuf_16
Xhold834 _6532_/Q VGND VGND VPWR VPWR hold834/X sky130_fd_sc_hd__bufbuf_16
X_3536_ _7049_/Q _5477_/A _4262_/A _6722_/Q _3535_/X VGND VGND VPWR VPWR _3546_/A
+ sky130_fd_sc_hd__a221o_4
X_6255_ _6550_/Q wire601/X _6293_/B1 _6723_/Q _6254_/X VGND VGND VPWR VPWR _6255_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_170_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5206_ wire753/A hold758/X _5206_/S VGND VGND VPWR VPWR _6810_/D sky130_fd_sc_hd__mux2_1
X_3467_ _3467_/A _3528_/B VGND VGND VPWR VPWR _4298_/A sky130_fd_sc_hd__nor2_8
X_3398_ _3398_/A _3398_/B _3398_/C _3398_/D VGND VGND VPWR VPWR _3415_/A sky130_fd_sc_hd__or4_1
X_6186_ _7043_/Q _6335_/B VGND VGND VPWR VPWR _6186_/X sky130_fd_sc_hd__and2_1
X_5137_ _5137_/A _5137_/B _5137_/C VGND VGND VPWR VPWR _5172_/B sky130_fd_sc_hd__or3_1
XFILLER_184_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5068_ _5069_/B _5068_/B _5067_/X VGND VGND VPWR VPWR _5132_/C sky130_fd_sc_hd__or3b_1
XFILLER_84_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4019_ hold478/X _5600_/A0 _4023_/S VGND VGND VPWR VPWR _4019_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold108 _6480_/Q VGND VGND VPWR VPWR hold108/X sky130_fd_sc_hd__bufbuf_16
X_4370_ _4484_/C VGND VGND VPWR VPWR _4370_/Y sky130_fd_sc_hd__inv_2
XFILLER_156_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold119 _3294_/X VGND VGND VPWR VPWR _3353_/B sky130_fd_sc_hd__bufbuf_16
XFILLER_125_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3321_ hold43/X hold95/X VGND VGND VPWR VPWR _5225_/B sky130_fd_sc_hd__or2_4
XFILLER_140_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _6893_/Q wire591/X _6179_/A2 _6861_/Q _6038_/X VGND VGND VPWR VPWR _6040_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _3260_/A VGND VGND VPWR VPWR _3314_/A sky130_fd_sc_hd__inv_2
XFILLER_112_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6942_ _7036_/CLK _6942_/D fanout869/X VGND VGND VPWR VPWR _6942_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6873_ _7128_/CLK _6873_/D _6421_/A VGND VGND VPWR VPWR _6873_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_81_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5824_ _7066_/Q _5669_/X _5698_/B _6986_/Q _5697_/X VGND VGND VPWR VPWR _5824_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5755_ _6879_/Q _5934_/B1 _5681_/X _6919_/Q _5754_/X VGND VGND VPWR VPWR _5763_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_175_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4706_ _5165_/A _4453_/Y _4695_/X _5166_/A VGND VGND VPWR VPWR _4706_/X sky130_fd_sc_hd__a31o_1
X_5686_ _6989_/Q _5684_/X wire691/X wire493/X VGND VGND VPWR VPWR _5686_/X sky130_fd_sc_hd__a22o_1
XFILLER_190_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4637_ _4636_/A _4844_/A _4591_/X _4635_/X VGND VGND VPWR VPWR _4637_/X sky130_fd_sc_hd__o211a_1
XFILLER_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold620 _7008_/Q VGND VGND VPWR VPWR hold620/X sky130_fd_sc_hd__bufbuf_16
Xhold642 _7112_/Q VGND VGND VPWR VPWR hold642/X sky130_fd_sc_hd__bufbuf_16
X_4568_ _4868_/A _4624_/B VGND VGND VPWR VPWR _4623_/A sky130_fd_sc_hd__nand2_2
XFILLER_116_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold631 _6851_/Q VGND VGND VPWR VPWR hold631/X sky130_fd_sc_hd__bufbuf_16
Xhold653 _6991_/Q VGND VGND VPWR VPWR hold653/X sky130_fd_sc_hd__bufbuf_16
X_4499_ _4553_/B _4507_/A _4499_/C VGND VGND VPWR VPWR _4586_/B sky130_fd_sc_hd__and3b_4
X_3519_ wire476/X _5558_/A _4124_/A _6603_/Q VGND VGND VPWR VPWR _3519_/X sky130_fd_sc_hd__a22o_1
XFILLER_104_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold675 _6615_/Q VGND VGND VPWR VPWR hold675/X sky130_fd_sc_hd__bufbuf_16
Xhold697 _6657_/Q VGND VGND VPWR VPWR hold697/X sky130_fd_sc_hd__bufbuf_16
Xhold686 _6655_/Q VGND VGND VPWR VPWR hold686/X sky130_fd_sc_hd__bufbuf_16
Xhold664 _7224_/Q VGND VGND VPWR VPWR hold664/X sky130_fd_sc_hd__bufbuf_16
X_6307_ _6288_/X _6294_/X _6306_/X _6357_/A2 _6532_/Q VGND VGND VPWR VPWR _6307_/X
+ sky130_fd_sc_hd__o32a_1
X_6238_ _6563_/Q wire590/X wire632/X _6589_/Q _6237_/X VGND VGND VPWR VPWR _6248_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6169_ _6986_/Q _6028_/X _6342_/B1 _6994_/Q _6168_/X VGND VGND VPWR VPWR _6170_/D
+ sky130_fd_sc_hd__a221o_2
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_43_csclk _6987_/CLK VGND VGND VPWR VPWR _6971_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_58_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7042_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_159_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3870_ _6463_/Q hold1/A _3874_/S VGND VGND VPWR VPWR _6464_/D sky130_fd_sc_hd__mux2_1
XFILLER_71_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5540_ _5540_/A _5576_/B VGND VGND VPWR VPWR _5548_/S sky130_fd_sc_hd__nand2_8
XFILLER_172_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5471_ wire780/X hold649/X _5476_/S VGND VGND VPWR VPWR _7039_/D sky130_fd_sc_hd__mux2_1
X_4422_ _4711_/A _4422_/B VGND VGND VPWR VPWR _4422_/Y sky130_fd_sc_hd__nand2_2
XFILLER_117_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7210_ _7210_/CLK _7210_/D VGND VGND VPWR VPWR _7210_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_160_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4353_ _4654_/A _4958_/A VGND VGND VPWR VPWR _4436_/B sky130_fd_sc_hd__and2_4
X_7141_ _7151_/CLK _7141_/D fanout880/X VGND VGND VPWR VPWR _7141_/Q sky130_fd_sc_hd__dfstp_1
X_7072_ _7072_/CLK _7072_/D fanout870/X VGND VGND VPWR VPWR _7072_/Q sky130_fd_sc_hd__dfrtp_2
X_3304_ _3314_/A _3304_/B VGND VGND VPWR VPWR _3304_/X sky130_fd_sc_hd__or2_4
X_4284_ _5249_/A0 hold486/X _4285_/S VGND VGND VPWR VPWR _6736_/D sky130_fd_sc_hd__mux2_1
X_3235_ _3235_/A VGND VGND VPWR VPWR _3235_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6023_ _6023_/A _6023_/B _6023_/C _6023_/D VGND VGND VPWR VPWR _6024_/D sky130_fd_sc_hd__or4_1
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6925_ _7151_/CLK _6925_/D fanout880/X VGND VGND VPWR VPWR _6925_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_82_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6856_ _7140_/CLK _6856_/D fanout862/X VGND VGND VPWR VPWR _6856_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_167_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5807_ _6857_/Q _5722_/B _5796_/X _5806_/X _6109_/S VGND VGND VPWR VPWR _5807_/X
+ sky130_fd_sc_hd__o221a_1
X_3999_ _6499_/Q _6410_/A0 _4003_/S VGND VGND VPWR VPWR _6499_/D sky130_fd_sc_hd__mux2_1
X_6787_ _6787_/CLK _6787_/D fanout850/X VGND VGND VPWR VPWR _6787_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_50_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire819 _3975_/B VGND VGND VPWR VPWR _3991_/S sky130_fd_sc_hd__buf_8
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5738_ _7094_/Q _5980_/A2 wire677/X _7078_/Q _5737_/X VGND VGND VPWR VPWR _5741_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_136_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length428 hold136/X VGND VGND VPWR VPWR wire427/A sky130_fd_sc_hd__buf_6
XFILLER_175_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5669_ _7165_/Q _5704_/B _5706_/B VGND VGND VPWR VPWR _5669_/X sky130_fd_sc_hd__and3_4
Xhold450 _5600_/X VGND VGND VPWR VPWR _7154_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_145_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold461 _5249_/X VGND VGND VPWR VPWR _6842_/D sky130_fd_sc_hd__bufbuf_16
Xhold472 _7076_/Q VGND VGND VPWR VPWR hold472/X sky130_fd_sc_hd__bufbuf_16
Xhold494 _6512_/Q VGND VGND VPWR VPWR hold494/X sky130_fd_sc_hd__bufbuf_16
Xhold483 _6510_/Q VGND VGND VPWR VPWR hold483/X sky130_fd_sc_hd__bufbuf_16
XFILLER_77_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_301 _5937_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_334 hold218/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_323 _4303_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_312 _3730_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_345 _5564_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_110_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4971_ _5130_/A _4971_/B _4970_/X VGND VGND VPWR VPWR _4971_/X sky130_fd_sc_hd__or3b_2
XFILLER_64_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6710_ _6712_/CLK _6710_/D fanout872/X VGND VGND VPWR VPWR _6710_/Q sky130_fd_sc_hd__dfstp_2
X_3922_ _6679_/Q _5606_/B VGND VGND VPWR VPWR _6678_/D sky130_fd_sc_hd__or2_1
XFILLER_149_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3853_ _3875_/B _6471_/Q _3853_/S VGND VGND VPWR VPWR _6471_/D sky130_fd_sc_hd__mux2_1
X_6641_ _6642_/CLK _6641_/D fanout856/X VGND VGND VPWR VPWR _6641_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_192_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6572_ _7210_/CLK _6572_/D VGND VGND VPWR VPWR _6572_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_9_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3784_ input11/X _3368_/Y _4286_/A _6738_/Q _3783_/X VGND VGND VPWR VPWR _3785_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5523_ _5532_/A0 wire493/X _5530_/S VGND VGND VPWR VPWR _7085_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5454_ wire769/X hold615/X _5458_/S VGND VGND VPWR VPWR _7024_/D sky130_fd_sc_hd__mux2_1
X_5385_ _5601_/A0 hold205/X _5386_/S VGND VGND VPWR VPWR _6963_/D sky130_fd_sc_hd__mux2_1
X_4405_ _4553_/A _4405_/B VGND VGND VPWR VPWR _4636_/A sky130_fd_sc_hd__or2_4
X_4336_ _4469_/A _4395_/D VGND VGND VPWR VPWR _4566_/A sky130_fd_sc_hd__nand2_8
XFILLER_160_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7124_ _7136_/CLK _7124_/D fanout871/X VGND VGND VPWR VPWR _7124_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_5_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7055_ _7128_/CLK _7055_/D _6421_/A VGND VGND VPWR VPWR _7055_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_140_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4267_ _6722_/Q _6411_/A0 _4267_/S VGND VGND VPWR VPWR _6722_/D sky130_fd_sc_hd__mux2_1
X_3218_ _3218_/A VGND VGND VPWR VPWR _3218_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6006_ _6035_/A _6018_/A _6035_/C VGND VGND VPWR VPWR _6022_/A sky130_fd_sc_hd__and3_4
XFILLER_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4198_ _5247_/A0 hold498/X _4201_/S VGND VGND VPWR VPWR _6660_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6908_ _6980_/CLK _6908_/D fanout878/X VGND VGND VPWR VPWR _6908_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6839_ _6842_/CLK _6839_/D fanout857/X VGND VGND VPWR VPWR _6839_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_183_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire616 _6031_/X VGND VGND VPWR VPWR wire616/X sky130_fd_sc_hd__buf_8
Xwire605 _5698_/Y VGND VGND VPWR VPWR _5722_/B sky130_fd_sc_hd__buf_8
XFILLER_10_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire627 _6012_/X VGND VGND VPWR VPWR wire627/X sky130_fd_sc_hd__buf_8
Xwire638 _6021_/C VGND VGND VPWR VPWR wire638/X sky130_fd_sc_hd__buf_8
Xwire649 _6027_/B VGND VGND VPWR VPWR wire649/X sky130_fd_sc_hd__buf_8
XFILLER_7_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold280 _6868_/Q VGND VGND VPWR VPWR hold280/X sky130_fd_sc_hd__bufbuf_16
XFILLER_151_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold291 _5314_/X VGND VGND VPWR VPWR _6900_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_104_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout760 wire763/A VGND VGND VPWR VPWR _4303_/A0 sky130_fd_sc_hd__buf_8
Xfanout771 wire773/A VGND VGND VPWR VPWR _5598_/A0 sky130_fd_sc_hd__buf_8
Xfanout793 hold38/A VGND VGND VPWR VPWR wire794/A sky130_fd_sc_hd__buf_8
XFILLER_172_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout782 hold7/X VGND VGND VPWR VPWR _5597_/A0 sky130_fd_sc_hd__buf_6
XFILLER_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_142 mgmt_gpio_in[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_120 _6480_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_131 mask_rev_in[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_175 _6395_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_164 wb_dat_i[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_153 spi_sck VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_186 _5581_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_197 wire475/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5170_ _4871_/A _4988_/A _4617_/A _4997_/B _4893_/A VGND VGND VPWR VPWR _5170_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4121_ hold838/X _6409_/A0 _4123_/S VGND VGND VPWR VPWR _6596_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4052_ hold832/X _6409_/A0 _4054_/S VGND VGND VPWR VPWR _6537_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput4 mask_rev_in[0] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_4
XFILLER_37_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4954_ _4636_/A _4986_/C _5005_/C _4591_/B VGND VGND VPWR VPWR _5075_/C sky130_fd_sc_hd__o22ai_4
XFILLER_91_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3905_ _6019_/A _6030_/A VGND VGND VPWR VPWR _3905_/X sky130_fd_sc_hd__or2_4
X_4885_ _4502_/A _4997_/A _4740_/X _4395_/D VGND VGND VPWR VPWR _5123_/D sky130_fd_sc_hd__o22a_1
XFILLER_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6624_ _6626_/CLK _6624_/D fanout873/X VGND VGND VPWR VPWR _6624_/Q sky130_fd_sc_hd__dfrtp_2
X_3836_ _3191_/Y _3840_/S _3825_/B hold59/A VGND VGND VPWR VPWR _3836_/X sky130_fd_sc_hd__o211a_1
XFILLER_118_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6555_ _7218_/CLK _6555_/D VGND VGND VPWR VPWR _6555_/Q sky130_fd_sc_hd__dfxtp_2
X_3767_ _6504_/Q _4004_/A _3765_/X _3766_/X VGND VGND VPWR VPWR _3767_/X sky130_fd_sc_hd__a211o_4
XFILLER_106_616 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5506_ _5578_/A0 _7070_/Q _5512_/S VGND VGND VPWR VPWR _7070_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6486_ _6668_/CLK _6486_/D _6441_/X VGND VGND VPWR VPWR _6486_/Q sky130_fd_sc_hd__dfrtp_2
X_3698_ _7094_/Q _5531_/A _4304_/A _6754_/Q _3675_/X VGND VGND VPWR VPWR _3699_/D
+ sky130_fd_sc_hd__a221o_1
Xoutput341 _7209_/Q VGND VGND VPWR VPWR wb_dat_o[30] sky130_fd_sc_hd__buf_8
XFILLER_133_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput330 _6559_/Q VGND VGND VPWR VPWR wb_dat_o[20] sky130_fd_sc_hd__buf_8
XFILLER_105_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5437_ _5572_/A0 hold519/X _5440_/S VGND VGND VPWR VPWR _7009_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5368_ wire742/X hold390/X _5368_/S VGND VGND VPWR VPWR _6948_/D sky130_fd_sc_hd__mux2_1
X_5299_ wire794/A _6886_/Q _5305_/S VGND VGND VPWR VPWR _6886_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7107_ _7107_/CLK _7107_/D fanout866/X VGND VGND VPWR VPWR _7107_/Q sky130_fd_sc_hd__dfrtp_2
X_4319_ _6765_/Q _6409_/A0 _4321_/S VGND VGND VPWR VPWR _6765_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7038_ _7129_/CLK _7038_/D fanout863/X VGND VGND VPWR VPWR _7038_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_47_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire413 _3338_/Y VGND VGND VPWR VPWR _5315_/A sky130_fd_sc_hd__buf_8
Xwire402 _3361_/Y VGND VGND VPWR VPWR _4234_/S sky130_fd_sc_hd__buf_8
Xwire424 _3325_/Y VGND VGND VPWR VPWR wire424/X sky130_fd_sc_hd__buf_8
XFILLER_167_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire457 _4402_/X VGND VGND VPWR VPWR _4995_/A sky130_fd_sc_hd__buf_8
Xwire435 wire436/X VGND VGND VPWR VPWR _5342_/A sky130_fd_sc_hd__buf_8
Xwire446 wire446/A VGND VGND VPWR VPWR _5558_/A sky130_fd_sc_hd__buf_8
Xwire479 _7109_/Q VGND VGND VPWR VPWR wire479/X sky130_fd_sc_hd__buf_6
XFILLER_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4670_ _4832_/B _4660_/X _4664_/X _4669_/X VGND VGND VPWR VPWR _4670_/X sky130_fd_sc_hd__o211a_1
XFILLER_119_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3621_ _6911_/Q wire424/X _3736_/A2 input45/X _3620_/X VGND VGND VPWR VPWR _3636_/A
+ sky130_fd_sc_hd__a221o_2
X_3552_ hold96/X _3552_/B VGND VGND VPWR VPWR _5218_/A sky130_fd_sc_hd__nor2_8
X_6340_ _6732_/Q wire603/X _6340_/B1 _6598_/Q _6339_/X VGND VGND VPWR VPWR _6343_/C
+ sky130_fd_sc_hd__a221o_4
XFILLER_142_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3483_ _7089_/Q _5522_/A _4118_/A _6598_/Q _3482_/X VGND VGND VPWR VPWR _3488_/C
+ sky130_fd_sc_hd__a221o_1
X_6271_ _6764_/Q wire649/X wire594/X _6719_/Q _6270_/X VGND VGND VPWR VPWR _6271_/X
+ sky130_fd_sc_hd__a221o_1
X_5222_ hold596/X wire769/X _5222_/S VGND VGND VPWR VPWR _6823_/D sky130_fd_sc_hd__mux2_1
X_5153_ _4737_/Y _5152_/X _4692_/C VGND VGND VPWR VPWR _5154_/B sky130_fd_sc_hd__o21a_2
XFILLER_111_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4104_ _6581_/Q wire350/X _4111_/S VGND VGND VPWR VPWR _6581_/D sky130_fd_sc_hd__mux2_1
XFILLER_111_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5084_ _5084_/A _5084_/B VGND VGND VPWR VPWR _5119_/B sky130_fd_sc_hd__or2_1
XFILLER_56_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4035_ _5595_/A0 hold665/X hold73/X VGND VGND VPWR VPWR _4035_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5986_ _6012_/A _6033_/C VGND VGND VPWR VPWR _6004_/A sky130_fd_sc_hd__nand2_8
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4937_ _5033_/A _5033_/B _5033_/C _5035_/C VGND VGND VPWR VPWR _4940_/C sky130_fd_sc_hd__or4_2
XANTENNA_31 _7144_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_20 _4244_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4868_ _4868_/A _4949_/B _4956_/B VGND VGND VPWR VPWR _5087_/D sky130_fd_sc_hd__and3_2
XFILLER_165_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_42 _4256_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6607_ _6623_/CLK _6607_/D fanout872/X VGND VGND VPWR VPWR _6607_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_53 _3562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3819_ _6482_/Q _6481_/Q _3828_/S _6483_/Q VGND VGND VPWR VPWR _3820_/C sky130_fd_sc_hd__a31o_1
XANTENNA_75 _3875_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_64 _3687_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_86 _5144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4799_ _4799_/A _4799_/B _5180_/A _4799_/D VGND VGND VPWR VPWR _4800_/D sky130_fd_sc_hd__or4_1
XANTENNA_97 _5871_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6538_ _6806_/CLK _6538_/D _6435_/A VGND VGND VPWR VPWR _6538_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6469_ _6668_/CLK _6469_/D _6424_/X VGND VGND VPWR VPWR _6469_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_133_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput193 _3214_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[26] sky130_fd_sc_hd__buf_8
Xoutput182 _3224_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[16] sky130_fd_sc_hd__buf_8
XFILLER_121_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput171 _3971_/X VGND VGND VPWR VPWR debug_in sky130_fd_sc_hd__buf_8
XFILLER_0_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5840_ _6883_/Q _5674_/X _5692_/X _7075_/Q VGND VGND VPWR VPWR _5840_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5771_ _6968_/Q _5691_/X wire665/X _6952_/Q VGND VGND VPWR VPWR _5771_/X sky130_fd_sc_hd__a22o_1
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4722_ _4722_/A _4722_/B _4368_/A VGND VGND VPWR VPWR _4812_/C sky130_fd_sc_hd__or3b_4
XFILLER_159_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4653_ _5164_/B _4832_/A VGND VGND VPWR VPWR _4653_/Y sky130_fd_sc_hd__nor2_2
Xinput40 mgmt_gpio_in[13] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__clkbuf_4
Xinput51 mgmt_gpio_in[23] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__buf_4
Xinput62 mgmt_gpio_in[33] VGND VGND VPWR VPWR input62/X sky130_fd_sc_hd__clkbuf_4
Xhold802 _4155_/X VGND VGND VPWR VPWR _6624_/D sky130_fd_sc_hd__bufbuf_16
X_4584_ _4584_/A _4740_/B VGND VGND VPWR VPWR _5005_/C sky130_fd_sc_hd__or2_4
Xinput73 pad_flash_io0_di VGND VGND VPWR VPWR _3964_/B sky130_fd_sc_hd__clkbuf_4
X_3604_ wire485/X _5531_/A _4322_/A _6771_/Q _3603_/X VGND VGND VPWR VPWR _3605_/D
+ sky130_fd_sc_hd__a221o_1
Xinput95 usr1_vcc_pwrgood VGND VGND VPWR VPWR wire836/A sky130_fd_sc_hd__buf_6
Xhold846 _6844_/Q VGND VGND VPWR VPWR hold846/X sky130_fd_sc_hd__bufbuf_16
Xinput84 spimemio_flash_csb VGND VGND VPWR VPWR wire843/A sky130_fd_sc_hd__buf_6
XFILLER_143_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold824 _6807_/Q VGND VGND VPWR VPWR hold824/X sky130_fd_sc_hd__bufbuf_16
Xhold813 _7051_/Q VGND VGND VPWR VPWR hold813/X sky130_fd_sc_hd__bufbuf_16
Xhold835 _7042_/Q VGND VGND VPWR VPWR hold835/X sky130_fd_sc_hd__bufbuf_16
X_3535_ input30/X _3283_/Y hold88/A _7129_/Q VGND VGND VPWR VPWR _3535_/X sky130_fd_sc_hd__a22o_1
X_6323_ _6766_/Q wire649/X wire594/X _6721_/Q _6322_/X VGND VGND VPWR VPWR _6323_/X
+ sky130_fd_sc_hd__a221o_1
X_6254_ _6718_/Q _6295_/B1 _6028_/X _6624_/Q VGND VGND VPWR VPWR _6254_/X sky130_fd_sc_hd__a22o_1
XFILLER_103_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3466_ _6961_/Q _3305_/Y _3763_/B1 _7137_/Q _3465_/X VGND VGND VPWR VPWR _3472_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_170_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5205_ _6411_/A0 _6809_/Q _5206_/S VGND VGND VPWR VPWR _6809_/D sky130_fd_sc_hd__mux2_1
X_3397_ input9/X _3320_/Y _5459_/A _7035_/Q _3392_/X VGND VGND VPWR VPWR _3398_/D
+ sky130_fd_sc_hd__a221o_4
X_6185_ _7194_/Q _5665_/Y _6183_/X _6184_/X VGND VGND VPWR VPWR _7194_/D sky130_fd_sc_hd__o22a_1
XFILLER_111_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5136_ _5136_/A _5136_/B _5136_/C _5136_/D VGND VGND VPWR VPWR _5137_/C sky130_fd_sc_hd__or4_1
XFILLER_57_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5067_ _4469_/A _4819_/A _4603_/B _4740_/B VGND VGND VPWR VPWR _5067_/X sky130_fd_sc_hd__a211o_2
XFILLER_84_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4018_ hold483/X _4017_/X _4024_/S VGND VGND VPWR VPWR _4018_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5969_ _6777_/Q wire694/X wire660/X _6608_/Q _5968_/X VGND VGND VPWR VPWR _5976_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_40_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold109 _3263_/X VGND VGND VPWR VPWR _3264_/B sky130_fd_sc_hd__bufbuf_16
XFILLER_171_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3320_ _5225_/A _3375_/B VGND VGND VPWR VPWR _3320_/Y sky130_fd_sc_hd__nor2_8
XFILLER_140_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ hold236/X hold117/X _3953_/A VGND VGND VPWR VPWR _3251_/X sky130_fd_sc_hd__mux2_8
XFILLER_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6941_ _7068_/CLK _6941_/D fanout878/X VGND VGND VPWR VPWR _6941_/Q sky130_fd_sc_hd__dfstp_4
X_6872_ _6930_/CLK _6872_/D fanout885/X VGND VGND VPWR VPWR _6872_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5823_ _7106_/Q _5857_/A2 wire692/A _6994_/Q _5822_/X VGND VGND VPWR VPWR _5826_/C
+ sky130_fd_sc_hd__a221o_1
X_5754_ _6959_/Q wire707/X wire680/X wire528/X VGND VGND VPWR VPWR _5754_/X sky130_fd_sc_hd__a22o_1
X_4705_ _5023_/B _4724_/B VGND VGND VPWR VPWR _5166_/A sky130_fd_sc_hd__nor2_2
XFILLER_147_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5685_ _7165_/Q _5707_/B _5701_/C VGND VGND VPWR VPWR _5685_/X sky130_fd_sc_hd__and3_4
XFILLER_108_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4636_ _4636_/A _4989_/A VGND VGND VPWR VPWR _5136_/B sky130_fd_sc_hd__nor2_2
Xhold621 _6944_/Q VGND VGND VPWR VPWR hold621/X sky130_fd_sc_hd__bufbuf_16
Xhold610 _7007_/Q VGND VGND VPWR VPWR hold610/X sky130_fd_sc_hd__bufbuf_16
XFILLER_190_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6306_ _6306_/A _6306_/B _6306_/C VGND VGND VPWR VPWR _6306_/X sky130_fd_sc_hd__or3_4
X_4567_ _4694_/A _4947_/B _6707_/Q VGND VGND VPWR VPWR _4567_/X sky130_fd_sc_hd__o21a_1
Xhold643 _6564_/Q VGND VGND VPWR VPWR hold643/X sky130_fd_sc_hd__bufbuf_16
Xhold654 _7140_/Q VGND VGND VPWR VPWR hold654/X sky130_fd_sc_hd__bufbuf_16
Xhold632 _5259_/X VGND VGND VPWR VPWR _6851_/D sky130_fd_sc_hd__bufbuf_16
Xhold665 _6522_/Q VGND VGND VPWR VPWR hold665/X sky130_fd_sc_hd__bufbuf_16
XFILLER_143_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4498_ _4986_/A _4745_/B VGND VGND VPWR VPWR _5119_/A sky130_fd_sc_hd__nor2_4
XFILLER_116_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3518_ _3543_/A _3733_/B VGND VGND VPWR VPWR _4124_/A sky130_fd_sc_hd__nor2_8
XFILLER_104_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold687 _7044_/Q VGND VGND VPWR VPWR hold687/X sky130_fd_sc_hd__bufbuf_16
Xhold676 _7100_/Q VGND VGND VPWR VPWR hold676/X sky130_fd_sc_hd__bufbuf_16
X_6237_ _6728_/Q wire604/X _6301_/B1 _6609_/Q VGND VGND VPWR VPWR _6237_/X sky130_fd_sc_hd__a22o_1
XFILLER_77_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3449_ wire907/X _3571_/A2 _5576_/A _7138_/Q _3448_/X VGND VGND VPWR VPWR _3450_/D
+ sky130_fd_sc_hd__a221o_4
Xhold698 _7222_/Q VGND VGND VPWR VPWR hold698/X sky130_fd_sc_hd__bufbuf_16
XFILLER_134_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6168_ _7074_/Q _6009_/X _6012_/X _6970_/Q VGND VGND VPWR VPWR _6168_/X sky130_fd_sc_hd__a22o_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5119_ _5119_/A _5119_/B _5119_/C VGND VGND VPWR VPWR _5135_/C sky130_fd_sc_hd__or3_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6099_ _7127_/Q wire598/X wire610/X wire519/X _6098_/X VGND VGND VPWR VPWR _6107_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A VGND VGND VPWR VPWR _7218_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_53_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5470_ _5578_/A0 _7038_/Q _5476_/S VGND VGND VPWR VPWR _7038_/D sky130_fd_sc_hd__mux2_1
X_4421_ _4728_/A _4671_/A VGND VGND VPWR VPWR _4702_/A sky130_fd_sc_hd__nor2_2
XFILLER_117_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4352_ _4352_/A _4352_/B _4352_/C VGND VGND VPWR VPWR _4529_/B sky130_fd_sc_hd__and3_4
X_7140_ _7140_/CLK _7140_/D fanout867/X VGND VGND VPWR VPWR _7140_/Q sky130_fd_sc_hd__dfrtp_2
X_4283_ _5498_/A0 _6735_/Q _4285_/S VGND VGND VPWR VPWR _6735_/D sky130_fd_sc_hd__mux2_1
XFILLER_125_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7071_ _7118_/CLK _7071_/D fanout869/X VGND VGND VPWR VPWR _7071_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_4_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3303_ _7028_/Q _3301_/Y _3302_/Y input28/X _3300_/X VGND VGND VPWR VPWR _3331_/A
+ sky130_fd_sc_hd__a221o_1
X_6022_ _6022_/A _6022_/B _6022_/C _6022_/D VGND VGND VPWR VPWR _6024_/C sky130_fd_sc_hd__or4_1
X_3234_ _6904_/Q VGND VGND VPWR VPWR _3234_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_58_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6924_ _6985_/CLK _6924_/D fanout878/X VGND VGND VPWR VPWR _6924_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_54_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6855_ _6996_/CLK _6855_/D fanout869/X VGND VGND VPWR VPWR _6855_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5806_ _5806_/A _5806_/B _5806_/C _5806_/D VGND VGND VPWR VPWR _5806_/X sky130_fd_sc_hd__or4_4
X_3998_ _6498_/Q _6409_/A0 _4003_/S VGND VGND VPWR VPWR _6498_/D sky130_fd_sc_hd__mux2_1
XFILLER_10_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6786_ _7225_/CLK _6786_/D fanout851/X VGND VGND VPWR VPWR _6786_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_148_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire809 _3241_/Y VGND VGND VPWR VPWR _5963_/B sky130_fd_sc_hd__buf_8
Xmax_length407 _3353_/Y VGND VGND VPWR VPWR _5288_/A sky130_fd_sc_hd__buf_6
X_5737_ _7014_/Q wire697/X wire662/X wire551/X VGND VGND VPWR VPWR _5737_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length418 _3736_/A2 VGND VGND VPWR VPWR _3571_/A2 sky130_fd_sc_hd__buf_6
Xmax_length429 wire430/X VGND VGND VPWR VPWR _3657_/A2 sky130_fd_sc_hd__buf_6
XFILLER_175_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5668_ _7163_/Q _7164_/Q VGND VGND VPWR VPWR _5706_/B sky130_fd_sc_hd__and2b_4
X_5599_ _5599_/A0 hold269/X hold66/X VGND VGND VPWR VPWR _7153_/D sky130_fd_sc_hd__mux2_1
XFILLER_151_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4619_ _4619_/A _4619_/B _4619_/C _4619_/D VGND VGND VPWR VPWR _4619_/X sky130_fd_sc_hd__and4_2
XFILLER_135_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold440 _6714_/Q VGND VGND VPWR VPWR hold440/X sky130_fd_sc_hd__bufbuf_16
Xhold451 _7066_/Q VGND VGND VPWR VPWR hold451/X sky130_fd_sc_hd__bufbuf_16
Xhold462 _6729_/Q VGND VGND VPWR VPWR hold462/X sky130_fd_sc_hd__bufbuf_16
Xhold495 _4022_/X VGND VGND VPWR VPWR _6512_/D sky130_fd_sc_hd__bufbuf_16
Xhold484 _4018_/X VGND VGND VPWR VPWR _6510_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_145_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold473 _6652_/Q VGND VGND VPWR VPWR hold473/X sky130_fd_sc_hd__bufbuf_16
XFILLER_77_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_324 wire763/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_302 _6856_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_313 wire594/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_335 hold409/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_346 hold59/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4970_ _5147_/A _4970_/B _4959_/A VGND VGND VPWR VPWR _4970_/X sky130_fd_sc_hd__or3b_1
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3921_ _3921_/A _3921_/B VGND VGND VPWR VPWR _5606_/B sky130_fd_sc_hd__nor2_1
XFILLER_32_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3852_ _6487_/Q _6486_/Q _6485_/Q _6664_/Q VGND VGND VPWR VPWR _3853_/S sky130_fd_sc_hd__or4b_1
X_6640_ _6642_/CLK _6640_/D fanout856/X VGND VGND VPWR VPWR _6640_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_177_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6571_ _7208_/CLK _6571_/D VGND VGND VPWR VPWR _6571_/Q sky130_fd_sc_hd__dfxtp_4
X_5522_ _5522_/A _5576_/B VGND VGND VPWR VPWR _5530_/S sky130_fd_sc_hd__nand2_8
X_3783_ _6989_/Q _5414_/A _5531_/A wire487/X VGND VGND VPWR VPWR _3783_/X sky130_fd_sc_hd__a22o_2
XFILLER_185_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5453_ wire780/X hold605/X _5458_/S VGND VGND VPWR VPWR _5453_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_42_csclk _6987_/CLK VGND VGND VPWR VPWR _6979_/CLK sky130_fd_sc_hd__clkbuf_8
X_5384_ _5600_/A0 hold453/X _5386_/S VGND VGND VPWR VPWR _6962_/D sky130_fd_sc_hd__mux2_1
X_4404_ _4553_/A _4405_/B VGND VGND VPWR VPWR _4845_/A sky130_fd_sc_hd__nor2_8
XFILLER_132_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4335_ _4707_/B _5050_/A VGND VGND VPWR VPWR _4728_/A sky130_fd_sc_hd__nand2_8
X_7123_ _7139_/CLK _7123_/D fanout867/X VGND VGND VPWR VPWR _7123_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_99_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7054_ _7153_/CLK _7054_/D fanout881/X VGND VGND VPWR VPWR _7054_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_140_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4266_ hold728/X _6410_/A0 _4267_/S VGND VGND VPWR VPWR _6721_/D sky130_fd_sc_hd__mux2_1
X_3217_ _3217_/A VGND VGND VPWR VPWR _3217_/Y sky130_fd_sc_hd__inv_2
X_6005_ _6014_/A _6010_/B VGND VGND VPWR VPWR _6025_/B sky130_fd_sc_hd__nor2_4
XFILLER_67_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_57_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7107_/CLK sky130_fd_sc_hd__clkbuf_8
X_4197_ wire799/A hold565/X _4201_/S VGND VGND VPWR VPWR _6659_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6907_ _6979_/CLK _6907_/D fanout878/X VGND VGND VPWR VPWR _6907_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_24_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6838_ _6842_/CLK _6838_/D fanout857/X VGND VGND VPWR VPWR _6838_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_168_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire606 _6037_/X VGND VGND VPWR VPWR _6335_/B sky130_fd_sc_hd__buf_8
XFILLER_136_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire639 _6021_/C VGND VGND VPWR VPWR wire639/X sky130_fd_sc_hd__buf_8
Xwire628 _6012_/X VGND VGND VPWR VPWR _6020_/D sky130_fd_sc_hd__buf_6
XFILLER_7_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6769_ _6771_/CLK _6769_/D fanout853/X VGND VGND VPWR VPWR _6769_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_109_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold270 _6971_/Q VGND VGND VPWR VPWR hold270/X sky130_fd_sc_hd__bufbuf_16
Xhold281 _5278_/X VGND VGND VPWR VPWR _6868_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_172_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold292 _7155_/Q VGND VGND VPWR VPWR hold292/X sky130_fd_sc_hd__bufbuf_16
XFILLER_2_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout772 hold83/A VGND VGND VPWR VPWR wire773/A sky130_fd_sc_hd__buf_6
Xfanout761 hold154/X VGND VGND VPWR VPWR hold155/A sky130_fd_sc_hd__buf_6
XFILLER_93_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_143 mgmt_gpio_in[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_110 _6835_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_121 _6473_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_132 mask_rev_in[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_176 _6384_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_165 wb_dat_i[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_154 spi_sdo VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_187 _5501_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_198 wire477/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4120_ hold535/X wire790/X _4123_/S VGND VGND VPWR VPWR _6595_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4051_ hold691/X _6408_/A0 _4054_/S VGND VGND VPWR VPWR _6536_/D sky130_fd_sc_hd__mux2_1
XFILLER_37_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput5 mask_rev_in[10] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4953_ _4953_/A _4965_/B VGND VGND VPWR VPWR _5068_/B sky130_fd_sc_hd__nor2_1
XFILLER_52_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3904_ _6012_/A _6037_/A VGND VGND VPWR VPWR _6030_/A sky130_fd_sc_hd__nand2_8
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4884_ _4898_/B _4756_/B _4623_/A VGND VGND VPWR VPWR _4907_/A sky130_fd_sc_hd__o21ai_2
X_6623_ _6623_/CLK _6623_/D fanout890/X VGND VGND VPWR VPWR _6623_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_32_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3835_ _3834_/X hold40/A _3840_/S VGND VGND VPWR VPWR _6479_/D sky130_fd_sc_hd__mux2_1
XFILLER_32_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6554_ _6554_/CLK _6554_/D fanout858/X VGND VGND VPWR VPWR _6554_/Q sky130_fd_sc_hd__dfrtp_2
X_3766_ _7005_/Q _5432_/A _4322_/A _6768_/Q VGND VGND VPWR VPWR _3766_/X sky130_fd_sc_hd__a22o_1
XFILLER_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6485_ _6668_/CLK _6485_/D _6440_/X VGND VGND VPWR VPWR _6485_/Q sky130_fd_sc_hd__dfrtp_2
X_5505_ _5532_/A0 _7069_/Q _5512_/S VGND VGND VPWR VPWR _7069_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5436_ wire769/X hold620/X _5440_/S VGND VGND VPWR VPWR _7008_/D sky130_fd_sc_hd__mux2_1
X_3697_ _6655_/Q _4190_/A _6406_/A _7222_/Q wire367/X VGND VGND VPWR VPWR _3699_/C
+ sky130_fd_sc_hd__a221o_2
XFILLER_160_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput342 _7210_/Q VGND VGND VPWR VPWR wb_dat_o[31] sky130_fd_sc_hd__buf_8
XFILLER_145_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput331 _6560_/Q VGND VGND VPWR VPWR wb_dat_o[21] sky130_fd_sc_hd__buf_8
Xoutput320 _6571_/Q VGND VGND VPWR VPWR wb_dat_o[11] sky130_fd_sc_hd__buf_8
XFILLER_99_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5367_ wire749/X hold492/X _5368_/S VGND VGND VPWR VPWR _5367_/X sky130_fd_sc_hd__mux2_1
X_5298_ _5595_/A0 _6885_/Q _5305_/S VGND VGND VPWR VPWR _6885_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7106_ _7107_/CLK _7106_/D fanout866/X VGND VGND VPWR VPWR _7106_/Q sky130_fd_sc_hd__dfrtp_2
X_4318_ hold712/X _6408_/A0 _4321_/S VGND VGND VPWR VPWR _6764_/D sky130_fd_sc_hd__mux2_1
X_4249_ _5602_/A0 hold314/X hold32/X VGND VGND VPWR VPWR _4249_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7037_ _7105_/CLK _7037_/D fanout861/X VGND VGND VPWR VPWR _7037_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_142_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire403 _3361_/Y VGND VGND VPWR VPWR _4232_/S sky130_fd_sc_hd__buf_8
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire458 _3945_/X VGND VGND VPWR VPWR wire458/X sky130_fd_sc_hd__buf_6
Xwire436 _3306_/Y VGND VGND VPWR VPWR wire436/X sky130_fd_sc_hd__buf_8
XFILLER_51_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire469 _7223_/Q VGND VGND VPWR VPWR wire469/X sky130_fd_sc_hd__clkbuf_8
XFILLER_109_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3620_ _7143_/Q _5585_/A _4280_/A _6735_/Q VGND VGND VPWR VPWR _3620_/X sky130_fd_sc_hd__a22o_1
XFILLER_128_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3551_ _3551_/A _5225_/B VGND VGND VPWR VPWR _3551_/Y sky130_fd_sc_hd__nor2_4
XFILLER_155_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3482_ wire500/X _3298_/Y _4082_/A _6567_/Q VGND VGND VPWR VPWR _3482_/X sky130_fd_sc_hd__a22o_1
X_6270_ _6551_/Q wire601/X wire580/X _6630_/Q VGND VGND VPWR VPWR _6270_/X sky130_fd_sc_hd__a22o_2
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5221_ hold768/X _5255_/A0 _5222_/S VGND VGND VPWR VPWR _6822_/D sky130_fd_sc_hd__mux2_1
X_5152_ _5062_/C _5050_/C _5041_/X _4668_/B VGND VGND VPWR VPWR _5152_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_111_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4103_ _6701_/Q _6362_/B VGND VGND VPWR VPWR _4111_/S sky130_fd_sc_hd__and2_4
XFILLER_110_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5083_ _5137_/A _5171_/B _5115_/A _5117_/A VGND VGND VPWR VPWR _5083_/X sky130_fd_sc_hd__or4_2
XFILLER_57_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4034_ _4034_/A _4241_/A _6421_/B hold31/X VGND VGND VPWR VPWR hold73/A sky130_fd_sc_hd__or4_4
XFILLER_65_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5985_ _7169_/Q _7168_/Q VGND VGND VPWR VPWR _6033_/C sky130_fd_sc_hd__nor2_8
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4936_ _4936_/A _4936_/B _4936_/C VGND VGND VPWR VPWR _5035_/C sky130_fd_sc_hd__or3_1
XFILLER_33_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_32 _7146_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4867_ _4818_/A _4740_/A _4452_/Y _4866_/X VGND VGND VPWR VPWR _4867_/X sky130_fd_sc_hd__a31o_1
XANTENNA_10 _6478_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 _6801_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_43 _4256_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6606_ _6747_/CLK _6606_/D fanout874/X VGND VGND VPWR VPWR _6606_/Q sky130_fd_sc_hd__dfstp_4
X_3818_ _6484_/Q _3840_/S _3817_/Y VGND VGND VPWR VPWR _6484_/D sky130_fd_sc_hd__a21o_1
XANTENNA_54 _3598_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_65 _3687_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 _4217_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4798_ _4798_/A _5022_/B _4798_/C _4798_/D VGND VGND VPWR VPWR _4799_/D sky130_fd_sc_hd__or4_1
XFILLER_119_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_87 _4763_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_98 _5871_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6537_ _6806_/CLK _6537_/D _6435_/A VGND VGND VPWR VPWR _6537_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_21_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3749_ _6965_/Q wire421/A _4154_/A _6624_/Q _3748_/X VGND VGND VPWR VPWR _3754_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6468_ _6668_/CLK _6468_/D _6423_/X VGND VGND VPWR VPWR _6468_/Q sky130_fd_sc_hd__dfrtp_2
X_6399_ _4236_/B _6399_/A2 _6399_/B1 _4238_/B _6398_/X VGND VGND VPWR VPWR _6399_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_133_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5419_ _5572_/A0 hold508/X _5422_/S VGND VGND VPWR VPWR _6993_/D sky130_fd_sc_hd__mux2_1
Xoutput194 _3213_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[27] sky130_fd_sc_hd__buf_8
Xoutput183 _3223_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[17] sky130_fd_sc_hd__buf_8
Xoutput172 _6825_/Q VGND VGND VPWR VPWR irq[0] sky130_fd_sc_hd__buf_8
XFILLER_153_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5770_ _3217_/A _5803_/B1 wire659/X _6936_/Q _5769_/X VGND VGND VPWR VPWR _5777_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4721_ _4818_/C _4724_/B _4238_/B VGND VGND VPWR VPWR _5003_/B sky130_fd_sc_hd__o21a_2
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4652_ _4758_/B _4652_/B VGND VGND VPWR VPWR _4832_/A sky130_fd_sc_hd__nand2_8
XFILLER_30_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput30 mask_rev_in[4] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__clkbuf_4
X_3603_ _3877_/C _4232_/S _4262_/A _6721_/Q _3602_/X VGND VGND VPWR VPWR _3603_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_190_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput52 mgmt_gpio_in[24] VGND VGND VPWR VPWR input52/X sky130_fd_sc_hd__clkbuf_4
XFILLER_162_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput41 mgmt_gpio_in[14] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__clkbuf_4
X_4583_ _4584_/A _4740_/B VGND VGND VPWR VPWR _4736_/B sky130_fd_sc_hd__nor2_8
Xinput63 mgmt_gpio_in[34] VGND VGND VPWR VPWR wire899/A sky130_fd_sc_hd__buf_6
XFILLER_116_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold803 _6798_/Q VGND VGND VPWR VPWR hold803/X sky130_fd_sc_hd__bufbuf_16
Xinput96 usr1_vdd_pwrgood VGND VGND VPWR VPWR wire835/A sky130_fd_sc_hd__buf_6
Xinput85 spimemio_flash_io0_do VGND VGND VPWR VPWR wire842/A sky130_fd_sc_hd__buf_6
XFILLER_115_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6322_ _6553_/Q wire601/X wire580/X _6632_/Q VGND VGND VPWR VPWR _6322_/X sky130_fd_sc_hd__a22o_4
Xhold814 _7050_/Q VGND VGND VPWR VPWR hold814/X sky130_fd_sc_hd__bufbuf_16
Xhold825 _6858_/Q VGND VGND VPWR VPWR hold825/X sky130_fd_sc_hd__bufbuf_16
Xinput74 pad_flash_io1_di VGND VGND VPWR VPWR _3965_/B sky130_fd_sc_hd__clkbuf_4
X_3534_ _3534_/A _5252_/A VGND VGND VPWR VPWR _4262_/A sky130_fd_sc_hd__nor2_8
Xhold836 _7082_/Q VGND VGND VPWR VPWR hold836/X sky130_fd_sc_hd__bufbuf_16
Xhold847 _6695_/Q VGND VGND VPWR VPWR hold847/X sky130_fd_sc_hd__bufbuf_16
XFILLER_89_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3465_ _6897_/Q _3352_/Y _4190_/A wire569/X VGND VGND VPWR VPWR _3465_/X sky130_fd_sc_hd__a22o_1
X_6253_ _6629_/Q wire580/X _6339_/B1 _6768_/Q VGND VGND VPWR VPWR _6253_/X sky130_fd_sc_hd__a22o_1
XFILLER_103_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5204_ _6410_/A0 hold708/X _5206_/S VGND VGND VPWR VPWR _6808_/D sky130_fd_sc_hd__mux2_1
X_3396_ wire532/X _5351_/A _5369_/A _6955_/Q _3387_/X VGND VGND VPWR VPWR _3398_/C
+ sky130_fd_sc_hd__a221o_4
X_6184_ _5611_/A _7193_/Q _5664_/X VGND VGND VPWR VPWR _6184_/X sky130_fd_sc_hd__a21o_1
XFILLER_97_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5135_ _5135_/A _5135_/B _5135_/C _5135_/D VGND VGND VPWR VPWR _5172_/A sky130_fd_sc_hd__or4_1
X_5066_ _5066_/A _5124_/B VGND VGND VPWR VPWR _5074_/A sky130_fd_sc_hd__nand2_1
XFILLER_96_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4017_ _6526_/Q hold150/X _4021_/S VGND VGND VPWR VPWR _4017_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5968_ _6732_/Q wire710/X wire689/X _6643_/Q VGND VGND VPWR VPWR _5968_/X sky130_fd_sc_hd__a22o_1
X_4919_ _4395_/D _4469_/Y _4656_/X _4796_/B _4412_/Y VGND VGND VPWR VPWR _5095_/B
+ sky130_fd_sc_hd__a311o_4
XFILLER_138_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5899_ _6625_/Q _5963_/B VGND VGND VPWR VPWR _5899_/X sky130_fd_sc_hd__or2_1
XFILLER_21_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_494 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ hold108/X _3845_/A hold235/X VGND VGND VPWR VPWR _3250_/X sky130_fd_sc_hd__a21bo_2
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6940_ _7156_/CLK _6940_/D fanout884/X VGND VGND VPWR VPWR _6940_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6871_ _7111_/CLK _6871_/D fanout875/X VGND VGND VPWR VPWR _6871_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_179_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5822_ _6882_/Q wire706/X _5855_/B1 _7034_/Q VGND VGND VPWR VPWR _5822_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5753_ _5753_/A _5753_/B _5753_/C _5753_/D VGND VGND VPWR VPWR _5753_/X sky130_fd_sc_hd__or4_2
XFILLER_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4704_ _4772_/A _4711_/C _4772_/C VGND VGND VPWR VPWR _4704_/X sky130_fd_sc_hd__and3_4
XFILLER_148_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5684_ _7165_/Q _5703_/B _5707_/B VGND VGND VPWR VPWR _5684_/X sky130_fd_sc_hd__and3_4
XFILLER_163_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4635_ _4996_/A _4844_/A _4631_/X _4633_/X _5144_/A VGND VGND VPWR VPWR _4635_/X
+ sky130_fd_sc_hd__o2111a_1
X_4566_ _4566_/A _4740_/B VGND VGND VPWR VPWR _4592_/B sky130_fd_sc_hd__or2_4
XFILLER_162_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold611 _5435_/X VGND VGND VPWR VPWR _7007_/D sky130_fd_sc_hd__bufbuf_16
Xhold600 _7016_/Q VGND VGND VPWR VPWR hold600/X sky130_fd_sc_hd__bufbuf_16
Xhold633 _6864_/Q VGND VGND VPWR VPWR hold633/X sky130_fd_sc_hd__bufbuf_16
Xhold622 _7056_/Q VGND VGND VPWR VPWR hold622/X sky130_fd_sc_hd__bufbuf_16
XFILLER_150_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6305_ _6305_/A _6305_/B _6305_/C _6305_/D VGND VGND VPWR VPWR _6306_/C sky130_fd_sc_hd__or4_1
X_3517_ _7009_/Q _5432_/A wire430/X _7065_/Q _3516_/X VGND VGND VPWR VPWR _3522_/C
+ sky130_fd_sc_hd__a221o_2
Xhold644 _6850_/Q VGND VGND VPWR VPWR hold644/X sky130_fd_sc_hd__bufbuf_16
XFILLER_171_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold666 _4035_/X VGND VGND VPWR VPWR _6522_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_143_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4497_ _5164_/B _4745_/B VGND VGND VPWR VPWR _5013_/A sky130_fd_sc_hd__nor2_4
XFILLER_104_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold688 _6771_/Q VGND VGND VPWR VPWR hold688/X sky130_fd_sc_hd__bufbuf_16
Xhold655 _5584_/X VGND VGND VPWR VPWR _7140_/D sky130_fd_sc_hd__bufbuf_16
Xhold677 _6688_/Q VGND VGND VPWR VPWR hold677/X sky130_fd_sc_hd__bufbuf_16
X_6236_ _6743_/Q wire598/X _6020_/D _6708_/Q VGND VGND VPWR VPWR _6248_/A sky130_fd_sc_hd__a22o_1
Xhold699 _6631_/Q VGND VGND VPWR VPWR hold699/X sky130_fd_sc_hd__bufbuf_16
X_3448_ wire504/X _5477_/A _5297_/A _6890_/Q VGND VGND VPWR VPWR _3448_/X sky130_fd_sc_hd__a22o_2
XFILLER_134_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3379_ _3379_/A _3379_/B _3379_/C VGND VGND VPWR VPWR _3379_/X sky130_fd_sc_hd__or3_2
X_6167_ wire475/X _6017_/Y _6030_/Y _7034_/Q _6166_/X VGND VGND VPWR VPWR _6170_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _5118_/A _5118_/B _5118_/C _5118_/D VGND VGND VPWR VPWR _5119_/C sky130_fd_sc_hd__or4_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6098_ _6887_/Q wire602/X wire581/X _7143_/Q _6097_/X VGND VGND VPWR VPWR _6098_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_85_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5049_ _4956_/C _4668_/B _5041_/X _4657_/B VGND VGND VPWR VPWR _5049_/X sky130_fd_sc_hd__a22o_1
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4420_ _4654_/A _4707_/B _5050_/A VGND VGND VPWR VPWR _4422_/B sky130_fd_sc_hd__and3_2
XFILLER_145_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4351_ _4351_/A _4351_/B _4351_/C _4351_/D VGND VGND VPWR VPWR _4352_/C sky130_fd_sc_hd__and4_1
XFILLER_125_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3302_ _3365_/A _5225_/A VGND VGND VPWR VPWR _3302_/Y sky130_fd_sc_hd__nor2_8
X_7070_ _7129_/CLK _7070_/D fanout863/X VGND VGND VPWR VPWR _7070_/Q sky130_fd_sc_hd__dfstp_4
X_4282_ wire790/X hold547/X _4285_/S VGND VGND VPWR VPWR _4282_/X sky130_fd_sc_hd__mux2_1
X_6021_ _6021_/A _6021_/B _6021_/C _6021_/D VGND VGND VPWR VPWR _6024_/B sky130_fd_sc_hd__or4_1
XFILLER_101_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3233_ _3233_/A VGND VGND VPWR VPWR _3233_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_1_csclk clkbuf_1_1_1_csclk/A VGND VGND VPWR VPWR clkbuf_2_3_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_104_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6923_ _6979_/CLK _6923_/D fanout878/X VGND VGND VPWR VPWR _6923_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_82_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6854_ _7036_/CLK _6854_/D fanout869/X VGND VGND VPWR VPWR _6854_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_168_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5805_ _6977_/Q _5676_/X wire691/X _7089_/Q _5804_/X VGND VGND VPWR VPWR _5806_/D
+ sky130_fd_sc_hd__a221o_2
X_3997_ _6497_/Q _6408_/A0 _4003_/S VGND VGND VPWR VPWR _6497_/D sky130_fd_sc_hd__mux2_1
X_6785_ _6787_/CLK _6785_/D fanout850/X VGND VGND VPWR VPWR _6785_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5736_ _6902_/Q _5814_/A2 _5725_/X _5735_/X VGND VGND VPWR VPWR _5736_/X sky130_fd_sc_hd__a211o_4
Xmax_length419 hold46/X VGND VGND VPWR VPWR _4209_/S sky130_fd_sc_hd__buf_6
XFILLER_148_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5667_ _7165_/Q _5703_/B _5704_/B VGND VGND VPWR VPWR _5667_/X sky130_fd_sc_hd__and3_4
XFILLER_108_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4618_ _4844_/A _4749_/C _4617_/A VGND VGND VPWR VPWR _4619_/D sky130_fd_sc_hd__a21o_1
XFILLER_190_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5598_ _5598_/A0 hold587/X hold66/X VGND VGND VPWR VPWR _7152_/D sky130_fd_sc_hd__mux2_1
XFILLER_135_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold463 hold511/X VGND VGND VPWR VPWR hold512/A sky130_fd_sc_hd__bufbuf_16
Xhold452 _6906_/Q VGND VGND VPWR VPWR hold452/X sky130_fd_sc_hd__bufbuf_16
Xhold430 _6610_/Q VGND VGND VPWR VPWR hold430/X sky130_fd_sc_hd__bufbuf_16
XFILLER_144_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4549_ _4987_/B _4624_/B _5114_/A _4548_/X VGND VGND VPWR VPWR _4549_/X sky130_fd_sc_hd__a211o_1
XFILLER_104_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold441 _6662_/Q VGND VGND VPWR VPWR hold441/X sky130_fd_sc_hd__bufbuf_16
Xhold474 _6874_/Q VGND VGND VPWR VPWR hold474/X sky130_fd_sc_hd__bufbuf_16
XFILLER_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold485 _7136_/Q VGND VGND VPWR VPWR hold485/X sky130_fd_sc_hd__bufbuf_16
Xhold496 _7072_/Q VGND VGND VPWR VPWR hold496/X sky130_fd_sc_hd__bufbuf_16
XFILLER_1_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6219_ _6219_/A _6219_/B _6219_/C _6219_/D VGND VGND VPWR VPWR _6219_/X sky130_fd_sc_hd__or4_1
X_7199_ _7220_/CLK _7199_/D fanout854/X VGND VGND VPWR VPWR _7199_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_57_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_314 wire616/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_303 _6740_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_325 _6410_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_336 hold502/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_347 wire548/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3920_ _5611_/A _3920_/B VGND VGND VPWR VPWR _3920_/Y sky130_fd_sc_hd__nand2_1
XFILLER_72_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3851_ _3797_/X _3898_/A _3850_/Y _6664_/Q VGND VGND VPWR VPWR _6472_/D sky130_fd_sc_hd__a211oi_2
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6570_ _7208_/CLK _6570_/D VGND VGND VPWR VPWR _6570_/Q sky130_fd_sc_hd__dfxtp_2
X_3782_ _7061_/Q _5495_/A _5540_/A _7101_/Q _3781_/X VGND VGND VPWR VPWR _3785_/C
+ sky130_fd_sc_hd__a221o_4
XFILLER_164_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5521_ wire739/X hold673/X _5521_/S VGND VGND VPWR VPWR _7084_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5452_ _5578_/A0 _7022_/Q _5458_/S VGND VGND VPWR VPWR _7022_/D sky130_fd_sc_hd__mux2_1
X_5383_ hold150/X hold227/X _5386_/S VGND VGND VPWR VPWR _6961_/D sky130_fd_sc_hd__mux2_1
X_4403_ _4671_/A _4617_/A VGND VGND VPWR VPWR _4847_/A sky130_fd_sc_hd__nor2_2
XFILLER_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7122_ _7122_/CLK _7122_/D fanout888/X VGND VGND VPWR VPWR _7122_/Q sky130_fd_sc_hd__dfrtp_2
X_4334_ _4707_/B _5050_/A VGND VGND VPWR VPWR _4696_/A sky130_fd_sc_hd__and2_4
XFILLER_141_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7053_ _7128_/CLK _7053_/D _6421_/A VGND VGND VPWR VPWR _7053_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_141_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4265_ hold760/X _5498_/A0 _4267_/S VGND VGND VPWR VPWR _4265_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6004_ _6004_/A _6014_/A VGND VGND VPWR VPWR _6023_/C sky130_fd_sc_hd__nor2_8
X_3216_ _3216_/A VGND VGND VPWR VPWR _3216_/Y sky130_fd_sc_hd__inv_2
X_4196_ _4196_/A _5242_/B VGND VGND VPWR VPWR _4201_/S sky130_fd_sc_hd__nand2_4
XFILLER_82_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6906_ _7154_/CLK _6906_/D fanout886/X VGND VGND VPWR VPWR _6906_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_70_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6837_ _6842_/CLK _6837_/D fanout857/X VGND VGND VPWR VPWR _6837_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_24_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire618 wire618/A VGND VGND VPWR VPWR wire618/X sky130_fd_sc_hd__buf_6
X_6768_ _6771_/CLK _6768_/D fanout853/X VGND VGND VPWR VPWR _6768_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_136_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5719_ _6917_/Q _5681_/X _5682_/X _7013_/Q _5677_/X VGND VGND VPWR VPWR _5720_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_109_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6699_ _7208_/CLK _6699_/D _6362_/B VGND VGND VPWR VPWR _6704_/D sky130_fd_sc_hd__dfrtp_2
XFILLER_40_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold271 _6953_/Q VGND VGND VPWR VPWR hold271/X sky130_fd_sc_hd__bufbuf_16
XFILLER_2_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold260 _5534_/X VGND VGND VPWR VPWR _7095_/D sky130_fd_sc_hd__bufbuf_16
Xhold293 _5601_/X VGND VGND VPWR VPWR _7155_/D sky130_fd_sc_hd__bufbuf_16
Xhold282 _6970_/Q VGND VGND VPWR VPWR hold282/X sky130_fd_sc_hd__bufbuf_16
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout740 hold21/X VGND VGND VPWR VPWR _5602_/A0 sky130_fd_sc_hd__buf_8
XFILLER_172_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout751 wire756/X VGND VGND VPWR VPWR wire753/A sky130_fd_sc_hd__buf_6
Xfanout795 hold36/X VGND VGND VPWR VPWR hold37/A sky130_fd_sc_hd__buf_8
XFILLER_92_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_100 _6009_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_133 _6508_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_122 _6476_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_111 debug_mode VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_166 wb_dat_i[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_144 mgmt_gpio_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_155 spi_sdoenb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_177 _6398_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_188 _6356_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_199 wire479/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length750 hold56/X VGND VGND VPWR VPWR hold57/A sky130_fd_sc_hd__buf_6
XFILLER_154_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length783 _5336_/A1 VGND VGND VPWR VPWR _5408_/A1 sky130_fd_sc_hd__buf_6
XFILLER_115_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4050_ hold743/X _6407_/A0 _4054_/S VGND VGND VPWR VPWR _6535_/D sky130_fd_sc_hd__mux2_1
Xinput6 mask_rev_in[11] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_4
XFILLER_37_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4952_ _4949_/A _4956_/A _4736_/B _4983_/B VGND VGND VPWR VPWR _5142_/B sky130_fd_sc_hd__a31o_2
XFILLER_17_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4883_ _4883_/A _4922_/A VGND VGND VPWR VPWR _4983_/B sky130_fd_sc_hd__or2_2
X_3903_ _7169_/Q _7168_/Q VGND VGND VPWR VPWR _6037_/A sky130_fd_sc_hd__and2b_4
XFILLER_189_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6622_ _6623_/CLK _6622_/D fanout872/X VGND VGND VPWR VPWR _6622_/Q sky130_fd_sc_hd__dfrtp_2
X_3834_ hold59/A _3845_/A _3827_/Y _3833_/X VGND VGND VPWR VPWR _3834_/X sky130_fd_sc_hd__a22o_1
XFILLER_32_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6553_ _6950_/CLK _6553_/D fanout875/X VGND VGND VPWR VPWR _6553_/Q sky130_fd_sc_hd__dfrtp_2
X_3765_ input4/X _3283_/Y _5441_/A _7013_/Q VGND VGND VPWR VPWR _3765_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6484_ _6668_/CLK _6484_/D _6439_/X VGND VGND VPWR VPWR _6484_/Q sky130_fd_sc_hd__dfrtp_1
X_5504_ _5504_/A _5576_/B VGND VGND VPWR VPWR _5512_/S sky130_fd_sc_hd__nand2_8
X_3696_ input21/X _3302_/Y _5441_/A _7014_/Q _3695_/X VGND VGND VPWR VPWR _3699_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_133_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5435_ wire780/X hold610/X _5440_/S VGND VGND VPWR VPWR _5435_/X sky130_fd_sc_hd__mux2_1
Xoutput310 _3952_/X VGND VGND VPWR VPWR serial_load sky130_fd_sc_hd__buf_8
Xoutput332 _6561_/Q VGND VGND VPWR VPWR wb_dat_o[22] sky130_fd_sc_hd__buf_8
Xoutput321 _6572_/Q VGND VGND VPWR VPWR wb_dat_o[12] sky130_fd_sc_hd__buf_8
Xoutput343 _6584_/Q VGND VGND VPWR VPWR wb_dat_o[3] sky130_fd_sc_hd__buf_8
XFILLER_120_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_662 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5366_ _5519_/A0 hold840/X _5368_/S VGND VGND VPWR VPWR _6946_/D sky130_fd_sc_hd__mux2_1
X_5297_ _5297_/A _5585_/B VGND VGND VPWR VPWR _5297_/Y sky130_fd_sc_hd__nand2_8
X_7105_ _7105_/CLK _7105_/D fanout862/X VGND VGND VPWR VPWR _7105_/Q sky130_fd_sc_hd__dfrtp_2
X_4317_ hold759/X _6407_/A0 _4321_/S VGND VGND VPWR VPWR _6763_/D sky130_fd_sc_hd__mux2_1
X_4248_ _5601_/A0 hold232/X hold32/X VGND VGND VPWR VPWR _4248_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7036_ _7036_/CLK _7036_/D fanout863/X VGND VGND VPWR VPWR _7036_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_83_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4179_ hold776/X _5234_/C _4183_/S VGND VGND VPWR VPWR _6644_/D sky130_fd_sc_hd__mux2_1
XFILLER_15_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire404 _3356_/Y VGND VGND VPWR VPWR _5351_/A sky130_fd_sc_hd__buf_8
XFILLER_11_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire437 _3305_/Y VGND VGND VPWR VPWR _5378_/A sky130_fd_sc_hd__buf_8
Xwire448 hold88/X VGND VGND VPWR VPWR hold89/A sky130_fd_sc_hd__buf_8
XFILLER_109_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire459 _3940_/X VGND VGND VPWR VPWR wire459/X sky130_fd_sc_hd__buf_6
XFILLER_152_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_41_csclk _6987_/CLK VGND VGND VPWR VPWR _6931_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_56_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7091_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_128_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3550_ _3549_/X _6794_/Q _3928_/A VGND VGND VPWR VPWR _6794_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3481_ _3534_/A _3543_/A VGND VGND VPWR VPWR _4082_/A sky130_fd_sc_hd__nor2_8
X_5220_ hold361/X _5578_/A0 _5222_/S VGND VGND VPWR VPWR _6821_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5151_ _5151_/A _5151_/B _5150_/X VGND VGND VPWR VPWR _5155_/B sky130_fd_sc_hd__or3b_1
X_5082_ _4581_/B _4987_/X _4950_/A _4411_/Y _4846_/X VGND VGND VPWR VPWR _5117_/A
+ sky130_fd_sc_hd__a2111o_4
XFILLER_111_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4102_ _4303_/A0 hold402/X _4102_/S VGND VGND VPWR VPWR _6580_/D sky130_fd_sc_hd__mux2_1
XFILLER_69_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4033_ _5602_/A0 hold298/X _4033_/S VGND VGND VPWR VPWR _4033_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5984_ _7188_/Q _6309_/S _5982_/X _5983_/X VGND VGND VPWR VPWR _7188_/D sky130_fd_sc_hd__o22a_1
XFILLER_24_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_7_0_csclk clkbuf_3_7_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_7_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
X_4935_ _4802_/A _5102_/D _4935_/C _4935_/D VGND VGND VPWR VPWR _4941_/C sky130_fd_sc_hd__nand4b_1
X_4866_ _5013_/A _4922_/A _5086_/A _4866_/D VGND VGND VPWR VPWR _4866_/X sky130_fd_sc_hd__or4_2
XANTENNA_22 _6808_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_11 _6484_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4797_ _5116_/A _4797_/B _4797_/C _4797_/D VGND VGND VPWR VPWR _4798_/D sky130_fd_sc_hd__or4_1
X_6605_ _6608_/CLK _6605_/D fanout858/X VGND VGND VPWR VPWR _6605_/Q sky130_fd_sc_hd__dfrtp_2
X_3817_ _3840_/S _3817_/B VGND VGND VPWR VPWR _3817_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_33 _7174_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_55 _3665_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_44 _3504_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_66 _3687_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3748_ _6609_/Q _4136_/A _4142_/A _6614_/Q VGND VGND VPWR VPWR _3748_/X sky130_fd_sc_hd__a22o_1
XANTENNA_88 _5056_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_99 _5927_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6536_ _6806_/CLK _6536_/D _6435_/A VGND VGND VPWR VPWR _6536_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_77 _4235_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3679_ _7118_/Q wire446/A _4160_/A _6630_/Q VGND VGND VPWR VPWR _3679_/X sky130_fd_sc_hd__a22o_1
X_6467_ _6668_/CLK _6467_/D _6422_/X VGND VGND VPWR VPWR _6467_/Q sky130_fd_sc_hd__dfrtp_2
X_6398_ _4236_/C _6398_/A2 _6398_/B1 _4236_/A VGND VGND VPWR VPWR _6398_/X sky130_fd_sc_hd__a22o_1
X_5418_ wire770/X hold422/X _5422_/S VGND VGND VPWR VPWR _6992_/D sky130_fd_sc_hd__mux2_1
Xoutput195 _3212_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[28] sky130_fd_sc_hd__buf_8
Xoutput184 _3222_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[18] sky130_fd_sc_hd__buf_8
X_5349_ _5601_/A0 hold346/X _5350_/S VGND VGND VPWR VPWR _6931_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput173 _3972_/X VGND VGND VPWR VPWR irq[1] sky130_fd_sc_hd__buf_8
XFILLER_87_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7019_ _7139_/CLK _7019_/D fanout865/X VGND VGND VPWR VPWR _7019_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4720_ _4706_/X _4713_/X _4917_/B VGND VGND VPWR VPWR _4720_/X sky130_fd_sc_hd__o21a_2
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4651_ _4728_/A _4651_/B VGND VGND VPWR VPWR _4652_/B sky130_fd_sc_hd__nor2_8
XFILLER_147_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3602_ _3204_/A _3346_/Y _4118_/A _6597_/Q VGND VGND VPWR VPWR _3602_/X sky130_fd_sc_hd__a22o_4
Xinput31 mask_rev_in[5] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__clkbuf_4
Xinput20 mask_rev_in[24] VGND VGND VPWR VPWR input20/X sky130_fd_sc_hd__clkbuf_4
Xinput42 mgmt_gpio_in[15] VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__clkbuf_4
Xinput53 mgmt_gpio_in[25] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__clkbuf_4
Xinput64 mgmt_gpio_in[35] VGND VGND VPWR VPWR input64/X sky130_fd_sc_hd__clkbuf_4
X_4582_ _4988_/A _4749_/C VGND VGND VPWR VPWR _5174_/A sky130_fd_sc_hd__nor2_1
Xinput97 usr2_vcc_pwrgood VGND VGND VPWR VPWR wire834/A sky130_fd_sc_hd__buf_6
Xinput86 spimemio_flash_io0_oeb VGND VGND VPWR VPWR wire841/A sky130_fd_sc_hd__buf_6
XFILLER_155_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3533_ _3533_/A _3533_/B _3533_/C VGND VGND VPWR VPWR _3547_/C sky130_fd_sc_hd__or3_1
Xwire790 wire790/A VGND VGND VPWR VPWR wire790/X sky130_fd_sc_hd__buf_8
Xhold815 _7106_/Q VGND VGND VPWR VPWR hold815/X sky130_fd_sc_hd__bufbuf_16
Xhold826 _5267_/X VGND VGND VPWR VPWR _6858_/D sky130_fd_sc_hd__bufbuf_16
Xhold804 _6824_/Q VGND VGND VPWR VPWR hold804/X sky130_fd_sc_hd__bufbuf_16
Xinput75 porb VGND VGND VPWR VPWR input75/X sky130_fd_sc_hd__clkbuf_4
Xhold837 _5519_/X VGND VGND VPWR VPWR _7082_/D sky130_fd_sc_hd__bufbuf_16
X_6321_ _6321_/A _6321_/B _6321_/C _6321_/D VGND VGND VPWR VPWR _6321_/X sky130_fd_sc_hd__or4_1
Xhold848 _7121_/Q VGND VGND VPWR VPWR hold848/X sky130_fd_sc_hd__bufbuf_16
XFILLER_143_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6252_ _6758_/Q _6337_/A2 _6252_/B1 _6753_/Q _6251_/X VGND VGND VPWR VPWR _6257_/C
+ sky130_fd_sc_hd__a221o_1
X_3464_ _3508_/A _3528_/B VGND VGND VPWR VPWR _4190_/A sky130_fd_sc_hd__nor2_8
XFILLER_131_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5203_ _6409_/A0 hold824/X _5206_/S VGND VGND VPWR VPWR _6807_/D sky130_fd_sc_hd__mux2_1
X_6183_ wire556/X _6060_/B _6170_/X _6182_/X _3197_/Y VGND VGND VPWR VPWR _6183_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_130_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3395_ wire553/X _3395_/A2 _5468_/A _7043_/Q _3394_/X VGND VGND VPWR VPWR _3398_/B
+ sky130_fd_sc_hd__a221o_1
X_5134_ _5077_/Y _5120_/X _5133_/Y _5112_/X VGND VGND VPWR VPWR _6782_/D sky130_fd_sc_hd__a211o_1
XFILLER_97_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5065_ _5065_/A _5130_/B VGND VGND VPWR VPWR _5124_/B sky130_fd_sc_hd__nor2_8
X_4016_ hold797/X _4015_/X _4024_/S VGND VGND VPWR VPWR _6509_/D sky130_fd_sc_hd__mux2_1
XFILLER_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5967_ _6567_/Q wire673/X wire653/X _6653_/Q VGND VGND VPWR VPWR _5967_/X sky130_fd_sc_hd__a22o_1
X_4918_ _5069_/B _5132_/A VGND VGND VPWR VPWR _5102_/D sky130_fd_sc_hd__nor2_4
XFILLER_193_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5898_ wire570/X wire657/X wire651/X _6759_/Q VGND VGND VPWR VPWR _5898_/X sky130_fd_sc_hd__a22o_1
XFILLER_32_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4849_ _4849_/A _5071_/A VGND VGND VPWR VPWR _5081_/B sky130_fd_sc_hd__or2_1
XFILLER_180_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6519_ _7147_/CLK _6519_/D fanout886/X VGND VGND VPWR VPWR _6519_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_146_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6870_ _7128_/CLK _6870_/D _6421_/A VGND VGND VPWR VPWR _6870_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_34_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5821_ _6962_/Q _5673_/X _5681_/X _6922_/Q _5820_/X VGND VGND VPWR VPWR _5826_/B
+ sky130_fd_sc_hd__a221o_4
XFILLER_34_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5752_ _6863_/Q wire667/X wire656/X wire530/X _5751_/X VGND VGND VPWR VPWR _5753_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_188_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4703_ _4773_/A _4930_/C _4773_/B VGND VGND VPWR VPWR _4772_/C sky130_fd_sc_hd__and3b_2
XFILLER_187_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5683_ _7165_/Q _5705_/B _5707_/C VGND VGND VPWR VPWR _5683_/X sky130_fd_sc_hd__and3_4
XFILLER_147_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4634_ _4845_/A _4634_/B VGND VGND VPWR VPWR _5144_/A sky130_fd_sc_hd__nand2_1
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4565_ _4566_/A _4740_/B VGND VGND VPWR VPWR _4565_/Y sky130_fd_sc_hd__nor2_8
Xhold601 _7048_/Q VGND VGND VPWR VPWR hold601/X sky130_fd_sc_hd__bufbuf_16
Xhold612 _6684_/Q VGND VGND VPWR VPWR hold612/X sky130_fd_sc_hd__bufbuf_16
XFILLER_190_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold623 _7000_/Q VGND VGND VPWR VPWR hold623/X sky130_fd_sc_hd__bufbuf_16
X_6304_ _6715_/Q wire640/X wire638/X _6547_/Q _6303_/X VGND VGND VPWR VPWR _6305_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3516_ _6772_/Q _4322_/A _5194_/A _6804_/Q VGND VGND VPWR VPWR _3516_/X sky130_fd_sc_hd__a22o_4
Xhold634 _6804_/Q VGND VGND VPWR VPWR hold634/X sky130_fd_sc_hd__bufbuf_16
Xhold645 _5258_/X VGND VGND VPWR VPWR _6850_/D sky130_fd_sc_hd__bufbuf_16
X_4496_ _4819_/B _4724_/A VGND VGND VPWR VPWR _4745_/B sky130_fd_sc_hd__or2_4
XFILLER_143_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold667 _7052_/Q VGND VGND VPWR VPWR hold667/X sky130_fd_sc_hd__bufbuf_16
Xhold656 _6761_/Q VGND VGND VPWR VPWR hold656/X sky130_fd_sc_hd__bufbuf_16
Xhold678 _6788_/Q VGND VGND VPWR VPWR hold678/X sky130_fd_sc_hd__bufbuf_16
XFILLER_134_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold689 _7092_/Q VGND VGND VPWR VPWR hold689/X sky130_fd_sc_hd__bufbuf_16
X_3447_ _7018_/Q _5441_/A _3369_/Y wire527/X _3446_/X VGND VGND VPWR VPWR _3450_/C
+ sky130_fd_sc_hd__a221o_1
X_6235_ _7196_/Q _5665_/Y _6233_/X _6234_/X VGND VGND VPWR VPWR _7196_/D sky130_fd_sc_hd__o22a_1
X_3378_ _3378_/A _3378_/B _3378_/C _3378_/D VGND VGND VPWR VPWR _3379_/C sky130_fd_sc_hd__or4_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6166_ _7002_/Q _5987_/Y _6191_/B1 _6922_/Q VGND VGND VPWR VPWR _6166_/X sky130_fd_sc_hd__a22o_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6097_ _7111_/Q wire650/X _6295_/B1 _7151_/Q VGND VGND VPWR VPWR _6097_/X sky130_fd_sc_hd__a22o_1
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5117_ _5117_/A _5117_/B VGND VGND VPWR VPWR _5120_/C sky130_fd_sc_hd__or2_2
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5048_ _5048_/A _5151_/B VGND VGND VPWR VPWR _5056_/A sky130_fd_sc_hd__or2_1
XFILLER_84_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6999_ _7129_/CLK _6999_/D fanout863/X VGND VGND VPWR VPWR _6999_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_159_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4350_ _4350_/A _4350_/B _4350_/C _4350_/D VGND VGND VPWR VPWR _4352_/B sky130_fd_sc_hd__and4_1
XFILLER_172_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3301_ _3505_/A hold63/X VGND VGND VPWR VPWR _3301_/Y sky130_fd_sc_hd__nor2_8
XFILLER_152_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4281_ _5487_/A0 hold806/X _4285_/S VGND VGND VPWR VPWR _6733_/D sky130_fd_sc_hd__mux2_1
XFILLER_140_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6020_ _6020_/A _6020_/B _6020_/C _6020_/D VGND VGND VPWR VPWR _6024_/A sky130_fd_sc_hd__or4_1
XFILLER_113_579 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3232_ _6920_/Q VGND VGND VPWR VPWR _3232_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6922_ _6979_/CLK _6922_/D fanout878/X VGND VGND VPWR VPWR _6922_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_82_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6853_ _6996_/CLK _6853_/D fanout869/X VGND VGND VPWR VPWR _6853_/Q sky130_fd_sc_hd__dfstp_1
X_5804_ _7065_/Q _5921_/A2 _5687_/X wire505/X VGND VGND VPWR VPWR _5804_/X sky130_fd_sc_hd__a22o_1
XFILLER_90_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6784_ _7210_/CLK _6784_/D wire915/A VGND VGND VPWR VPWR _6784_/Q sky130_fd_sc_hd__dfrtp_2
X_3996_ _6496_/Q _6407_/A0 _4003_/S VGND VGND VPWR VPWR _6496_/D sky130_fd_sc_hd__mux2_1
X_5735_ _6910_/Q wire699/X wire666/X _6862_/Q _5726_/X VGND VGND VPWR VPWR _5735_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5666_ _7161_/Q _7162_/Q VGND VGND VPWR VPWR _5704_/B sky130_fd_sc_hd__and2b_4
Xmax_length409 _3352_/Y VGND VGND VPWR VPWR _3582_/B1 sky130_fd_sc_hd__buf_6
X_4617_ _4617_/A _4617_/B VGND VGND VPWR VPWR _4617_/Y sky130_fd_sc_hd__nor2_2
X_5597_ _5597_/A0 hold247/X hold66/X VGND VGND VPWR VPWR _5597_/X sky130_fd_sc_hd__mux2_1
Xhold420 _7123_/Q VGND VGND VPWR VPWR hold420/X sky130_fd_sc_hd__bufbuf_16
XFILLER_190_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold442 _6894_/Q VGND VGND VPWR VPWR hold442/X sky130_fd_sc_hd__bufbuf_16
Xhold453 _6962_/Q VGND VGND VPWR VPWR hold453/X sky130_fd_sc_hd__bufbuf_16
Xhold431 _4138_/X VGND VGND VPWR VPWR _6610_/D sky130_fd_sc_hd__bufbuf_16
X_4548_ _5081_/A _4849_/A _4548_/C _4548_/D VGND VGND VPWR VPWR _4548_/X sky130_fd_sc_hd__or4_1
XFILLER_116_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold475 _6914_/Q VGND VGND VPWR VPWR hold475/X sky130_fd_sc_hd__bufbuf_16
Xhold464 hold513/X VGND VGND VPWR VPWR hold514/A sky130_fd_sc_hd__bufbuf_16
XFILLER_131_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4479_ _4775_/A _4636_/A VGND VGND VPWR VPWR _4766_/A sky130_fd_sc_hd__nor2_2
XFILLER_104_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold486 _6736_/Q VGND VGND VPWR VPWR hold486/X sky130_fd_sc_hd__bufbuf_16
XFILLER_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6218_ _6988_/Q _6028_/X _6034_/Y _6996_/Q _6217_/X VGND VGND VPWR VPWR _6219_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_58_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold497 _6635_/Q VGND VGND VPWR VPWR hold497/X sky130_fd_sc_hd__bufbuf_16
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7198_ _7220_/CLK _7198_/D fanout854/X VGND VGND VPWR VPWR _7198_/Q sky130_fd_sc_hd__dfrtp_1
X_6149_ wire539/X wire600/X wire646/X _6937_/Q _6148_/X VGND VGND VPWR VPWR _6156_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_304 _7122_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_315 wire632/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_326 _5598_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_348 _4303_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_337 hold555/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3850_ _6470_/Q _3797_/X _6472_/Q VGND VGND VPWR VPWR _3850_/Y sky130_fd_sc_hd__a21oi_1
X_3781_ input20/X _3302_/Y _3320_/Y input34/X VGND VGND VPWR VPWR _3781_/X sky130_fd_sc_hd__a22o_2
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5520_ wire746/X hold737/X _5521_/S VGND VGND VPWR VPWR _7083_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5451_ wire802/X _7021_/Q _5458_/S VGND VGND VPWR VPWR _7021_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4402_ _4553_/B _4410_/C _4513_/A VGND VGND VPWR VPWR _4402_/X sky130_fd_sc_hd__or3_2
X_5382_ wire773/A hold329/X _5386_/S VGND VGND VPWR VPWR _5382_/X sky130_fd_sc_hd__mux2_1
X_7121_ _7133_/CLK _7121_/D fanout883/X VGND VGND VPWR VPWR _7121_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_160_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4333_ _6411_/A0 hold614/X _4333_/S VGND VGND VPWR VPWR _6777_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7052_ _7140_/CLK _7052_/D fanout865/X VGND VGND VPWR VPWR _7052_/Q sky130_fd_sc_hd__dfrtp_2
X_4264_ hold764/X _6408_/A0 _4267_/S VGND VGND VPWR VPWR _4264_/X sky130_fd_sc_hd__mux2_1
X_3215_ _7056_/Q VGND VGND VPWR VPWR _3215_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6003_ _6037_/B _6033_/C _6018_/A VGND VGND VPWR VPWR _6021_/C sky130_fd_sc_hd__and3_4
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4195_ _6411_/A0 hold597/X _4195_/S VGND VGND VPWR VPWR _4195_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6905_ _6951_/CLK _6905_/D _6421_/A VGND VGND VPWR VPWR _6905_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_82_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6836_ _6980_/CLK _6836_/D fanout878/X VGND VGND VPWR VPWR _6836_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_24_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6767_ _7223_/CLK _6767_/D fanout850/X VGND VGND VPWR VPWR _6767_/Q sky130_fd_sc_hd__dfrtp_2
X_3979_ wire903/X hold512/X _3993_/S VGND VGND VPWR VPWR _3979_/X sky130_fd_sc_hd__mux2_8
X_5718_ wire509/X _5803_/B1 wire670/X _6925_/Q _5717_/X VGND VGND VPWR VPWR _5720_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_10_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6698_ _7220_/CLK _6698_/D _6362_/B VGND VGND VPWR VPWR _6698_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_156_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5649_ _7170_/Q _5654_/A VGND VGND VPWR VPWR _5649_/Y sky130_fd_sc_hd__nor2_1
XFILLER_151_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold261 _7218_/Q VGND VGND VPWR VPWR hold261/X sky130_fd_sc_hd__bufbuf_16
XFILLER_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold250 _6907_/Q VGND VGND VPWR VPWR hold250/X sky130_fd_sc_hd__bufbuf_16
XFILLER_104_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold294 _7060_/Q VGND VGND VPWR VPWR hold294/X sky130_fd_sc_hd__bufbuf_16
Xhold283 _7004_/Q VGND VGND VPWR VPWR hold283/X sky130_fd_sc_hd__bufbuf_16
Xhold272 _6969_/Q VGND VGND VPWR VPWR hold272/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout741 hold263/X VGND VGND VPWR VPWR hold264/A sky130_fd_sc_hd__buf_6
Xfanout774 hold81/X VGND VGND VPWR VPWR hold82/A sky130_fd_sc_hd__buf_8
Xfanout785 hold11/X VGND VGND VPWR VPWR hold12/A sky130_fd_sc_hd__buf_8
XFILLER_93_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_101 _6029_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_134 _6508_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_112 debug_oeb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_123 _6457_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_167 wb_sel_i[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_156 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_145 pad_flash_io0_di VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_178 _6393_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_189 _5741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_1_1_1_csclk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_182_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length762 hold156/X VGND VGND VPWR VPWR _5572_/A0 sky130_fd_sc_hd__buf_8
Xmax_length784 _5597_/A0 VGND VGND VPWR VPWR _5336_/A1 sky130_fd_sc_hd__buf_8
XFILLER_123_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput7 mask_rev_in[12] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_4
XFILLER_64_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4951_ _4949_/B _4536_/B _4959_/A _4903_/A VGND VGND VPWR VPWR _5148_/A sky130_fd_sc_hd__a31o_1
XFILLER_17_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4882_ _4736_/B _4692_/C _4657_/B _4581_/B _4581_/A VGND VGND VPWR VPWR _4903_/C
+ sky130_fd_sc_hd__a32o_2
X_3902_ _7166_/Q _7167_/Q VGND VGND VPWR VPWR _6012_/A sky130_fd_sc_hd__and2b_4
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6621_ _6621_/CLK _6621_/D fanout872/X VGND VGND VPWR VPWR _6621_/Q sky130_fd_sc_hd__dfstp_4
X_3833_ hold59/A _6477_/Q hold40/A VGND VGND VPWR VPWR _3833_/X sky130_fd_sc_hd__a21o_1
X_6552_ _6950_/CLK _6552_/D fanout874/X VGND VGND VPWR VPWR _6552_/Q sky130_fd_sc_hd__dfstp_2
X_3764_ _3764_/A _3764_/B _3764_/C _3764_/D VGND VGND VPWR VPWR _3764_/X sky130_fd_sc_hd__or4_4
XFILLER_185_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5503_ wire742/X hold370/X _5503_/S VGND VGND VPWR VPWR _7068_/D sky130_fd_sc_hd__mux2_1
X_3695_ _7070_/Q _5504_/A _4292_/A _6744_/Q VGND VGND VPWR VPWR _3695_/X sky130_fd_sc_hd__a22o_1
X_6483_ _6668_/CLK _6483_/D _6438_/X VGND VGND VPWR VPWR _6483_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_10_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5434_ _5578_/A0 _7006_/Q _5440_/S VGND VGND VPWR VPWR _7006_/D sky130_fd_sc_hd__mux2_1
Xoutput300 _6489_/Q VGND VGND VPWR VPWR pll_trim[9] sky130_fd_sc_hd__buf_8
XFILLER_133_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput333 _6562_/Q VGND VGND VPWR VPWR wb_dat_o[23] sky130_fd_sc_hd__buf_8
XFILLER_126_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput322 _6573_/Q VGND VGND VPWR VPWR wb_dat_o[13] sky130_fd_sc_hd__buf_8
Xoutput344 _6585_/Q VGND VGND VPWR VPWR wb_dat_o[4] sky130_fd_sc_hd__buf_8
Xoutput311 _3951_/X VGND VGND VPWR VPWR serial_resetn sky130_fd_sc_hd__buf_8
Xclkbuf_3_3_0_csclk clkbuf_3_3_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_3_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
X_5365_ _5572_/A0 hold477/X _5365_/S VGND VGND VPWR VPWR _6945_/D sky130_fd_sc_hd__mux2_1
X_7104_ _7140_/CLK _7104_/D fanout865/X VGND VGND VPWR VPWR _7104_/Q sky130_fd_sc_hd__dfrtp_2
X_5296_ _5602_/A0 hold356/X _5296_/S VGND VGND VPWR VPWR _6884_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4316_ _4316_/A _6406_/B VGND VGND VPWR VPWR _4321_/S sky130_fd_sc_hd__and2_4
X_4247_ hold3/X hold847/X hold32/X VGND VGND VPWR VPWR hold4/A sky130_fd_sc_hd__mux2_1
X_7035_ _7042_/CLK _7035_/D fanout865/X VGND VGND VPWR VPWR _7035_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4178_ _4178_/A _5242_/B VGND VGND VPWR VPWR _4183_/S sky130_fd_sc_hd__and2_4
XFILLER_67_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_23_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6819_ _7103_/CLK _6819_/D fanout861/X VGND VGND VPWR VPWR _6819_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_11_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire427 wire427/A VGND VGND VPWR VPWR _4025_/A sky130_fd_sc_hd__buf_8
XFILLER_109_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire438 wire438/A VGND VGND VPWR VPWR wire438/X sky130_fd_sc_hd__buf_8
XFILLER_11_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3480_ _3543_/A _5252_/B VGND VGND VPWR VPWR _4118_/A sky130_fd_sc_hd__nor2_8
XFILLER_170_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5150_ _4947_/B _4832_/B _5050_/C _4832_/A _4835_/X VGND VGND VPWR VPWR _5150_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5081_ _5081_/A _5081_/B _5081_/C _4623_/A VGND VGND VPWR VPWR _5115_/A sky130_fd_sc_hd__or4b_4
X_4101_ hold83/X _6579_/Q _4102_/S VGND VGND VPWR VPWR _4101_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4032_ _5601_/A0 hold225/X _4033_/S VGND VGND VPWR VPWR _4032_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5983_ wire824/X _7187_/Q wire381/X VGND VGND VPWR VPWR _5983_/X sky130_fd_sc_hd__a21o_1
XFILLER_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4934_ _4398_/Y _5023_/B _5062_/C _4933_/Y VGND VGND VPWR VPWR _4935_/C sky130_fd_sc_hd__o22a_2
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4865_ _5118_/B _4865_/B _4865_/C VGND VGND VPWR VPWR _4866_/D sky130_fd_sc_hd__or3_1
XANTENNA_12 _6486_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 _6823_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4796_ _5140_/B _4796_/B _4796_/C _4796_/D VGND VGND VPWR VPWR _4797_/D sky130_fd_sc_hd__or4_1
X_6604_ _6950_/CLK _6604_/D fanout874/X VGND VGND VPWR VPWR _6604_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_45 _3516_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_34 _7187_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3816_ _3255_/X _3256_/Y _3820_/B VGND VGND VPWR VPWR _3817_/B sky130_fd_sc_hd__mux2_1
XANTENNA_56 _3654_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3747_ _6861_/Q wire439/X _5306_/A _6893_/Q _3746_/X VGND VGND VPWR VPWR _3754_/A
+ sky130_fd_sc_hd__a221o_2
XANTENNA_67 _3693_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6535_ _6806_/CLK _6535_/D _6435_/A VGND VGND VPWR VPWR _6535_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_89 _5234_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_78 _4235_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6466_ _3938_/A1 _6466_/D _6421_/X VGND VGND VPWR VPWR hold19/A sky130_fd_sc_hd__dfrtp_4
XFILLER_173_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3678_ _6831_/Q _5227_/A _4298_/A _6749_/Q VGND VGND VPWR VPWR _3678_/X sky130_fd_sc_hd__a22o_1
X_6397_ _6396_/X _7217_/Q _6400_/S VGND VGND VPWR VPWR _7217_/D sky130_fd_sc_hd__mux2_1
X_5417_ wire780/X hold653/X _5422_/S VGND VGND VPWR VPWR _6991_/D sky130_fd_sc_hd__mux2_1
Xoutput185 _3221_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[19] sky130_fd_sc_hd__buf_8
X_5348_ _5600_/A0 hold426/X _5350_/S VGND VGND VPWR VPWR _6930_/D sky130_fd_sc_hd__mux2_1
Xoutput174 _3973_/X VGND VGND VPWR VPWR irq[2] sky130_fd_sc_hd__buf_8
Xoutput196 _3211_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[29] sky130_fd_sc_hd__buf_8
XFILLER_101_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5279_ _5279_/A _5594_/B VGND VGND VPWR VPWR _5287_/S sky130_fd_sc_hd__nand2_8
XFILLER_87_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7018_ _7139_/CLK _7018_/D fanout868/X VGND VGND VPWR VPWR _7018_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_101_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4650_ _4722_/B _4650_/B VGND VGND VPWR VPWR _5062_/B sky130_fd_sc_hd__or2_4
XFILLER_175_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput10 mask_rev_in[15] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__clkbuf_4
X_3601_ _7024_/Q _3301_/Y _4328_/A _6776_/Q _3561_/X VGND VGND VPWR VPWR _3605_/C
+ sky130_fd_sc_hd__a221o_1
Xinput21 mask_rev_in[25] VGND VGND VPWR VPWR input21/X sky130_fd_sc_hd__clkbuf_4
X_4581_ _4581_/A _4581_/B VGND VGND VPWR VPWR _4612_/B sky130_fd_sc_hd__nand2_1
Xinput43 mgmt_gpio_in[16] VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__clkbuf_4
Xinput54 mgmt_gpio_in[26] VGND VGND VPWR VPWR input54/X sky130_fd_sc_hd__clkbuf_4
XFILLER_128_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6320_ _6627_/Q _6028_/X _6342_/B1 _6726_/Q _6319_/X VGND VGND VPWR VPWR _6321_/D
+ sky130_fd_sc_hd__a221o_2
Xinput32 mask_rev_in[6] VGND VGND VPWR VPWR input32/X sky130_fd_sc_hd__clkbuf_4
Xinput98 usr2_vdd_pwrgood VGND VGND VPWR VPWR wire833/A sky130_fd_sc_hd__buf_6
Xinput87 spimemio_flash_io1_do VGND VGND VPWR VPWR wire840/A sky130_fd_sc_hd__buf_6
XFILLER_155_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput65 mgmt_gpio_in[36] VGND VGND VPWR VPWR _7228_/A sky130_fd_sc_hd__buf_6
X_3532_ wire484/X _5531_/A _4097_/A _6580_/Q _3530_/X VGND VGND VPWR VPWR _3533_/C
+ sky130_fd_sc_hd__a221o_1
Xwire780 wire780/A VGND VGND VPWR VPWR wire780/X sky130_fd_sc_hd__buf_8
Xhold805 _5224_/X VGND VGND VPWR VPWR _6824_/D sky130_fd_sc_hd__bufbuf_16
Xhold827 _7138_/Q VGND VGND VPWR VPWR hold827/X sky130_fd_sc_hd__bufbuf_16
Xhold816 _7090_/Q VGND VGND VPWR VPWR hold816/X sky130_fd_sc_hd__bufbuf_16
Xinput76 qspi_enabled VGND VGND VPWR VPWR wire845/A sky130_fd_sc_hd__buf_6
Xhold849 _7147_/Q VGND VGND VPWR VPWR hold849/X sky130_fd_sc_hd__bufbuf_16
X_6251_ _6619_/Q wire623/X wire611/X _6738_/Q VGND VGND VPWR VPWR _6251_/X sky130_fd_sc_hd__a22o_1
X_3463_ wire539/X _3338_/Y _4256_/A _6717_/Q _3461_/X VGND VGND VPWR VPWR _3472_/B
+ sky130_fd_sc_hd__a221o_1
Xhold838 _6596_/Q VGND VGND VPWR VPWR hold838/X sky130_fd_sc_hd__bufbuf_16
XFILLER_170_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6182_ _6306_/A _6182_/B _6182_/C VGND VGND VPWR VPWR _6182_/X sky130_fd_sc_hd__or3_4
XFILLER_115_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5202_ _6408_/A0 _6806_/Q _5206_/S VGND VGND VPWR VPWR _6806_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3394_ _7059_/Q wire438/X wire450/X wire521/X VGND VGND VPWR VPWR _3394_/X sky130_fd_sc_hd__a22o_1
X_5133_ _5133_/A _5133_/B VGND VGND VPWR VPWR _5133_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5064_ _4949_/C _4748_/A _4657_/B _4903_/C _4846_/B VGND VGND VPWR VPWR _5130_/B
+ sky130_fd_sc_hd__a311o_4
XFILLER_97_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4015_ hold562/X _5598_/A0 _4021_/S VGND VGND VPWR VPWR _4015_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5966_ _6613_/Q wire657/X wire651/X _6762_/Q VGND VGND VPWR VPWR _5981_/B sky130_fd_sc_hd__a22o_1
XFILLER_12_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4917_ _4917_/A _4917_/B _5003_/C VGND VGND VPWR VPWR _5102_/C sky130_fd_sc_hd__and3_4
X_5897_ _6645_/Q wire690/X _5964_/B1 _6600_/Q VGND VGND VPWR VPWR _5897_/X sky130_fd_sc_hd__a22o_1
XFILLER_178_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4848_ _4845_/A _4634_/B _4920_/A VGND VGND VPWR VPWR _5136_/C sky130_fd_sc_hd__a21o_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4779_ _4724_/B _4757_/B _5081_/A VGND VGND VPWR VPWR _4799_/A sky130_fd_sc_hd__o21bai_1
X_6518_ _7152_/CLK _6518_/D fanout886/X VGND VGND VPWR VPWR _6518_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_180_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6449_ _6455_/A _6455_/B VGND VGND VPWR VPWR _6449_/X sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_40_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _6930_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_122_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_0_0_csclk clkbuf_2_1_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_1_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_102_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_55_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _6992_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_56_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5820_ _6970_/Q _5691_/X wire665/X _6954_/Q VGND VGND VPWR VPWR _5820_/X sky130_fd_sc_hd__a22o_1
X_5751_ _7031_/Q wire686/X wire675/X _7079_/Q VGND VGND VPWR VPWR _5751_/X sky130_fd_sc_hd__a22o_2
XFILLER_62_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4702_ _4702_/A _4702_/B VGND VGND VPWR VPWR _4773_/B sky130_fd_sc_hd__or2_1
XFILLER_147_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5682_ _7165_/Q _5702_/B _5707_/C VGND VGND VPWR VPWR _5682_/X sky130_fd_sc_hd__and3_4
XFILLER_175_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4633_ _4986_/A _4996_/A VGND VGND VPWR VPWR _4633_/X sky130_fd_sc_hd__or2_2
X_4564_ _4564_/A _4672_/A VGND VGND VPWR VPWR _4740_/B sky130_fd_sc_hd__nand2_8
Xhold602 _6976_/Q VGND VGND VPWR VPWR hold602/X sky130_fd_sc_hd__bufbuf_16
XFILLER_118_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold624 _7096_/Q VGND VGND VPWR VPWR hold624/X sky130_fd_sc_hd__bufbuf_16
X_6303_ wire568/X wire647/X wire632/X _6591_/Q VGND VGND VPWR VPWR _6303_/X sky130_fd_sc_hd__a22o_1
XFILLER_128_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3515_ _5234_/A hold87/X VGND VGND VPWR VPWR _5194_/A sky130_fd_sc_hd__nor2_8
Xhold635 _6767_/Q VGND VGND VPWR VPWR hold635/X sky130_fd_sc_hd__bufbuf_16
Xhold613 _4227_/X VGND VGND VPWR VPWR _6684_/D sky130_fd_sc_hd__bufbuf_16
X_4495_ _4651_/B _4707_/B _5050_/A VGND VGND VPWR VPWR _4724_/A sky130_fd_sc_hd__or3b_4
Xhold668 _6546_/Q VGND VGND VPWR VPWR hold668/X sky130_fd_sc_hd__bufbuf_16
Xhold657 _7012_/Q VGND VGND VPWR VPWR hold657/X sky130_fd_sc_hd__bufbuf_16
Xhold646 _6492_/Q VGND VGND VPWR VPWR hold646/X sky130_fd_sc_hd__bufbuf_16
X_6234_ _5611_/A _7195_/Q _5664_/X VGND VGND VPWR VPWR _6234_/X sky130_fd_sc_hd__a21o_1
Xhold679 _6663_/Q VGND VGND VPWR VPWR hold679/X sky130_fd_sc_hd__bufbuf_16
X_3446_ wire535/X _3306_/Y _5200_/A _6810_/Q VGND VGND VPWR VPWR _3446_/X sky130_fd_sc_hd__a22o_1
X_3377_ _3377_/A _3377_/B _3377_/C _3377_/D VGND VGND VPWR VPWR _3378_/D sky130_fd_sc_hd__or4_2
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ _7018_/Q wire575/X _6037_/X _7042_/Q _6162_/X VGND VGND VPWR VPWR _6170_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5116_ _5116_/A _5116_/B _5116_/C _4881_/A VGND VGND VPWR VPWR _5117_/B sky130_fd_sc_hd__or4b_4
X_6096_ _7079_/Q _6211_/B _6091_/X _6093_/X _6095_/X VGND VGND VPWR VPWR _6096_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_57_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5047_ _5047_/A _5047_/B _5047_/C _5047_/D VGND VGND VPWR VPWR _5151_/B sky130_fd_sc_hd__or4_2
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6998_ _7140_/CLK _6998_/D fanout862/X VGND VGND VPWR VPWR _6998_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_41_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5949_ _6548_/Q wire706/X wire686/X _6771_/Q VGND VGND VPWR VPWR _5949_/X sky130_fd_sc_hd__a22o_1
XFILLER_53_586 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3300_ wire499/X wire438/X _5414_/A _6996_/Q VGND VGND VPWR VPWR _3300_/X sky130_fd_sc_hd__a22o_2
X_4280_ _4280_/A _5378_/B VGND VGND VPWR VPWR _4285_/S sky130_fd_sc_hd__nand2_8
XFILLER_125_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3231_ _6928_/Q VGND VGND VPWR VPWR _3231_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6921_ _6981_/CLK _6921_/D fanout878/X VGND VGND VPWR VPWR _6921_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_81_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6852_ _6992_/CLK _6852_/D fanout868/X VGND VGND VPWR VPWR _6852_/Q sky130_fd_sc_hd__dfrtp_1
X_5803_ wire480/X _5857_/A2 _5803_/B1 _7041_/Q _5802_/X VGND VGND VPWR VPWR _5806_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_90_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6783_ _7210_/CLK _6783_/D wire915/A VGND VGND VPWR VPWR _6783_/Q sky130_fd_sc_hd__dfrtp_2
X_3995_ _3995_/A _6406_/B VGND VGND VPWR VPWR _4003_/S sky130_fd_sc_hd__and2_4
XFILLER_148_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5734_ _5734_/A _5734_/B _5734_/C _5734_/D VGND VGND VPWR VPWR _5734_/X sky130_fd_sc_hd__or4_1
XFILLER_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5665_ _5665_/A _5665_/B VGND VGND VPWR VPWR _5665_/Y sky130_fd_sc_hd__nor2_8
XFILLER_148_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4616_ _4502_/A _4997_/A _5123_/C _4881_/A VGND VGND VPWR VPWR _4619_/C sky130_fd_sc_hd__o211a_1
Xhold410 _4212_/X VGND VGND VPWR VPWR _6673_/D sky130_fd_sc_hd__bufbuf_16
X_5596_ hold38/X _7150_/Q hold66/X VGND VGND VPWR VPWR hold67/A sky130_fd_sc_hd__mux2_1
XFILLER_151_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold432 _6898_/Q VGND VGND VPWR VPWR hold432/X sky130_fd_sc_hd__bufbuf_16
Xhold443 _6878_/Q VGND VGND VPWR VPWR hold443/X sky130_fd_sc_hd__bufbuf_16
X_4547_ _4986_/B _4988_/A VGND VGND VPWR VPWR _4548_/D sky130_fd_sc_hd__nor2_1
XFILLER_116_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold454 _6727_/Q VGND VGND VPWR VPWR hold454/X sky130_fd_sc_hd__bufbuf_16
Xhold421 _5565_/X VGND VGND VPWR VPWR _7123_/D sky130_fd_sc_hd__bufbuf_16
Xhold465 hold465/A VGND VGND VPWR VPWR hold465/X sky130_fd_sc_hd__bufbuf_16
X_4478_ _4707_/B _4478_/B _4478_/C VGND VGND VPWR VPWR _4844_/B sky130_fd_sc_hd__or3_4
XFILLER_143_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold487 _6726_/Q VGND VGND VPWR VPWR hold487/X sky130_fd_sc_hd__bufbuf_16
Xhold476 _6489_/Q VGND VGND VPWR VPWR hold476/X sky130_fd_sc_hd__bufbuf_16
XFILLER_104_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6217_ _7076_/Q _6009_/X wire627/X _6972_/Q VGND VGND VPWR VPWR _6217_/X sky130_fd_sc_hd__a22o_1
XFILLER_77_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold498 _6660_/Q VGND VGND VPWR VPWR hold498/X sky130_fd_sc_hd__bufbuf_16
X_3429_ _7042_/Q _5468_/A _5423_/A _7002_/Q _3428_/X VGND VGND VPWR VPWR _3450_/B
+ sky130_fd_sc_hd__a221o_1
X_7197_ _7220_/CLK _7197_/D fanout856/X VGND VGND VPWR VPWR _7197_/Q sky130_fd_sc_hd__dfrtp_4
X_6148_ _6953_/Q wire637/X wire635/X _6929_/Q VGND VGND VPWR VPWR _6148_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6079_ wire555/X wire585/X wire618/A _7046_/Q _6078_/X VGND VGND VPWR VPWR _6082_/C
+ sky130_fd_sc_hd__a221o_4
XFILLER_57_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_305 mgmt_gpio_in[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_316 wire647/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_349 _5598_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_338 hold578/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_327 _6408_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3780_ _6805_/Q _5200_/A _4166_/A _6634_/Q _3779_/X VGND VGND VPWR VPWR _3785_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5450_ _5450_/A _5576_/B VGND VGND VPWR VPWR _5458_/S sky130_fd_sc_hd__nand2_8
XFILLER_173_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4401_ _4553_/B _4410_/C _4513_/A VGND VGND VPWR VPWR _4575_/B sky130_fd_sc_hd__nor3_4
XFILLER_117_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5381_ _5597_/A0 hold287/X _5386_/S VGND VGND VPWR VPWR _6959_/D sky130_fd_sc_hd__mux2_1
X_7120_ _7147_/CLK _7120_/D fanout888/X VGND VGND VPWR VPWR _7120_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_113_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A VGND VGND VPWR VPWR _7210_/CLK sky130_fd_sc_hd__clkbuf_8
X_4332_ _6410_/A0 hold669/X _4333_/S VGND VGND VPWR VPWR _6776_/D sky130_fd_sc_hd__mux2_1
XFILLER_140_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4263_ hold594/X wire799/A _4267_/S VGND VGND VPWR VPWR _6718_/D sky130_fd_sc_hd__mux2_1
X_7051_ _7140_/CLK _7051_/D fanout865/X VGND VGND VPWR VPWR _7051_/Q sky130_fd_sc_hd__dfrtp_2
X_3214_ _3214_/A VGND VGND VPWR VPWR _3214_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6002_ _6019_/A _6010_/B VGND VGND VPWR VPWR _6002_/Y sky130_fd_sc_hd__nor2_2
X_4194_ _6410_/A0 hold697/X _4195_/S VGND VGND VPWR VPWR _6657_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6904_ _7152_/CLK _6904_/D fanout882/X VGND VGND VPWR VPWR _6904_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6835_ _6980_/CLK _6835_/D fanout878/X VGND VGND VPWR VPWR _6835_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3978_ _3978_/A _6406_/B VGND VGND VPWR VPWR _3994_/S sky130_fd_sc_hd__and2_4
X_6766_ _7223_/CLK _6766_/D fanout850/X VGND VGND VPWR VPWR _6766_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_164_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5717_ _6909_/Q _5680_/X _5931_/A2 _6869_/Q VGND VGND VPWR VPWR _5717_/X sky130_fd_sc_hd__a22o_1
Xwire609 _6111_/B VGND VGND VPWR VPWR _6211_/B sky130_fd_sc_hd__buf_8
X_6697_ _7133_/CLK _6697_/D fanout882/X VGND VGND VPWR VPWR _6697_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5648_ _7170_/Q _5648_/B _6035_/A VGND VGND VPWR VPWR _5654_/B sky130_fd_sc_hd__and3_1
X_5579_ _5579_/A0 hold792/X _5580_/S VGND VGND VPWR VPWR _7135_/D sky130_fd_sc_hd__mux2_1
Xhold262 _3993_/X VGND VGND VPWR VPWR hold20/A sky130_fd_sc_hd__bufbuf_16
Xhold240 _6865_/Q VGND VGND VPWR VPWR hold240/X sky130_fd_sc_hd__bufbuf_16
XFILLER_123_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold251 _6689_/Q VGND VGND VPWR VPWR wire821/A sky130_fd_sc_hd__bufbuf_16
Xhold295 _5494_/X VGND VGND VPWR VPWR _7060_/D sky130_fd_sc_hd__bufbuf_16
Xhold284 _5431_/X VGND VGND VPWR VPWR _7004_/D sky130_fd_sc_hd__bufbuf_16
Xhold273 _6955_/Q VGND VGND VPWR VPWR hold273/X sky130_fd_sc_hd__bufbuf_16
XFILLER_132_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout720 _5242_/B VGND VGND VPWR VPWR _6406_/B sky130_fd_sc_hd__buf_8
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout764 hold154/X VGND VGND VPWR VPWR _5599_/A0 sky130_fd_sc_hd__buf_8
XFILLER_172_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout797 wire799/A VGND VGND VPWR VPWR _6407_/A0 sky130_fd_sc_hd__buf_8
XFILLER_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_102 _6029_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_113 debug_oeb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_124 mask_rev_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_157 wb_adr_i[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_135 mgmt_gpio_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_146 pad_flash_io0_di VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_168 input92/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_179 _3929_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length730 wire729/A VGND VGND VPWR VPWR fanout724/A sky130_fd_sc_hd__buf_6
Xmax_length752 wire753/X VGND VGND VPWR VPWR _5519_/A0 sky130_fd_sc_hd__buf_6
XFILLER_182_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput8 mask_rev_in[13] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4950_ _4950_/A _4950_/B _4950_/C VGND VGND VPWR VPWR _5129_/B sky130_fd_sc_hd__or3_4
XFILLER_64_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4881_ _4881_/A _4881_/B VGND VGND VPWR VPWR _4905_/B sky130_fd_sc_hd__nand2_1
X_3901_ _7170_/Q _7171_/Q VGND VGND VPWR VPWR _6019_/A sky130_fd_sc_hd__nand2b_4
X_6620_ _6621_/CLK _6620_/D fanout873/X VGND VGND VPWR VPWR _6620_/Q sky130_fd_sc_hd__dfrtp_2
X_3832_ _3831_/X _6480_/Q _3840_/S VGND VGND VPWR VPWR _6480_/D sky130_fd_sc_hd__mux2_1
XFILLER_158_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6551_ _6554_/CLK _6551_/D fanout858/X VGND VGND VPWR VPWR _6551_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3763_ _6885_/Q _5297_/A _3763_/B1 _7133_/Q _3738_/X VGND VGND VPWR VPWR _3764_/D
+ sky130_fd_sc_hd__a221o_1
X_5502_ _5547_/A0 hold811/X _5502_/S VGND VGND VPWR VPWR _7067_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6482_ _6668_/CLK _6482_/D _6437_/X VGND VGND VPWR VPWR _6482_/Q sky130_fd_sc_hd__dfrtp_2
X_3694_ _6812_/Q _5207_/A _3365_/Y _7134_/Q _3678_/X VGND VGND VPWR VPWR _3699_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5433_ wire802/X _7005_/Q _5440_/S VGND VGND VPWR VPWR _5433_/X sky130_fd_sc_hd__mux2_1
Xoutput301 _6820_/Q VGND VGND VPWR VPWR pwr_ctrl_out[0] sky130_fd_sc_hd__buf_8
XFILLER_161_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput334 _7203_/Q VGND VGND VPWR VPWR wb_dat_o[24] sky130_fd_sc_hd__buf_8
X_5364_ wire773/X hold621/X _5368_/S VGND VGND VPWR VPWR _6944_/D sky130_fd_sc_hd__mux2_1
Xoutput323 _6574_/Q VGND VGND VPWR VPWR wb_dat_o[14] sky130_fd_sc_hd__buf_8
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput312 _3970_/X VGND VGND VPWR VPWR spi_sdi sky130_fd_sc_hd__buf_8
XFILLER_126_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput345 _6586_/Q VGND VGND VPWR VPWR wb_dat_o[5] sky130_fd_sc_hd__buf_8
X_7103_ _7103_/CLK _7103_/D fanout861/X VGND VGND VPWR VPWR _7103_/Q sky130_fd_sc_hd__dfrtp_2
X_4315_ hold651/X _6411_/A0 _4315_/S VGND VGND VPWR VPWR _6762_/D sky130_fd_sc_hd__mux2_1
X_5295_ _5601_/A0 _6883_/Q _5296_/S VGND VGND VPWR VPWR _5295_/X sky130_fd_sc_hd__mux2_1
X_4246_ _5599_/A0 hold310/X hold32/X VGND VGND VPWR VPWR _4246_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7034_ _7042_/CLK _7034_/D fanout865/X VGND VGND VPWR VPWR _7034_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_67_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4177_ hold652/X _6411_/A0 _4177_/S VGND VGND VPWR VPWR _6643_/D sky130_fd_sc_hd__mux2_1
XFILLER_82_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6818_ _7103_/CLK _6818_/D fanout861/X VGND VGND VPWR VPWR _6818_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_23_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire406 _3353_/Y VGND VGND VPWR VPWR wire406/X sky130_fd_sc_hd__buf_8
XFILLER_149_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire439 wire439/A VGND VGND VPWR VPWR wire439/X sky130_fd_sc_hd__buf_8
Xwire417 _3334_/Y VGND VGND VPWR VPWR _5468_/A sky130_fd_sc_hd__buf_8
X_6749_ _7225_/CLK _6749_/D fanout851/X VGND VGND VPWR VPWR _6749_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_109_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length582 _6252_/B1 VGND VGND VPWR VPWR _6339_/A2 sky130_fd_sc_hd__buf_6
XFILLER_6_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4100_ _5498_/A0 hold755/X _4102_/S VGND VGND VPWR VPWR _6578_/D sky130_fd_sc_hd__mux2_1
X_5080_ _4586_/B _4987_/X _4850_/X _4617_/Y _4798_/A VGND VGND VPWR VPWR _5171_/B
+ sky130_fd_sc_hd__a2111o_4
XFILLER_110_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4031_ _5600_/A0 hold468/X _4033_/S VGND VGND VPWR VPWR _6519_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5982_ _6534_/Q _5722_/B _5976_/X _5981_/X _6308_/S VGND VGND VPWR VPWR _5982_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_64_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4933_ _5165_/A _4933_/B VGND VGND VPWR VPWR _4933_/Y sky130_fd_sc_hd__nand2_1
XFILLER_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_13 _6517_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4864_ _4648_/B _5164_/B _4638_/X VGND VGND VPWR VPWR _4865_/C sky130_fd_sc_hd__o21ai_2
XFILLER_60_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_24 _6864_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6603_ _6747_/CLK _6603_/D fanout874/X VGND VGND VPWR VPWR _6603_/Q sky130_fd_sc_hd__dfrtp_2
X_4795_ _4772_/A _5165_/A _4428_/C _4794_/X VGND VGND VPWR VPWR _4796_/D sky130_fd_sc_hd__a31o_1
XANTENNA_46 _4124_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_57 _3687_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3815_ _6483_/Q _6482_/Q _6481_/Q _3828_/S VGND VGND VPWR VPWR _3820_/B sky130_fd_sc_hd__nand4_2
XANTENNA_35 _3255_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_79 _4238_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3746_ _6941_/Q wire401/X _4268_/A _6723_/Q VGND VGND VPWR VPWR _3746_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_68 _3693_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6534_ _7225_/CLK _6534_/D fanout850/X VGND VGND VPWR VPWR _6534_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_180_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6465_ _3938_/A1 _6465_/D _6420_/X VGND VGND VPWR VPWR _6465_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3677_ _6489_/Q _3978_/A _4322_/A _6769_/Q _3676_/X VGND VGND VPWR VPWR _3717_/A
+ sky130_fd_sc_hd__a221o_2
X_5416_ _5578_/A0 hold438/X _5422_/S VGND VGND VPWR VPWR _6990_/D sky130_fd_sc_hd__mux2_1
X_6396_ _4236_/C _6396_/A2 _6396_/B1 _4238_/B _6395_/X VGND VGND VPWR VPWR _6396_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5347_ hold150/X hold242/X _5350_/S VGND VGND VPWR VPWR _6929_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput175 wire442/X VGND VGND VPWR VPWR mgmt_gpio_oeb[0] sky130_fd_sc_hd__buf_8
Xoutput186 _3946_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[1] sky130_fd_sc_hd__buf_8
X_5278_ _5602_/A0 hold280/X _5278_/S VGND VGND VPWR VPWR _5278_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput197 _3237_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[2] sky130_fd_sc_hd__buf_8
X_4229_ hold584/X _4228_/X _4235_/S VGND VGND VPWR VPWR _4229_/X sky130_fd_sc_hd__mux2_1
X_7017_ _7095_/CLK _7017_/D fanout863/X VGND VGND VPWR VPWR _7017_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_101_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout380 _5664_/X VGND VGND VPWR VPWR wire381/A sky130_fd_sc_hd__buf_8
XFILLER_19_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4580_ _4581_/B _4634_/B _4536_/X _4581_/A VGND VGND VPWR VPWR _4612_/A sky130_fd_sc_hd__a22oi_4
XFILLER_174_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3600_ _6756_/Q _4304_/A _4049_/A _6538_/Q _3560_/X VGND VGND VPWR VPWR _3605_/B
+ sky130_fd_sc_hd__a221o_2
Xinput11 mask_rev_in[16] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__clkbuf_4
XFILLER_30_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput22 mask_rev_in[26] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__clkbuf_4
Xinput55 mgmt_gpio_in[27] VGND VGND VPWR VPWR input55/X sky130_fd_sc_hd__clkbuf_8
XFILLER_174_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput44 mgmt_gpio_in[17] VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__clkbuf_4
XFILLER_162_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3531_ _3543_/A _3539_/B VGND VGND VPWR VPWR _4097_/A sky130_fd_sc_hd__nor2_8
Xwire770 wire770/A VGND VGND VPWR VPWR wire770/X sky130_fd_sc_hd__buf_8
Xinput33 mask_rev_in[7] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__clkbuf_4
XFILLER_183_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput88 spimemio_flash_io1_oeb VGND VGND VPWR VPWR wire839/A sky130_fd_sc_hd__buf_6
Xhold806 _6733_/Q VGND VGND VPWR VPWR hold806/X sky130_fd_sc_hd__bufbuf_16
Xinput66 mgmt_gpio_in[37] VGND VGND VPWR VPWR wire897/A sky130_fd_sc_hd__buf_6
XFILLER_128_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold828 _6829_/Q VGND VGND VPWR VPWR hold828/X sky130_fd_sc_hd__bufbuf_16
XFILLER_6_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold817 _5528_/X VGND VGND VPWR VPWR _7090_/D sky130_fd_sc_hd__bufbuf_16
Xinput77 ser_tx VGND VGND VPWR VPWR input77/X sky130_fd_sc_hd__clkbuf_4
Xinput99 wb_adr_i[0] VGND VGND VPWR VPWR _4672_/A sky130_fd_sc_hd__buf_8
XFILLER_143_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3462_ _3540_/A hold45/X VGND VGND VPWR VPWR _4256_/A sky130_fd_sc_hd__nor2_8
X_6250_ _6594_/Q _6340_/B1 _6036_/Y _6748_/Q _6249_/X VGND VGND VPWR VPWR _6257_/B
+ sky130_fd_sc_hd__a221o_1
Xhold839 _6755_/Q VGND VGND VPWR VPWR hold839/X sky130_fd_sc_hd__bufbuf_16
X_6181_ _6181_/A _6181_/B _6181_/C _6181_/D VGND VGND VPWR VPWR _6182_/C sky130_fd_sc_hd__or4_1
XFILLER_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3393_ _6963_/Q _3305_/Y _5576_/A _7139_/Q _3390_/X VGND VGND VPWR VPWR _3398_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5201_ _6407_/A0 hold754/X _5206_/S VGND VGND VPWR VPWR _6805_/D sky130_fd_sc_hd__mux2_1
X_5132_ _5132_/A _5133_/A _5132_/C VGND VGND VPWR VPWR _5143_/B sky130_fd_sc_hd__or3_2
XFILLER_96_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5063_ _4505_/X _5062_/B _4963_/Y _5062_/X _4612_/C VGND VGND VPWR VPWR _5066_/A
+ sky130_fd_sc_hd__o2111a_4
XFILLER_111_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4014_ hold385/X _4013_/X _4024_/S VGND VGND VPWR VPWR _4014_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5965_ _6742_/Q wire700/X wire679/X _7225_/Q VGND VGND VPWR VPWR _5981_/A sky130_fd_sc_hd__a22o_1
XFILLER_40_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4916_ _6779_/Q _4239_/X _4807_/X _4915_/X VGND VGND VPWR VPWR _6779_/D sky130_fd_sc_hd__o22a_1
X_5896_ _7184_/Q _6309_/S _5895_/X VGND VGND VPWR VPWR _7184_/D sky130_fd_sc_hd__o21a_1
X_4847_ _4847_/A _5174_/A VGND VGND VPWR VPWR _5171_/A sky130_fd_sc_hd__or2_2
XFILLER_32_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4778_ _5165_/A _4778_/B VGND VGND VPWR VPWR _5033_/C sky130_fd_sc_hd__and2_1
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6517_ _7152_/CLK _6517_/D fanout886/X VGND VGND VPWR VPWR _6517_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_174_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3729_ _3728_/X _6791_/Q _3928_/A VGND VGND VPWR VPWR _6791_/D sky130_fd_sc_hd__mux2_1
XFILLER_106_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6448_ _6455_/A _6455_/B VGND VGND VPWR VPWR _6448_/X sky130_fd_sc_hd__and2_1
X_6379_ _6378_/X _7211_/Q _6400_/S VGND VGND VPWR VPWR _7211_/D sky130_fd_sc_hd__mux2_1
XFILLER_164_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5750_ _6895_/Q wire672/X _5749_/X VGND VGND VPWR VPWR _5753_/C sky130_fd_sc_hd__a21o_1
XFILLER_97_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4701_ _5050_/A _4711_/A _4707_/B VGND VGND VPWR VPWR _4702_/B sky130_fd_sc_hd__a21oi_1
X_5681_ _5864_/B _5702_/B _5706_/B VGND VGND VPWR VPWR _5681_/X sky130_fd_sc_hd__and3_4
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4632_ _4996_/A _4989_/A VGND VGND VPWR VPWR _5078_/B sky130_fd_sc_hd__nor2_2
XFILLER_190_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4563_ _4763_/B _4980_/A _4559_/X _4980_/B _4367_/X VGND VGND VPWR VPWR _4563_/X
+ sky130_fd_sc_hd__o41a_2
Xhold603 _7040_/Q VGND VGND VPWR VPWR hold603/X sky130_fd_sc_hd__bufbuf_16
X_4494_ _4501_/A _4648_/B VGND VGND VPWR VPWR _4494_/Y sky130_fd_sc_hd__nor2_4
X_6302_ wire572/X wire585/X wire618/X _6641_/Q _6301_/X VGND VGND VPWR VPWR _6305_/C
+ sky130_fd_sc_hd__a221o_1
X_3514_ _3514_/A _3732_/B VGND VGND VPWR VPWR _4322_/A sky130_fd_sc_hd__nor2_8
Xhold614 _6777_/Q VGND VGND VPWR VPWR hold614/X sky130_fd_sc_hd__bufbuf_16
Xhold636 _6999_/Q VGND VGND VPWR VPWR hold636/X sky130_fd_sc_hd__bufbuf_16
Xhold625 _6789_/Q VGND VGND VPWR VPWR hold625/X sky130_fd_sc_hd__bufbuf_16
XFILLER_171_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold647 _6511_/Q VGND VGND VPWR VPWR hold647/X sky130_fd_sc_hd__bufbuf_16
XFILLER_116_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold658 _7108_/Q VGND VGND VPWR VPWR hold658/X sky130_fd_sc_hd__bufbuf_16
XFILLER_6_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold669 _6776_/Q VGND VGND VPWR VPWR hold669/X sky130_fd_sc_hd__bufbuf_16
X_6233_ _6860_/Q _6060_/B _6219_/X _6232_/X _3197_/Y VGND VGND VPWR VPWR _6233_/X
+ sky130_fd_sc_hd__o221a_1
X_3445_ _7010_/Q _5432_/A _3325_/Y wire536/X _3444_/X VGND VGND VPWR VPWR _3451_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_170_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3376_ _6876_/Q _3425_/B1 _5369_/A _6956_/Q _3373_/X VGND VGND VPWR VPWR _3377_/D
+ sky130_fd_sc_hd__a221o_4
X_6164_ _7026_/Q wire589/X wire615/X _7090_/Q _6163_/X VGND VGND VPWR VPWR _6170_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6095_ _6983_/Q _6028_/X _6342_/B1 _6991_/Q _6094_/X VGND VGND VPWR VPWR _6095_/X
+ sky130_fd_sc_hd__a221o_1
X_5115_ _5115_/A _5115_/B VGND VGND VPWR VPWR _5137_/B sky130_fd_sc_hd__or2_1
XFILLER_57_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5046_ _5046_/A _5108_/A _5154_/A VGND VGND VPWR VPWR _5057_/A sky130_fd_sc_hd__or3_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6997_ _7140_/CLK _6997_/D fanout862/X VGND VGND VPWR VPWR _6997_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_26_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5948_ _6622_/Q wire707/X _5681_/X _6597_/Q _5947_/X VGND VGND VPWR VPWR _5953_/B
+ sky130_fd_sc_hd__a221o_4
XFILLER_43_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5879_ _6634_/Q _5973_/A2 wire694/X _6773_/Q VGND VGND VPWR VPWR _5879_/X sky130_fd_sc_hd__a22o_1
XFILLER_193_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3230_ _6936_/Q VGND VGND VPWR VPWR _3230_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6920_ _7068_/CLK _6920_/D fanout878/X VGND VGND VPWR VPWR _6920_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_94_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6851_ _6851_/CLK _6851_/D _6447_/A VGND VGND VPWR VPWR _6851_/Q sky130_fd_sc_hd__dfrtp_1
X_5802_ _6913_/Q wire699/X wire666/X _6865_/Q VGND VGND VPWR VPWR _5802_/X sky130_fd_sc_hd__a22o_4
XFILLER_62_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6782_ _7190_/CLK _6782_/D wire915/A VGND VGND VPWR VPWR _6782_/Q sky130_fd_sc_hd__dfrtp_2
X_3994_ _6495_/Q wire739/X _3994_/S VGND VGND VPWR VPWR _6495_/D sky130_fd_sc_hd__mux2_1
X_5733_ _6974_/Q wire702/X _5702_/X _6886_/Q _5732_/X VGND VGND VPWR VPWR _5734_/D
+ sky130_fd_sc_hd__a221o_4
XFILLER_176_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5664_ _5665_/A _5665_/B VGND VGND VPWR VPWR _5664_/X sky130_fd_sc_hd__or2_4
X_5595_ _5595_/A0 hold726/X hold66/X VGND VGND VPWR VPWR _7149_/D sky130_fd_sc_hd__mux2_1
X_4615_ _4846_/B _4615_/B _4615_/C VGND VGND VPWR VPWR _4619_/B sky130_fd_sc_hd__and3b_1
XFILLER_129_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_54_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7082_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_191_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold400 _5554_/X VGND VGND VPWR VPWR _7113_/D sky130_fd_sc_hd__bufbuf_16
X_4546_ _4850_/A _5022_/A _4546_/C _4546_/D VGND VGND VPWR VPWR _4548_/C sky130_fd_sc_hd__or4_1
Xhold411 _6849_/Q VGND VGND VPWR VPWR hold411/X sky130_fd_sc_hd__bufbuf_16
Xhold433 _7058_/Q VGND VGND VPWR VPWR hold433/X sky130_fd_sc_hd__bufbuf_16
Xhold444 _5290_/X VGND VGND VPWR VPWR _6878_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_150_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold422 _6992_/Q VGND VGND VPWR VPWR hold422/X sky130_fd_sc_hd__bufbuf_16
Xhold466 _4242_/X VGND VGND VPWR VPWR _6690_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_171_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4477_ _4603_/B _4749_/C VGND VGND VPWR VPWR _4883_/A sky130_fd_sc_hd__nor2_1
XFILLER_89_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold455 _4273_/X VGND VGND VPWR VPWR _6727_/D sky130_fd_sc_hd__bufbuf_16
Xhold477 _6945_/Q VGND VGND VPWR VPWR hold477/X sky130_fd_sc_hd__bufbuf_16
X_6216_ _7124_/Q _6252_/B1 wire579/X _7036_/Q _6215_/X VGND VGND VPWR VPWR _6219_/C
+ sky130_fd_sc_hd__a221o_2
Xhold488 _4272_/X VGND VGND VPWR VPWR _6726_/D sky130_fd_sc_hd__bufbuf_16
Xclkbuf_leaf_69_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7118_/CLK sky130_fd_sc_hd__clkbuf_8
X_3428_ input31/X _3283_/Y _3335_/Y _6493_/Q VGND VGND VPWR VPWR _3428_/X sky130_fd_sc_hd__a22o_2
X_7196_ _7196_/CLK _7196_/D fanout868/X VGND VGND VPWR VPWR _7196_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout913 wire915/A VGND VGND VPWR VPWR _6362_/B sky130_fd_sc_hd__buf_8
Xhold499 _7074_/Q VGND VGND VPWR VPWR hold499/X sky130_fd_sc_hd__bufbuf_16
X_3359_ _3505_/A _3375_/B VGND VGND VPWR VPWR _5441_/A sky130_fd_sc_hd__nor2_8
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6147_ _7129_/Q wire597/X wire611/X _7009_/Q wire441/X VGND VGND VPWR VPWR _6157_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_100_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6078_ _7102_/Q wire712/X wire625/X _6942_/Q VGND VGND VPWR VPWR _6078_/X sky130_fd_sc_hd__a22o_1
XFILLER_57_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5029_ _4414_/B _4711_/C _4704_/X _4802_/A _4932_/B VGND VGND VPWR VPWR _5101_/A
+ sky130_fd_sc_hd__a2111o_1
XANTENNA_306 _6828_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_328 _5595_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_339 hold617/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_317 wire649/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4400_ _4400_/A _4513_/A VGND VGND VPWR VPWR _4617_/A sky130_fd_sc_hd__or2_4
X_5380_ hold38/X _6958_/Q _5386_/S VGND VGND VPWR VPWR _6958_/D sky130_fd_sc_hd__mux2_1
XFILLER_126_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4331_ _6409_/A0 _6775_/Q _4333_/S VGND VGND VPWR VPWR _6775_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4262_ _4262_/A _5242_/B VGND VGND VPWR VPWR _4267_/S sky130_fd_sc_hd__and2_4
X_7050_ _7140_/CLK _7050_/D fanout865/X VGND VGND VPWR VPWR _7050_/Q sky130_fd_sc_hd__dfrtp_2
X_3213_ _3213_/A VGND VGND VPWR VPWR _3213_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6001_ _6037_/A _6032_/A VGND VGND VPWR VPWR _6010_/B sky130_fd_sc_hd__nand2_8
XFILLER_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4193_ _6409_/A0 _6656_/Q _4195_/S VGND VGND VPWR VPWR _6656_/D sky130_fd_sc_hd__mux2_1
X_6903_ _7111_/CLK _6903_/D _6421_/A VGND VGND VPWR VPWR _6903_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_63_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6834_ _6980_/CLK hold8/X fanout878/X VGND VGND VPWR VPWR _6834_/Q sky130_fd_sc_hd__dfrtp_2
X_6765_ _7223_/CLK _6765_/D fanout848/X VGND VGND VPWR VPWR _6765_/Q sky130_fd_sc_hd__dfstp_4
X_3977_ hold140/X hold252/X hold69/X VGND VGND VPWR VPWR hold70/A sky130_fd_sc_hd__o21ai_4
XFILLER_50_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5716_ _6861_/Q wire667/A wire653/A wire503/X _5686_/X VGND VGND VPWR VPWR _5720_/B
+ sky130_fd_sc_hd__a221o_1
X_6696_ _7133_/CLK _6696_/D fanout882/X VGND VGND VPWR VPWR _6696_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_164_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5647_ _7169_/Q _5635_/B _5645_/Y _5646_/X VGND VGND VPWR VPWR _7169_/D sky130_fd_sc_hd__a31o_1
XFILLER_191_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5578_ _5578_/A0 hold396/X _5580_/S VGND VGND VPWR VPWR _7134_/D sky130_fd_sc_hd__mux2_1
X_4529_ _4529_/A _4529_/B _4529_/C VGND VGND VPWR VPWR _4533_/B sky130_fd_sc_hd__and3_4
Xhold241 _7065_/Q VGND VGND VPWR VPWR hold241/X sky130_fd_sc_hd__bufbuf_16
XFILLER_117_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold230 _6711_/Q VGND VGND VPWR VPWR hold230/X sky130_fd_sc_hd__bufbuf_16
Xhold252 _3975_/B VGND VGND VPWR VPWR hold252/X sky130_fd_sc_hd__bufbuf_16
Xhold263 hold20/X VGND VGND VPWR VPWR hold263/X sky130_fd_sc_hd__bufbuf_16
Xhold296 _6747_/Q VGND VGND VPWR VPWR hold296/X sky130_fd_sc_hd__bufbuf_16
Xhold285 _6887_/Q VGND VGND VPWR VPWR hold285/X sky130_fd_sc_hd__bufbuf_16
Xhold274 _6889_/Q VGND VGND VPWR VPWR hold274/X sky130_fd_sc_hd__bufbuf_16
XFILLER_104_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout721 fanout724/A VGND VGND VPWR VPWR _5242_/B sky130_fd_sc_hd__buf_8
Xfanout765 hold154/X VGND VGND VPWR VPWR hold150/A sky130_fd_sc_hd__buf_8
Xfanout754 wire758/X VGND VGND VPWR VPWR _5600_/A0 sky130_fd_sc_hd__buf_8
Xfanout743 wire749/X VGND VGND VPWR VPWR wire746/A sky130_fd_sc_hd__buf_6
XFILLER_86_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7179_ _7196_/CLK _7179_/D fanout869/X VGND VGND VPWR VPWR _7179_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout776 _5579_/A0 VGND VGND VPWR VPWR _6409_/A0 sky130_fd_sc_hd__buf_8
XFILLER_105_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout798 wire802/A VGND VGND VPWR VPWR wire799/A sky130_fd_sc_hd__buf_8
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_114 debug_out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_125 mask_rev_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_103 _6072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_158 wb_adr_i[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_136 mgmt_gpio_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_147 pad_flash_io1_di VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_169 input81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput9 mask_rev_in[14] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4880_ _4875_/A _4588_/X _4593_/Y VGND VGND VPWR VPWR _4962_/A sky130_fd_sc_hd__o21ai_2
X_3900_ _6707_/Q _3883_/X _6702_/Q VGND VGND VPWR VPWR _6707_/D sky130_fd_sc_hd__a21o_1
XFILLER_177_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3831_ hold40/A _3845_/A _3824_/B _3830_/X VGND VGND VPWR VPWR _3831_/X sky130_fd_sc_hd__a22o_1
X_6550_ _6950_/CLK _6550_/D fanout874/X VGND VGND VPWR VPWR _6550_/Q sky130_fd_sc_hd__dfrtp_2
X_3762_ _6917_/Q _5333_/A _4292_/A _6743_/Q _3737_/X VGND VGND VPWR VPWR _3764_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5501_ _5600_/A0 hold451/X _5501_/S VGND VGND VPWR VPWR _7066_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3693_ _3693_/A _3693_/B _3693_/C _3693_/D VGND VGND VPWR VPWR _3727_/B sky130_fd_sc_hd__or4_2
XFILLER_9_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6481_ _6668_/CLK _6481_/D _6436_/X VGND VGND VPWR VPWR _6481_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_146_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5432_ _5432_/A _5576_/B VGND VGND VPWR VPWR _5440_/S sky130_fd_sc_hd__nand2_8
Xoutput313 wire807/X VGND VGND VPWR VPWR spimemio_flash_io0_di sky130_fd_sc_hd__buf_8
XFILLER_160_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput335 _7204_/Q VGND VGND VPWR VPWR wb_dat_o[25] sky130_fd_sc_hd__buf_8
Xoutput324 _6575_/Q VGND VGND VPWR VPWR wb_dat_o[15] sky130_fd_sc_hd__buf_8
X_5363_ wire786/X hold210/X _5365_/S VGND VGND VPWR VPWR _5363_/X sky130_fd_sc_hd__mux2_1
Xoutput302 _6821_/Q VGND VGND VPWR VPWR pwr_ctrl_out[1] sky130_fd_sc_hd__buf_8
XFILLER_160_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput346 _6587_/Q VGND VGND VPWR VPWR wb_dat_o[6] sky130_fd_sc_hd__buf_8
X_7102_ _7103_/CLK _7102_/D fanout861/X VGND VGND VPWR VPWR _7102_/Q sky130_fd_sc_hd__dfstp_4
X_4314_ hold656/X _6410_/A0 _4315_/S VGND VGND VPWR VPWR _6761_/D sky130_fd_sc_hd__mux2_1
X_5294_ _5600_/A0 hold507/X _5296_/S VGND VGND VPWR VPWR _6882_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4245_ _5598_/A0 hold626/X hold32/X VGND VGND VPWR VPWR _4245_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7033_ _7118_/CLK _7033_/D fanout869/X VGND VGND VPWR VPWR _7033_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_19_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4176_ hold709/X _6410_/A0 _4177_/S VGND VGND VPWR VPWR _6642_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6817_ _7103_/CLK _6817_/D fanout861/X VGND VGND VPWR VPWR _6817_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_167_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6748_ _6752_/CLK _6748_/D fanout857/X VGND VGND VPWR VPWR _6748_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6679_ _7194_/CLK _6679_/D fanout866/X VGND VGND VPWR VPWR _6679_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_151_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length583 _6017_/Y VGND VGND VPWR VPWR _6252_/B1 sky130_fd_sc_hd__buf_6
XFILLER_6_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4030_ hold150/X hold218/X _4033_/S VGND VGND VPWR VPWR _6518_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5981_ _5981_/A _5981_/B _5981_/C _5981_/D VGND VGND VPWR VPWR _5981_/X sky130_fd_sc_hd__or4_2
XFILLER_64_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4932_ _4932_/A _4932_/B _4932_/C VGND VGND VPWR VPWR _4940_/B sky130_fd_sc_hd__or3_1
XANTENNA_14 _6518_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6602_ _6950_/CLK _6602_/D fanout874/X VGND VGND VPWR VPWR _6602_/Q sky130_fd_sc_hd__dfrtp_2
X_4863_ _5118_/A _4863_/B _4863_/C _5084_/A VGND VGND VPWR VPWR _4865_/B sky130_fd_sc_hd__or4_1
XANTENNA_25 _5278_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4794_ _5165_/A _4793_/Y _4791_/X _5035_/B VGND VGND VPWR VPWR _4794_/X sky130_fd_sc_hd__a211o_1
XFILLER_119_702 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_47 _3522_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_36 hold97/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3814_ _6480_/Q _3830_/B VGND VGND VPWR VPWR _3828_/S sky130_fd_sc_hd__and2_2
XFILLER_20_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_69 _3709_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 _3687_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3745_ wire493/X _5522_/A _5459_/A wire511/X VGND VGND VPWR VPWR _3745_/X sky130_fd_sc_hd__a22o_1
X_6533_ _7225_/CLK _6533_/D fanout856/X VGND VGND VPWR VPWR _6533_/Q sky130_fd_sc_hd__dfstp_4
X_6464_ _3938_/A1 _6464_/D _6419_/X VGND VGND VPWR VPWR hold1/A sky130_fd_sc_hd__dfrtp_2
XFILLER_161_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3676_ input35/X _3320_/Y _4049_/A _6536_/Q VGND VGND VPWR VPWR _3676_/X sky130_fd_sc_hd__a22o_1
X_5415_ wire802/X _6989_/Q _5422_/S VGND VGND VPWR VPWR _6989_/D sky130_fd_sc_hd__mux2_1
X_6395_ _4236_/B _6395_/A2 _6395_/B1 _4236_/A VGND VGND VPWR VPWR _6395_/X sky130_fd_sc_hd__a22o_1
X_5346_ _5598_/A0 hold561/X _5350_/S VGND VGND VPWR VPWR _6928_/D sky130_fd_sc_hd__mux2_1
Xoutput176 _3230_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[10] sky130_fd_sc_hd__buf_8
XFILLER_99_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput187 _3220_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[20] sky130_fd_sc_hd__buf_8
Xoutput198 _3210_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[30] sky130_fd_sc_hd__buf_8
XFILLER_153_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5277_ _5601_/A0 hold212/X _5278_/S VGND VGND VPWR VPWR _5277_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7016_ _7132_/CLK _7016_/D fanout863/X VGND VGND VPWR VPWR _7016_/Q sky130_fd_sc_hd__dfrtp_2
X_4228_ hold411/X wire763/X _4234_/S VGND VGND VPWR VPWR _4228_/X sky130_fd_sc_hd__mux2_1
X_4159_ hold379/X _5599_/A0 _4159_/S VGND VGND VPWR VPWR _6628_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_1_0_mgmt_gpio_in[4] clkbuf_2_1_0_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR _6668_/CLK
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_19_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput12 mask_rev_in[17] VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__clkbuf_4
XFILLER_190_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput45 mgmt_gpio_in[18] VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__buf_4
X_3530_ _6633_/Q _4160_/A _4112_/A _6593_/Q VGND VGND VPWR VPWR _3530_/X sky130_fd_sc_hd__a22o_1
Xinput34 mask_rev_in[8] VGND VGND VPWR VPWR input34/X sky130_fd_sc_hd__clkbuf_4
Xinput23 mask_rev_in[27] VGND VGND VPWR VPWR input23/X sky130_fd_sc_hd__clkbuf_4
Xinput89 spimemio_flash_io2_do VGND VGND VPWR VPWR input89/X sky130_fd_sc_hd__clkbuf_4
XFILLER_155_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput56 mgmt_gpio_in[28] VGND VGND VPWR VPWR wire905/A sky130_fd_sc_hd__buf_6
XFILLER_128_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold818 _7026_/Q VGND VGND VPWR VPWR hold818/X sky130_fd_sc_hd__bufbuf_16
Xhold807 _6787_/Q VGND VGND VPWR VPWR hold807/X sky130_fd_sc_hd__bufbuf_16
Xinput78 spi_csb VGND VGND VPWR VPWR input78/X sky130_fd_sc_hd__clkbuf_4
Xinput67 mgmt_gpio_in[3] VGND VGND VPWR VPWR wire896/A sky130_fd_sc_hd__buf_6
XFILLER_182_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold829 _5231_/X VGND VGND VPWR VPWR _6829_/D sky130_fd_sc_hd__bufbuf_16
X_3461_ _6767_/Q _4316_/A _4328_/A _6777_/Q VGND VGND VPWR VPWR _3461_/X sky130_fd_sc_hd__a22o_4
XFILLER_170_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6180_ _7066_/Q wire648/X wire633/X _6914_/Q _6161_/X VGND VGND VPWR VPWR _6181_/D
+ sky130_fd_sc_hd__a221o_1
X_5200_ _5200_/A _6406_/B VGND VGND VPWR VPWR _5206_/S sky130_fd_sc_hd__nand2_4
X_3392_ _7091_/Q _5522_/A _5441_/A _7019_/Q VGND VGND VPWR VPWR _3392_/X sky130_fd_sc_hd__a22o_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5131_ _5131_/A _5146_/A _5143_/A VGND VGND VPWR VPWR _5133_/B sky130_fd_sc_hd__nor3_1
XFILLER_69_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5062_ _5062_/A _5062_/B _5062_/C VGND VGND VPWR VPWR _5062_/X sky130_fd_sc_hd__or3_1
X_4013_ _6524_/Q _5248_/A0 _4021_/S VGND VGND VPWR VPWR _4013_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5964_ _6648_/Q wire690/X _5964_/B1 _6603_/Q VGND VGND VPWR VPWR _5964_/X sky130_fd_sc_hd__a22o_1
X_4915_ _4367_/X _4867_/X _4914_/X VGND VGND VPWR VPWR _4915_/X sky130_fd_sc_hd__a21o_1
X_5895_ wire824/X _7183_/Q wire381/X _5894_/X VGND VGND VPWR VPWR _5895_/X sky130_fd_sc_hd__a211o_1
XFILLER_33_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4846_ _5033_/A _4846_/B VGND VGND VPWR VPWR _4846_/X sky130_fd_sc_hd__or2_2
XFILLER_138_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6516_ _7152_/CLK _6516_/D fanout882/X VGND VGND VPWR VPWR _6516_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_165_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4777_ _4772_/A _5165_/B _4698_/Y VGND VGND VPWR VPWR _4778_/B sky130_fd_sc_hd__a21o_1
XFILLER_21_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3728_ _3727_/X _6790_/Q _3857_/C VGND VGND VPWR VPWR _3728_/X sky130_fd_sc_hd__mux2_1
X_6447_ _6447_/A _6447_/B VGND VGND VPWR VPWR _6447_/X sky130_fd_sc_hd__and2_1
X_3659_ _6775_/Q _4328_/A _4172_/A _6641_/Q VGND VGND VPWR VPWR _3659_/X sky130_fd_sc_hd__a22o_1
X_6378_ _4236_/C _6378_/A2 _6378_/B1 _4238_/B _6377_/X VGND VGND VPWR VPWR _6378_/X
+ sky130_fd_sc_hd__a221o_1
X_5329_ hold150/X hold246/X _5332_/S VGND VGND VPWR VPWR _6913_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4700_ _4422_/Y _4423_/X _4424_/Y _4414_/B VGND VGND VPWR VPWR _4930_/C sky130_fd_sc_hd__o2bb2a_2
X_5680_ _5864_/B _5705_/B _5707_/C VGND VGND VPWR VPWR _5680_/X sky130_fd_sc_hd__and3_4
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4631_ _4995_/A _4844_/A _4575_/Y _4627_/X _4630_/Y VGND VGND VPWR VPWR _4631_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_30_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4562_ _4819_/B _4562_/B VGND VGND VPWR VPWR _4980_/B sky130_fd_sc_hd__nor2_8
XFILLER_128_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold626 _6693_/Q VGND VGND VPWR VPWR hold626/X sky130_fd_sc_hd__bufbuf_16
Xwire590 wire591/X VGND VGND VPWR VPWR wire590/X sky130_fd_sc_hd__buf_6
X_6301_ _6636_/Q wire711/X _6301_/B1 _6611_/Q VGND VGND VPWR VPWR _6301_/X sky130_fd_sc_hd__a22o_1
X_4493_ _4648_/B _5164_/B VGND VGND VPWR VPWR _4840_/A sky130_fd_sc_hd__nor2_1
X_3513_ wire905/X wire427/A _4049_/A _6539_/Q _3512_/X VGND VGND VPWR VPWR _3522_/B
+ sky130_fd_sc_hd__a221o_1
Xhold615 _7024_/Q VGND VGND VPWR VPWR hold615/X sky130_fd_sc_hd__bufbuf_16
Xhold604 _5472_/X VGND VGND VPWR VPWR _7040_/D sky130_fd_sc_hd__bufbuf_16
Xhold648 _4020_/X VGND VGND VPWR VPWR _6511_/D sky130_fd_sc_hd__bufbuf_16
Xhold637 _6936_/Q VGND VGND VPWR VPWR hold637/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3444_ input25/X _3302_/Y _3320_/Y input8/X VGND VGND VPWR VPWR _3444_/X sky130_fd_sc_hd__a22o_2
Xhold659 _6815_/Q VGND VGND VPWR VPWR hold659/X sky130_fd_sc_hd__bufbuf_16
X_6232_ _6232_/A _6232_/B _6232_/C VGND VGND VPWR VPWR _6232_/X sky130_fd_sc_hd__or3_1
XFILLER_112_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3375_ _3540_/A _3375_/B VGND VGND VPWR VPWR _5369_/A sky130_fd_sc_hd__nor2_8
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6163_ _7138_/Q wire642/X _6212_/B1 _7098_/Q VGND VGND VPWR VPWR _6163_/X sky130_fd_sc_hd__a22o_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5114_ _5114_/A _5114_/B _5114_/C _5114_/D VGND VGND VPWR VPWR _5115_/B sky130_fd_sc_hd__or4_1
X_6094_ _7071_/Q _6009_/X wire627/X wire528/X VGND VGND VPWR VPWR _6094_/X sky130_fd_sc_hd__a22o_1
XFILLER_69_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _4758_/B _5042_/Y _5016_/C _5035_/A VGND VGND VPWR VPWR _5154_/A sky130_fd_sc_hd__a211o_2
XFILLER_27_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6996_ _6996_/CLK _6996_/D fanout869/X VGND VGND VPWR VPWR _6996_/Q sky130_fd_sc_hd__dfrtp_2
X_5947_ _6711_/Q wire680/X wire664/X _6617_/Q VGND VGND VPWR VPWR _5947_/X sky130_fd_sc_hd__a22o_1
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5878_ _6659_/Q _5974_/A2 wire700/X _6738_/Q _5877_/X VGND VGND VPWR VPWR _5883_/B
+ sky130_fd_sc_hd__a221o_1
X_4829_ _4736_/B _4657_/B _4697_/Y _4828_/Y VGND VGND VPWR VPWR _4829_/X sky130_fd_sc_hd__a211o_1
XFILLER_166_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1 hold1/A VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__bufbuf_16
XFILLER_94_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6850_ _6994_/CLK _6850_/D fanout870/X VGND VGND VPWR VPWR _6850_/Q sky130_fd_sc_hd__dfrtp_4
X_5801_ _7017_/Q _5682_/X wire653/A wire500/X _5800_/X VGND VGND VPWR VPWR _5806_/B
+ sky130_fd_sc_hd__a221o_1
X_6781_ _7190_/CLK _6781_/D wire915/A VGND VGND VPWR VPWR _6781_/Q sky130_fd_sc_hd__dfrtp_2
X_3993_ hold19/X hold261/X _3993_/S VGND VGND VPWR VPWR _3993_/X sky130_fd_sc_hd__mux2_4
X_5732_ wire498/X _5921_/A2 wire671/X _6982_/Q _5697_/X VGND VGND VPWR VPWR _5732_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_50_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_1_mgmt_gpio_in[4] clkbuf_1_1_1_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR clkbuf_2_3_0_mgmt_gpio_in[4]/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_13_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5663_ _5663_/A _5663_/B VGND VGND VPWR VPWR _5663_/Y sky130_fd_sc_hd__nor2_2
XFILLER_30_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5594_ hold65/X _5594_/B VGND VGND VPWR VPWR hold66/A sky130_fd_sc_hd__nand2_8
X_4614_ _4997_/A _4844_/A VGND VGND VPWR VPWR _4615_/C sky130_fd_sc_hd__or2_1
XFILLER_163_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4545_ _4500_/A _4622_/B _4772_/A _4399_/Y _4847_/A VGND VGND VPWR VPWR _4546_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_129_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold401 _6752_/Q VGND VGND VPWR VPWR hold401/X sky130_fd_sc_hd__bufbuf_16
Xhold445 _6862_/Q VGND VGND VPWR VPWR hold445/X sky130_fd_sc_hd__bufbuf_16
XFILLER_190_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold434 _7130_/Q VGND VGND VPWR VPWR hold434/X sky130_fd_sc_hd__bufbuf_16
XFILLER_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold423 _7001_/Q VGND VGND VPWR VPWR hold423/X sky130_fd_sc_hd__bufbuf_16
Xhold412 _5257_/X VGND VGND VPWR VPWR _6849_/D sky130_fd_sc_hd__bufbuf_16
Xhold478 _6527_/Q VGND VGND VPWR VPWR hold478/X sky130_fd_sc_hd__bufbuf_16
X_4476_ _4558_/B _4584_/A VGND VGND VPWR VPWR _4749_/C sky130_fd_sc_hd__or2_4
XFILLER_89_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold456 _6543_/Q VGND VGND VPWR VPWR hold456/X sky130_fd_sc_hd__bufbuf_16
Xhold467 _6854_/Q VGND VGND VPWR VPWR hold467/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6215_ _7004_/Q wire604/X _6022_/D _6924_/Q VGND VGND VPWR VPWR _6215_/X sky130_fd_sc_hd__a22o_2
XFILLER_89_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3427_ _6816_/Q _5207_/A _5459_/A _7034_/Q wire369/X VGND VGND VPWR VPWR _3450_/A
+ sky130_fd_sc_hd__a221o_1
Xhold489 _6852_/Q VGND VGND VPWR VPWR hold489/X sky130_fd_sc_hd__bufbuf_16
Xfanout914 input164/X VGND VGND VPWR VPWR wire915/A sky130_fd_sc_hd__buf_8
X_7195_ _7196_/CLK _7195_/D fanout868/A VGND VGND VPWR VPWR _7195_/Q sky130_fd_sc_hd__dfrtp_4
X_6146_ _6889_/Q wire602/X wire581/X _7145_/Q _6145_/X VGND VGND VPWR VPWR _6146_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3358_ _5252_/A hold87/X VGND VGND VPWR VPWR hold88/A sky130_fd_sc_hd__nor2_8
XFILLER_97_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6077_ _6870_/Q wire593/X wire591/X _6894_/Q _6076_/X VGND VGND VPWR VPWR _6082_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_100_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3289_ hold42/X hold86/X VGND VGND VPWR VPWR _3343_/A sky130_fd_sc_hd__nand2_2
XANTENNA_307 wb_dat_i[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5028_ _5180_/C _5028_/B _5098_/B _5163_/B VGND VGND VPWR VPWR _5036_/A sky130_fd_sc_hd__or4_2
XFILLER_66_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_318 wire673/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_329 _3972_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6979_ _6979_/CLK _6979_/D fanout884/X VGND VGND VPWR VPWR _6979_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_186_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4330_ _6408_/A0 hold703/X _4333_/S VGND VGND VPWR VPWR _6774_/D sky130_fd_sc_hd__mux2_1
X_4261_ hold300/X _5599_/A0 _4261_/S VGND VGND VPWR VPWR _6717_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3212_ _7080_/Q VGND VGND VPWR VPWR _3212_/Y sky130_fd_sc_hd__inv_2
X_6000_ _6037_/B _6035_/A _6018_/A VGND VGND VPWR VPWR _6023_/B sky130_fd_sc_hd__and3_4
XFILLER_86_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4192_ _6408_/A0 hold686/X _4195_/S VGND VGND VPWR VPWR _6655_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6902_ _7128_/CLK _6902_/D _6421_/A VGND VGND VPWR VPWR _6902_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_54_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6833_ _6833_/CLK _6833_/D fanout873/X VGND VGND VPWR VPWR _6833_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6764_ _7223_/CLK _6764_/D fanout850/X VGND VGND VPWR VPWR _6764_/Q sky130_fd_sc_hd__dfrtp_2
X_3976_ hold140/X hold252/X hold69/X VGND VGND VPWR VPWR _3976_/X sky130_fd_sc_hd__o21a_1
XFILLER_50_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6695_ _7133_/CLK hold4/X fanout881/X VGND VGND VPWR VPWR _6695_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5715_ _6965_/Q wire680/X wire659/X _6933_/Q _5714_/X VGND VGND VPWR VPWR _5720_/A
+ sky130_fd_sc_hd__a221o_1
X_5646_ _6679_/Q _6037_/A _6037_/B VGND VGND VPWR VPWR _5646_/X sky130_fd_sc_hd__and3_1
XFILLER_163_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5577_ _5595_/A0 _7133_/Q _5581_/S VGND VGND VPWR VPWR _7133_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold220 _4146_/X VGND VGND VPWR VPWR _6617_/D sky130_fd_sc_hd__bufbuf_16
X_4528_ _4444_/B _4958_/B VGND VGND VPWR VPWR _4949_/B sky130_fd_sc_hd__and2b_4
Xhold242 _6929_/Q VGND VGND VPWR VPWR hold242/X sky130_fd_sc_hd__bufbuf_16
XFILLER_132_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold231 _4254_/X VGND VGND VPWR VPWR _6711_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_104_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold253 _3976_/X VGND VGND VPWR VPWR hold253/X sky130_fd_sc_hd__bufbuf_16
Xhold275 _7055_/Q VGND VGND VPWR VPWR hold275/X sky130_fd_sc_hd__bufbuf_16
Xhold286 _6892_/Q VGND VGND VPWR VPWR hold286/X sky130_fd_sc_hd__bufbuf_16
Xhold264 hold264/A VGND VGND VPWR VPWR hold21/A sky130_fd_sc_hd__bufbuf_16
XFILLER_131_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4459_ _4694_/A _4989_/A VGND VGND VPWR VPWR _4763_/B sky130_fd_sc_hd__nor2_1
Xfanout733 _4719_/C VGND VGND VPWR VPWR _4692_/C sky130_fd_sc_hd__buf_8
Xhold297 _4297_/X VGND VGND VPWR VPWR _6747_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_77_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout722 _5459_/B VGND VGND VPWR VPWR _5576_/B sky130_fd_sc_hd__buf_8
Xfanout755 hold25/X VGND VGND VPWR VPWR hold26/A sky130_fd_sc_hd__buf_6
XFILLER_131_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7178_ _7196_/CLK _7178_/D fanout869/X VGND VGND VPWR VPWR _7178_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_58_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout766 _5249_/A0 VGND VGND VPWR VPWR _6410_/A0 sky130_fd_sc_hd__buf_8
X_6129_ _3209_/A wire711/X _6022_/B _6944_/Q VGND VGND VPWR VPWR _6129_/X sky130_fd_sc_hd__a22o_2
Xfanout777 wire786/X VGND VGND VPWR VPWR wire780/A sky130_fd_sc_hd__buf_6
XFILLER_85_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout788 wire790/X VGND VGND VPWR VPWR _6408_/A0 sky130_fd_sc_hd__buf_8
XFILLER_100_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_104 _6082_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_115 _6938_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_137 mgmt_gpio_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_148 porb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_126 mask_rev_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_159 wb_adr_i[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length787 hold13/X VGND VGND VPWR VPWR _5248_/A0 sky130_fd_sc_hd__buf_6
XFILLER_6_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_53_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _6994_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_29_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_68_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7036_/CLK sky130_fd_sc_hd__clkbuf_8
X_3830_ _6480_/Q _3830_/B VGND VGND VPWR VPWR _3830_/X sky130_fd_sc_hd__or2_1
XFILLER_158_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3761_ _6909_/Q wire424/X _4160_/A _6629_/Q _3736_/X VGND VGND VPWR VPWR _3764_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_60_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5500_ hold150/X hold241/X _5501_/S VGND VGND VPWR VPWR _7065_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6480_ _6668_/CLK _6480_/D _6435_/X VGND VGND VPWR VPWR _6480_/Q sky130_fd_sc_hd__dfrtp_2
X_3692_ _6640_/Q _4172_/A _3551_/Y wire835/X _3669_/X VGND VGND VPWR VPWR _3693_/D
+ sky130_fd_sc_hd__a221o_2
X_5431_ _5602_/A0 hold283/X _5431_/S VGND VGND VPWR VPWR _5431_/X sky130_fd_sc_hd__mux2_1
Xoutput314 wire806/X VGND VGND VPWR VPWR spimemio_flash_io1_di sky130_fd_sc_hd__buf_8
Xoutput325 _6555_/Q VGND VGND VPWR VPWR wb_dat_o[16] sky130_fd_sc_hd__buf_8
X_5362_ _5578_/A0 _6942_/Q _5368_/S VGND VGND VPWR VPWR _6942_/D sky130_fd_sc_hd__mux2_1
Xoutput303 _6822_/Q VGND VGND VPWR VPWR pwr_ctrl_out[2] sky130_fd_sc_hd__buf_8
Xoutput336 _7205_/Q VGND VGND VPWR VPWR wb_dat_o[26] sky130_fd_sc_hd__buf_8
Xoutput347 _6588_/Q VGND VGND VPWR VPWR wb_dat_o[7] sky130_fd_sc_hd__buf_8
X_7101_ _7103_/CLK _7101_/D fanout861/X VGND VGND VPWR VPWR _7101_/Q sky130_fd_sc_hd__dfstp_2
X_4313_ _6760_/Q _6409_/A0 _4315_/S VGND VGND VPWR VPWR _6760_/D sky130_fd_sc_hd__mux2_1
X_5293_ hold150/X hold245/X _5296_/S VGND VGND VPWR VPWR _6881_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7032_ _7095_/CLK _7032_/D fanout865/X VGND VGND VPWR VPWR _7032_/Q sky130_fd_sc_hd__dfrtp_2
X_4244_ _5248_/A0 hold214/X hold32/X VGND VGND VPWR VPWR _4244_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4175_ _6641_/Q _6409_/A0 _4177_/S VGND VGND VPWR VPWR _6641_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6816_ _7103_/CLK _6816_/D fanout861/X VGND VGND VPWR VPWR _6816_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6747_ _6747_/CLK _6747_/D _6420_/A VGND VGND VPWR VPWR _6747_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire408 _3352_/Y VGND VGND VPWR VPWR _5306_/A sky130_fd_sc_hd__buf_8
X_3959_ _6474_/Q _3959_/B VGND VGND VPWR VPWR _3960_/A sky130_fd_sc_hd__nand2b_4
XFILLER_164_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6678_ _7194_/CLK _6678_/D fanout866/X VGND VGND VPWR VPWR _6678_/Q sky130_fd_sc_hd__dfrtp_2
X_5629_ _7163_/Q _5629_/B VGND VGND VPWR VPWR _5633_/B sky130_fd_sc_hd__or2_2
XFILLER_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length540 _6904_/Q VGND VGND VPWR VPWR _3581_/A1 sky130_fd_sc_hd__buf_6
XFILLER_41_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length595 _6021_/B VGND VGND VPWR VPWR _6295_/B1 sky130_fd_sc_hd__buf_6
Xmax_length584 _6017_/Y VGND VGND VPWR VPWR _6023_/D sky130_fd_sc_hd__buf_6
XFILLER_69_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5980_ _6789_/Q _5980_/A2 wire675/X wire569/X _5979_/X VGND VGND VPWR VPWR _5981_/D
+ sky130_fd_sc_hd__a221o_1
X_4931_ _4735_/B _4494_/Y _4957_/A _4930_/X VGND VGND VPWR VPWR _4932_/C sky130_fd_sc_hd__a211o_4
XFILLER_80_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4862_ _4735_/B _4486_/B _4554_/A _4554_/X VGND VGND VPWR VPWR _5084_/A sky130_fd_sc_hd__a31o_4
XFILLER_60_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6601_ _6950_/CLK _6601_/D fanout874/X VGND VGND VPWR VPWR _6601_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_60_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3813_ hold40/A hold59/A _6477_/Q VGND VGND VPWR VPWR _3830_/B sky130_fd_sc_hd__and3_1
XFILLER_193_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_15 _6519_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 _6874_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4793_ _4793_/A VGND VGND VPWR VPWR _4793_/Y sky130_fd_sc_hd__inv_2
XANTENNA_37 hold97/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 _3522_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_59 _3687_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3744_ _6488_/Q _3978_/A _3730_/X _5223_/A VGND VGND VPWR VPWR _3744_/X sky130_fd_sc_hd__a22o_1
X_6532_ _7225_/CLK _6532_/D fanout856/X VGND VGND VPWR VPWR _6532_/Q sky130_fd_sc_hd__dfrtp_2
X_6463_ _3938_/A1 _6463_/D _6418_/X VGND VGND VPWR VPWR _6463_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_146_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3675_ _7126_/Q hold88/A _4232_/S input47/X VGND VGND VPWR VPWR _3675_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5414_ _5414_/A _5576_/B VGND VGND VPWR VPWR _5422_/S sky130_fd_sc_hd__nand2_8
X_6394_ _6393_/X hold23/A _6400_/S VGND VGND VPWR VPWR _7216_/D sky130_fd_sc_hd__mux2_1
X_5345_ _5498_/A0 hold744/X _5350_/S VGND VGND VPWR VPWR _6927_/D sky130_fd_sc_hd__mux2_1
Xoutput177 _3229_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[11] sky130_fd_sc_hd__buf_8
Xoutput199 _3209_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[31] sky130_fd_sc_hd__buf_8
Xoutput188 _3219_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[21] sky130_fd_sc_hd__buf_8
X_5276_ wire758/X _6866_/Q _5278_/S VGND VGND VPWR VPWR _5276_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7015_ _7134_/CLK _7015_/D fanout864/X VGND VGND VPWR VPWR _7015_/Q sky130_fd_sc_hd__dfrtp_2
X_4227_ hold612/X _4226_/X _4235_/S VGND VGND VPWR VPWR _4227_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4158_ hold255/X hold83/X _4159_/S VGND VGND VPWR VPWR _6627_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4089_ _6568_/Q wire350/X _4096_/S VGND VGND VPWR VPWR _6568_/D sky130_fd_sc_hd__mux2_1
XFILLER_15_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput13 mask_rev_in[18] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__clkbuf_4
Xinput46 mgmt_gpio_in[19] VGND VGND VPWR VPWR wire908/A sky130_fd_sc_hd__clkbuf_4
XFILLER_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput35 mask_rev_in[9] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__clkbuf_4
Xinput24 mask_rev_in[28] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__clkbuf_4
Xhold808 _6669_/Q VGND VGND VPWR VPWR hold808/X sky130_fd_sc_hd__bufbuf_16
Xwire794 wire794/A VGND VGND VPWR VPWR wire794/X sky130_fd_sc_hd__buf_6
Xinput57 mgmt_gpio_in[29] VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__clkbuf_4
XFILLER_143_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput68 mgmt_gpio_in[5] VGND VGND VPWR VPWR wire895/A sky130_fd_sc_hd__buf_6
Xinput79 spi_enabled VGND VGND VPWR VPWR _3970_/B sky130_fd_sc_hd__buf_4
Xhold819 _7011_/Q VGND VGND VPWR VPWR hold819/X sky130_fd_sc_hd__bufbuf_16
XFILLER_143_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3460_ _3514_/A hold44/X VGND VGND VPWR VPWR _4328_/A sky130_fd_sc_hd__nor2_8
XFILLER_170_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3391_ _7027_/Q _3301_/Y _5540_/A _7107_/Q VGND VGND VPWR VPWR _3391_/X sky130_fd_sc_hd__a22o_1
X_5130_ _5130_/A _5130_/B _5130_/C _4970_/X VGND VGND VPWR VPWR _5175_/B sky130_fd_sc_hd__or4b_4
XFILLER_111_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5061_ _5132_/A _5133_/A VGND VGND VPWR VPWR _5061_/Y sky130_fd_sc_hd__nor2_1
X_4012_ hold350/X _4011_/X _4024_/S VGND VGND VPWR VPWR _4012_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5963_ _6628_/Q _5963_/B VGND VGND VPWR VPWR _5963_/X sky130_fd_sc_hd__or2_1
XFILLER_53_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4914_ _5003_/B _4838_/X _4913_/X _4567_/X _5156_/A VGND VGND VPWR VPWR _4914_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_52_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5894_ _6530_/Q _5722_/B _5883_/X _5893_/X _6308_/S VGND VGND VPWR VPWR _5894_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4845_ _4845_/A _4845_/B VGND VGND VPWR VPWR _4863_/B sky130_fd_sc_hd__and2_2
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4776_ _4776_/A _4776_/B VGND VGND VPWR VPWR _5165_/B sky130_fd_sc_hd__nor2_2
XFILLER_148_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6515_ _7096_/CLK _6515_/D fanout882/X VGND VGND VPWR VPWR _6515_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_146_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3727_ _3727_/A _3727_/B _3727_/C _3727_/D VGND VGND VPWR VPWR _3727_/X sky130_fd_sc_hd__or4_4
XFILLER_180_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3658_ _7111_/Q hold97/A _5261_/A _6855_/Q _3657_/X VGND VGND VPWR VPWR _3664_/C
+ sky130_fd_sc_hd__a221o_4
X_6446_ _6446_/A _6447_/B VGND VGND VPWR VPWR _6446_/X sky130_fd_sc_hd__and2_1
X_6377_ _4236_/B _6377_/A2 _6377_/B1 _4236_/A VGND VGND VPWR VPWR _6377_/X sky130_fd_sc_hd__a22o_1
X_3589_ input23/X _3302_/Y _5459_/A _7032_/Q _3553_/X VGND VGND VPWR VPWR _3593_/A
+ sky130_fd_sc_hd__a221o_2
X_5328_ _5598_/A0 hold568/X _5332_/S VGND VGND VPWR VPWR _6912_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5259_ _5259_/A0 hold631/X _5260_/S VGND VGND VPWR VPWR _5259_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4630_ _5079_/B VGND VGND VPWR VPWR _4630_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4561_ _4562_/B VGND VGND VPWR VPWR _4561_/Y sky130_fd_sc_hd__inv_2
X_6300_ _6542_/Q wire592/X wire590/X _6565_/Q _6299_/X VGND VGND VPWR VPWR _6305_/B
+ sky130_fd_sc_hd__a221o_1
Xhold627 _4245_/X VGND VGND VPWR VPWR _6693_/D sky130_fd_sc_hd__bufbuf_16
X_4492_ _4566_/A _4663_/B VGND VGND VPWR VPWR _4687_/A sky130_fd_sc_hd__or2_4
Xwire591 _6025_/B VGND VGND VPWR VPWR wire591/X sky130_fd_sc_hd__buf_8
X_3512_ _7081_/Q _3638_/B1 _4142_/A _6618_/Q VGND VGND VPWR VPWR _3512_/X sky130_fd_sc_hd__a22o_1
Xwire580 _6021_/D VGND VGND VPWR VPWR wire580/X sky130_fd_sc_hd__buf_8
XFILLER_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold605 _7023_/Q VGND VGND VPWR VPWR hold605/X sky130_fd_sc_hd__bufbuf_16
Xhold616 _7225_/Q VGND VGND VPWR VPWR hold616/X sky130_fd_sc_hd__bufbuf_16
XFILLER_170_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold638 _6880_/Q VGND VGND VPWR VPWR hold638/X sky130_fd_sc_hd__bufbuf_16
X_6231_ _6231_/A _6231_/B _6231_/C _6231_/D VGND VGND VPWR VPWR _6232_/C sky130_fd_sc_hd__or4_4
X_3443_ wire538/X _3443_/A2 _5513_/A _7082_/Q _3430_/X VGND VGND VPWR VPWR _3451_/B
+ sky130_fd_sc_hd__a221o_1
Xhold649 _7039_/Q VGND VGND VPWR VPWR hold649/X sky130_fd_sc_hd__bufbuf_16
XFILLER_103_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _7082_/Q _6211_/B VGND VGND VPWR VPWR _6162_/X sky130_fd_sc_hd__and2_1
X_5113_ _4871_/A _4989_/A _4995_/A VGND VGND VPWR VPWR _5114_/D sky130_fd_sc_hd__a21oi_1
XFILLER_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3374_ _3543_/A hold87/X VGND VGND VPWR VPWR _3374_/Y sky130_fd_sc_hd__nor2_8
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6093_ _7119_/Q _6252_/B1 wire579/X _7031_/Q _6092_/X VGND VGND VPWR VPWR _6093_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _4745_/A _4756_/B _5050_/C _4757_/B _5043_/X VGND VGND VPWR VPWR _5108_/A
+ sky130_fd_sc_hd__o221ai_2
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6995_ _7072_/CLK _6995_/D fanout870/X VGND VGND VPWR VPWR _6995_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5946_ _6776_/Q wire694/X wire660/X _6607_/Q _5945_/X VGND VGND VPWR VPWR _5953_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5877_ _6748_/Q _5979_/A2 wire667/X _6535_/Q VGND VGND VPWR VPWR _5877_/X sky130_fd_sc_hd__a22o_1
X_4828_ _4687_/A _4898_/B _5147_/B VGND VGND VPWR VPWR _4828_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_139_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4759_ _5062_/B _4739_/X _4753_/X _4733_/X VGND VGND VPWR VPWR _4759_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6429_ _6446_/A _6447_/B VGND VGND VPWR VPWR _6429_/X sky130_fd_sc_hd__and2_1
XFILLER_108_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2 hold2/A VGND VGND VPWR VPWR hold2/X sky130_fd_sc_hd__bufbuf_16
XFILLER_94_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_618 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5800_ _6937_/Q wire659/X _5799_/X wire671/X VGND VGND VPWR VPWR _5800_/X sky130_fd_sc_hd__a22o_1
X_6780_ _7218_/CLK _6780_/D wire915/A VGND VGND VPWR VPWR _6780_/Q sky130_fd_sc_hd__dfrtp_2
X_3992_ _6494_/Q _5547_/A0 _3994_/S VGND VGND VPWR VPWR _6494_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5731_ _7102_/Q _5973_/A2 wire692/X _6990_/Q _5730_/X VGND VGND VPWR VPWR _5734_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_188_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5662_ _6832_/Q _5626_/A _6680_/Q _3918_/X _5661_/X VGND VGND VPWR VPWR _7175_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4613_ _4997_/A _4617_/B VGND VGND VPWR VPWR _4950_/A sky130_fd_sc_hd__nor2_2
X_5593_ _5602_/A0 hold357/X _5593_/S VGND VGND VPWR VPWR _5593_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4544_ _4987_/B _4586_/B _4542_/X _4543_/X VGND VGND VPWR VPWR _4546_/C sky130_fd_sc_hd__a211o_1
XFILLER_144_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold402 _6580_/Q VGND VGND VPWR VPWR hold402/X sky130_fd_sc_hd__bufbuf_16
Xhold435 _7146_/Q VGND VGND VPWR VPWR hold435/X sky130_fd_sc_hd__bufbuf_16
XFILLER_144_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold413 _7139_/Q VGND VGND VPWR VPWR hold413/X sky130_fd_sc_hd__bufbuf_16
Xhold424 _6848_/Q VGND VGND VPWR VPWR hold424/X sky130_fd_sc_hd__bufbuf_16
Xhold468 _6519_/Q VGND VGND VPWR VPWR hold468/X sky130_fd_sc_hd__bufbuf_16
Xhold446 _6600_/Q VGND VGND VPWR VPWR hold446/X sky130_fd_sc_hd__bufbuf_16
Xhold457 _6978_/Q VGND VGND VPWR VPWR hold457/X sky130_fd_sc_hd__bufbuf_16
X_4475_ _4558_/B _4584_/A VGND VGND VPWR VPWR _4634_/B sky130_fd_sc_hd__nor2_8
XFILLER_89_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6214_ _7020_/Q wire575/X _6335_/B _7044_/Q _6211_/X VGND VGND VPWR VPWR _6219_/B
+ sky130_fd_sc_hd__a221o_1
X_3426_ _7058_/Q wire438/X _5549_/A _7114_/Q VGND VGND VPWR VPWR _3426_/X sky130_fd_sc_hd__a22o_2
Xhold479 _4040_/X VGND VGND VPWR VPWR _6527_/D sky130_fd_sc_hd__bufbuf_16
X_7194_ _7194_/CLK _7194_/D fanout868/A VGND VGND VPWR VPWR _7194_/Q sky130_fd_sc_hd__dfrtp_4
X_6145_ _7113_/Q wire650/X _6295_/B1 _7153_/Q VGND VGND VPWR VPWR _6145_/X sky130_fd_sc_hd__a22o_1
XFILLER_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3357_ _7108_/Q _5540_/A _3683_/B1 wire531/X _3354_/X VGND VGND VPWR VPWR _3377_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ _6958_/Q wire624/X wire613/X _7054_/Q VGND VGND VPWR VPWR _6076_/X sky130_fd_sc_hd__a22o_1
XFILLER_112_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5027_ _4758_/C _4684_/Y _4941_/B _4653_/Y _4386_/Y VGND VGND VPWR VPWR _5163_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3288_ hold94/X hold61/X VGND VGND VPWR VPWR hold95/A sky130_fd_sc_hd__nand2b_4
XFILLER_173_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_308 input72/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_319 wire739/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6978_ _7154_/CLK _6978_/D fanout884/X VGND VGND VPWR VPWR _6978_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_179_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5929_ _6646_/Q wire690/X wire653/X _6651_/Q _5928_/X VGND VGND VPWR VPWR _5937_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_186_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4260_ _6716_/Q hold83/A _4261_/S VGND VGND VPWR VPWR hold78/A sky130_fd_sc_hd__mux2_1
XFILLER_140_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3211_ _3211_/A VGND VGND VPWR VPWR _3211_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4191_ _6407_/A0 hold780/X _4195_/S VGND VGND VPWR VPWR _6654_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6901_ _6969_/CLK _6901_/D fanout880/X VGND VGND VPWR VPWR _6901_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_63_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6832_ _7107_/CLK _6832_/D fanout867/X VGND VGND VPWR VPWR _6832_/Q sky130_fd_sc_hd__dfrtp_2
X_6763_ _7223_/CLK _6763_/D fanout850/X VGND VGND VPWR VPWR _6763_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3975_ hold68/X _3975_/B VGND VGND VPWR VPWR hold69/A sky130_fd_sc_hd__nand2b_2
X_6694_ _7145_/CLK _6694_/D fanout881/X VGND VGND VPWR VPWR _6694_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5714_ _6981_/Q wire671/X wire656/X _6941_/Q _5697_/X VGND VGND VPWR VPWR _5714_/X
+ sky130_fd_sc_hd__a221o_1
X_5645_ _5648_/B _6035_/A VGND VGND VPWR VPWR _5645_/Y sky130_fd_sc_hd__nand2_1
XFILLER_176_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold210 _6943_/Q VGND VGND VPWR VPWR hold210/X sky130_fd_sc_hd__bufbuf_16
X_5576_ _5576_/A _5576_/B VGND VGND VPWR VPWR _5584_/S sky130_fd_sc_hd__nand2_4
XFILLER_191_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold232 _6696_/Q VGND VGND VPWR VPWR hold232/X sky130_fd_sc_hd__bufbuf_16
Xhold221 _7131_/Q VGND VGND VPWR VPWR hold221/X sky130_fd_sc_hd__bufbuf_16
Xhold243 _6841_/Q VGND VGND VPWR VPWR hold243/X sky130_fd_sc_hd__bufbuf_16
XFILLER_144_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4527_ _4986_/A _4648_/B VGND VGND VPWR VPWR _4805_/A sky130_fd_sc_hd__nor2_1
X_4458_ _4558_/B _4818_/B VGND VGND VPWR VPWR _4617_/B sky130_fd_sc_hd__or2_4
Xhold276 _6863_/Q VGND VGND VPWR VPWR hold276/X sky130_fd_sc_hd__bufbuf_16
Xhold287 _6959_/Q VGND VGND VPWR VPWR hold287/X sky130_fd_sc_hd__bufbuf_16
Xhold265 _4023_/X VGND VGND VPWR VPWR hold265/X sky130_fd_sc_hd__bufbuf_16
XFILLER_132_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold254 _4164_/X VGND VGND VPWR VPWR _6632_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_104_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold298 _6521_/Q VGND VGND VPWR VPWR hold298/X sky130_fd_sc_hd__bufbuf_16
XFILLER_132_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout723 _5585_/B VGND VGND VPWR VPWR _5594_/B sky130_fd_sc_hd__bufbuf_16
X_3409_ wire542/X _3582_/B1 _5227_/A _3385_/X VGND VGND VPWR VPWR _3409_/X sky130_fd_sc_hd__a22o_2
X_7177_ _7190_/CLK _7177_/D fanout869/X VGND VGND VPWR VPWR _7177_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_49_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6128_ wire550/X wire593/X wire591/X _3235_/A _6127_/X VGND VGND VPWR VPWR _6131_/C
+ sky130_fd_sc_hd__a221o_1
X_4389_ _4507_/A _4851_/B VGND VGND VPWR VPWR _4405_/B sky130_fd_sc_hd__nand2_8
XFILLER_131_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout767 wire770/A VGND VGND VPWR VPWR _5249_/A0 sky130_fd_sc_hd__buf_8
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout789 wire796/X VGND VGND VPWR VPWR wire790/A sky130_fd_sc_hd__buf_6
XFILLER_85_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6059_ _6059_/A _6059_/B _6059_/C _6059_/D VGND VGND VPWR VPWR _6059_/X sky130_fd_sc_hd__or4_4
XFILLER_73_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_116 _6738_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_105 _6157_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_138 mgmt_gpio_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_149 porb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_127 mask_rev_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length744 wire746/X VGND VGND VPWR VPWR _5547_/A0 sky130_fd_sc_hd__buf_6
XFILLER_182_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3760_ _7117_/Q _5558_/A _5245_/A input61/X _3741_/X VGND VGND VPWR VPWR _3764_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_192_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5430_ _5601_/A0 hold223/X _5431_/S VGND VGND VPWR VPWR _5430_/X sky130_fd_sc_hd__mux2_1
X_3691_ wire498/X wire430/X _4130_/A _6605_/Q _3671_/X VGND VGND VPWR VPWR _3693_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput315 _7228_/X VGND VGND VPWR VPWR spimemio_flash_io2_di sky130_fd_sc_hd__buf_8
XFILLER_161_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5361_ hold465/X _6941_/Q _5368_/S VGND VGND VPWR VPWR _6941_/D sky130_fd_sc_hd__mux2_1
Xoutput326 _6556_/Q VGND VGND VPWR VPWR wb_dat_o[17] sky130_fd_sc_hd__buf_8
Xoutput304 _6823_/Q VGND VGND VPWR VPWR pwr_ctrl_out[3] sky130_fd_sc_hd__buf_8
X_5292_ _5598_/A0 hold638/X _5296_/S VGND VGND VPWR VPWR _6880_/D sky130_fd_sc_hd__mux2_1
Xoutput337 _7206_/Q VGND VGND VPWR VPWR wb_dat_o[27] sky130_fd_sc_hd__buf_8
XFILLER_114_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput348 _6568_/Q VGND VGND VPWR VPWR wb_dat_o[8] sky130_fd_sc_hd__buf_8
X_4312_ hold690/X _6408_/A0 _4315_/S VGND VGND VPWR VPWR _6759_/D sky130_fd_sc_hd__mux2_1
X_7100_ _7132_/CLK _7100_/D fanout863/X VGND VGND VPWR VPWR _7100_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_141_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4243_ hold38/A hold841/X hold32/X VGND VGND VPWR VPWR hold33/A sky130_fd_sc_hd__mux2_1
X_7031_ _7118_/CLK _7031_/D fanout869/X VGND VGND VPWR VPWR _7031_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_59_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4174_ hold745/X _6408_/A0 _4177_/S VGND VGND VPWR VPWR _6640_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6815_ _6815_/CLK _6815_/D fanout861/X VGND VGND VPWR VPWR _6815_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_23_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6746_ _6951_/CLK _6746_/D _6420_/A VGND VGND VPWR VPWR _6746_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_51_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3958_ _6473_/Q _6446_/A VGND VGND VPWR VPWR _3958_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3889_ _4368_/A _4722_/A VGND VGND VPWR VPWR _4346_/S sky130_fd_sc_hd__and2_2
XFILLER_137_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6677_ _7194_/CLK _6677_/D fanout868/X VGND VGND VPWR VPWR _6677_/Q sky130_fd_sc_hd__dfstp_4
X_5628_ _5663_/B _5702_/B _5705_/B _7162_/Q _5621_/X VGND VGND VPWR VPWR _7162_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_164_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5559_ _5595_/A0 _7117_/Q _5564_/S VGND VGND VPWR VPWR _7117_/D sky130_fd_sc_hd__mux2_1
X_7229_ _7229_/A VGND VGND VPWR VPWR _7229_/X sky130_fd_sc_hd__buf_2
XFILLER_74_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_1_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A VGND VGND VPWR VPWR _7208_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_54_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire910 wire910/A VGND VGND VPWR VPWR _3202_/A sky130_fd_sc_hd__buf_6
XFILLER_167_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length574 _6036_/Y VGND VGND VPWR VPWR _6139_/A2 sky130_fd_sc_hd__buf_6
XFILLER_157_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4930_ _4426_/A _4707_/A _4930_/C _4930_/D VGND VGND VPWR VPWR _4930_/X sky130_fd_sc_hd__and4bb_2
XFILLER_64_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4861_ _4376_/Y _4845_/B _5136_/C _4859_/X _4860_/X VGND VGND VPWR VPWR _4863_/C
+ sky130_fd_sc_hd__a2111o_1
XFILLER_33_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6600_ _6950_/CLK _6600_/D fanout874/X VGND VGND VPWR VPWR _6600_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_60_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3812_ _6664_/Q _3812_/B VGND VGND VPWR VPWR _3840_/S sky130_fd_sc_hd__nand2b_4
XFILLER_33_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_27 _5358_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_16 _6519_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4792_ _4775_/A _4776_/A _4776_/B _5147_/B _4745_/A VGND VGND VPWR VPWR _4793_/A
+ sky130_fd_sc_hd__o32a_1
XANTENNA_38 _3377_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_49 _3533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3743_ _7037_/Q _3334_/Y _5216_/A _6819_/Q VGND VGND VPWR VPWR _3743_/X sky130_fd_sc_hd__a22o_1
X_6531_ _7225_/CLK _6531_/D fanout856/X VGND VGND VPWR VPWR _6531_/Q sky130_fd_sc_hd__dfrtp_2
X_6462_ _3938_/A1 _6462_/D _6417_/X VGND VGND VPWR VPWR _6462_/Q sky130_fd_sc_hd__dfrtp_2
X_3674_ _7150_/Q hold65/A _5245_/A input62/X VGND VGND VPWR VPWR _3674_/X sky130_fd_sc_hd__a22o_4
XFILLER_146_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6393_ _4236_/C _6393_/A2 _6393_/B1 _4238_/B _6392_/X VGND VGND VPWR VPWR _6393_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5413_ hold582/X wire739/A _5413_/S VGND VGND VPWR VPWR _5413_/X sky130_fd_sc_hd__mux2_1
X_5344_ hold38/X hold249/X _5350_/S VGND VGND VPWR VPWR _6926_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput189 _3218_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[22] sky130_fd_sc_hd__buf_8
X_5275_ hold150/X hold240/X _5278_/S VGND VGND VPWR VPWR _6865_/D sky130_fd_sc_hd__mux2_1
Xoutput178 _3228_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[12] sky130_fd_sc_hd__buf_8
XFILLER_99_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7014_ _7134_/CLK _7014_/D fanout864/X VGND VGND VPWR VPWR _7014_/Q sky130_fd_sc_hd__dfstp_2
X_4226_ hold424/X wire770/X _4234_/S VGND VGND VPWR VPWR _4226_/X sky130_fd_sc_hd__mux2_1
X_4157_ hold545/X _5336_/A1 _4159_/S VGND VGND VPWR VPWR _6626_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4088_ _6700_/Q _6362_/B VGND VGND VPWR VPWR _4096_/S sky130_fd_sc_hd__and2_4
XFILLER_55_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6729_ _6771_/CLK _6729_/D fanout854/X VGND VGND VPWR VPWR _6729_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_164_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_67_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7129_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_120_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput14 mask_rev_in[19] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__clkbuf_4
Xinput36 mgmt_gpio_in[0] VGND VGND VPWR VPWR wire911/A sky130_fd_sc_hd__buf_6
Xinput25 mask_rev_in[29] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__clkbuf_4
Xhold809 _4204_/X VGND VGND VPWR VPWR _6669_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_183_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire773 wire773/A VGND VGND VPWR VPWR wire773/X sky130_fd_sc_hd__buf_6
XFILLER_128_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput69 mgmt_gpio_in[6] VGND VGND VPWR VPWR input69/X sky130_fd_sc_hd__clkbuf_4
Xinput47 mgmt_gpio_in[1] VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__clkbuf_4
Xinput58 mgmt_gpio_in[2] VGND VGND VPWR VPWR wire904/A sky130_fd_sc_hd__buf_6
XFILLER_182_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3390_ _6891_/Q _5297_/A _5405_/A _6987_/Q VGND VGND VPWR VPWR _3390_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5060_ _5060_/A _5060_/B VGND VGND VPWR VPWR _5133_/A sky130_fd_sc_hd__or2_2
XFILLER_69_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4011_ _6523_/Q hold38/A _4021_/S VGND VGND VPWR VPWR _4011_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5962_ _7187_/Q _6309_/S _5961_/X VGND VGND VPWR VPWR _7187_/D sky130_fd_sc_hd__o21a_1
X_4913_ _4978_/B _4913_/B _4913_/C _5069_/C VGND VGND VPWR VPWR _4913_/X sky130_fd_sc_hd__or4_1
X_5893_ _5893_/A _5893_/B _5893_/C _5893_/D VGND VGND VPWR VPWR _5893_/X sky130_fd_sc_hd__or4_4
XFILLER_33_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4844_ _4844_/A _4844_/B VGND VGND VPWR VPWR _5086_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4775_ _4775_/A _4927_/B VGND VGND VPWR VPWR _5099_/B sky130_fd_sc_hd__nor2_1
X_6514_ _7096_/CLK _6514_/D fanout882/X VGND VGND VPWR VPWR _6514_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_119_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3726_ _3726_/A _3726_/B _3726_/C _3726_/D VGND VGND VPWR VPWR _3727_/D sky130_fd_sc_hd__or4_1
XFILLER_174_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3657_ _7063_/Q _3657_/A2 _5531_/A wire486/X VGND VGND VPWR VPWR _3657_/X sky130_fd_sc_hd__a22o_1
X_6445_ _6447_/A _6447_/B VGND VGND VPWR VPWR _6445_/X sky130_fd_sc_hd__and2_1
X_6376_ _6376_/A _6376_/B _6376_/C _6374_/X VGND VGND VPWR VPWR _6400_/S sky130_fd_sc_hd__or4b_4
XFILLER_164_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3588_ _3588_/A _3588_/B _3588_/C _3588_/D VGND VGND VPWR VPWR _3606_/A sky130_fd_sc_hd__or4_4
X_5327_ _5498_/A0 hold715/X _5332_/S VGND VGND VPWR VPWR _6911_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5258_ _5519_/A0 hold644/X _5260_/S VGND VGND VPWR VPWR _5258_/X sky130_fd_sc_hd__mux2_1
X_4209_ hold626/X _5598_/A0 _4209_/S VGND VGND VPWR VPWR _4209_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5189_ _6410_/A0 hold678/X _5190_/S VGND VGND VPWR VPWR _6788_/D sky130_fd_sc_hd__mux2_1
XFILLER_29_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4560_ _4812_/A _4697_/A VGND VGND VPWR VPWR _4562_/B sky130_fd_sc_hd__or2_4
XFILLER_128_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold617 _6517_/Q VGND VGND VPWR VPWR hold617/X sky130_fd_sc_hd__bufbuf_16
Xwire570 _6610_/Q VGND VGND VPWR VPWR wire570/X sky130_fd_sc_hd__buf_6
X_4491_ _5004_/A _4659_/A VGND VGND VPWR VPWR _4648_/B sky130_fd_sc_hd__nand2_8
Xwire581 _6021_/D VGND VGND VPWR VPWR wire581/X sky130_fd_sc_hd__buf_8
Xwire592 _6023_/C VGND VGND VPWR VPWR wire592/X sky130_fd_sc_hd__buf_8
X_3511_ _3540_/A _3528_/B VGND VGND VPWR VPWR _4142_/A sky130_fd_sc_hd__nor2_8
XFILLER_7_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold606 _5453_/X VGND VGND VPWR VPWR _7023_/D sky130_fd_sc_hd__bufbuf_16
X_3442_ _7146_/Q _5585_/A _5369_/A _6954_/Q _3441_/X VGND VGND VPWR VPWR _3451_/A
+ sky130_fd_sc_hd__a221o_4
X_6230_ wire525/X wire641/X wire639/X _6884_/Q _6229_/X VGND VGND VPWR VPWR _6231_/D
+ sky130_fd_sc_hd__a221o_1
Xhold628 _6920_/Q VGND VGND VPWR VPWR hold628/X sky130_fd_sc_hd__bufbuf_16
Xhold639 _6732_/Q VGND VGND VPWR VPWR hold639/X sky130_fd_sc_hd__bufbuf_16
X_6161_ _6978_/Q wire641/X wire639/X _6882_/Q VGND VGND VPWR VPWR _6161_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3373_ _7124_/Q wire446/A _3739_/B1 _6988_/Q VGND VGND VPWR VPWR _3373_/X sky130_fd_sc_hd__a22o_1
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5112_ _6782_/Q _5156_/A _5038_/Y _5111_/X _5103_/X VGND VGND VPWR VPWR _5112_/X
+ sky130_fd_sc_hd__a221o_2
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ _6999_/Q wire604/X _6140_/B1 _6919_/Q VGND VGND VPWR VPWR _6092_/X sky130_fd_sc_hd__a22o_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _4818_/A _4566_/A _4756_/B _4893_/B VGND VGND VPWR VPWR _5043_/X sky130_fd_sc_hd__o31a_1
XFILLER_84_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_wbbd_sck _7219_/Q VGND VGND VPWR VPWR clkbuf_0_wbbd_sck/X sky130_fd_sc_hd__clkbuf_8
X_6994_ _6994_/CLK _6994_/D fanout870/X VGND VGND VPWR VPWR _6994_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_80_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5945_ _6731_/Q wire710/X wire689/X _6642_/Q VGND VGND VPWR VPWR _5945_/X sky130_fd_sc_hd__a22o_1
XFILLER_40_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5876_ _6785_/Q _5926_/A2 wire656/X _6609_/Q _5875_/X VGND VGND VPWR VPWR _5883_/A
+ sky130_fd_sc_hd__a221o_4
XFILLER_80_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4827_ _4827_/A _5013_/B _5047_/C _4826_/X VGND VGND VPWR VPWR _4834_/B sky130_fd_sc_hd__or4b_2
XFILLER_193_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4758_ _4758_/A _4758_/B _4758_/C VGND VGND VPWR VPWR _5105_/A sky130_fd_sc_hd__and3_1
XFILLER_147_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3709_ _3709_/A _3709_/B _3709_/C _3709_/D VGND VGND VPWR VPWR _3709_/X sky130_fd_sc_hd__or4_4
XFILLER_146_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4689_ _4717_/B VGND VGND VPWR VPWR _4689_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_108_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6428_ _6446_/A _6447_/B VGND VGND VPWR VPWR _6428_/X sky130_fd_sc_hd__and2_1
XFILLER_88_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6359_ _7201_/Q _6309_/S _6357_/X _6358_/X VGND VGND VPWR VPWR _7201_/D sky130_fd_sc_hd__o22a_1
XFILLER_102_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold3 hold3/A VGND VGND VPWR VPWR hold3/X sky130_fd_sc_hd__bufbuf_16
XFILLER_121_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3991_ hold196/X _7217_/Q _3991_/S VGND VGND VPWR VPWR _3991_/X sky130_fd_sc_hd__mux2_4
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5730_ wire546/X wire706/X wire686/X _7030_/Q VGND VGND VPWR VPWR _5730_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5661_ _6677_/Q _5659_/C _7175_/Q VGND VGND VPWR VPWR _5661_/X sky130_fd_sc_hd__a21o_1
XFILLER_30_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4612_ _4612_/A _4612_/B _4612_/C _4612_/D VGND VGND VPWR VPWR _4615_/B sky130_fd_sc_hd__and4_2
XFILLER_163_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5592_ hold57/X hold849/X _5593_/S VGND VGND VPWR VPWR hold58/A sky130_fd_sc_hd__mux2_1
XFILLER_175_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4543_ _4772_/A _4409_/Y _4412_/Y _5116_/A VGND VGND VPWR VPWR _4543_/X sky130_fd_sc_hd__a211o_1
XFILLER_144_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold436 _6938_/Q VGND VGND VPWR VPWR hold436/X sky130_fd_sc_hd__bufbuf_16
XFILLER_143_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold403 _7033_/Q VGND VGND VPWR VPWR hold403/X sky130_fd_sc_hd__bufbuf_16
Xhold425 _5256_/X VGND VGND VPWR VPWR _6848_/D sky130_fd_sc_hd__bufbuf_16
Xhold414 _6648_/Q VGND VGND VPWR VPWR hold414/X sky130_fd_sc_hd__bufbuf_16
Xhold458 _5402_/X VGND VGND VPWR VPWR _6978_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_131_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4474_ _4949_/A _4956_/A VGND VGND VPWR VPWR _4603_/B sky130_fd_sc_hd__nand2_8
Xhold447 _6637_/Q VGND VGND VPWR VPWR hold447/X sky130_fd_sc_hd__bufbuf_16
Xhold469 _6769_/Q VGND VGND VPWR VPWR hold469/X sky130_fd_sc_hd__bufbuf_16
X_6213_ _7028_/Q wire589/X wire615/X _7092_/Q _6212_/X VGND VGND VPWR VPWR _6219_/A
+ sky130_fd_sc_hd__a221o_2
Xfanout916 _4665_/A VGND VGND VPWR VPWR _4707_/B sky130_fd_sc_hd__buf_8
XFILLER_131_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3425_ wire533/X _3683_/B1 _3425_/B1 wire547/X VGND VGND VPWR VPWR _3425_/X sky130_fd_sc_hd__a22o_1
X_7193_ _7196_/CLK _7193_/D fanout870/X VGND VGND VPWR VPWR _7193_/Q sky130_fd_sc_hd__dfrtp_4
X_6144_ _6144_/A _6144_/B _6144_/C _6144_/D VGND VGND VPWR VPWR _6144_/X sky130_fd_sc_hd__or4_4
X_3356_ _3540_/A hold87/X VGND VGND VPWR VPWR _3356_/Y sky130_fd_sc_hd__nor2_8
XFILLER_58_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6075_ _6902_/Q wire600/X wire645/X _6934_/Q _6074_/X VGND VGND VPWR VPWR _6082_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_85_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3287_ input33/X _3283_/Y _5522_/A _7092_/Q VGND VGND VPWR VPWR _3287_/X sky130_fd_sc_hd__a22o_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5026_ _5164_/A _4990_/A _4926_/X _5025_/X VGND VGND VPWR VPWR _5098_/B sky130_fd_sc_hd__o211ai_4
XFILLER_100_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_309 _3957_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6977_ _6980_/CLK _6977_/D fanout889/X VGND VGND VPWR VPWR _6977_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5928_ _6636_/Q _5973_/A2 wire694/X _6775_/Q VGND VGND VPWR VPWR _5928_/X sky130_fd_sc_hd__a22o_1
XFILLER_53_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5859_ _6916_/Q _5680_/X _5689_/X _6908_/Q VGND VGND VPWR VPWR _5859_/X sky130_fd_sc_hd__a22o_1
XFILLER_154_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3210_ _7096_/Q VGND VGND VPWR VPWR _3210_/Y sky130_fd_sc_hd__inv_2
X_4190_ _4190_/A _6406_/B VGND VGND VPWR VPWR _4195_/S sky130_fd_sc_hd__nand2_4
XFILLER_79_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6900_ _7152_/CLK _6900_/D fanout886/X VGND VGND VPWR VPWR _6900_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_63_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6831_ _7091_/CLK _6831_/D fanout866/X VGND VGND VPWR VPWR _6831_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3974_ _6707_/Q _3974_/B VGND VGND VPWR VPWR _6699_/D sky130_fd_sc_hd__and2_1
X_6762_ _6787_/CLK _6762_/D fanout848/X VGND VGND VPWR VPWR _6762_/Q sky130_fd_sc_hd__dfrtp_2
X_6693_ _7122_/CLK _6693_/D fanout887/X VGND VGND VPWR VPWR _6693_/Q sky130_fd_sc_hd__dfrtp_1
X_5713_ _6901_/Q _5689_/X _5710_/X _5712_/X VGND VGND VPWR VPWR _5713_/X sky130_fd_sc_hd__a211o_4
X_5644_ _7169_/Q _7168_/Q VGND VGND VPWR VPWR _6035_/A sky130_fd_sc_hd__and2_4
XFILLER_191_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold200 hold56/X VGND VGND VPWR VPWR hold200/X sky130_fd_sc_hd__bufbuf_16
XFILLER_163_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold211 _5363_/X VGND VGND VPWR VPWR _6943_/D sky130_fd_sc_hd__bufbuf_16
X_5575_ wire739/A hold470/X _5575_/S VGND VGND VPWR VPWR _5575_/X sky130_fd_sc_hd__mux2_1
Xhold244 _5248_/X VGND VGND VPWR VPWR _6841_/D sky130_fd_sc_hd__bufbuf_16
Xhold233 _4248_/X VGND VGND VPWR VPWR _6696_/D sky130_fd_sc_hd__bufbuf_16
Xhold222 _5574_/X VGND VGND VPWR VPWR _7131_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_144_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4526_ _4749_/C _4965_/A VGND VGND VPWR VPWR _4557_/C sky130_fd_sc_hd__nor2_1
XFILLER_2_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4457_ _4558_/B _4818_/B VGND VGND VPWR VPWR _4868_/A sky130_fd_sc_hd__nor2_8
Xhold277 _6876_/Q VGND VGND VPWR VPWR hold277/X sky130_fd_sc_hd__bufbuf_16
XFILLER_171_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold266 _4024_/X VGND VGND VPWR VPWR _6513_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_116_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold255 _6627_/Q VGND VGND VPWR VPWR hold255/X sky130_fd_sc_hd__bufbuf_16
Xhold299 _4033_/X VGND VGND VPWR VPWR _6521_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_172_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold288 _6964_/Q VGND VGND VPWR VPWR hold288/X sky130_fd_sc_hd__bufbuf_16
Xfanout713 _4588_/X VGND VGND VPWR VPWR _4898_/B sky130_fd_sc_hd__buf_8
Xfanout724 fanout724/A VGND VGND VPWR VPWR _5236_/B sky130_fd_sc_hd__buf_8
X_3408_ _6859_/Q _5261_/A _3571_/A2 wire906/X _3407_/X VGND VGND VPWR VPWR _3414_/A
+ sky130_fd_sc_hd__a221o_1
X_7176_ _7190_/CLK _7176_/D fanout869/X VGND VGND VPWR VPWR _7176_/Q sky130_fd_sc_hd__dfrtp_4
X_4388_ _4478_/C _4388_/B VGND VGND VPWR VPWR _4851_/B sky130_fd_sc_hd__and2_4
X_6127_ _6960_/Q wire624/X wire613/X _7056_/Q VGND VGND VPWR VPWR _6127_/X sky130_fd_sc_hd__a22o_1
Xfanout735 _4687_/A VGND VGND VPWR VPWR _5164_/B sky130_fd_sc_hd__buf_8
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout768 wire775/X VGND VGND VPWR VPWR wire770/A sky130_fd_sc_hd__buf_6
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ _3505_/A _5225_/B VGND VGND VPWR VPWR _5459_/A sky130_fd_sc_hd__nor2_8
X_6058_ _6306_/A _6058_/B _6058_/C VGND VGND VPWR VPWR _6059_/D sky130_fd_sc_hd__or3_2
XANTENNA_106 _6178_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5009_ _5004_/A _4469_/Y _4652_/B _4494_/Y VGND VGND VPWR VPWR _5105_/B sky130_fd_sc_hd__a31o_1
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_117 _7133_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_139 mgmt_gpio_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_128 mask_rev_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length734 _4692_/C VGND VGND VPWR VPWR _4758_/B sky130_fd_sc_hd__buf_8
XFILLER_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length778 wire780/X VGND VGND VPWR VPWR _5579_/A0 sky130_fd_sc_hd__buf_6
Xmax_length745 wire746/X VGND VGND VPWR VPWR _5259_/A0 sky130_fd_sc_hd__buf_6
XFILLER_146_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3690_ _6910_/Q wire424/X _5297_/A _6886_/Q _3689_/X VGND VGND VPWR VPWR _3693_/B
+ sky130_fd_sc_hd__a221o_4
XFILLER_118_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput316 _7229_/X VGND VGND VPWR VPWR spimemio_flash_io3_di sky130_fd_sc_hd__buf_8
XFILLER_99_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput305 _3730_/X VGND VGND VPWR VPWR reset sky130_fd_sc_hd__buf_8
X_5360_ _5360_/A _5576_/B VGND VGND VPWR VPWR _5365_/S sky130_fd_sc_hd__nand2_4
X_5291_ _5498_/A0 hold714/X _5296_/S VGND VGND VPWR VPWR _6879_/D sky130_fd_sc_hd__mux2_1
XFILLER_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput338 _7207_/Q VGND VGND VPWR VPWR wb_dat_o[28] sky130_fd_sc_hd__buf_8
XFILLER_126_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput327 _6557_/Q VGND VGND VPWR VPWR wb_dat_o[18] sky130_fd_sc_hd__buf_8
Xoutput349 _6569_/Q VGND VGND VPWR VPWR wb_dat_o[9] sky130_fd_sc_hd__buf_8
X_4311_ hold779/X _6407_/A0 _4315_/S VGND VGND VPWR VPWR _6758_/D sky130_fd_sc_hd__mux2_1
X_4242_ hold465/X hold842/X hold32/X VGND VGND VPWR VPWR _4242_/X sky130_fd_sc_hd__mux2_1
X_7030_ _7140_/CLK _7030_/D fanout862/X VGND VGND VPWR VPWR _7030_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_141_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4173_ hold793/X _6407_/A0 _4177_/S VGND VGND VPWR VPWR _6639_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6814_ _6815_/CLK _6814_/D fanout855/X VGND VGND VPWR VPWR _6814_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_51_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6745_ _6951_/CLK _6745_/D _6420_/A VGND VGND VPWR VPWR _6745_/Q sky130_fd_sc_hd__dfstp_4
X_3957_ wire844/X _3957_/A1 _6473_/Q VGND VGND VPWR VPWR _3957_/X sky130_fd_sc_hd__mux2_1
X_6676_ _7133_/CLK _6676_/D fanout882/X VGND VGND VPWR VPWR _6676_/Q sky130_fd_sc_hd__dfrtp_2
X_3888_ _4350_/C _4350_/D _4349_/A _4349_/B VGND VGND VPWR VPWR _3895_/C sky130_fd_sc_hd__or4_2
XFILLER_176_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5627_ _6677_/Q _5663_/B VGND VGND VPWR VPWR _5635_/B sky130_fd_sc_hd__nand2_4
X_5558_ _5558_/A _5594_/B VGND VGND VPWR VPWR _5564_/S sky130_fd_sc_hd__nand2_8
XFILLER_132_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4509_ _4996_/A _4775_/A VGND VGND VPWR VPWR _4920_/B sky130_fd_sc_hd__nor2_1
XFILLER_3_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5489_ _5597_/A0 hold275/X _5494_/S VGND VGND VPWR VPWR _7055_/D sky130_fd_sc_hd__mux2_1
X_7228_ _7228_/A VGND VGND VPWR VPWR _7228_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_116_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7159_ _7194_/CLK _7159_/D fanout866/X VGND VGND VPWR VPWR _7159_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire900 wire900/A VGND VGND VPWR VPWR wire900/X sky130_fd_sc_hd__buf_6
XFILLER_167_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire911 wire911/A VGND VGND VPWR VPWR _3971_/A sky130_fd_sc_hd__buf_6
XFILLER_182_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length586 _6025_/D VGND VGND VPWR VPWR _6179_/A2 sky130_fd_sc_hd__buf_6
XFILLER_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4860_ _4575_/B _4845_/B _5079_/B _5079_/A VGND VGND VPWR VPWR _4860_/X sky130_fd_sc_hd__a211o_1
X_3811_ _6666_/Q _3843_/B _3898_/B _3845_/A VGND VGND VPWR VPWR _3812_/B sky130_fd_sc_hd__a31o_2
XFILLER_32_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_28 _7096_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4791_ _4772_/A _5165_/A _4772_/C _4936_/A VGND VGND VPWR VPWR _4791_/X sky130_fd_sc_hd__a31o_1
XANTENNA_39 _3398_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_17 _6535_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6530_ _7225_/CLK _6530_/D fanout850/X VGND VGND VPWR VPWR _6530_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_186_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3742_ input52/X _4025_/A hold65/A _7149_/Q VGND VGND VPWR VPWR _3742_/X sky130_fd_sc_hd__a22o_4
XFILLER_13_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6461_ _3938_/A1 _6461_/D _6416_/X VGND VGND VPWR VPWR hold5/A sky130_fd_sc_hd__dfrtp_2
X_3673_ _5225_/A hold63/X VGND VGND VPWR VPWR _5191_/A sky130_fd_sc_hd__nor2_4
X_6392_ _4236_/B _6392_/A2 _6392_/B1 _4236_/A VGND VGND VPWR VPWR _6392_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5412_ hold783/X wire746/A _5413_/S VGND VGND VPWR VPWR _6987_/D sky130_fd_sc_hd__mux2_1
X_5343_ _5595_/A0 _6925_/Q _5350_/S VGND VGND VPWR VPWR _6925_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5274_ _5598_/A0 hold633/X _5278_/S VGND VGND VPWR VPWR _6864_/D sky130_fd_sc_hd__mux2_1
Xoutput179 _3227_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[13] sky130_fd_sc_hd__buf_8
XFILLER_102_616 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7013_ _7134_/CLK _7013_/D fanout861/X VGND VGND VPWR VPWR _7013_/Q sky130_fd_sc_hd__dfstp_4
X_4225_ hold756/X _4224_/X _4235_/S VGND VGND VPWR VPWR _4225_/X sky130_fd_sc_hd__mux2_1
X_4156_ hold693/X wire794/X _4159_/S VGND VGND VPWR VPWR _6625_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4087_ hold328/X _5599_/A0 _4087_/S VGND VGND VPWR VPWR _6567_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4989_ _4989_/A _4989_/B VGND VGND VPWR VPWR _5121_/C sky130_fd_sc_hd__nor2_1
XFILLER_183_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6728_ _6787_/CLK _6728_/D fanout854/X VGND VGND VPWR VPWR _6728_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6659_ _6752_/CLK _6659_/D fanout857/X VGND VGND VPWR VPWR _6659_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_191_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput37 mgmt_gpio_in[10] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__clkbuf_4
Xinput15 mask_rev_in[1] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__clkbuf_4
Xinput26 mask_rev_in[2] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__clkbuf_4
XFILLER_183_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput48 mgmt_gpio_in[20] VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__clkbuf_4
XFILLER_143_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput59 mgmt_gpio_in[30] VGND VGND VPWR VPWR wire901/A sky130_fd_sc_hd__buf_6
Xwire763 wire763/A VGND VGND VPWR VPWR wire763/X sky130_fd_sc_hd__buf_8
Xwire796 hold36/X VGND VGND VPWR VPWR wire796/X sky130_fd_sc_hd__buf_8
Xmax_length372 _6060_/B VGND VGND VPWR VPWR _6357_/A2 sky130_fd_sc_hd__buf_8
Xmax_length394 _3374_/Y VGND VGND VPWR VPWR _3425_/B1 sky130_fd_sc_hd__buf_6
XFILLER_6_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4010_ hold810/X _4009_/X _4024_/S VGND VGND VPWR VPWR _6506_/D sky130_fd_sc_hd__mux2_1
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5961_ wire824/X _7186_/Q wire381/X _5960_/X VGND VGND VPWR VPWR _5961_/X sky130_fd_sc_hd__a211o_2
X_4912_ _4965_/B _4898_/B _4603_/B VGND VGND VPWR VPWR _5069_/C sky130_fd_sc_hd__a21oi_1
X_5892_ _6768_/Q wire686/X wire678/X _7221_/Q _5891_/X VGND VGND VPWR VPWR _5893_/D
+ sky130_fd_sc_hd__a221o_4
XFILLER_178_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4843_ _5023_/A _4986_/C VGND VGND VPWR VPWR _4845_/B sky130_fd_sc_hd__nand2_8
X_4774_ _4774_/A _4776_/B _4774_/C _4930_/C VGND VGND VPWR VPWR _4927_/B sky130_fd_sc_hd__or4b_4
XFILLER_193_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6513_ _7156_/CLK _6513_/D fanout880/X VGND VGND VPWR VPWR _6513_/Q sky130_fd_sc_hd__dfrtp_4
X_3725_ _3725_/A _3725_/B _3725_/C _3725_/D VGND VGND VPWR VPWR _3726_/D sky130_fd_sc_hd__or4_1
XFILLER_173_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6444_ _6447_/A _6447_/B VGND VGND VPWR VPWR _6444_/X sky130_fd_sc_hd__and2_1
XFILLER_161_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3656_ wire519/X _5432_/A _5441_/A _7015_/Q _3655_/X VGND VGND VPWR VPWR _3664_/B
+ sky130_fd_sc_hd__a221o_1
X_6375_ _6402_/A2 _6372_/A _4236_/C VGND VGND VPWR VPWR _6376_/B sky130_fd_sc_hd__a21boi_1
X_3587_ _3587_/A _3587_/B _3587_/C _3587_/D VGND VGND VPWR VPWR _3588_/D sky130_fd_sc_hd__or4_1
X_5326_ wire794/A _6910_/Q _5332_/S VGND VGND VPWR VPWR _6910_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5257_ wire763/X hold411/X _5260_/S VGND VGND VPWR VPWR _5257_/X sky130_fd_sc_hd__mux2_1
X_4208_ hold407/X _4207_/X _4218_/S VGND VGND VPWR VPWR _4208_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5188_ _6409_/A0 hold807/X _5190_/S VGND VGND VPWR VPWR _6787_/D sky130_fd_sc_hd__mux2_1
X_4139_ _5498_/A0 _6611_/Q _4141_/S VGND VGND VPWR VPWR _6611_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3510_ _5234_/A _3510_/B VGND VGND VPWR VPWR _4049_/A sky130_fd_sc_hd__nor2_8
Xwire560 _6787_/Q VGND VGND VPWR VPWR wire560/X sky130_fd_sc_hd__buf_6
X_4490_ _4651_/B _4746_/A VGND VGND VPWR VPWR _4819_/D sky130_fd_sc_hd__or2_2
XFILLER_128_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire593 _6023_/C VGND VGND VPWR VPWR wire593/X sky130_fd_sc_hd__buf_8
XFILLER_7_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold618 _7103_/Q VGND VGND VPWR VPWR hold618/X sky130_fd_sc_hd__bufbuf_16
Xhold607 _6832_/Q VGND VGND VPWR VPWR hold607/X sky130_fd_sc_hd__bufbuf_16
Xwire571 _6596_/Q VGND VGND VPWR VPWR wire571/X sky130_fd_sc_hd__buf_6
Xhold629 _6952_/Q VGND VGND VPWR VPWR hold629/X sky130_fd_sc_hd__bufbuf_16
XFILLER_143_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3441_ _6970_/Q _3327_/Y _4234_/S wire895/A VGND VGND VPWR VPWR _3441_/X sky130_fd_sc_hd__a22o_4
XFILLER_143_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3372_ hold96/X _3540_/A VGND VGND VPWR VPWR _3372_/Y sky130_fd_sc_hd__nor2_1
X_6160_ _7193_/Q _5665_/Y _6159_/X VGND VGND VPWR VPWR _7193_/D sky130_fd_sc_hd__o21a_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5111_ _5157_/B _5155_/A _5178_/B _5156_/C VGND VGND VPWR VPWR _5111_/X sky130_fd_sc_hd__or4_4
XFILLER_69_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6091_ _7015_/Q _6036_/Y _6139_/B1 _7039_/Q VGND VGND VPWR VPWR _6091_/X sky130_fd_sc_hd__a22o_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _4745_/A _5062_/C _4734_/X VGND VGND VPWR VPWR _5042_/Y sky130_fd_sc_hd__o21ai_2
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_51_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _7072_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_53_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6993_ _7129_/CLK _6993_/D fanout863/X VGND VGND VPWR VPWR _6993_/Q sky130_fd_sc_hd__dfrtp_2
X_5944_ _6647_/Q wire690/X _5964_/B1 _6602_/Q VGND VGND VPWR VPWR _5944_/X sky130_fd_sc_hd__a22o_2
XFILLER_80_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5875_ _6713_/Q wire702/X _5702_/X _6550_/Q VGND VGND VPWR VPWR _5875_/X sky130_fd_sc_hd__a22o_1
XFILLER_178_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4826_ _4562_/B _5062_/B _4725_/Y _4823_/X _4825_/X VGND VGND VPWR VPWR _4826_/X
+ sky130_fd_sc_hd__o2111a_1
Xclkbuf_leaf_66_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7135_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_147_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4757_ _4965_/B _4757_/B VGND VGND VPWR VPWR _5174_/B sky130_fd_sc_hd__nor2_1
XFILLER_119_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4688_ _4728_/A _4690_/A _5062_/B VGND VGND VPWR VPWR _4717_/B sky130_fd_sc_hd__or3_4
XFILLER_107_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3708_ _6650_/Q _4184_/A _3543_/Y _6541_/Q _3680_/X VGND VGND VPWR VPWR _3709_/D
+ sky130_fd_sc_hd__a221o_4
XFILLER_146_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3639_ input22/X _3302_/Y _4286_/A _6740_/Q VGND VGND VPWR VPWR _3639_/X sky130_fd_sc_hd__a22o_1
X_6427_ _6455_/A _6455_/B VGND VGND VPWR VPWR _6427_/X sky130_fd_sc_hd__and2_1
XFILLER_162_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6358_ wire824/X _7200_/Q wire381/X VGND VGND VPWR VPWR _6358_/X sky130_fd_sc_hd__a21o_1
XFILLER_191_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5309_ _5498_/A0 hold721/X _5314_/S VGND VGND VPWR VPWR _6895_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_606 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6289_ wire563/X wire575/X _6335_/B _6775_/Q VGND VGND VPWR VPWR _6289_/X sky130_fd_sc_hd__a22o_1
XFILLER_102_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_19_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _6951_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_16_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold4 hold4/A VGND VGND VPWR VPWR hold4/X sky130_fd_sc_hd__bufbuf_16
XFILLER_79_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3990_ _6493_/Q wire753/X _3994_/S VGND VGND VPWR VPWR _6493_/D sky130_fd_sc_hd__mux2_1
XFILLER_35_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5660_ _7158_/Q _5659_/X _5658_/S _7174_/Q VGND VGND VPWR VPWR _7174_/D sky130_fd_sc_hd__a2bb2o_1
X_4611_ _4875_/A _5005_/C _4610_/Y _4564_/A _4593_/Y VGND VGND VPWR VPWR _4612_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_175_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5591_ _5600_/A0 hold435/X _5593_/S VGND VGND VPWR VPWR _7146_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4542_ _5033_/A _4542_/B _4542_/C _4542_/D VGND VGND VPWR VPWR _4542_/X sky130_fd_sc_hd__or4_1
XFILLER_128_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold415 _6675_/Q VGND VGND VPWR VPWR hold415/X sky130_fd_sc_hd__bufbuf_16
X_4473_ _4525_/A _4572_/A VGND VGND VPWR VPWR _4956_/A sky130_fd_sc_hd__nor2_8
Xhold426 _6930_/Q VGND VGND VPWR VPWR hold426/X sky130_fd_sc_hd__bufbuf_16
XFILLER_143_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold404 _6593_/Q VGND VGND VPWR VPWR hold404/X sky130_fd_sc_hd__bufbuf_16
Xwire390 _4262_/A VGND VGND VPWR VPWR wire390/X sky130_fd_sc_hd__buf_6
X_3424_ _6962_/Q _5378_/A _5306_/A _6898_/Q VGND VGND VPWR VPWR _3424_/X sky130_fd_sc_hd__a22o_1
Xhold437 _5357_/X VGND VGND VPWR VPWR _6938_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_144_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold448 _6608_/Q VGND VGND VPWR VPWR hold448/X sky130_fd_sc_hd__bufbuf_16
X_6212_ _7140_/Q wire642/X _6212_/B1 _7100_/Q VGND VGND VPWR VPWR _6212_/X sky130_fd_sc_hd__a22o_1
Xhold459 _6597_/Q VGND VGND VPWR VPWR hold459/X sky130_fd_sc_hd__bufbuf_16
XFILLER_143_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7192_ _7196_/CLK _7192_/D fanout869/X VGND VGND VPWR VPWR _7192_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_98_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6143_ _6985_/Q _6028_/X _6034_/Y _6993_/Q _6142_/X VGND VGND VPWR VPWR _6144_/D
+ sky130_fd_sc_hd__a221o_1
X_3355_ _3508_/A _3355_/B VGND VGND VPWR VPWR _5540_/A sky130_fd_sc_hd__nor2_8
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _6950_/Q wire637/X wire635/X _6926_/Q VGND VGND VPWR VPWR _6074_/X sky130_fd_sc_hd__a22o_1
X_3286_ _3508_/A hold63/X VGND VGND VPWR VPWR _5522_/A sky130_fd_sc_hd__nor2_8
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5025_ _5164_/B _4756_/B _4746_/X _4724_/B VGND VGND VPWR VPWR _5025_/X sky130_fd_sc_hd__o22a_2
XFILLER_85_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6976_ _6979_/CLK _6976_/D fanout884/X VGND VGND VPWR VPWR _6976_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5927_ _5927_/A _5927_/B _5927_/C _5927_/D VGND VGND VPWR VPWR _5927_/X sky130_fd_sc_hd__or4_4
XFILLER_81_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5858_ wire552/X _5700_/X _5857_/X VGND VGND VPWR VPWR _5861_/C sky130_fd_sc_hd__a21o_1
XFILLER_22_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4809_ _4697_/A _5005_/C _4746_/X VGND VGND VPWR VPWR _4809_/X sky130_fd_sc_hd__a21o_1
XFILLER_119_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5789_ _6881_/Q _5674_/X wire673/X _6897_/Q _5788_/X VGND VGND VPWR VPWR _5796_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6830_ _7107_/CLK _6830_/D fanout866/X VGND VGND VPWR VPWR _6830_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6761_ _6806_/CLK _6761_/D fanout848/X VGND VGND VPWR VPWR _6761_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5712_ _6877_/Q _5934_/B1 _5690_/X wire487/X _5711_/X VGND VGND VPWR VPWR _5712_/X
+ sky130_fd_sc_hd__a221o_2
X_3973_ _6838_/Q _3973_/B VGND VGND VPWR VPWR _3973_/X sky130_fd_sc_hd__and2_4
XFILLER_188_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6692_ _7122_/CLK _6692_/D fanout887/X VGND VGND VPWR VPWR _6692_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5643_ _7168_/Q _5648_/B _5642_/Y VGND VGND VPWR VPWR _7168_/D sky130_fd_sc_hd__a21oi_1
X_5574_ _5601_/A0 hold221/X hold91/X VGND VGND VPWR VPWR _5574_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4525_ _4525_/A _4572_/A _4538_/A VGND VGND VPWR VPWR _4965_/A sky130_fd_sc_hd__or3b_4
Xhold201 _5331_/X VGND VGND VPWR VPWR _6915_/D sky130_fd_sc_hd__bufbuf_16
Xhold212 _6867_/Q VGND VGND VPWR VPWR hold212/X sky130_fd_sc_hd__bufbuf_16
Xhold223 _7003_/Q VGND VGND VPWR VPWR hold223/X sky130_fd_sc_hd__bufbuf_16
XFILLER_132_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold234 _6481_/Q VGND VGND VPWR VPWR _3249_/B sky130_fd_sc_hd__bufbuf_16
Xhold245 _6881_/Q VGND VGND VPWR VPWR hold245/X sky130_fd_sc_hd__bufbuf_16
Xhold278 _6529_/Q VGND VGND VPWR VPWR hold278/X sky130_fd_sc_hd__bufbuf_16
Xhold267 _6977_/Q VGND VGND VPWR VPWR hold267/X sky130_fd_sc_hd__bufbuf_16
X_4456_ _4469_/A _4558_/B VGND VGND VPWR VPWR _4844_/A sky130_fd_sc_hd__or2_4
Xhold256 _6923_/Q VGND VGND VPWR VPWR hold256/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4387_ _4958_/A _4408_/A VGND VGND VPWR VPWR _4513_/A sky130_fd_sc_hd__or2_4
Xhold289 _7111_/Q VGND VGND VPWR VPWR hold289/X sky130_fd_sc_hd__bufbuf_16
X_3407_ _7075_/Q _5504_/A _3324_/Y _6923_/Q VGND VGND VPWR VPWR _3407_/X sky130_fd_sc_hd__a22o_1
X_7175_ _7194_/CLK _7175_/D fanout867/X VGND VGND VPWR VPWR _7175_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout747 hold200/X VGND VGND VPWR VPWR _5601_/A0 sky130_fd_sc_hd__buf_8
X_6126_ _6904_/Q wire600/X wire646/X _6936_/Q _6125_/X VGND VGND VPWR VPWR _6132_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_86_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3338_ _3353_/B _5225_/B VGND VGND VPWR VPWR _3338_/Y sky130_fd_sc_hd__nor2_8
XFILLER_105_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6057_ _6057_/A _6057_/B _6057_/C _6057_/D VGND VGND VPWR VPWR _6058_/C sky130_fd_sc_hd__or4_1
XFILLER_100_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3269_ hold60/X hold165/X _3953_/A VGND VGND VPWR VPWR _3269_/X sky130_fd_sc_hd__mux2_8
X_5008_ _5008_/A _5008_/B VGND VGND VPWR VPWR _5012_/A sky130_fd_sc_hd__nand2_1
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_107 _6196_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 _7153_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_129 mask_rev_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6959_ _7111_/CLK _6959_/D _6421_/A VGND VGND VPWR VPWR _6959_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_10_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length779 wire780/X VGND VGND VPWR VPWR _5255_/A0 sky130_fd_sc_hd__buf_6
XFILLER_146_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold790 _6563_/Q VGND VGND VPWR VPWR hold790/X sky130_fd_sc_hd__bufbuf_16
XFILLER_122_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput306 _3969_/X VGND VGND VPWR VPWR ser_rx sky130_fd_sc_hd__buf_8
Xoutput317 _7202_/Q VGND VGND VPWR VPWR wb_ack_o sky130_fd_sc_hd__buf_8
X_5290_ wire794/A hold443/X _5296_/S VGND VGND VPWR VPWR _5290_/X sky130_fd_sc_hd__mux2_1
Xoutput339 _7208_/Q VGND VGND VPWR VPWR wb_dat_o[29] sky130_fd_sc_hd__buf_8
XFILLER_126_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput328 _6558_/Q VGND VGND VPWR VPWR wb_dat_o[19] sky130_fd_sc_hd__buf_8
XFILLER_113_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4310_ _4310_/A _6406_/B VGND VGND VPWR VPWR _4315_/S sky130_fd_sc_hd__and2_4
X_4241_ _4241_/A hold45/X _6421_/B hold31/X VGND VGND VPWR VPWR hold32/A sky130_fd_sc_hd__or4_4
XFILLER_114_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4172_ _4172_/A _6406_/B VGND VGND VPWR VPWR _4177_/S sky130_fd_sc_hd__and2_4
XFILLER_121_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6813_ _6815_/CLK _6813_/D fanout855/X VGND VGND VPWR VPWR _6813_/Q sky130_fd_sc_hd__dfstp_4
X_3956_ _6474_/Q _6446_/A VGND VGND VPWR VPWR _3956_/Y sky130_fd_sc_hd__nor2_1
X_6744_ _6744_/CLK _6744_/D wire860/X VGND VGND VPWR VPWR _6744_/Q sky130_fd_sc_hd__dfrtp_2
X_6675_ _7133_/CLK _6675_/D fanout882/X VGND VGND VPWR VPWR _6675_/Q sky130_fd_sc_hd__dfrtp_2
X_3887_ _4349_/C _4349_/D _3887_/C input116/X VGND VGND VPWR VPWR _3895_/B sky130_fd_sc_hd__or4b_4
X_5626_ _5626_/A _6679_/Q VGND VGND VPWR VPWR _5654_/A sky130_fd_sc_hd__nor2_4
XFILLER_191_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5557_ hold366/X _5602_/A0 _5557_/S VGND VGND VPWR VPWR _5557_/X sky130_fd_sc_hd__mux2_1
X_5488_ hold38/X _7054_/Q _5494_/S VGND VGND VPWR VPWR _7054_/D sky130_fd_sc_hd__mux2_1
X_4508_ _4711_/A _4581_/B VGND VGND VPWR VPWR _5033_/A sky130_fd_sc_hd__and2_2
XFILLER_132_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4439_ _4774_/A _4593_/A VGND VGND VPWR VPWR _4525_/A sky130_fd_sc_hd__or2_4
XFILLER_132_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7227_ _7227_/A VGND VGND VPWR VPWR _7227_/X sky130_fd_sc_hd__buf_2
XFILLER_160_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7158_ _7194_/CLK _7158_/D fanout867/X VGND VGND VPWR VPWR _7158_/Q sky130_fd_sc_hd__dfrtp_2
X_6109_ _7190_/Q _6108_/X _6109_/S VGND VGND VPWR VPWR _6109_/X sky130_fd_sc_hd__mux2_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7089_ _7095_/CLK _7089_/D fanout862/X VGND VGND VPWR VPWR _7089_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire901 wire901/A VGND VGND VPWR VPWR wire901/X sky130_fd_sc_hd__buf_6
Xwire912 wire912/A VGND VGND VPWR VPWR wire912/X sky130_fd_sc_hd__buf_6
XFILLER_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length576 _6034_/Y VGND VGND VPWR VPWR _6293_/B1 sky130_fd_sc_hd__buf_6
XFILLER_170_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4790_ _4692_/C _4758_/C _4668_/B _4411_/Y VGND VGND VPWR VPWR _4796_/C sky130_fd_sc_hd__a31o_1
XFILLER_82_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3810_ _6467_/Q _3810_/B VGND VGND VPWR VPWR _3898_/B sky130_fd_sc_hd__nand2_1
XANTENNA_29 _7120_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_18 _4208_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3741_ _6901_/Q _5315_/A _5585_/A _7141_/Q VGND VGND VPWR VPWR _3741_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6460_ _3938_/A1 _6460_/D _6415_/X VGND VGND VPWR VPWR hold49/A sky130_fd_sc_hd__dfrtp_2
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3672_ _3672_/A _5234_/A VGND VGND VPWR VPWR _5242_/A sky130_fd_sc_hd__nor2_4
X_6391_ _6390_/X _7215_/Q _6400_/S VGND VGND VPWR VPWR _7215_/D sky130_fd_sc_hd__mux2_1
X_5411_ hold534/X wire757/X _5413_/S VGND VGND VPWR VPWR _6986_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5342_ _5342_/A _5594_/B VGND VGND VPWR VPWR _5350_/S sky130_fd_sc_hd__nand2_8
XFILLER_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5273_ _5597_/A0 hold276/X _5278_/S VGND VGND VPWR VPWR _6863_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7012_ _7140_/CLK _7012_/D fanout865/X VGND VGND VPWR VPWR _7012_/Q sky130_fd_sc_hd__dfrtp_2
X_4224_ hold571/X _5255_/A0 _4234_/S VGND VGND VPWR VPWR _4224_/X sky130_fd_sc_hd__mux2_1
X_4155_ hold801/X _5487_/A0 _4159_/S VGND VGND VPWR VPWR _4155_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4086_ _6566_/Q hold83/X _4087_/S VGND VGND VPWR VPWR _4086_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4988_ _4988_/A _4997_/B VGND VGND VPWR VPWR _5081_/C sky130_fd_sc_hd__nor2_4
XFILLER_11_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3939_ _6506_/Q wire896/A _3939_/S VGND VGND VPWR VPWR _3939_/X sky130_fd_sc_hd__mux2_2
X_6727_ _6727_/CLK _6727_/D wire860/X VGND VGND VPWR VPWR _6727_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_176_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6658_ _6806_/CLK _6658_/D fanout848/X VGND VGND VPWR VPWR _6658_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_137_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5609_ _5617_/A _5609_/B _5609_/C VGND VGND VPWR VPWR _7157_/D sky130_fd_sc_hd__and3_1
X_6589_ _6591_/CLK _6589_/D fanout873/X VGND VGND VPWR VPWR _6589_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire731 _3895_/Y VGND VGND VPWR VPWR _3915_/B sky130_fd_sc_hd__buf_6
XFILLER_155_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire742 hold21/X VGND VGND VPWR VPWR wire742/X sky130_fd_sc_hd__buf_8
XFILLER_128_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput16 mask_rev_in[20] VGND VGND VPWR VPWR input16/X sky130_fd_sc_hd__buf_4
Xinput27 mask_rev_in[30] VGND VGND VPWR VPWR input27/X sky130_fd_sc_hd__clkbuf_4
XFILLER_182_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire775 hold81/X VGND VGND VPWR VPWR wire775/X sky130_fd_sc_hd__buf_6
Xinput49 mgmt_gpio_in[21] VGND VGND VPWR VPWR wire907/A sky130_fd_sc_hd__buf_6
Xwire786 hold13/X VGND VGND VPWR VPWR wire786/X sky130_fd_sc_hd__buf_8
Xinput38 mgmt_gpio_in[11] VGND VGND VPWR VPWR wire910/A sky130_fd_sc_hd__buf_6
XFILLER_109_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire753 wire753/A VGND VGND VPWR VPWR wire753/X sky130_fd_sc_hd__buf_8
Xmax_length395 _5405_/A VGND VGND VPWR VPWR _3739_/B1 sky130_fd_sc_hd__buf_6
Xmax_length384 _5566_/S VGND VGND VPWR VPWR _5565_/S sky130_fd_sc_hd__buf_6
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5960_ _6533_/Q _5722_/B _5953_/X _5959_/X _6308_/S VGND VGND VPWR VPWR _5960_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_53_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4911_ _4983_/B _4911_/B _4976_/A _4911_/D VGND VGND VPWR VPWR _4913_/C sky130_fd_sc_hd__or4_1
X_5891_ _6545_/Q wire706/X wire651/A _6758_/Q VGND VGND VPWR VPWR _5891_/X sky130_fd_sc_hd__a22o_1
X_4842_ _4554_/A _5087_/A _4554_/B _4507_/A VGND VGND VPWR VPWR _4842_/X sky130_fd_sc_hd__a22o_4
XANTENNA_290 _6805_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4773_ _4773_/A _4773_/B VGND VGND VPWR VPWR _4776_/B sky130_fd_sc_hd__or2_4
XFILLER_119_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6512_ _6931_/CLK _6512_/D fanout885/X VGND VGND VPWR VPWR _6512_/Q sky130_fd_sc_hd__dfrtp_1
X_3724_ _6714_/Q _4256_/A _4118_/A _6595_/Q _3723_/X VGND VGND VPWR VPWR _3725_/D
+ sky130_fd_sc_hd__a221o_4
XFILLER_174_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6443_ _6455_/A _6455_/B VGND VGND VPWR VPWR _6443_/X sky130_fd_sc_hd__and2_1
X_3655_ _6991_/Q _5414_/A _4310_/A _6760_/Q VGND VGND VPWR VPWR _3655_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6374_ _6372_/A _6374_/A2 wire817/X VGND VGND VPWR VPWR _6374_/X sky130_fd_sc_hd__a21bo_1
X_3586_ _6976_/Q _5396_/A _5245_/A input64/X _3585_/X VGND VGND VPWR VPWR _3587_/D
+ sky130_fd_sc_hd__a221o_4
XFILLER_161_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5325_ _5595_/A0 _6909_/Q _5332_/S VGND VGND VPWR VPWR _6909_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5256_ wire770/X hold424/X _5260_/S VGND VGND VPWR VPWR _5256_/X sky130_fd_sc_hd__mux2_1
X_4207_ hold214/X _5248_/A0 _4209_/S VGND VGND VPWR VPWR _4207_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5187_ _6408_/A0 hold695/X _5190_/S VGND VGND VPWR VPWR _5187_/X sky130_fd_sc_hd__mux2_1
X_4138_ wire794/A hold430/X _4141_/S VGND VGND VPWR VPWR _4138_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4069_ _5247_/A0 hold570/X _4072_/S VGND VGND VPWR VPWR _6551_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire550 _6872_/Q VGND VGND VPWR VPWR wire550/X sky130_fd_sc_hd__buf_6
XFILLER_183_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire594 _6002_/Y VGND VGND VPWR VPWR wire594/X sky130_fd_sc_hd__buf_6
Xhold608 _5235_/X VGND VGND VPWR VPWR _6832_/D sky130_fd_sc_hd__bufbuf_16
Xwire572 _6537_/Q VGND VGND VPWR VPWR wire572/X sky130_fd_sc_hd__buf_6
Xwire561 _6786_/Q VGND VGND VPWR VPWR wire561/X sky130_fd_sc_hd__buf_6
XFILLER_171_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3440_ _7098_/Q _5531_/A _5360_/A _6946_/Q _3439_/X VGND VGND VPWR VPWR _3452_/C
+ sky130_fd_sc_hd__a221o_1
Xhold619 _5543_/X VGND VGND VPWR VPWR _7103_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_112_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3371_ _3668_/A _3552_/B VGND VGND VPWR VPWR _3371_/Y sky130_fd_sc_hd__nor2_4
X_5110_ _5004_/A _4469_/Y _4659_/A _5099_/A _5046_/A VGND VGND VPWR VPWR _5156_/C
+ sky130_fd_sc_hd__a311o_2
XFILLER_97_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6090_ wire515/X wire589/X wire615/X _7087_/Q _6088_/X VGND VGND VPWR VPWR _6090_/X
+ sky130_fd_sc_hd__a221o_2
X_5041_ _4469_/A _4470_/B _4565_/Y VGND VGND VPWR VPWR _5041_/X sky130_fd_sc_hd__a21o_2
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_wb_clk_i wb_clk_i VGND VGND VPWR VPWR clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_8
XFILLER_93_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6992_ _6992_/CLK _6992_/D fanout868/X VGND VGND VPWR VPWR _6992_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_179_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5943_ _6566_/Q wire673/X wire653/X _6652_/Q VGND VGND VPWR VPWR _5959_/A sky130_fd_sc_hd__a22o_1
XFILLER_179_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5874_ _7183_/Q _6110_/S _5872_/X _5873_/X VGND VGND VPWR VPWR _7183_/D sky130_fd_sc_hd__o22a_1
XFILLER_33_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4825_ _4898_/B _4728_/X _4746_/X _5164_/B _4824_/X VGND VGND VPWR VPWR _4825_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_193_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4756_ _4965_/B _4756_/B VGND VGND VPWR VPWR _5071_/B sky130_fd_sc_hd__nor2_1
XFILLER_175_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4687_ _4687_/A _4832_/C VGND VGND VPWR VPWR _5095_/A sky130_fd_sc_hd__nor2_4
X_3707_ _6950_/Q _5369_/A wire391/X wire561/X _3706_/X VGND VGND VPWR VPWR _3709_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3638_ _7031_/Q _5459_/A _3638_/B1 _7079_/Q _3637_/X VGND VGND VPWR VPWR _3645_/A
+ sky130_fd_sc_hd__a221o_4
X_6426_ _6446_/A _6447_/B VGND VGND VPWR VPWR _6426_/X sky130_fd_sc_hd__and2_1
XFILLER_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3569_ _6928_/Q wire436/X _3567_/X _3568_/X VGND VGND VPWR VPWR _3588_/B sky130_fd_sc_hd__a211o_1
XFILLER_68_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6357_ _6534_/Q _6357_/A2 _6356_/X _6308_/S VGND VGND VPWR VPWR _6357_/X sky130_fd_sc_hd__o211a_2
X_5308_ wire794/A hold442/X _5314_/S VGND VGND VPWR VPWR _6894_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6288_ _6760_/Q wire589/X _6337_/B1 _6646_/Q _6287_/X VGND VGND VPWR VPWR _6288_/X
+ sky130_fd_sc_hd__a221o_1
X_5239_ hold7/X _6834_/Q _5241_/S VGND VGND VPWR VPWR hold8/A sky130_fd_sc_hd__mux2_1
XFILLER_102_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold5 hold5/A VGND VGND VPWR VPWR hold5/X sky130_fd_sc_hd__bufbuf_16
XFILLER_75_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4610_ _4536_/B _4537_/X _4735_/B _4740_/A _4949_/B VGND VGND VPWR VPWR _4610_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_175_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5590_ _5599_/A0 hold303/X _5593_/S VGND VGND VPWR VPWR _5590_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4541_ _5023_/A _4871_/A _4997_/A VGND VGND VPWR VPWR _4542_/D sky130_fd_sc_hd__a21oi_1
XFILLER_128_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4472_ _4707_/B _4534_/B VGND VGND VPWR VPWR _4949_/A sky130_fd_sc_hd__nor2_8
Xhold416 _6462_/Q VGND VGND VPWR VPWR hold75/A sky130_fd_sc_hd__bufbuf_16
XFILLER_144_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold427 _7137_/Q VGND VGND VPWR VPWR hold427/X sky130_fd_sc_hd__bufbuf_16
Xhold405 _6544_/Q VGND VGND VPWR VPWR hold405/X sky130_fd_sc_hd__bufbuf_16
Xwire391 _5185_/A VGND VGND VPWR VPWR wire391/X sky130_fd_sc_hd__buf_6
Xhold449 _7154_/Q VGND VGND VPWR VPWR hold449/X sky130_fd_sc_hd__bufbuf_16
XFILLER_143_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7191_ _7196_/CLK _7191_/D fanout869/X VGND VGND VPWR VPWR _7191_/Q sky130_fd_sc_hd__dfrtp_1
X_3423_ _7188_/Q _6829_/Q _6831_/Q VGND VGND VPWR VPWR _3423_/X sky130_fd_sc_hd__mux2_8
X_6211_ _7084_/Q _6211_/B VGND VGND VPWR VPWR _6211_/X sky130_fd_sc_hd__and2_1
Xhold438 _6990_/Q VGND VGND VPWR VPWR hold438/X sky130_fd_sc_hd__bufbuf_16
X_6142_ _7073_/Q _6009_/X wire627/X _6969_/Q VGND VGND VPWR VPWR _6142_/X sky130_fd_sc_hd__a22o_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3354_ wire541/X _3582_/B1 _3353_/Y _6884_/Q VGND VGND VPWR VPWR _3354_/X sky130_fd_sc_hd__a22o_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3285_ hold62/X hold43/X VGND VGND VPWR VPWR hold63/A sky130_fd_sc_hd__or2_4
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ _7126_/Q wire597/X wire611/X _7006_/Q _6072_/X VGND VGND VPWR VPWR _6083_/B
+ sky130_fd_sc_hd__a221o_1
X_5024_ _5024_/A _5035_/B _5024_/C _5035_/D VGND VGND VPWR VPWR _5028_/B sky130_fd_sc_hd__or4_2
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6975_ _7111_/CLK _6975_/D fanout875/X VGND VGND VPWR VPWR _6975_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5926_ wire560/X _5926_/A2 _5964_/B1 _6601_/Q _5925_/X VGND VGND VPWR VPWR _5927_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5857_ _7108_/Q _5857_/A2 _5706_/X wire499/X VGND VGND VPWR VPWR _5857_/X sky130_fd_sc_hd__a22o_1
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4808_ _4808_/A _5069_/B VGND VGND VPWR VPWR _5037_/A sky130_fd_sc_hd__or2_2
X_5788_ _7009_/Q wire701/X wire692/X _6993_/Q VGND VGND VPWR VPWR _5788_/X sky130_fd_sc_hd__a22o_1
XFILLER_182_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4739_ _4714_/B _5147_/C _4738_/Y _4734_/X _4505_/X VGND VGND VPWR VPWR _4739_/X
+ sky130_fd_sc_hd__o2111a_2
XFILLER_147_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6409_ _6409_/A0 hold812/X _6411_/S VGND VGND VPWR VPWR _7223_/D sky130_fd_sc_hd__mux2_1
XFILLER_1_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_50_csclk clkbuf_3_3_0_csclk/X VGND VGND VPWR VPWR _6996_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_65_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7134_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_82_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6760_ _6787_/CLK _6760_/D fanout854/X VGND VGND VPWR VPWR _6760_/Q sky130_fd_sc_hd__dfstp_4
X_5711_ wire520/X _5678_/X _5702_/X _6885_/Q VGND VGND VPWR VPWR _5711_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3972_ _6837_/Q _3972_/B VGND VGND VPWR VPWR _3972_/X sky130_fd_sc_hd__and2_4
X_6691_ _6930_/CLK hold33/X fanout887/X VGND VGND VPWR VPWR _6691_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5642_ _7168_/Q _5635_/B _5648_/B VGND VGND VPWR VPWR _5642_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_176_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5573_ _5600_/A0 hold434/X hold91/X VGND VGND VPWR VPWR _7130_/D sky130_fd_sc_hd__mux2_1
Xhold202 _6875_/Q VGND VGND VPWR VPWR hold202/X sky130_fd_sc_hd__bufbuf_16
X_4524_ _4988_/A _4671_/A VGND VGND VPWR VPWR _4849_/A sky130_fd_sc_hd__nor2_2
Xhold213 _5277_/X VGND VGND VPWR VPWR _6867_/D sky130_fd_sc_hd__bufbuf_16
Xhold224 _5430_/X VGND VGND VPWR VPWR _7003_/D sky130_fd_sc_hd__bufbuf_16
Xclkbuf_leaf_18_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _6950_/CLK sky130_fd_sc_hd__clkbuf_8
Xhold235 _3249_/Y VGND VGND VPWR VPWR hold235/X sky130_fd_sc_hd__bufbuf_16
Xhold246 _6913_/Q VGND VGND VPWR VPWR hold246/X sky130_fd_sc_hd__bufbuf_16
Xhold268 _6922_/Q VGND VGND VPWR VPWR hold268/X sky130_fd_sc_hd__bufbuf_16
X_4455_ _4694_/A _4745_/A VGND VGND VPWR VPWR _4808_/A sky130_fd_sc_hd__nor2_2
XFILLER_104_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold257 _7087_/Q VGND VGND VPWR VPWR hold257/X sky130_fd_sc_hd__bufbuf_16
Xhold279 _4042_/X VGND VGND VPWR VPWR _6529_/D sky130_fd_sc_hd__bufbuf_16
X_4386_ _4996_/A _5164_/A VGND VGND VPWR VPWR _4386_/Y sky130_fd_sc_hd__nor2_1
XFILLER_132_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3406_ _6907_/Q _3443_/A2 _3726_/A _3403_/X _3405_/X VGND VGND VPWR VPWR _3415_/C
+ sky130_fd_sc_hd__a2111o_1
X_7174_ _7194_/CLK _7174_/D fanout866/X VGND VGND VPWR VPWR _7174_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout748 hold198/X VGND VGND VPWR VPWR hold199/A sky130_fd_sc_hd__buf_6
X_6125_ _6952_/Q wire637/X wire635/X _6928_/Q VGND VGND VPWR VPWR _6125_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3337_ _6818_/Q _5207_/A _3336_/X VGND VGND VPWR VPWR _3378_/A sky130_fd_sc_hd__a21o_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout759 _4303_/A0 VGND VGND VPWR VPWR _6411_/A0 sky130_fd_sc_hd__buf_8
X_6056_ _6933_/Q wire646/X wire593/X _6869_/Q _6055_/X VGND VGND VPWR VPWR _6057_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_105_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ hold59/X _6477_/Q _3845_/A VGND VGND VPWR VPWR hold60/A sky130_fd_sc_hd__mux2_1
X_5007_ _4707_/B _4746_/B _5050_/C _4745_/A _4648_/B VGND VGND VPWR VPWR _5008_/B
+ sky130_fd_sc_hd__o32a_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3199_ _6680_/Q VGND VGND VPWR VPWR _5659_/C sky130_fd_sc_hd__inv_2
XFILLER_39_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_108 _6293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_119 _6908_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6958_ _7111_/CLK _6958_/D fanout875/X VGND VGND VPWR VPWR _6958_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_157_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6889_ _6969_/CLK _6889_/D fanout880/X VGND VGND VPWR VPWR _6889_/Q sky130_fd_sc_hd__dfrtp_2
X_5909_ _6714_/Q wire702/X _5702_/X _6551_/Q _5908_/X VGND VGND VPWR VPWR _5910_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_167_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length703 _5857_/A2 VGND VGND VPWR VPWR _5973_/A2 sky130_fd_sc_hd__buf_6
XFILLER_10_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold791 _6629_/Q VGND VGND VPWR VPWR hold791/X sky130_fd_sc_hd__bufbuf_16
Xhold780 _6654_/Q VGND VGND VPWR VPWR hold780/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput307 _3920_/B VGND VGND VPWR VPWR serial_clock sky130_fd_sc_hd__buf_8
XFILLER_141_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput329 _6582_/Q VGND VGND VPWR VPWR wb_dat_o[1] sky130_fd_sc_hd__buf_8
Xoutput318 _6581_/Q VGND VGND VPWR VPWR wb_dat_o[0] sky130_fd_sc_hd__buf_8
XFILLER_4_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4240_ _6360_/A _3953_/A _6704_/Q _4237_/X _4239_/X VGND VGND VPWR VPWR _6689_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4171_ _4303_/A0 hold397/X _4171_/S VGND VGND VPWR VPWR _6638_/D sky130_fd_sc_hd__mux2_1
XFILLER_122_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6812_ _7103_/CLK _6812_/D fanout861/X VGND VGND VPWR VPWR _6812_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_168_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6743_ _6951_/CLK _6743_/D _6421_/A VGND VGND VPWR VPWR _6743_/Q sky130_fd_sc_hd__dfrtp_2
X_3955_ wire843/X _3877_/C _6474_/Q VGND VGND VPWR VPWR _3955_/X sky130_fd_sc_hd__mux2_8
X_6674_ _7133_/CLK hold48/X fanout881/X VGND VGND VPWR VPWR _6674_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3886_ _4351_/A _4351_/B _3886_/C VGND VGND VPWR VPWR _3895_/A sky130_fd_sc_hd__or3_4
XFILLER_137_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5625_ _7162_/Q _7161_/Q VGND VGND VPWR VPWR _5705_/B sky130_fd_sc_hd__and2_4
X_5556_ hold301/X _5601_/A0 _5557_/S VGND VGND VPWR VPWR _5556_/X sky130_fd_sc_hd__mux2_1
X_5487_ _5487_/A0 hold775/X _5494_/S VGND VGND VPWR VPWR _7053_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4507_ _4507_/A _4711_/A _4659_/A VGND VGND VPWR VPWR _4920_/A sky130_fd_sc_hd__and3_4
XFILLER_132_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4438_ _4722_/A _4438_/B VGND VGND VPWR VPWR _4593_/A sky130_fd_sc_hd__xor2_4
XFILLER_160_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4369_ _4529_/A _4650_/B VGND VGND VPWR VPWR _4484_/C sky130_fd_sc_hd__nand2_8
X_7157_ _7194_/CLK _7157_/D fanout866/X VGND VGND VPWR VPWR _7157_/Q sky130_fd_sc_hd__dfrtp_2
X_6108_ _6090_/X _6096_/X _6107_/X _6357_/A2 _6855_/Q VGND VGND VPWR VPWR _6108_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7088_ _7132_/CLK _7088_/D fanout863/X VGND VGND VPWR VPWR _7088_/Q sky130_fd_sc_hd__dfrtp_2
X_6039_ _6877_/Q wire639/X wire624/X _6957_/Q VGND VGND VPWR VPWR _6039_/X sky130_fd_sc_hd__a22o_1
XFILLER_86_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire902 wire904/A VGND VGND VPWR VPWR _3875_/B sky130_fd_sc_hd__buf_8
XFILLER_155_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length577 _6034_/Y VGND VGND VPWR VPWR _6342_/B1 sky130_fd_sc_hd__buf_6
XFILLER_142_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length588 _6010_/Y VGND VGND VPWR VPWR _6337_/A2 sky130_fd_sc_hd__buf_6
XFILLER_123_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_19 _4208_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3740_ _6933_/Q _5351_/A _5279_/A _6869_/Q VGND VGND VPWR VPWR _3740_/X sky130_fd_sc_hd__a22o_2
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3671_ _6739_/Q _4286_/A _5194_/A _6801_/Q VGND VGND VPWR VPWR _3671_/X sky130_fd_sc_hd__a22o_4
X_6390_ _4236_/C _6390_/A2 _6390_/B1 _4236_/A _6389_/X VGND VGND VPWR VPWR _6390_/X
+ sky130_fd_sc_hd__a221o_1
X_5410_ hold349/X hold150/X _5413_/S VGND VGND VPWR VPWR _6985_/D sky130_fd_sc_hd__mux2_1
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5341_ hold382/X wire742/X _5341_/S VGND VGND VPWR VPWR _5341_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5272_ wire794/A hold445/X _5278_/S VGND VGND VPWR VPWR _6862_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7011_ _7042_/CLK _7011_/D fanout865/X VGND VGND VPWR VPWR _7011_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_141_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4223_ hold738/X _4222_/X _4235_/S VGND VGND VPWR VPWR _4223_/X sky130_fd_sc_hd__mux2_1
X_4154_ _4154_/A _4154_/B VGND VGND VPWR VPWR _4159_/S sky130_fd_sc_hd__and2_4
X_4085_ hold549/X _5336_/A1 _4087_/S VGND VGND VPWR VPWR _6565_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4987_ _4987_/A _4987_/B _4992_/B VGND VGND VPWR VPWR _4987_/X sky130_fd_sc_hd__or3_4
X_6726_ _6736_/CLK _6726_/D wire860/X VGND VGND VPWR VPWR _6726_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3938_ _6507_/Q _3938_/A1 _3938_/S VGND VGND VPWR VPWR _3938_/X sky130_fd_sc_hd__mux2_1
X_3869_ hold1/A _6465_/Q _3874_/S VGND VGND VPWR VPWR _6465_/D sky130_fd_sc_hd__mux2_1
X_6657_ _6787_/CLK _6657_/D fanout848/X VGND VGND VPWR VPWR _6657_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_176_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5608_ _7157_/Q _5615_/D VGND VGND VPWR VPWR _5609_/C sky130_fd_sc_hd__or2_1
X_6588_ _7208_/CLK _6588_/D VGND VGND VPWR VPWR _6588_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_192_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5539_ wire739/X hold676/X _5539_/S VGND VGND VPWR VPWR _7100_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_690 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7209_ _7210_/CLK _7209_/D VGND VGND VPWR VPWR _7209_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_587 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire710 _5667_/X VGND VGND VPWR VPWR wire710/X sky130_fd_sc_hd__buf_8
Xwire732 _3859_/Y VGND VGND VPWR VPWR _3874_/S sky130_fd_sc_hd__buf_8
XFILLER_10_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput28 mask_rev_in[31] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__clkbuf_4
Xinput17 mask_rev_in[21] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__clkbuf_4
XFILLER_167_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput39 mgmt_gpio_in[12] VGND VGND VPWR VPWR wire909/A sky130_fd_sc_hd__buf_6
XFILLER_155_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5890_ _6619_/Q wire707/X wire675/A _6654_/Q _5889_/X VGND VGND VPWR VPWR _5893_/C
+ sky130_fd_sc_hd__a221o_1
X_4910_ _5128_/A _5075_/B _4910_/C VGND VGND VPWR VPWR _4911_/D sky130_fd_sc_hd__or3_1
XFILLER_93_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4841_ _4412_/Y _5123_/C VGND VGND VPWR VPWR _5116_/B sky130_fd_sc_hd__nand2b_2
XANTENNA_291 _6913_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_280 hold475/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4772_ _4772_/A _5165_/A _4772_/C VGND VGND VPWR VPWR _4936_/B sky130_fd_sc_hd__and3_1
XFILLER_159_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6511_ _7156_/CLK _6511_/D fanout882/X VGND VGND VPWR VPWR _6511_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_158_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3723_ _6577_/Q _4097_/A _5242_/A _6838_/Q VGND VGND VPWR VPWR _3723_/X sky130_fd_sc_hd__a22o_2
XFILLER_146_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3654_ _3654_/A _3654_/B _3654_/C _3654_/D VGND VGND VPWR VPWR _3664_/A sky130_fd_sc_hd__or4_1
X_6442_ _6446_/A _6447_/B VGND VGND VPWR VPWR _6442_/X sky130_fd_sc_hd__and2_1
XFILLER_173_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6373_ _4236_/A _6371_/Y _6372_/Y _4236_/B VGND VGND VPWR VPWR _6376_/C sky130_fd_sc_hd__a22o_1
XFILLER_161_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3585_ _6553_/Q _3473_/Y _4136_/A _6612_/Q VGND VGND VPWR VPWR _3585_/X sky130_fd_sc_hd__a22o_4
XFILLER_115_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_0_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A VGND VGND VPWR VPWR _7220_/CLK sky130_fd_sc_hd__clkbuf_8
X_5324_ _5324_/A _5594_/B VGND VGND VPWR VPWR _5332_/S sky130_fd_sc_hd__nand2_8
XFILLER_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5255_ _5255_/A0 hold571/X _5260_/S VGND VGND VPWR VPWR _5255_/X sky130_fd_sc_hd__mux2_1
X_4206_ hold323/X _4205_/X _4218_/S VGND VGND VPWR VPWR _4206_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5186_ _6407_/A0 hold784/X _5190_/S VGND VGND VPWR VPWR _6785_/D sky130_fd_sc_hd__mux2_1
X_4137_ _5487_/A0 hold767/X _4141_/S VGND VGND VPWR VPWR _6609_/D sky130_fd_sc_hd__mux2_1
X_4068_ _5487_/A0 hold773/X _4072_/S VGND VGND VPWR VPWR _6550_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6709_ _6712_/CLK _6709_/D fanout872/X VGND VGND VPWR VPWR _6709_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_152_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire551 _6870_/Q VGND VGND VPWR VPWR wire551/X sky130_fd_sc_hd__buf_6
XFILLER_128_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire573 _6404_/X VGND VGND VPWR VPWR wire573/X sky130_fd_sc_hd__buf_6
XFILLER_116_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold609 _7032_/Q VGND VGND VPWR VPWR hold609/X sky130_fd_sc_hd__bufbuf_16
Xwire562 _6765_/Q VGND VGND VPWR VPWR wire562/X sky130_fd_sc_hd__buf_6
XFILLER_143_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3370_ input19/X _3368_/Y _3369_/Y wire525/X _3366_/X VGND VGND VPWR VPWR _3377_/C
+ sky130_fd_sc_hd__a221o_2
XFILLER_151_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _4565_/Y _4689_/Y _4817_/C _5039_/X VGND VGND VPWR VPWR _5048_/A sky130_fd_sc_hd__a211o_2
XFILLER_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6991_ _7135_/CLK _6991_/D fanout864/X VGND VGND VPWR VPWR _6991_/Q sky130_fd_sc_hd__dfrtp_2
X_5942_ _6627_/Q _5963_/B VGND VGND VPWR VPWR _5942_/X sky130_fd_sc_hd__or2_1
XFILLER_93_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5873_ _5611_/A _7182_/Q wire381/A VGND VGND VPWR VPWR _5873_/X sky130_fd_sc_hd__a21o_1
X_4824_ _5164_/B _4756_/B _4746_/X _4898_/B VGND VGND VPWR VPWR _4824_/X sky130_fd_sc_hd__o22a_1
XFILLER_21_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4755_ _4898_/B _4757_/B VGND VGND VPWR VPWR _4893_/B sky130_fd_sc_hd__or2_4
XFILLER_21_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3706_ _6870_/Q _5279_/A _4124_/A _6600_/Q VGND VGND VPWR VPWR _3706_/X sky130_fd_sc_hd__a22o_1
X_4686_ _4724_/B _4832_/C VGND VGND VPWR VPWR _5022_/B sky130_fd_sc_hd__nor2_1
XFILLER_107_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3637_ _7071_/Q _5504_/A _4178_/A _6646_/Q VGND VGND VPWR VPWR _3637_/X sky130_fd_sc_hd__a22o_1
X_6425_ _6455_/A _6425_/B VGND VGND VPWR VPWR _6425_/X sky130_fd_sc_hd__and2_1
XFILLER_161_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3568_ _6602_/Q _4124_/A _4112_/A _6592_/Q _3555_/X VGND VGND VPWR VPWR _3568_/X
+ sky130_fd_sc_hd__a221o_4
X_6356_ _6356_/A _6356_/B _6356_/C _6356_/D VGND VGND VPWR VPWR _6356_/X sky130_fd_sc_hd__or4_2
X_5307_ _5595_/A0 _6893_/Q _5314_/S VGND VGND VPWR VPWR _6893_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3499_ input7/X _3320_/Y _5200_/A _6809_/Q _3498_/X VGND VGND VPWR VPWR _3504_/C
+ sky130_fd_sc_hd__a221o_4
X_6287_ wire567/X wire642/X wire630/X wire560/X VGND VGND VPWR VPWR _6287_/X sky130_fd_sc_hd__a22o_1
X_5238_ _5238_/A _5594_/B VGND VGND VPWR VPWR _5241_/S sky130_fd_sc_hd__nand2_2
XFILLER_69_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5169_ _5169_/A _5169_/B _5169_/C VGND VGND VPWR VPWR _6783_/D sky130_fd_sc_hd__or3_1
XFILLER_29_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__1132_ clkbuf_0__1132_/X VGND VGND VPWR VPWR _6367_/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_193_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold6 hold6/A VGND VGND VPWR VPWR hold6/X sky130_fd_sc_hd__bufbuf_16
XFILLER_59_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4540_ _5140_/A _5140_/B _4520_/X VGND VGND VPWR VPWR _4542_/C sky130_fd_sc_hd__or3b_1
XFILLER_128_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold417 hold75/X VGND VGND VPWR VPWR hold417/X sky130_fd_sc_hd__bufbuf_16
XFILLER_183_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4471_ _4818_/B _4663_/B VGND VGND VPWR VPWR _4697_/A sky130_fd_sc_hd__or2_4
XFILLER_129_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire370 _3404_/X VGND VGND VPWR VPWR wire370/X sky130_fd_sc_hd__buf_6
Xwire381 wire381/A VGND VGND VPWR VPWR wire381/X sky130_fd_sc_hd__buf_8
XFILLER_7_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire392 _3384_/Y VGND VGND VPWR VPWR _5227_/A sky130_fd_sc_hd__buf_8
Xhold406 _6598_/Q VGND VGND VPWR VPWR hold406/X sky130_fd_sc_hd__bufbuf_16
XFILLER_143_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold439 _6554_/Q VGND VGND VPWR VPWR hold439/X sky130_fd_sc_hd__bufbuf_16
Xhold428 _5581_/X VGND VGND VPWR VPWR _7137_/D sky130_fd_sc_hd__bufbuf_16
X_7190_ _7190_/CLK _7190_/D fanout869/X VGND VGND VPWR VPWR _7190_/Q sky130_fd_sc_hd__dfrtp_1
X_3422_ _5234_/A _3543_/B VGND VGND VPWR VPWR _5200_/A sky130_fd_sc_hd__nor2_8
X_6210_ _7195_/Q _5665_/Y _6209_/X VGND VGND VPWR VPWR _7195_/D sky130_fd_sc_hd__o21a_1
X_6141_ wire476/X _6252_/B1 wire579/X _7033_/Q _6140_/X VGND VGND VPWR VPWR _6144_/C
+ sky130_fd_sc_hd__a221o_2
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _3365_/A _3353_/B VGND VGND VPWR VPWR _3353_/Y sky130_fd_sc_hd__nor2_8
X_6072_ _6886_/Q wire602/X wire581/X _7142_/Q _6062_/X VGND VGND VPWR VPWR _6072_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_112_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3284_ _3421_/A _3284_/B VGND VGND VPWR VPWR hold43/A sky130_fd_sc_hd__or2_4
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5023_ _5023_/A _5023_/B VGND VGND VPWR VPWR _5035_/D sky130_fd_sc_hd__nor2_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6974_ _6974_/CLK _6974_/D fanout875/X VGND VGND VPWR VPWR _6974_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_80_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5925_ wire572/X wire667/A wire665/X _6616_/Q VGND VGND VPWR VPWR _5925_/X sky130_fd_sc_hd__a22o_1
XFILLER_110_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5856_ _7100_/Q _5856_/A2 wire660/X wire531/X _5855_/X VGND VGND VPWR VPWR _5861_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_166_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4807_ _4980_/B _4980_/C _5132_/A _4806_/X _4917_/B VGND VGND VPWR VPWR _4807_/X
+ sky130_fd_sc_hd__o41a_2
X_5787_ _7179_/Q _6110_/S _5785_/X _5786_/X VGND VGND VPWR VPWR _7179_/D sky130_fd_sc_hd__o22a_1
X_4738_ _4758_/A _4758_/C _4737_/Y VGND VGND VPWR VPWR _4738_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_107_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4669_ _4697_/A _4687_/A _4724_/B _4886_/B VGND VGND VPWR VPWR _4669_/X sky130_fd_sc_hd__a31o_1
XFILLER_147_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6408_ _6408_/A0 hold698/X _6411_/S VGND VGND VPWR VPWR _7222_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6339_ _6757_/Q _6339_/A2 _6339_/B1 _6772_/Q VGND VGND VPWR VPWR _6339_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3971_ _3971_/A input1/X VGND VGND VPWR VPWR _3971_/X sky130_fd_sc_hd__and2_2
X_5710_ _6957_/Q wire707/X _5695_/X VGND VGND VPWR VPWR _5710_/X sky130_fd_sc_hd__a21o_1
XFILLER_188_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6690_ _6930_/CLK _6690_/D fanout887/X VGND VGND VPWR VPWR _6690_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5641_ _5663_/B _6012_/A _6032_/A _5621_/X _7167_/Q VGND VGND VPWR VPWR _7167_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_31_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5572_ _5572_/A0 hold503/X _5575_/S VGND VGND VPWR VPWR _5572_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4523_ _4671_/A _4990_/A VGND VGND VPWR VPWR _5114_/A sky130_fd_sc_hd__nor2_4
Xclkbuf_1_0_1_csclk clkbuf_1_0_1_csclk/A VGND VGND VPWR VPWR clkbuf_2_1_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
Xhold225 _6520_/Q VGND VGND VPWR VPWR hold225/X sky130_fd_sc_hd__bufbuf_16
Xhold203 _6939_/Q VGND VGND VPWR VPWR hold203/X sky130_fd_sc_hd__bufbuf_16
Xhold214 _6692_/Q VGND VGND VPWR VPWR hold214/X sky130_fd_sc_hd__bufbuf_16
Xhold269 _7153_/Q VGND VGND VPWR VPWR hold269/X sky130_fd_sc_hd__bufbuf_16
Xhold247 _7151_/Q VGND VGND VPWR VPWR hold247/X sky130_fd_sc_hd__bufbuf_16
X_4454_ _4584_/A _4663_/B VGND VGND VPWR VPWR _4745_/A sky130_fd_sc_hd__or2_4
XFILLER_132_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold236 _3250_/X VGND VGND VPWR VPWR hold236/X sky130_fd_sc_hd__bufbuf_16
Xhold258 _5525_/X VGND VGND VPWR VPWR _7087_/D sky130_fd_sc_hd__bufbuf_16
X_4385_ _5023_/A _4871_/A VGND VGND VPWR VPWR _5164_/A sky130_fd_sc_hd__and2_4
XFILLER_132_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3405_ _7011_/Q _5432_/A _3995_/A _6502_/Q wire370/X VGND VGND VPWR VPWR _3405_/X
+ sky130_fd_sc_hd__a221o_4
X_7173_ _7194_/CLK _7173_/D fanout867/X VGND VGND VPWR VPWR _7173_/Q sky130_fd_sc_hd__dfrtp_2
X_6124_ _3206_/A wire598/X wire610/X _3221_/A _6123_/X VGND VGND VPWR VPWR _6132_/B
+ sky130_fd_sc_hd__a221o_1
Xfanout738 wire742/X VGND VGND VPWR VPWR wire739/A sky130_fd_sc_hd__buf_8
XFILLER_86_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout727 hold141/X VGND VGND VPWR VPWR hold142/A sky130_fd_sc_hd__buf_6
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3336_ _7044_/Q _5468_/A _3335_/Y _6495_/Q VGND VGND VPWR VPWR _3336_/X sky130_fd_sc_hd__a22o_1
XFILLER_112_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6055_ _6909_/Q wire632/X wire579/X wire511/X VGND VGND VPWR VPWR _6055_/X sky130_fd_sc_hd__a22o_2
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _4832_/A _4728_/X _5050_/C VGND VGND VPWR VPWR _5008_/A sky130_fd_sc_hd__a21o_1
XFILLER_100_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3267_ hold42/X _3284_/B VGND VGND VPWR VPWR _3267_/Y sky130_fd_sc_hd__nand2_2
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3198_ _6677_/Q VGND VGND VPWR VPWR _5626_/A sky130_fd_sc_hd__inv_2
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_109 _6306_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6957_ _7153_/CLK _6957_/D fanout882/X VGND VGND VPWR VPWR _6957_/Q sky130_fd_sc_hd__dfstp_4
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6888_ _7154_/CLK _6888_/D fanout886/X VGND VGND VPWR VPWR _6888_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_167_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5908_ _6660_/Q _5974_/A2 wire671/X _5899_/X VGND VGND VPWR VPWR _5908_/X sky130_fd_sc_hd__a22o_1
XFILLER_14_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5839_ _5839_/A _5839_/B _5839_/C _5839_/D VGND VGND VPWR VPWR _5839_/X sky130_fd_sc_hd__or4_4
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length704 _5675_/X VGND VGND VPWR VPWR _5857_/A2 sky130_fd_sc_hd__buf_6
Xmax_length726 _5236_/B VGND VGND VPWR VPWR _4154_/B sky130_fd_sc_hd__buf_8
XFILLER_14_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold770 _6713_/Q VGND VGND VPWR VPWR hold770/X sky130_fd_sc_hd__bufbuf_16
XFILLER_150_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold781 _6687_/Q VGND VGND VPWR VPWR hold781/X sky130_fd_sc_hd__bufbuf_16
Xhold792 _7135_/Q VGND VGND VPWR VPWR hold792/X sky130_fd_sc_hd__bufbuf_16
XFILLER_77_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput308 _3423_/X VGND VGND VPWR VPWR serial_data_1 sky130_fd_sc_hd__buf_8
XFILLER_114_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput319 _6570_/Q VGND VGND VPWR VPWR wb_dat_o[10] sky130_fd_sc_hd__buf_8
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4170_ _5249_/A0 hold447/X _4171_/S VGND VGND VPWR VPWR _6637_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6811_ _6815_/CLK _6811_/D fanout855/X VGND VGND VPWR VPWR _6811_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_35_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6742_ _6806_/CLK _6742_/D _6435_/A VGND VGND VPWR VPWR _6742_/Q sky130_fd_sc_hd__dfrtp_2
X_3954_ _3953_/A _3954_/A2 _6455_/B _3953_/Y VGND VGND VPWR VPWR _3954_/X sky130_fd_sc_hd__a22o_2
X_6673_ _7133_/CLK _6673_/D fanout881/X VGND VGND VPWR VPWR _6673_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_188_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3885_ _4351_/C _4351_/D _4350_/A _4350_/B VGND VGND VPWR VPWR _3886_/C sky130_fd_sc_hd__or4_1
XFILLER_176_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5624_ _6679_/Q _5702_/B VGND VGND VPWR VPWR _5629_/B sky130_fd_sc_hd__nand2_1
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5555_ hold505/X _5600_/A0 _5557_/S VGND VGND VPWR VPWR _5555_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4506_ _4502_/A _4749_/C _5164_/B _4812_/A VGND VGND VPWR VPWR _4506_/X sky130_fd_sc_hd__a31o_1
X_5486_ _5486_/A _5594_/B VGND VGND VPWR VPWR _5486_/Y sky130_fd_sc_hd__nand2_8
X_4437_ _4529_/B _4529_/C VGND VGND VPWR VPWR _4438_/B sky130_fd_sc_hd__nand2_4
X_7225_ _7225_/CLK _7225_/D fanout850/X VGND VGND VPWR VPWR _7225_/Q sky130_fd_sc_hd__dfrtp_2
X_7156_ _7156_/CLK _7156_/D fanout889/X VGND VGND VPWR VPWR _7156_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_116_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4368_ _4368_/A _4722_/A VGND VGND VPWR VPWR _4650_/B sky130_fd_sc_hd__or2_4
X_6107_ _6306_/A _6107_/B _6107_/C VGND VGND VPWR VPWR _6107_/X sky130_fd_sc_hd__or3_4
XFILLER_86_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4299_ wire799/A hold560/X _4303_/S VGND VGND VPWR VPWR _6748_/D sky130_fd_sc_hd__mux2_1
X_3319_ _3367_/A hold95/X VGND VGND VPWR VPWR _3375_/B sky130_fd_sc_hd__or2_4
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7087_ _7129_/CLK _7087_/D fanout863/X VGND VGND VPWR VPWR _7087_/Q sky130_fd_sc_hd__dfrtp_2
X_6038_ wire487/X wire631/X wire616/X wire493/X VGND VGND VPWR VPWR _6038_/X sky130_fd_sc_hd__a22o_2
XFILLER_100_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire903 wire904/X VGND VGND VPWR VPWR wire903/X sky130_fd_sc_hd__buf_6
XFILLER_10_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length523 hold623/X VGND VGND VPWR VPWR wire522/A sky130_fd_sc_hd__buf_6
XFILLER_108_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_64_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7103_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_41_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length545 _6880_/Q VGND VGND VPWR VPWR _3194_/A sky130_fd_sc_hd__buf_6
XFILLER_108_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length578 wire579/X VGND VGND VPWR VPWR _6339_/B1 sky130_fd_sc_hd__buf_6
XFILLER_150_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_79_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6806_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_123_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_17_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _6747_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3670_ wire555/X _3295_/Y _3327_/Y wire529/X VGND VGND VPWR VPWR _3670_/X sky130_fd_sc_hd__a22o_1
XFILLER_40_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5340_ hold256/X hold57/X _5341_/S VGND VGND VPWR VPWR _6923_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5271_ _5595_/A0 _6861_/Q _5278_/S VGND VGND VPWR VPWR _6861_/D sky130_fd_sc_hd__mux2_1
XFILLER_126_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7010_ _7107_/CLK _7010_/D fanout865/X VGND VGND VPWR VPWR _7010_/Q sky130_fd_sc_hd__dfrtp_2
X_4222_ hold550/X _6408_/A0 _4232_/S VGND VGND VPWR VPWR _4222_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4153_ hold327/X _5599_/A0 _4153_/S VGND VGND VPWR VPWR _6623_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4084_ hold643/X wire794/X _4087_/S VGND VGND VPWR VPWR _6564_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4986_ _4986_/A _4986_/B _4986_/C VGND VGND VPWR VPWR _4997_/B sky130_fd_sc_hd__and3_4
XFILLER_63_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6725_ _6833_/CLK _6725_/D fanout873/X VGND VGND VPWR VPWR _6725_/Q sky130_fd_sc_hd__dfstp_4
X_3937_ _6508_/Q wire904/X _3939_/S VGND VGND VPWR VPWR _3937_/X sky130_fd_sc_hd__mux2_2
XFILLER_137_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3868_ _6465_/Q hold19/A _3874_/S VGND VGND VPWR VPWR _6466_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6656_ _6787_/CLK _6656_/D fanout854/X VGND VGND VPWR VPWR _6656_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_191_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5607_ _7157_/Q _5615_/D VGND VGND VPWR VPWR _5609_/B sky130_fd_sc_hd__nand2_1
X_3799_ _6486_/Q _3801_/B VGND VGND VPWR VPWR _3802_/A sky130_fd_sc_hd__nand2_1
X_6587_ _7208_/CLK _6587_/D VGND VGND VPWR VPWR _6587_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5538_ wire746/X hold736/X _5538_/S VGND VGND VPWR VPWR _7099_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7208_ _7208_/CLK _7208_/D VGND VGND VPWR VPWR _7208_/Q sky130_fd_sc_hd__dfxtp_4
X_5469_ wire802/X hold552/X _5476_/S VGND VGND VPWR VPWR _7037_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7139_ _7139_/CLK _7139_/D fanout868/X VGND VGND VPWR VPWR _7139_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_101_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire700 wire701/X VGND VGND VPWR VPWR wire700/X sky130_fd_sc_hd__buf_8
XFILLER_183_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire711 _5653_/X VGND VGND VPWR VPWR wire711/X sky130_fd_sc_hd__buf_8
Xinput18 mask_rev_in[22] VGND VGND VPWR VPWR input18/X sky130_fd_sc_hd__clkbuf_4
Xinput29 mask_rev_in[3] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__clkbuf_4
XFILLER_10_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire799 wire799/A VGND VGND VPWR VPWR _5234_/C sky130_fd_sc_hd__buf_6
XFILLER_184_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_270 _6670_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4840_ _4840_/A _4957_/A VGND VGND VPWR VPWR _5046_/A sky130_fd_sc_hd__or2_2
XFILLER_45_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_281 hold575/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_292 _3331_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6510_ _6931_/CLK _6510_/D fanout885/X VGND VGND VPWR VPWR _6510_/Q sky130_fd_sc_hd__dfrtp_2
X_4771_ _4986_/B _5031_/B VGND VGND VPWR VPWR _4806_/B sky130_fd_sc_hd__nor2_1
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3722_ _7030_/Q _5459_/A _5423_/A _6998_/Q _3721_/X VGND VGND VPWR VPWR _3725_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6441_ _6446_/A _6447_/B VGND VGND VPWR VPWR _6441_/X sky130_fd_sc_hd__and2_1
X_3653_ _7087_/Q _5522_/A _3978_/A _6490_/Q _3652_/X VGND VGND VPWR VPWR _3654_/D
+ sky130_fd_sc_hd__a221o_1
X_6372_ _6372_/A _6372_/B VGND VGND VPWR VPWR _6372_/Y sky130_fd_sc_hd__nand2_1
X_5323_ wire742/X hold309/X _5323_/S VGND VGND VPWR VPWR _6908_/D sky130_fd_sc_hd__mux2_1
X_3584_ input55/X wire427/A _4154_/A _6627_/Q _3583_/X VGND VGND VPWR VPWR _3587_/C
+ sky130_fd_sc_hd__a221o_4
XFILLER_142_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5254_ _6408_/A0 hold550/X _5260_/S VGND VGND VPWR VPWR _5254_/X sky130_fd_sc_hd__mux2_1
X_4205_ _6691_/Q hold38/A _4209_/S VGND VGND VPWR VPWR _4205_/X sky130_fd_sc_hd__mux2_1
X_5185_ _5185_/A _6406_/B VGND VGND VPWR VPWR _5190_/S sky130_fd_sc_hd__nand2_4
X_4136_ _4136_/A _5378_/B VGND VGND VPWR VPWR _4141_/S sky130_fd_sc_hd__nand2_4
Xclkbuf_3_6_0_csclk clkbuf_3_7_0_csclk/A VGND VGND VPWR VPWR _6987_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_113_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4067_ _4067_/A _4154_/B VGND VGND VPWR VPWR _4067_/Y sky130_fd_sc_hd__nand2_8
XFILLER_71_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4969_ _4949_/B _4571_/Y _4959_/A _4905_/B VGND VGND VPWR VPWR _4973_/C sky130_fd_sc_hd__a31o_2
X_6708_ _6708_/CLK _6708_/D fanout873/X VGND VGND VPWR VPWR _6708_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_137_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6639_ _6642_/CLK _6639_/D fanout856/X VGND VGND VPWR VPWR _6639_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire541 _6900_/Q VGND VGND VPWR VPWR wire541/X sky130_fd_sc_hd__buf_6
Xwire530 _6943_/Q VGND VGND VPWR VPWR wire530/X sky130_fd_sc_hd__buf_6
Xwire552 _6868_/Q VGND VGND VPWR VPWR wire552/X sky130_fd_sc_hd__buf_8
XFILLER_171_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire585 _6014_/Y VGND VGND VPWR VPWR wire585/X sky130_fd_sc_hd__buf_8
XFILLER_7_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire563 _6750_/Q VGND VGND VPWR VPWR wire563/X sky130_fd_sc_hd__buf_6
XFILLER_155_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire596 _6002_/Y VGND VGND VPWR VPWR _6021_/B sky130_fd_sc_hd__buf_8
XFILLER_143_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6990_ _7118_/CLK _6990_/D fanout869/X VGND VGND VPWR VPWR _6990_/Q sky130_fd_sc_hd__dfstp_2
X_5941_ _6592_/Q _5977_/A2 wire667/X _6538_/Q VGND VGND VPWR VPWR _5941_/X sky130_fd_sc_hd__a22o_1
XFILLER_93_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5872_ _6860_/Q _5698_/Y _5861_/X _5871_/X _6109_/S VGND VGND VPWR VPWR _5872_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4823_ _5164_/B _5017_/A _4756_/B _4898_/B VGND VGND VPWR VPWR _4823_/X sky130_fd_sc_hd__o22a_2
XFILLER_61_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4754_ _4898_/B _4754_/B VGND VGND VPWR VPWR _4950_/B sky130_fd_sc_hd__nor2_4
X_3705_ _6894_/Q _5306_/A _4136_/A _6610_/Q _3704_/X VGND VGND VPWR VPWR _3709_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4685_ _4685_/A _4746_/B VGND VGND VPWR VPWR _5017_/A sky130_fd_sc_hd__or2_4
XFILLER_161_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3636_ _3636_/A _3636_/B _3636_/C _3636_/D VGND VGND VPWR VPWR _3665_/A sky130_fd_sc_hd__or4_4
X_6424_ _6455_/A _6455_/B VGND VGND VPWR VPWR _6424_/X sky130_fd_sc_hd__and2_1
X_3567_ _3233_/A wire424/X _5387_/A _6968_/Q _3554_/X VGND VGND VPWR VPWR _3567_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_108_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6355_ _6355_/A _6355_/B _6355_/C _6355_/D VGND VGND VPWR VPWR _6356_/D sky130_fd_sc_hd__or4_1
X_5306_ _5306_/A _5594_/B VGND VGND VPWR VPWR _5314_/S sky130_fd_sc_hd__nand2_8
X_6286_ _6616_/Q wire636/X wire634/X _6601_/Q VGND VGND VPWR VPWR _6286_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5237_ _5487_/A0 hold798/X _5237_/S VGND VGND VPWR VPWR _6833_/D sky130_fd_sc_hd__mux2_1
X_3498_ _6993_/Q _5414_/A _6406_/A _7225_/Q VGND VGND VPWR VPWR _3498_/X sky130_fd_sc_hd__a22o_2
X_5168_ _6783_/Q _5156_/A _5155_/X _5158_/Y _5167_/X VGND VGND VPWR VPWR _5169_/C
+ sky130_fd_sc_hd__a221o_2
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5099_ _5099_/A _5099_/B _5099_/C VGND VGND VPWR VPWR _5101_/C sky130_fd_sc_hd__or3_1
X_4119_ hold641/X wire799/A _4123_/S VGND VGND VPWR VPWR _6594_/D sky130_fd_sc_hd__mux2_1
XFILLER_140_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold7 hold7/A VGND VGND VPWR VPWR hold7/X sky130_fd_sc_hd__bufbuf_16
XFILLER_121_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire360 _5521_/S VGND VGND VPWR VPWR _5517_/S sky130_fd_sc_hd__buf_4
X_4470_ _4740_/A _4470_/B VGND VGND VPWR VPWR _5005_/A sky130_fd_sc_hd__nand2_4
Xhold418 _3985_/X VGND VGND VPWR VPWR hold80/A sky130_fd_sc_hd__bufbuf_16
Xhold407 _6671_/Q VGND VGND VPWR VPWR hold407/X sky130_fd_sc_hd__bufbuf_16
Xwire371 _6082_/X VGND VGND VPWR VPWR _6083_/C sky130_fd_sc_hd__buf_4
XFILLER_143_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire382 hold90/X VGND VGND VPWR VPWR _5575_/S sky130_fd_sc_hd__buf_6
XFILLER_128_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire393 _3374_/Y VGND VGND VPWR VPWR _5279_/A sky130_fd_sc_hd__buf_8
XFILLER_171_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold429 _6633_/Q VGND VGND VPWR VPWR hold429/X sky130_fd_sc_hd__bufbuf_16
X_3421_ _3421_/A _3421_/B _3421_/C VGND VGND VPWR VPWR _3543_/B sky130_fd_sc_hd__or3_4
XFILLER_171_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6140_ _7001_/Q wire604/X _6140_/B1 _6921_/Q VGND VGND VPWR VPWR _6140_/X sky130_fd_sc_hd__a22o_1
X_3352_ hold63/X _3543_/A VGND VGND VPWR VPWR _3352_/Y sky130_fd_sc_hd__nor2_4
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6071_ _6071_/A _6071_/B _6071_/C _6071_/D VGND VGND VPWR VPWR _6071_/X sky130_fd_sc_hd__or4_1
X_3283_ _5225_/A _3534_/A VGND VGND VPWR VPWR _3283_/Y sky130_fd_sc_hd__nor2_8
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _5022_/A _5022_/B _5022_/C _5022_/D VGND VGND VPWR VPWR _5180_/C sky130_fd_sc_hd__or4_2
XFILLER_100_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6973_ _6974_/CLK _6973_/D fanout875/X VGND VGND VPWR VPWR _6973_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5924_ wire571/X _5681_/X _5923_/X VGND VGND VPWR VPWR _5927_/C sky130_fd_sc_hd__a21o_1
XFILLER_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5855_ _7020_/Q wire697/X _5855_/B1 _7036_/Q VGND VGND VPWR VPWR _5855_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4806_ _5142_/A _4806_/B _5099_/B _4806_/D VGND VGND VPWR VPWR _4806_/X sky130_fd_sc_hd__or4_1
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5786_ _5611_/A _7178_/Q wire381/A VGND VGND VPWR VPWR _5786_/X sky130_fd_sc_hd__a21o_1
X_4737_ _4898_/B _5062_/C VGND VGND VPWR VPWR _4737_/Y sky130_fd_sc_hd__nor2_4
XFILLER_147_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4668_ _4692_/C _4668_/B VGND VGND VPWR VPWR _4886_/B sky130_fd_sc_hd__nand2_8
XFILLER_135_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3619_ wire528/X wire421/A wire401/X wire530/X VGND VGND VPWR VPWR _3619_/X sky130_fd_sc_hd__a22o_1
XFILLER_79_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6407_ _6407_/A0 hold766/X _6411_/S VGND VGND VPWR VPWR _7221_/D sky130_fd_sc_hd__mux2_1
XFILLER_162_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4599_ _4622_/B _4868_/A VGND VGND VPWR VPWR _4893_/A sky130_fd_sc_hd__nand2_2
XFILLER_103_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6338_ wire569/X _6311_/B _6036_/Y _6752_/Q _6335_/X VGND VGND VPWR VPWR _6343_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6269_ _6269_/A _6269_/B _6269_/C _6269_/D VGND VGND VPWR VPWR _6269_/X sky130_fd_sc_hd__or4_1
XFILLER_88_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_3_0_csclk clkbuf_2_3_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_7_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_28_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3970_ _3970_/A _3970_/B VGND VGND VPWR VPWR _3970_/X sky130_fd_sc_hd__and2_2
XFILLER_16_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5640_ _7167_/Q _7166_/Q VGND VGND VPWR VPWR _6032_/A sky130_fd_sc_hd__and2b_4
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5571_ hold83/A _7128_/Q hold91/X VGND VGND VPWR VPWR hold92/A sky130_fd_sc_hd__mux2_1
X_4522_ _5023_/A _4871_/A _4617_/A VGND VGND VPWR VPWR _5022_/A sky130_fd_sc_hd__a21oi_2
XFILLER_116_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold226 _4032_/X VGND VGND VPWR VPWR _6520_/D sky130_fd_sc_hd__bufbuf_16
Xhold204 _5358_/X VGND VGND VPWR VPWR _6939_/D sky130_fd_sc_hd__bufbuf_16
Xhold215 _4244_/X VGND VGND VPWR VPWR _6692_/D sky130_fd_sc_hd__bufbuf_16
X_4453_ _4584_/A _4663_/B VGND VGND VPWR VPWR _4453_/Y sky130_fd_sc_hd__nor2_8
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold248 _5597_/X VGND VGND VPWR VPWR _7151_/D sky130_fd_sc_hd__bufbuf_16
X_3404_ _7115_/Q _5549_/A hold65/A _7155_/Q VGND VGND VPWR VPWR _3404_/X sky130_fd_sc_hd__a22o_4
XFILLER_144_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold259 _7095_/Q VGND VGND VPWR VPWR hold259/X sky130_fd_sc_hd__bufbuf_16
Xhold237 _3251_/X VGND VGND VPWR VPWR hold237/X sky130_fd_sc_hd__bufbuf_16
X_4384_ _5031_/A _4584_/A VGND VGND VPWR VPWR _4871_/A sky130_fd_sc_hd__or2_4
X_7172_ _7194_/CLK _7172_/D fanout866/X VGND VGND VPWR VPWR _7172_/Q sky130_fd_sc_hd__dfrtp_1
X_6123_ _6888_/Q wire602/X wire581/X _7144_/Q _6122_/X VGND VGND VPWR VPWR _6123_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3335_ _5225_/A hold96/X VGND VGND VPWR VPWR _3335_/Y sky130_fd_sc_hd__nor2_4
XFILLER_140_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6054_ _6925_/Q wire634/X _6010_/Y _7021_/Q _6053_/X VGND VGND VPWR VPWR _6057_/C
+ sky130_fd_sc_hd__a221o_4
XFILLER_100_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3266_ _3953_/A hold174/X hold110/X VGND VGND VPWR VPWR _3266_/Y sky130_fd_sc_hd__a21oi_4
X_5005_ _5005_/A _5062_/A _5005_/C VGND VGND VPWR VPWR _5050_/C sky130_fd_sc_hd__and3_4
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3197_ _5611_/A VGND VGND VPWR VPWR _3197_/Y sky130_fd_sc_hd__inv_8
XFILLER_26_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6956_ _6980_/CLK hold22/X fanout878/X VGND VGND VPWR VPWR _6956_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5907_ _6635_/Q _5973_/A2 wire692/X _6724_/Q _5906_/X VGND VGND VPWR VPWR _5910_/C
+ sky130_fd_sc_hd__a221o_1
X_6887_ _7111_/CLK _6887_/D fanout881/X VGND VGND VPWR VPWR _6887_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_14_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5838_ _6963_/Q _5673_/X _5699_/X _6931_/Q _5837_/X VGND VGND VPWR VPWR _5839_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_167_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length705 _5674_/X VGND VGND VPWR VPWR _5934_/B1 sky130_fd_sc_hd__buf_6
X_5769_ wire522/A _5667_/X _5687_/X _3216_/A VGND VGND VPWR VPWR _5769_/X sky130_fd_sc_hd__a22o_1
XFILLER_135_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold760 _6720_/Q VGND VGND VPWR VPWR hold760/X sky130_fd_sc_hd__bufbuf_16
XFILLER_122_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold771 _6753_/Q VGND VGND VPWR VPWR hold771/X sky130_fd_sc_hd__bufbuf_16
Xhold782 _4233_/X VGND VGND VPWR VPWR _6687_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_150_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold793 _6639_/Q VGND VGND VPWR VPWR hold793/X sky130_fd_sc_hd__bufbuf_16
XFILLER_162_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput309 _3385_/X VGND VGND VPWR VPWR serial_data_2 sky130_fd_sc_hd__buf_8
XFILLER_5_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6810_ _6810_/CLK _6810_/D fanout853/X VGND VGND VPWR VPWR _6810_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_63_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6741_ _6806_/CLK _6741_/D _6435_/A VGND VGND VPWR VPWR _6741_/Q sky130_fd_sc_hd__dfrtp_2
X_3953_ _3953_/A _3953_/B VGND VGND VPWR VPWR _3953_/Y sky130_fd_sc_hd__nor2_2
XFILLER_50_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6672_ _7122_/CLK _6672_/D fanout887/X VGND VGND VPWR VPWR _6672_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_31_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3884_ _6472_/Q _6456_/Q _6425_/B VGND VGND VPWR VPWR _3974_/B sky130_fd_sc_hd__o21ai_4
XFILLER_149_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5623_ _7162_/Q _7161_/Q VGND VGND VPWR VPWR _5702_/B sky130_fd_sc_hd__nor2_8
X_5554_ hold399/X _5599_/A0 _5557_/S VGND VGND VPWR VPWR _5554_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4505_ _4812_/A _4687_/A VGND VGND VPWR VPWR _4505_/X sky130_fd_sc_hd__or2_4
XFILLER_160_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5485_ hold667/X wire739/X _5485_/S VGND VGND VPWR VPWR _7052_/D sky130_fd_sc_hd__mux2_1
X_4436_ _4696_/A _4436_/B _4446_/B VGND VGND VPWR VPWR _4529_/C sky130_fd_sc_hd__and3_4
XFILLER_116_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7224_ _7225_/CLK _7224_/D fanout850/X VGND VGND VPWR VPWR _7224_/Q sky130_fd_sc_hd__dfrtp_2
X_7155_ _7155_/CLK _7155_/D fanout884/X VGND VGND VPWR VPWR _7155_/Q sky130_fd_sc_hd__dfrtp_2
X_4367_ _4728_/A _4478_/B _4502_/A _4236_/B VGND VGND VPWR VPWR _4367_/X sky130_fd_sc_hd__o31a_4
XFILLER_116_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6106_ _6106_/A _6106_/B _6106_/C _6106_/D VGND VGND VPWR VPWR _6107_/C sky130_fd_sc_hd__or4_2
XFILLER_86_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3318_ _6860_/Q _5261_/A wire430/X _7068_/Q VGND VGND VPWR VPWR _3318_/X sky130_fd_sc_hd__a22o_1
XFILLER_112_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7086_ _7129_/CLK _7086_/D fanout863/X VGND VGND VPWR VPWR _7086_/Q sky130_fd_sc_hd__dfstp_4
X_4298_ _4298_/A _6406_/B VGND VGND VPWR VPWR _4303_/S sky130_fd_sc_hd__nand2_4
XFILLER_132_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6037_ _6037_/A _6037_/B _6037_/C VGND VGND VPWR VPWR _6037_/X sky130_fd_sc_hd__and3_4
X_3249_ _3845_/A _3249_/B VGND VGND VPWR VPWR _3249_/Y sky130_fd_sc_hd__nand2b_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6939_ _7147_/CLK _6939_/D fanout888/X VGND VGND VPWR VPWR _6939_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire915 wire915/A VGND VGND VPWR VPWR wire915/X sky130_fd_sc_hd__buf_8
Xwire904 wire904/A VGND VGND VPWR VPWR wire904/X sky130_fd_sc_hd__buf_8
XFILLER_155_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0_csclk _3954_/X VGND VGND VPWR VPWR clkbuf_0_csclk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_150_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold590 _6996_/Q VGND VGND VPWR VPWR hold590/X sky130_fd_sc_hd__bufbuf_16
XFILLER_173_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_1_0_1_csclk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5270_ _5270_/A _5594_/B VGND VGND VPWR VPWR _5270_/Y sky130_fd_sc_hd__nand2_8
XFILLER_141_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4221_ hold734/X _4220_/X _4235_/S VGND VGND VPWR VPWR _4221_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4152_ hold194/X hold83/X _4153_/S VGND VGND VPWR VPWR _6622_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4083_ hold790/X _5487_/A0 _4087_/S VGND VGND VPWR VPWR _6563_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4985_ _4507_/A _5004_/B _4842_/X VGND VGND VPWR VPWR _4985_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_177_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6724_ _6724_/CLK _6724_/D wire860/X VGND VGND VPWR VPWR _6724_/Q sky130_fd_sc_hd__dfrtp_2
X_3936_ _6842_/Q input81/X _3970_/B VGND VGND VPWR VPWR _3936_/X sky130_fd_sc_hd__mux2_4
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_2_0_csclk clkbuf_3_3_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_2_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_137_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6655_ _6806_/CLK _6655_/D fanout848/X VGND VGND VPWR VPWR _6655_/Q sky130_fd_sc_hd__dfrtp_2
X_3867_ _3875_/B _3864_/B _3861_/B _6467_/Q _3866_/X VGND VGND VPWR VPWR _6467_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_192_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5606_ _6680_/Q _5606_/B _5665_/B VGND VGND VPWR VPWR _5617_/A sky130_fd_sc_hd__or3_2
X_3798_ _6664_/Q _3797_/X _6485_/Q VGND VGND VPWR VPWR _3801_/B sky130_fd_sc_hd__o21a_1
X_6586_ _7208_/CLK _6586_/D VGND VGND VPWR VPWR _6586_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_191_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5537_ wire753/X hold822/X _5538_/S VGND VGND VPWR VPWR _7098_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7207_ _7210_/CLK _7207_/D VGND VGND VPWR VPWR _7207_/Q sky130_fd_sc_hd__dfxtp_4
X_5468_ _5468_/A _5576_/B VGND VGND VPWR VPWR _5476_/S sky130_fd_sc_hd__nand2_8
X_4419_ _4707_/B _4773_/A VGND VGND VPWR VPWR _4426_/A sky130_fd_sc_hd__nand2_1
X_5399_ hold724/X _5498_/A0 _5404_/S VGND VGND VPWR VPWR _6975_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7138_ _7139_/CLK _7138_/D fanout867/X VGND VGND VPWR VPWR _7138_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_143_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7069_ _7132_/CLK _7069_/D fanout863/X VGND VGND VPWR VPWR _7069_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_47_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire701 _5678_/X VGND VGND VPWR VPWR wire701/X sky130_fd_sc_hd__buf_8
Xwire712 _5653_/X VGND VGND VPWR VPWR wire712/X sky130_fd_sc_hd__buf_8
Xinput19 mask_rev_in[23] VGND VGND VPWR VPWR input19/X sky130_fd_sc_hd__clkbuf_4
XFILLER_183_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire756 wire757/X VGND VGND VPWR VPWR wire756/X sky130_fd_sc_hd__buf_6
XFILLER_182_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length398 _5576_/A VGND VGND VPWR VPWR _3763_/B1 sky130_fd_sc_hd__buf_6
XFILLER_2_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_260 _3202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_282 hold575/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_271 hold514/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_293 _3522_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4770_ _5087_/A _5087_/C _5165_/A VGND VGND VPWR VPWR _5035_/B sky130_fd_sc_hd__o21a_2
XFILLER_158_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3721_ _6497_/Q _3995_/A _4262_/A _6719_/Q VGND VGND VPWR VPWR _3721_/X sky130_fd_sc_hd__a22o_2
XFILLER_174_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3652_ wire482/X _5540_/A _3551_/Y wire834/X VGND VGND VPWR VPWR _3652_/X sky130_fd_sc_hd__a22o_1
X_6440_ _6446_/A _6447_/B VGND VGND VPWR VPWR _6440_/X sky130_fd_sc_hd__and2_1
X_6371_ _6372_/A _6371_/B VGND VGND VPWR VPWR _6371_/Y sky130_fd_sc_hd__nand2_1
XFILLER_173_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3583_ _7128_/Q _3583_/A2 _4160_/A _6632_/Q VGND VGND VPWR VPWR _3583_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5322_ hold57/X hold250/X _5323_/S VGND VGND VPWR VPWR _6907_/D sky130_fd_sc_hd__mux2_1
XFILLER_5_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5253_ _6407_/A0 hold543/X _5260_/S VGND VGND VPWR VPWR _5253_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4204_ hold808/X _4203_/X _4218_/S VGND VGND VPWR VPWR _4204_/X sky130_fd_sc_hd__mux2_1
X_5184_ _5184_/A _5184_/B VGND VGND VPWR VPWR _6784_/D sky130_fd_sc_hd__or2_1
X_4135_ _4303_/A0 hold448/X _4135_/S VGND VGND VPWR VPWR _6608_/D sky130_fd_sc_hd__mux2_1
XFILLER_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_63_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7105_/CLK sky130_fd_sc_hd__clkbuf_8
X_4066_ _5599_/A0 hold336/X _4066_/S VGND VGND VPWR VPWR _6549_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_78_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6810_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_24_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4968_ _4537_/X _4959_/A _4959_/B _4906_/B VGND VGND VPWR VPWR _5071_/D sky130_fd_sc_hd__a31o_2
X_4899_ _4965_/A _4899_/B VGND VGND VPWR VPWR _4976_/A sky130_fd_sc_hd__nor2_1
X_6707_ _7210_/CLK _6707_/D _6362_/B VGND VGND VPWR VPWR _6707_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3919_ _6832_/Q _5626_/A _3918_/X VGND VGND VPWR VPWR _6677_/D sky130_fd_sc_hd__o21ai_1
XFILLER_165_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6638_ _6752_/CLK _6638_/D fanout857/X VGND VGND VPWR VPWR _6638_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_137_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6569_ _7208_/CLK _6569_/D VGND VGND VPWR VPWR _6569_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_16_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _6844_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_145_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire531 _6940_/Q VGND VGND VPWR VPWR wire531/X sky130_fd_sc_hd__buf_6
XFILLER_156_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire542 _6899_/Q VGND VGND VPWR VPWR wire542/X sky130_fd_sc_hd__buf_6
XFILLER_11_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire520 _7005_/Q VGND VGND VPWR VPWR wire520/X sky130_fd_sc_hd__buf_6
Xwire564 _6747_/Q VGND VGND VPWR VPWR wire564/X sky130_fd_sc_hd__buf_6
XFILLER_156_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire553 _6867_/Q VGND VGND VPWR VPWR wire553/X sky130_fd_sc_hd__buf_6
Xwire575 _6036_/Y VGND VGND VPWR VPWR wire575/X sky130_fd_sc_hd__buf_8
XFILLER_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire597 _6023_/A VGND VGND VPWR VPWR wire597/X sky130_fd_sc_hd__buf_8
XFILLER_170_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5940_ _7186_/Q _6309_/S _5938_/X _5939_/X VGND VGND VPWR VPWR _7186_/D sky130_fd_sc_hd__o22a_1
XFILLER_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5871_ _5871_/A _5871_/B _5871_/C _5871_/D VGND VGND VPWR VPWR _5871_/X sky130_fd_sc_hd__or4_1
XFILLER_34_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4822_ _4956_/C _4684_/Y _4653_/Y VGND VGND VPWR VPWR _5047_/C sky130_fd_sc_hd__a21o_1
X_4753_ _4753_/A _4753_/B _4753_/C _4753_/D VGND VGND VPWR VPWR _4753_/X sky130_fd_sc_hd__and4_2
X_3704_ wire546/X wire406/X _4148_/A _6620_/Q VGND VGND VPWR VPWR _3704_/X sky130_fd_sc_hd__a22o_2
X_4684_ _4685_/A _4746_/B VGND VGND VPWR VPWR _4684_/Y sky130_fd_sc_hd__nor2_2
XFILLER_146_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6423_ _6455_/A _6455_/B VGND VGND VPWR VPWR _6423_/X sky130_fd_sc_hd__and2_1
X_3635_ _3635_/A _3635_/B _3635_/C _3635_/D VGND VGND VPWR VPWR _3636_/D sky130_fd_sc_hd__or4_1
XFILLER_134_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3566_ _6936_/Q _3356_/Y _4256_/A _6716_/Q VGND VGND VPWR VPWR _3588_/A sky130_fd_sc_hd__a22o_2
X_6354_ _6717_/Q wire640/X wire638/X _6549_/Q _6353_/X VGND VGND VPWR VPWR _6355_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5305_ _5602_/A0 hold286/X _5305_/S VGND VGND VPWR VPWR _6892_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6285_ _7198_/Q _6309_/S _6284_/X VGND VGND VPWR VPWR _7198_/D sky130_fd_sc_hd__o21a_1
X_3497_ _3508_/A _3520_/B VGND VGND VPWR VPWR _6406_/A sky130_fd_sc_hd__nor2_8
XFILLER_130_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5236_ _5236_/A _5236_/B VGND VGND VPWR VPWR _5237_/S sky130_fd_sc_hd__nand2_1
XFILLER_124_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5167_ _5101_/B _5163_/X _5166_/X _5161_/X VGND VGND VPWR VPWR _5167_/X sky130_fd_sc_hd__o31a_2
XFILLER_69_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5098_ _5098_/A _5098_/B _5098_/C VGND VGND VPWR VPWR _5101_/B sky130_fd_sc_hd__or3_2
XFILLER_84_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4118_ _4118_/A _5242_/B VGND VGND VPWR VPWR _4123_/S sky130_fd_sc_hd__and2_4
XFILLER_56_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4049_ _4049_/A _6406_/B VGND VGND VPWR VPWR _4054_/S sky130_fd_sc_hd__and2_4
XFILLER_44_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold8 hold8/A VGND VGND VPWR VPWR hold8/X sky130_fd_sc_hd__bufbuf_16
XFILLER_87_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire350 _3794_/X VGND VGND VPWR VPWR wire350/X sky130_fd_sc_hd__buf_6
Xhold408 _4208_/X VGND VGND VPWR VPWR _6671_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_171_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire383 hold90/X VGND VGND VPWR VPWR hold91/A sky130_fd_sc_hd__buf_8
Xwire361 _5503_/S VGND VGND VPWR VPWR _5501_/S sky130_fd_sc_hd__buf_8
XFILLER_128_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3420_ _4241_/A _3539_/B VGND VGND VPWR VPWR _5245_/A sky130_fd_sc_hd__nor2_8
XFILLER_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold419 _4278_/X VGND VGND VPWR VPWR _6731_/D sky130_fd_sc_hd__bufbuf_16
X_3351_ _7004_/Q wire450/X hold65/A _7156_/Q _3348_/X VGND VGND VPWR VPWR _3351_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6070_ _6982_/Q _6028_/X _6342_/B1 _6990_/Q _6069_/X VGND VGND VPWR VPWR _6071_/D
+ sky130_fd_sc_hd__a221o_1
X_3282_ _3367_/A _3383_/C VGND VGND VPWR VPWR _3534_/A sky130_fd_sc_hd__or2_4
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5021_ _6780_/Q _4239_/X _4979_/X _5020_/X VGND VGND VPWR VPWR _6780_/D sky130_fd_sc_hd__o22a_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6972_ _6980_/CLK _6972_/D fanout889/X VGND VGND VPWR VPWR _6972_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5923_ _6591_/Q _5977_/A2 _5923_/B1 _6641_/Q VGND VGND VPWR VPWR _5923_/X sky130_fd_sc_hd__a22o_1
XFILLER_53_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5854_ _6964_/Q _5673_/X _5676_/X wire525/X _5853_/X VGND VGND VPWR VPWR _5861_/A
+ sky130_fd_sc_hd__a221o_4
XFILLER_167_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4805_ _4805_/A _4805_/B _4805_/C _4638_/X VGND VGND VPWR VPWR _4806_/D sky130_fd_sc_hd__or4b_1
XFILLER_22_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5785_ _6856_/Q _5698_/Y _5777_/X _5784_/X _3197_/Y VGND VGND VPWR VPWR _5785_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_9_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4736_ _4748_/A _4736_/B VGND VGND VPWR VPWR _5147_/C sky130_fd_sc_hd__nor2_4
XFILLER_119_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4667_ _5050_/A _4714_/B VGND VGND VPWR VPWR _5147_/B sky130_fd_sc_hd__or2_4
XFILLER_174_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3618_ _6606_/Q _4130_/A _4082_/A _6565_/Q VGND VGND VPWR VPWR _3618_/X sky130_fd_sc_hd__a22o_1
X_6406_ _6406_/A _6406_/B VGND VGND VPWR VPWR _6411_/S sky130_fd_sc_hd__nand2_4
X_4598_ _4997_/A _4749_/C VGND VGND VPWR VPWR _4846_/B sky130_fd_sc_hd__nor2_4
XFILLER_122_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6337_ _6762_/Q _6337_/A2 _6337_/B1 _6648_/Q _6336_/X VGND VGND VPWR VPWR _6343_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3549_ _4108_/A1 _6793_/Q _3857_/C VGND VGND VPWR VPWR _3549_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6268_ _6625_/Q _6028_/X _6342_/B1 _6724_/Q _6267_/X VGND VGND VPWR VPWR _6269_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6199_ _6907_/Q _6021_/A wire646/X wire532/X _6198_/X VGND VGND VPWR VPWR _6206_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5219_ wire559/X _5532_/A0 _5222_/S VGND VGND VPWR VPWR _6820_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5570_ hold13/X _7127_/Q hold91/A VGND VGND VPWR VPWR hold14/A sky130_fd_sc_hd__mux2_1
XFILLER_157_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4521_ _4871_/A _4617_/A VGND VGND VPWR VPWR _4798_/A sky130_fd_sc_hd__nor2_2
XFILLER_129_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold205 _6963_/Q VGND VGND VPWR VPWR hold205/X sky130_fd_sc_hd__bufbuf_16
XFILLER_172_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold216 _7062_/Q VGND VGND VPWR VPWR hold216/X sky130_fd_sc_hd__bufbuf_16
X_4452_ _4694_/A VGND VGND VPWR VPWR _4452_/Y sky130_fd_sc_hd__inv_2
Xhold227 _6961_/Q VGND VGND VPWR VPWR hold227/X sky130_fd_sc_hd__bufbuf_16
Xhold249 _6926_/Q VGND VGND VPWR VPWR hold249/X sky130_fd_sc_hd__bufbuf_16
XFILLER_144_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3403_ wire473/X hold89/A _3425_/B1 _6875_/Q VGND VGND VPWR VPWR _3403_/X sky130_fd_sc_hd__a22o_1
Xhold238 _3260_/A VGND VGND VPWR VPWR _3309_/A sky130_fd_sc_hd__bufbuf_16
XFILLER_171_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4383_ _5031_/A _4584_/A VGND VGND VPWR VPWR _4500_/A sky130_fd_sc_hd__nor2_8
XFILLER_131_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7171_ _3949_/A1 _7171_/D fanout871/X VGND VGND VPWR VPWR _7171_/Q sky130_fd_sc_hd__dfrtp_2
X_6122_ _7112_/Q wire650/X _6021_/B _7152_/Q VGND VGND VPWR VPWR _6122_/X sky130_fd_sc_hd__a22o_1
XFILLER_124_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3334_ _3505_/A _3355_/B VGND VGND VPWR VPWR _3334_/Y sky130_fd_sc_hd__nor2_4
XFILLER_105_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6053_ _6949_/Q wire636/X _6009_/X _7069_/Q VGND VGND VPWR VPWR _6053_/X sky130_fd_sc_hd__a22o_1
XFILLER_100_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__1132_ _3548_/X VGND VGND VPWR VPWR clkbuf_0__1132_/X sky130_fd_sc_hd__clkbuf_8
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3265_ _3953_/A hold174/X hold110/X VGND VGND VPWR VPWR _3265_/X sky130_fd_sc_hd__a21o_4
X_5004_ _5004_/A _5004_/B VGND VGND VPWR VPWR _5037_/B sky130_fd_sc_hd__and2_2
XFILLER_85_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3196_ _6666_/Q VGND VGND VPWR VPWR _3196_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6955_ _6971_/CLK _6955_/D fanout879/X VGND VGND VPWR VPWR _6955_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_121_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5906_ _6546_/Q wire706/X wire686/X _6769_/Q VGND VGND VPWR VPWR _5906_/X sky130_fd_sc_hd__a22o_1
XFILLER_167_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6886_ _7111_/CLK _6886_/D fanout880/X VGND VGND VPWR VPWR _6886_/Q sky130_fd_sc_hd__dfstp_4
X_5837_ _7003_/Q _5667_/X _5681_/X _6923_/Q VGND VGND VPWR VPWR _5837_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5768_ _3211_/A _5685_/X _5699_/X _6928_/Q VGND VGND VPWR VPWR _5768_/X sky130_fd_sc_hd__a22o_1
XFILLER_10_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4719_ _4690_/A _4719_/B _4719_/C VGND VGND VPWR VPWR _4719_/X sky130_fd_sc_hd__and3b_4
XFILLER_154_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5699_ _5864_/B _5706_/B _5707_/B VGND VGND VPWR VPWR _5699_/X sky130_fd_sc_hd__and3_4
XFILLER_162_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold772 _6604_/Q VGND VGND VPWR VPWR hold772/X sky130_fd_sc_hd__bufbuf_16
Xhold761 _4265_/X VGND VGND VPWR VPWR _6720_/D sky130_fd_sc_hd__bufbuf_16
Xhold750 _6672_/Q VGND VGND VPWR VPWR hold750/X sky130_fd_sc_hd__bufbuf_16
XFILLER_122_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold794 _6576_/Q VGND VGND VPWR VPWR hold794/X sky130_fd_sc_hd__bufbuf_16
Xhold783 _6987_/Q VGND VGND VPWR VPWR hold783/X sky130_fd_sc_hd__bufbuf_16
XFILLER_39_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6740_ _6810_/CLK _6740_/D fanout853/X VGND VGND VPWR VPWR _6740_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_189_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3952_ _7174_/Q _6827_/Q _6831_/Q VGND VGND VPWR VPWR _3952_/X sky130_fd_sc_hd__mux2_2
X_6671_ _7122_/CLK _6671_/D fanout887/X VGND VGND VPWR VPWR _6671_/Q sky130_fd_sc_hd__dfrtp_2
X_3883_ _6472_/Q _6456_/Q _6425_/B VGND VGND VPWR VPWR _3883_/X sky130_fd_sc_hd__o21a_2
XFILLER_149_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5622_ _6679_/Q _5620_/Y _7161_/Q VGND VGND VPWR VPWR _7161_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5553_ hold642/X _5598_/A0 _5557_/S VGND VGND VPWR VPWR _7112_/D sky130_fd_sc_hd__mux2_1
XFILLER_136_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4504_ _4812_/A _5164_/B VGND VGND VPWR VPWR _5087_/B sky130_fd_sc_hd__nor2_1
XFILLER_117_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5484_ hold813/X _5547_/A0 _5485_/S VGND VGND VPWR VPWR _7051_/D sky130_fd_sc_hd__mux2_1
X_4435_ _4696_/A _4446_/B VGND VGND VPWR VPWR _4440_/B sky130_fd_sc_hd__nand2_8
XFILLER_172_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7223_ _7223_/CLK _7223_/D fanout850/X VGND VGND VPWR VPWR _7223_/Q sky130_fd_sc_hd__dfstp_1
X_7154_ _7154_/CLK _7154_/D fanout886/X VGND VGND VPWR VPWR _7154_/Q sky130_fd_sc_hd__dfrtp_2
X_4366_ _4364_/A _4364_/B _4388_/B VGND VGND VPWR VPWR _4553_/B sky130_fd_sc_hd__o21bai_4
XFILLER_160_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6105_ _6863_/Q _6025_/D wire618/X wire507/X _6104_/X VGND VGND VPWR VPWR _6106_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_113_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3317_ _3508_/A hold87/X VGND VGND VPWR VPWR _5495_/A sky130_fd_sc_hd__nor2_8
X_4297_ _5599_/A0 hold296/X _4297_/S VGND VGND VPWR VPWR _4297_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7085_ _7105_/CLK _7085_/D fanout862/X VGND VGND VPWR VPWR _7085_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_100_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6036_ _6036_/A _6036_/B VGND VGND VPWR VPWR _6036_/Y sky130_fd_sc_hd__nor2_8
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3248_ _6487_/Q _6486_/Q _6485_/Q VGND VGND VPWR VPWR _3857_/C sky130_fd_sc_hd__or3_4
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6938_ _7147_/CLK _6938_/D fanout888/X VGND VGND VPWR VPWR _6938_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6869_ _7153_/CLK _6869_/D fanout881/X VGND VGND VPWR VPWR _6869_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_167_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire905 wire905/A VGND VGND VPWR VPWR wire905/X sky130_fd_sc_hd__buf_6
XFILLER_22_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length514 _7024_/Q VGND VGND VPWR VPWR wire513/A sky130_fd_sc_hd__buf_6
XFILLER_41_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold580 _6917_/Q VGND VGND VPWR VPWR hold580/X sky130_fd_sc_hd__bufbuf_16
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold591 _5422_/X VGND VGND VPWR VPWR _6996_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_131_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4220_ hold543/X _6407_/A0 _4232_/S VGND VGND VPWR VPWR _4220_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4151_ hold700/X _5408_/A1 _4153_/S VGND VGND VPWR VPWR _6621_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4082_ _4082_/A _4154_/B VGND VGND VPWR VPWR _4087_/S sky130_fd_sc_hd__and2_4
XFILLER_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4984_ _4871_/A _4749_/C _4812_/A VGND VGND VPWR VPWR _5004_/B sky130_fd_sc_hd__a21oi_4
XFILLER_51_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6723_ _6833_/CLK _6723_/D fanout873/X VGND VGND VPWR VPWR _6723_/Q sky130_fd_sc_hd__dfrtp_2
X_3935_ _6840_/Q input78/X _3970_/B VGND VGND VPWR VPWR _3935_/X sky130_fd_sc_hd__mux2_4
XFILLER_32_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6654_ _6787_/CLK _6654_/D fanout853/X VGND VGND VPWR VPWR _6654_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_32_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5605_ _5615_/D VGND VGND VPWR VPWR _5605_/Y sky130_fd_sc_hd__inv_2
X_3866_ _6664_/Q _3866_/B VGND VGND VPWR VPWR _3866_/X sky130_fd_sc_hd__and2b_1
XFILLER_176_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3797_ _6667_/Q _6666_/Q VGND VGND VPWR VPWR _3797_/X sky130_fd_sc_hd__or2_4
X_6585_ _7220_/CLK _6585_/D VGND VGND VPWR VPWR _6585_/Q sky130_fd_sc_hd__dfxtp_2
X_5536_ hold150/X hold179/X _5536_/S VGND VGND VPWR VPWR _5536_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5467_ wire739/A hold573/X _5467_/S VGND VGND VPWR VPWR _7036_/D sky130_fd_sc_hd__mux2_1
X_4418_ _5050_/A _4711_/A VGND VGND VPWR VPWR _4773_/A sky130_fd_sc_hd__xor2_4
XFILLER_133_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7206_ _7208_/CLK _7206_/D VGND VGND VPWR VPWR _7206_/Q sky130_fd_sc_hd__dfxtp_4
X_5398_ _6974_/Q wire794/A _5404_/S VGND VGND VPWR VPWR _6974_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4349_ _4349_/A _4349_/B _4349_/C _4349_/D VGND VGND VPWR VPWR _4352_/A sky130_fd_sc_hd__and4_1
XFILLER_143_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7137_ _7137_/CLK _7137_/D fanout871/X VGND VGND VPWR VPWR _7137_/Q sky130_fd_sc_hd__dfrtp_2
X_7068_ _7068_/CLK _7068_/D fanout879/X VGND VGND VPWR VPWR _7068_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_101_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout378 _5665_/Y VGND VGND VPWR VPWR _6110_/S sky130_fd_sc_hd__buf_8
XFILLER_74_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6019_ _6019_/A _6036_/B VGND VGND VPWR VPWR _6021_/D sky130_fd_sc_hd__nor2_8
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire702 _5676_/X VGND VGND VPWR VPWR wire702/X sky130_fd_sc_hd__buf_8
XFILLER_155_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire757 wire758/X VGND VGND VPWR VPWR wire757/X sky130_fd_sc_hd__buf_6
Xwire746 wire746/A VGND VGND VPWR VPWR wire746/X sky130_fd_sc_hd__buf_8
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout890 fanout891/X VGND VGND VPWR VPWR fanout890/X sky130_fd_sc_hd__buf_8
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_261 _3202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_250 _5532_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_283 hold575/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_272 hold465/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_294 _3606_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3720_ _6990_/Q _5414_/A _3368_/Y input12/X _3679_/X VGND VGND VPWR VPWR _3725_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_13_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3651_ _6532_/Q _4043_/A _4166_/A _6636_/Q _3650_/X VGND VGND VPWR VPWR _3654_/C
+ sky130_fd_sc_hd__a221o_4
XFILLER_146_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3582_ _6920_/Q _3582_/A2 _3582_/B1 _3235_/A _3581_/X VGND VGND VPWR VPWR _3587_/B
+ sky130_fd_sc_hd__a221o_1
X_6370_ _7210_/Q wire353/X _6370_/S VGND VGND VPWR VPWR _7210_/D sky130_fd_sc_hd__mux2_1
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5321_ _5600_/A0 hold452/X _5323_/S VGND VGND VPWR VPWR _6906_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5252_ _5252_/A _5252_/B _5252_/C hold71/X VGND VGND VPWR VPWR _5260_/S sky130_fd_sc_hd__or4_4
XFILLER_130_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4203_ _6690_/Q _5595_/A0 _4209_/S VGND VGND VPWR VPWR _4203_/X sky130_fd_sc_hd__mux2_1
X_5183_ _5143_/Y _5146_/Y _5175_/X _5182_/X VGND VGND VPWR VPWR _5184_/B sky130_fd_sc_hd__a31o_1
XFILLER_87_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4134_ hold83/X _6607_/Q _4135_/S VGND VGND VPWR VPWR _4134_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4065_ hold83/X _6548_/Q _4066_/S VGND VGND VPWR VPWR _6548_/D sky130_fd_sc_hd__mux2_1
XFILLER_36_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4967_ _4956_/C _4719_/X _4959_/X _4571_/Y _4628_/Y VGND VGND VPWR VPWR _5073_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_51_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4898_ _4965_/A _4898_/B VGND VGND VPWR VPWR _4911_/B sky130_fd_sc_hd__nor2_1
X_6706_ _7208_/CLK _6706_/D _6362_/B VGND VGND VPWR VPWR _6706_/Q sky130_fd_sc_hd__dfrtp_2
X_3918_ _5659_/C _3918_/B VGND VGND VPWR VPWR _3918_/X sky130_fd_sc_hd__or2_1
XFILLER_192_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6637_ _6752_/CLK _6637_/D fanout857/X VGND VGND VPWR VPWR _6637_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3849_ _3196_/Y _6668_/Q _3859_/B _6473_/Q VGND VGND VPWR VPWR _6473_/D sky130_fd_sc_hd__a31o_1
X_6568_ _7210_/CLK _6568_/D VGND VGND VPWR VPWR _6568_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_22_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5519_ _5519_/A0 hold836/X _5521_/S VGND VGND VPWR VPWR _5519_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6499_ _6810_/CLK _6499_/D fanout853/X VGND VGND VPWR VPWR _6499_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_160_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire532 _6939_/Q VGND VGND VPWR VPWR wire532/X sky130_fd_sc_hd__buf_6
Xwire521 _7003_/Q VGND VGND VPWR VPWR wire521/X sky130_fd_sc_hd__buf_6
XFILLER_7_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire510 _7032_/Q VGND VGND VPWR VPWR _3218_/A sky130_fd_sc_hd__buf_8
XFILLER_183_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire565 _6746_/Q VGND VGND VPWR VPWR wire565/X sky130_fd_sc_hd__buf_6
Xwire554 _6864_/Q VGND VGND VPWR VPWR _3238_/A sky130_fd_sc_hd__buf_6
Xwire543 _6896_/Q VGND VGND VPWR VPWR _3235_/A sky130_fd_sc_hd__buf_6
XFILLER_143_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire598 _6023_/A VGND VGND VPWR VPWR wire598/X sky130_fd_sc_hd__buf_8
Xwire587 _6014_/Y VGND VGND VPWR VPWR _6025_/D sky130_fd_sc_hd__buf_8
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5870_ _6972_/Q _5691_/X _5699_/X _6932_/Q _5869_/X VGND VGND VPWR VPWR _5871_/D
+ sky130_fd_sc_hd__a221o_4
XFILLER_92_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4821_ _5119_/A _5135_/A VGND VGND VPWR VPWR _5013_/B sky130_fd_sc_hd__or2_4
XFILLER_73_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4752_ _4592_/B _5147_/C _4756_/B VGND VGND VPWR VPWR _4753_/D sky130_fd_sc_hd__a21o_1
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3703_ _6926_/Q _5342_/A _5396_/A _6974_/Q _3702_/X VGND VGND VPWR VPWR _3709_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4683_ _4745_/A _4832_/B VGND VGND VPWR VPWR _5151_/A sky130_fd_sc_hd__nor2_1
X_3634_ _6863_/Q wire439/X _5306_/A _6895_/Q _3633_/X VGND VGND VPWR VPWR _3635_/D
+ sky130_fd_sc_hd__a221o_1
X_6422_ _6455_/A _6455_/B VGND VGND VPWR VPWR _6422_/X sky130_fd_sc_hd__and2_1
XFILLER_146_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6353_ _6663_/Q wire647/X wire632/X _6593_/Q VGND VGND VPWR VPWR _6353_/X sky130_fd_sc_hd__a22o_1
X_3565_ _7016_/Q _5441_/A _4274_/A _6731_/Q VGND VGND VPWR VPWR _3565_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5304_ _5601_/A0 hold229/X _5305_/S VGND VGND VPWR VPWR _6891_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3496_ input24/X _3302_/Y _5360_/A _6945_/Q _3495_/X VGND VGND VPWR VPWR _3504_/B
+ sky130_fd_sc_hd__a221o_4
X_6284_ wire824/X _7197_/Q wire381/X _6283_/X VGND VGND VPWR VPWR _6284_/X sky130_fd_sc_hd__a211o_2
XFILLER_130_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5235_ hold607/X _5227_/A _5576_/B _5234_/X VGND VGND VPWR VPWR _5235_/X sky130_fd_sc_hd__o211a_1
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5166_ _5166_/A _5166_/B _5166_/C _4935_/C VGND VGND VPWR VPWR _5166_/X sky130_fd_sc_hd__or4b_4
XFILLER_69_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5097_ _5164_/A _4995_/A _5096_/X VGND VGND VPWR VPWR _5098_/C sky130_fd_sc_hd__o21ai_1
X_4117_ _4303_/A0 hold404/X _4117_/S VGND VGND VPWR VPWR _6593_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4048_ _6534_/Q _6411_/A0 _4048_/S VGND VGND VPWR VPWR _6534_/D sky130_fd_sc_hd__mux2_1
XFILLER_140_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5999_ _6019_/A _6004_/A VGND VGND VPWR VPWR _6023_/A sky130_fd_sc_hd__nor2_8
XFILLER_184_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput290 _6818_/Q VGND VGND VPWR VPWR pll_trim[23] sky130_fd_sc_hd__buf_8
Xhold9 hold9/A VGND VGND VPWR VPWR hold9/X sky130_fd_sc_hd__bufbuf_16
XFILLER_181_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire351 _3452_/X VGND VGND VPWR VPWR wire351/X sky130_fd_sc_hd__buf_6
Xhold409 _6673_/Q VGND VGND VPWR VPWR hold409/X sky130_fd_sc_hd__bufbuf_16
Xwire373 _6027_/X VGND VGND VPWR VPWR _6060_/B sky130_fd_sc_hd__buf_8
Xclkbuf_leaf_62_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7140_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_7_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire362 _5502_/S VGND VGND VPWR VPWR _5503_/S sky130_fd_sc_hd__buf_6
XFILLER_152_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3350_ hold63/X _5252_/A VGND VGND VPWR VPWR hold64/A sky130_fd_sc_hd__nor2_4
XFILLER_152_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_77_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6787_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5020_ _5102_/C _4946_/X _5002_/X _5019_/X VGND VGND VPWR VPWR _5020_/X sky130_fd_sc_hd__a211o_1
X_3281_ _3281_/A _3281_/B VGND VGND VPWR VPWR _3383_/C sky130_fd_sc_hd__nand2_2
XFILLER_3_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6971_ _6971_/CLK _6971_/D fanout879/X VGND VGND VPWR VPWR _6971_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_93_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5922_ _6715_/Q wire702/X _5682_/X wire563/X _5921_/X VGND VGND VPWR VPWR _5927_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_15_csclk _6708_/CLK VGND VGND VPWR VPWR _6720_/CLK sky130_fd_sc_hd__clkbuf_8
X_5853_ _6924_/Q _5681_/X wire651/A _7028_/Q VGND VGND VPWR VPWR _5853_/X sky130_fd_sc_hd__a22o_1
XFILLER_110_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4804_ _4654_/A _4958_/A _4702_/A _4711_/C _4803_/X VGND VGND VPWR VPWR _4805_/C
+ sky130_fd_sc_hd__a41o_4
X_5784_ _5784_/A _5784_/B _5784_/C VGND VGND VPWR VPWR _5784_/X sky130_fd_sc_hd__or3_4
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4735_ _4735_/A _4735_/B _4566_/A VGND VGND VPWR VPWR _4735_/X sky130_fd_sc_hd__or3b_4
XFILLER_159_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4666_ _5050_/A _4714_/B VGND VGND VPWR VPWR _4668_/B sky130_fd_sc_hd__nor2_8
XFILLER_119_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3617_ _6887_/Q _5297_/A wire406/X _6879_/Q VGND VGND VPWR VPWR _3617_/X sky130_fd_sc_hd__a22o_1
X_4597_ _4648_/B _4947_/B VGND VGND VPWR VPWR _4957_/A sky130_fd_sc_hd__nor2_8
X_6405_ hold68/A _6704_/Q _4239_/X wire573/X VGND VGND VPWR VPWR _7220_/D sky130_fd_sc_hd__o31a_1
XFILLER_134_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3548_ _3548_/A _3548_/B _3548_/C VGND VGND VPWR VPWR _3548_/X sky130_fd_sc_hd__or3_2
X_6336_ _6737_/Q wire643/X wire630/X _6789_/Q VGND VGND VPWR VPWR _6336_/X sky130_fd_sc_hd__a22o_1
XFILLER_103_524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3479_ wire548/X _3374_/Y _4148_/A _6623_/Q _3477_/X VGND VGND VPWR VPWR _3488_/B
+ sky130_fd_sc_hd__a221o_1
X_6267_ _7222_/Q _6009_/X wire627/X _6709_/Q VGND VGND VPWR VPWR _6267_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6198_ _6955_/Q wire637/X wire635/X _6931_/Q VGND VGND VPWR VPWR _6198_/X sky130_fd_sc_hd__a22o_1
XFILLER_69_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5218_ _5218_/A _5576_/B VGND VGND VPWR VPWR _5222_/S sky130_fd_sc_hd__and2_4
XFILLER_28_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5149_ _5146_/A _5146_/B _5175_/C _5143_/Y VGND VGND VPWR VPWR _5169_/B sky130_fd_sc_hd__o31a_2
XFILLER_151_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4520_ _4370_/Y _4503_/Y _4506_/X _4484_/B _4533_/A VGND VGND VPWR VPWR _4520_/X
+ sky130_fd_sc_hd__a2111o_1
Xhold217 _6516_/Q VGND VGND VPWR VPWR hold217/X sky130_fd_sc_hd__bufbuf_16
X_4451_ _4525_/A _4590_/A VGND VGND VPWR VPWR _4694_/A sky130_fd_sc_hd__or2_4
Xhold206 _6899_/Q VGND VGND VPWR VPWR hold206/X sky130_fd_sc_hd__bufbuf_16
XFILLER_171_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold228 _7059_/Q VGND VGND VPWR VPWR hold228/X sky130_fd_sc_hd__bufbuf_16
Xhold239 _5295_/X VGND VGND VPWR VPWR _6883_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_132_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3402_ _6883_/Q _5288_/A _5360_/A _6947_/Q _3401_/X VGND VGND VPWR VPWR _3415_/B
+ sky130_fd_sc_hd__a221o_1
X_7170_ _3949_/A1 _7170_/D fanout871/X VGND VGND VPWR VPWR _7170_/Q sky130_fd_sc_hd__dfstp_4
X_4382_ _4469_/A _4819_/A VGND VGND VPWR VPWR _4584_/A sky130_fd_sc_hd__nand2_8
XFILLER_124_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6121_ _6121_/A _6121_/B _6121_/C _6121_/D VGND VGND VPWR VPWR _6121_/X sky130_fd_sc_hd__or4_2
XFILLER_98_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ _5225_/A _3510_/B VGND VGND VPWR VPWR _5207_/A sky130_fd_sc_hd__nor2_8
X_6052_ _6901_/Q wire600/X _6295_/B1 _7149_/Q _6051_/X VGND VGND VPWR VPWR _6057_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_140_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3264_ _3953_/A _3264_/B VGND VGND VPWR VPWR _3264_/X sky130_fd_sc_hd__and2b_4
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _5003_/A _5003_/B _5003_/C VGND VGND VPWR VPWR _5003_/X sky130_fd_sc_hd__and3_1
XFILLER_66_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3195_ _6704_/Q VGND VGND VPWR VPWR _3916_/A sky130_fd_sc_hd__clkinv_8
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6954_ _6979_/CLK _6954_/D fanout885/X VGND VGND VPWR VPWR _6954_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_121_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5905_ _6620_/Q wire707/X _5681_/X _6595_/Q _5904_/X VGND VGND VPWR VPWR _5910_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_81_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6885_ _7153_/CLK _6885_/D fanout881/X VGND VGND VPWR VPWR _6885_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_167_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5836_ _6971_/Q _5691_/X _5835_/X VGND VGND VPWR VPWR _5839_/C sky130_fd_sc_hd__a21o_1
X_5767_ _3235_/A wire674/X _5812_/B1 _7056_/Q VGND VGND VPWR VPWR _5767_/X sky130_fd_sc_hd__a22o_1
X_4718_ _4745_/A _4757_/B VGND VGND VPWR VPWR _5178_/A sky130_fd_sc_hd__nor2_2
XFILLER_108_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5698_ _5864_/B _5698_/B VGND VGND VPWR VPWR _5698_/Y sky130_fd_sc_hd__nand2_8
XFILLER_190_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4649_ _4722_/B _4650_/B VGND VGND VPWR VPWR _4719_/C sky130_fd_sc_hd__nor2_4
XFILLER_135_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold751 _4210_/X VGND VGND VPWR VPWR _6672_/D sky130_fd_sc_hd__bufbuf_16
Xhold773 _6550_/Q VGND VGND VPWR VPWR hold773/X sky130_fd_sc_hd__bufbuf_16
Xhold762 _7035_/Q VGND VGND VPWR VPWR hold762/X sky130_fd_sc_hd__bufbuf_16
Xhold740 _7019_/Q VGND VGND VPWR VPWR hold740/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold795 _6545_/Q VGND VGND VPWR VPWR hold795/X sky130_fd_sc_hd__bufbuf_16
XFILLER_103_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6319_ _7224_/Q _6009_/X wire627/X _6711_/Q VGND VGND VPWR VPWR _6319_/X sky130_fd_sc_hd__a22o_1
Xhold784 _6785_/Q VGND VGND VPWR VPWR hold784/X sky130_fd_sc_hd__bufbuf_16
XFILLER_162_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3951_ _7172_/Q _6828_/Q _6831_/Q VGND VGND VPWR VPWR _3951_/X sky130_fd_sc_hd__mux2_2
XFILLER_51_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6670_ _6930_/CLK _6670_/D fanout887/X VGND VGND VPWR VPWR _6670_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3882_ _7173_/Q _6826_/Q _6831_/Q VGND VGND VPWR VPWR _3920_/B sky130_fd_sc_hd__mux2_8
XFILLER_188_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5621_ _6677_/Q _6679_/Q VGND VGND VPWR VPWR _5621_/X sky130_fd_sc_hd__or2_2
X_5552_ hold289/X _5597_/A0 _5557_/S VGND VGND VPWR VPWR _7111_/D sky130_fd_sc_hd__mux2_1
XFILLER_157_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4503_ _5087_/A VGND VGND VPWR VPWR _4503_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5483_ hold814/X wire753/X _5485_/S VGND VGND VPWR VPWR _7050_/D sky130_fd_sc_hd__mux2_1
X_4434_ _4735_/A _4672_/A _4469_/A _4395_/D VGND VGND VPWR VPWR _4446_/B sky130_fd_sc_hd__o211a_4
XFILLER_6_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7222_ _7225_/CLK _7222_/D fanout850/X VGND VGND VPWR VPWR _7222_/Q sky130_fd_sc_hd__dfrtp_2
X_7153_ _7153_/CLK _7153_/D fanout881/X VGND VGND VPWR VPWR _7153_/Q sky130_fd_sc_hd__dfrtp_2
X_4365_ _4707_/B _4364_/B _4340_/B VGND VGND VPWR VPWR _4388_/B sky130_fd_sc_hd__o21a_1
XFILLER_98_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6104_ wire482/X wire711/X _6301_/B1 wire530/X VGND VGND VPWR VPWR _6104_/X sky130_fd_sc_hd__a22o_1
XFILLER_113_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3316_ _3421_/A hold86/X hold95/X VGND VGND VPWR VPWR hold87/A sky130_fd_sc_hd__or3_4
X_7084_ _7132_/CLK _7084_/D fanout868/X VGND VGND VPWR VPWR _7084_/Q sky130_fd_sc_hd__dfrtp_2
X_4296_ hold83/X hold208/X _4297_/S VGND VGND VPWR VPWR _4296_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6035_ _6035_/A _6037_/C _6035_/C VGND VGND VPWR VPWR _6111_/B sky130_fd_sc_hd__and3_4
XFILLER_58_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3247_ _4707_/B VGND VGND VPWR VPWR _4655_/A sky130_fd_sc_hd__inv_6
XFILLER_100_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6937_ _7133_/CLK _6937_/D fanout883/X VGND VGND VPWR VPWR _6937_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6868_ _7152_/CLK _6868_/D fanout886/X VGND VGND VPWR VPWR _6868_/Q sky130_fd_sc_hd__dfrtp_2
Xwire917 _4735_/A VGND VGND VPWR VPWR _4818_/A sky130_fd_sc_hd__buf_8
XFILLER_179_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire906 wire906/A VGND VGND VPWR VPWR wire906/X sky130_fd_sc_hd__buf_6
X_5819_ _7042_/Q wire694/X wire660/X wire533/X _5810_/X VGND VGND VPWR VPWR _5826_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_10_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6799_ _6806_/CLK _6799_/D _6435_/A VGND VGND VPWR VPWR _6799_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold581 _6981_/Q VGND VGND VPWR VPWR hold581/X sky130_fd_sc_hd__bufbuf_16
Xhold570 _6551_/Q VGND VGND VPWR VPWR hold570/X sky130_fd_sc_hd__bufbuf_16
XFILLER_2_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold592 _6839_/Q VGND VGND VPWR VPWR hold592/X sky130_fd_sc_hd__bufbuf_16
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4150_ hold683/X wire794/X _4153_/S VGND VGND VPWR VPWR _6620_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4081_ _6562_/Q wire353/X _4081_/S VGND VGND VPWR VPWR _6562_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4983_ _5013_/A _4983_/B VGND VGND VPWR VPWR _5135_/B sky130_fd_sc_hd__or2_2
XFILLER_189_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3934_ _6839_/Q input80/X _3970_/B VGND VGND VPWR VPWR _3934_/X sky130_fd_sc_hd__mux2_2
X_6722_ _7223_/CLK _6722_/D fanout851/X VGND VGND VPWR VPWR _6722_/Q sky130_fd_sc_hd__dfstp_4
X_6653_ _6752_/CLK _6653_/D fanout857/X VGND VGND VPWR VPWR _6653_/Q sky130_fd_sc_hd__dfrtp_2
X_3865_ _3866_/B _3865_/B VGND VGND VPWR VPWR _6468_/D sky130_fd_sc_hd__xnor2_1
X_5604_ _5611_/A _6680_/Q _6679_/Q _3920_/Y VGND VGND VPWR VPWR _5615_/D sky130_fd_sc_hd__o31a_4
XFILLER_191_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6584_ _7208_/CLK _6584_/D VGND VGND VPWR VPWR _6584_/Q sky130_fd_sc_hd__dfxtp_2
X_3796_ _6790_/Q _3928_/A wire350/X _3795_/Y VGND VGND VPWR VPWR _6790_/D sky130_fd_sc_hd__a22o_1
XFILLER_157_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5535_ _5598_/A0 hold624/X _5536_/S VGND VGND VPWR VPWR _7096_/D sky130_fd_sc_hd__mux2_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5466_ _5547_/A0 hold762/X _5467_/S VGND VGND VPWR VPWR _7035_/D sky130_fd_sc_hd__mux2_1
X_4417_ _4650_/B _4416_/B _4415_/X VGND VGND VPWR VPWR _5165_/A sky130_fd_sc_hd__a21oi_4
XFILLER_160_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7205_ _7208_/CLK _7205_/D VGND VGND VPWR VPWR _7205_/Q sky130_fd_sc_hd__dfxtp_4
X_5397_ _6973_/Q hold465/X _5404_/S VGND VGND VPWR VPWR _6973_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4348_ _4368_/A _4722_/B VGND VGND VPWR VPWR _4774_/A sky130_fd_sc_hd__or2_4
X_7136_ _7136_/CLK _7136_/D fanout871/X VGND VGND VPWR VPWR _7136_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_59_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7067_ _7140_/CLK _7067_/D fanout865/X VGND VGND VPWR VPWR _7067_/Q sky130_fd_sc_hd__dfrtp_2
X_4279_ _6411_/A0 hold639/X _4279_/S VGND VGND VPWR VPWR _6732_/D sky130_fd_sc_hd__mux2_1
XFILLER_100_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6018_ _6018_/A _6035_/C _6032_/C VGND VGND VPWR VPWR _6022_/D sky130_fd_sc_hd__and3_4
XFILLER_74_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire714 _5062_/A VGND VGND VPWR VPWR _4965_/B sky130_fd_sc_hd__buf_8
Xwire725 _4154_/B VGND VGND VPWR VPWR _5378_/B sky130_fd_sc_hd__buf_8
XFILLER_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire758 hold27/X VGND VGND VPWR VPWR wire758/X sky130_fd_sc_hd__buf_8
Xwire736 _4502_/A VGND VGND VPWR VPWR _4986_/A sky130_fd_sc_hd__buf_8
XFILLER_109_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire769 wire770/X VGND VGND VPWR VPWR wire769/X sky130_fd_sc_hd__buf_8
XFILLER_182_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout880 fanout889/X VGND VGND VPWR VPWR fanout880/X sky130_fd_sc_hd__buf_8
XFILLER_92_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout891 input75/X VGND VGND VPWR VPWR fanout891/X sky130_fd_sc_hd__buf_8
XFILLER_133_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_251 _5963_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_240 _5259_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_262 wire912/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_284 hold575/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_273 hold465/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_295 _3785_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3650_ input13/X _3368_/Y _5238_/A _6834_/Q VGND VGND VPWR VPWR _3650_/X sky130_fd_sc_hd__a22o_4
XFILLER_127_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3581_ _3581_/A1 _5315_/A _4097_/A _6579_/Q VGND VGND VPWR VPWR _3581_/X sky130_fd_sc_hd__a22o_2
X_5320_ _5599_/A0 hold352/X _5323_/S VGND VGND VPWR VPWR _5320_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5251_ hold27/X hold846/X _5251_/S VGND VGND VPWR VPWR hold28/A sky130_fd_sc_hd__mux2_1
XFILLER_142_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4202_ hold45/X _6421_/B _4007_/X hold46/X _5594_/B VGND VGND VPWR VPWR _4218_/S
+ sky130_fd_sc_hd__o221a_4
XFILLER_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5182_ _6784_/Q _5156_/A _5158_/Y _5178_/X _5181_/X VGND VGND VPWR VPWR _5182_/X
+ sky130_fd_sc_hd__a221o_1
X_4133_ _5498_/A0 _6606_/Q _4135_/S VGND VGND VPWR VPWR _6606_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4064_ _5408_/A1 hold685/X _4066_/S VGND VGND VPWR VPWR _6547_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4966_ _4443_/X _4536_/B _4959_/A _4909_/B VGND VGND VPWR VPWR _5145_/B sky130_fd_sc_hd__a31o_2
X_6705_ _7210_/CLK _6705_/D _6362_/B VGND VGND VPWR VPWR _6705_/Q sky130_fd_sc_hd__dfrtp_2
X_4897_ _5003_/A _4897_/B VGND VGND VPWR VPWR _4913_/B sky130_fd_sc_hd__nand2_1
X_3917_ _6457_/Q _3192_/Y _6664_/Q _3843_/B _6665_/Q VGND VGND VPWR VPWR _6665_/D
+ sky130_fd_sc_hd__a41o_1
XFILLER_20_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6636_ _6752_/CLK _6636_/D fanout857/X VGND VGND VPWR VPWR _6636_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_22_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3848_ _6474_/Q _6459_/Q _3848_/S VGND VGND VPWR VPWR _6474_/D sky130_fd_sc_hd__mux2_1
XFILLER_164_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6567_ _6623_/CLK _6567_/D fanout890/X VGND VGND VPWR VPWR _6567_/Q sky130_fd_sc_hd__dfrtp_2
X_3779_ _7175_/Q _3384_/Y _6406_/A _7221_/Q VGND VGND VPWR VPWR _3779_/X sky130_fd_sc_hd__a22o_1
XFILLER_192_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5518_ hold156/X hold852/X _5521_/S VGND VGND VPWR VPWR _5518_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6498_ _6810_/CLK _6498_/D fanout853/X VGND VGND VPWR VPWR _6498_/Q sky130_fd_sc_hd__dfstp_4
X_5449_ wire739/X hold672/X _5449_/S VGND VGND VPWR VPWR _7020_/D sky130_fd_sc_hd__mux2_1
XFILLER_120_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7119_ _7119_/CLK _7119_/D fanout871/X VGND VGND VPWR VPWR _7119_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f_wbbd_sck clkbuf_0_wbbd_sck/X VGND VGND VPWR VPWR _6401_/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_179_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire500 _7057_/Q VGND VGND VPWR VPWR wire500/X sky130_fd_sc_hd__buf_6
XFILLER_8_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire533 _6938_/Q VGND VGND VPWR VPWR wire533/X sky130_fd_sc_hd__buf_6
Xwire522 wire522/A VGND VGND VPWR VPWR wire522/X sky130_fd_sc_hd__buf_6
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire511 _7029_/Q VGND VGND VPWR VPWR wire511/X sky130_fd_sc_hd__buf_6
Xwire555 _6862_/Q VGND VGND VPWR VPWR wire555/X sky130_fd_sc_hd__buf_6
Xwire544 _6888_/Q VGND VGND VPWR VPWR _3236_/A sky130_fd_sc_hd__buf_6
XFILLER_7_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire566 _6740_/Q VGND VGND VPWR VPWR wire566/X sky130_fd_sc_hd__buf_6
XFILLER_171_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire599 _6021_/A VGND VGND VPWR VPWR wire599/X sky130_fd_sc_hd__buf_6
XFILLER_170_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4820_ _5003_/C _4820_/B VGND VGND VPWR VPWR _4827_/A sky130_fd_sc_hd__nand2_1
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751_ _4754_/B _4735_/X _5123_/B _4935_/D _5144_/B VGND VGND VPWR VPWR _4753_/C
+ sky130_fd_sc_hd__o2111a_1
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3702_ _6902_/Q _5315_/A _4061_/A _6546_/Q VGND VGND VPWR VPWR _3702_/X sky130_fd_sc_hd__a22o_1
XFILLER_147_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4682_ _4697_/A _4832_/B VGND VGND VPWR VPWR _4682_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6421_ _6421_/A _6421_/B VGND VGND VPWR VPWR _6421_/X sky130_fd_sc_hd__and2_1
XFILLER_147_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3633_ _7127_/Q hold89/A _3763_/B1 _7135_/Q VGND VGND VPWR VPWR _3633_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6352_ _6539_/Q wire585/X _6352_/B1 _6643_/Q _6351_/X VGND VGND VPWR VPWR _6355_/C
+ sky130_fd_sc_hd__a221o_1
X_3564_ wire522/X _5423_/A _4310_/A _6761_/Q VGND VGND VPWR VPWR _3564_/X sky130_fd_sc_hd__a22o_1
X_5303_ wire758/X _6890_/Q _5305_/S VGND VGND VPWR VPWR _5303_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3495_ _6732_/Q _4274_/A _4196_/A _6663_/Q VGND VGND VPWR VPWR _3495_/X sky130_fd_sc_hd__a22o_4
X_6283_ _6531_/Q _6357_/A2 _6269_/X _6282_/X _6308_/S VGND VGND VPWR VPWR _6283_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_130_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5234_ _5234_/A _5234_/B _5234_/C VGND VGND VPWR VPWR _5234_/X sky130_fd_sc_hd__or3_4
X_5165_ _5165_/A _5165_/B _5165_/C VGND VGND VPWR VPWR _5166_/B sky130_fd_sc_hd__and3_1
XFILLER_69_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4116_ hold83/X hold158/X _4117_/S VGND VGND VPWR VPWR _4116_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5096_ _5164_/B _5017_/A _4756_/B _4724_/B VGND VGND VPWR VPWR _5096_/X sky130_fd_sc_hd__o22a_1
XFILLER_84_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4047_ _6533_/Q _6410_/A0 _4048_/S VGND VGND VPWR VPWR _6533_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5998_ _6019_/A _6037_/B _6033_/C VGND VGND VPWR VPWR _5998_/X sky130_fd_sc_hd__and3b_4
XFILLER_52_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4949_ _4949_/A _4949_/B _4949_/C _4959_/A VGND VGND VPWR VPWR _4950_/C sky130_fd_sc_hd__and4_1
XFILLER_149_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6619_ _6621_/CLK _6619_/D fanout872/X VGND VGND VPWR VPWR _6619_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput280 _6494_/Q VGND VGND VPWR VPWR pll_trim[14] sky130_fd_sc_hd__buf_8
XFILLER_121_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput291 _6504_/Q VGND VGND VPWR VPWR pll_trim[24] sky130_fd_sc_hd__buf_8
XFILLER_87_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire352 _3415_/X VGND VGND VPWR VPWR wire352/X sky130_fd_sc_hd__buf_8
Xwire363 _5365_/S VGND VGND VPWR VPWR _5368_/S sky130_fd_sc_hd__buf_8
Xwire374 _6232_/A VGND VGND VPWR VPWR _6356_/A sky130_fd_sc_hd__buf_6
Xwire385 _5564_/S VGND VGND VPWR VPWR _5566_/S sky130_fd_sc_hd__buf_8
XFILLER_109_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire396 _3372_/Y VGND VGND VPWR VPWR _5405_/A sky130_fd_sc_hd__buf_8
XFILLER_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3280_ _5225_/A VGND VGND VPWR VPWR _3280_/Y sky130_fd_sc_hd__inv_2
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6970_ _6971_/CLK _6970_/D fanout879/X VGND VGND VPWR VPWR _6970_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_93_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5921_ wire568/X _5921_/A2 _5684_/X _6725_/Q VGND VGND VPWR VPWR _5921_/X sky130_fd_sc_hd__a22o_1
XFILLER_93_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5852_ _7182_/Q _6110_/S _5850_/X _5851_/X VGND VGND VPWR VPWR _7182_/D sky130_fd_sc_hd__o22a_1
XFILLER_34_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4803_ _4654_/A _4958_/A _5165_/A _4702_/A _4704_/X VGND VGND VPWR VPWR _4803_/X
+ sky130_fd_sc_hd__a41o_1
X_5783_ _6944_/Q wire656/A _5707_/X _3219_/A _5782_/X VGND VGND VPWR VPWR _5784_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4734_ _4724_/A _4724_/B _4503_/Y VGND VGND VPWR VPWR _4734_/X sky130_fd_sc_hd__o21a_1
XFILLER_119_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4665_ _4665_/A _4696_/B VGND VGND VPWR VPWR _4714_/B sky130_fd_sc_hd__nand2_8
XFILLER_175_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6404_ wire813/X _4238_/B _6374_/X _6403_/X _6372_/A VGND VGND VPWR VPWR _6404_/X
+ sky130_fd_sc_hd__a32o_4
X_3616_ _6959_/Q _5378_/A _5396_/A _6975_/Q VGND VGND VPWR VPWR _3616_/X sky130_fd_sc_hd__a22o_1
X_4596_ _4745_/B _4947_/B VGND VGND VPWR VPWR _5135_/A sky130_fd_sc_hd__nor2_8
XFILLER_127_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3547_ _3547_/A _3547_/B _3547_/C _3547_/D VGND VGND VPWR VPWR _3548_/C sky130_fd_sc_hd__or4_2
X_6335_ _6777_/Q _6335_/B VGND VGND VPWR VPWR _6335_/X sky130_fd_sc_hd__and2_1
XFILLER_130_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3478_ _3534_/A _3540_/A VGND VGND VPWR VPWR _4148_/A sky130_fd_sc_hd__nor2_8
X_6266_ _6754_/Q _6339_/A2 _6339_/B1 _6769_/Q _6265_/X VGND VGND VPWR VPWR _6269_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5217_ wire802/X hold524/X _5217_/S VGND VGND VPWR VPWR _6819_/D sky130_fd_sc_hd__mux2_1
X_6197_ wire473/X wire597/X _6033_/X _7011_/Q _6196_/X VGND VGND VPWR VPWR _6207_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_185_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5148_ _5148_/A _5148_/B _5066_/A _4612_/A VGND VGND VPWR VPWR _5175_/C sky130_fd_sc_hd__or4bb_4
XFILLER_151_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5079_ _5079_/A _5079_/B _5079_/C VGND VGND VPWR VPWR _5137_/A sky130_fd_sc_hd__or3_1
XFILLER_28_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold207 _5313_/X VGND VGND VPWR VPWR _6899_/D sky130_fd_sc_hd__bufbuf_16
X_4450_ _4572_/A _4572_/B VGND VGND VPWR VPWR _4590_/A sky130_fd_sc_hd__or2_1
Xhold218 _6518_/Q VGND VGND VPWR VPWR hold218/X sky130_fd_sc_hd__bufbuf_16
Xhold229 _6891_/Q VGND VGND VPWR VPWR hold229/X sky130_fd_sc_hd__bufbuf_16
X_4381_ _4395_/D _4987_/B VGND VGND VPWR VPWR _5023_/A sky130_fd_sc_hd__nand2_8
X_3401_ wire526/X _3369_/Y _3399_/X _3400_/X VGND VGND VPWR VPWR _3401_/X sky130_fd_sc_hd__a211o_4
X_6120_ _6984_/Q _6028_/X _6293_/B1 _3223_/A _6119_/X VGND VGND VPWR VPWR _6121_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_98_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3332_ _3383_/C _3343_/A VGND VGND VPWR VPWR _3510_/B sky130_fd_sc_hd__or2_4
XFILLER_140_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6051_ _7125_/Q wire598/X _6020_/D _6965_/Q VGND VGND VPWR VPWR _6051_/X sky130_fd_sc_hd__a22o_1
XFILLER_98_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ hold108/X hold40/X _3845_/A VGND VGND VPWR VPWR _3263_/X sky130_fd_sc_hd__mux2_1
X_5002_ _5084_/B _5001_/X _5121_/A VGND VGND VPWR VPWR _5002_/X sky130_fd_sc_hd__o21ba_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3194_ _3194_/A VGND VGND VPWR VPWR _3194_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6953_ _6969_/CLK _6953_/D fanout880/X VGND VGND VPWR VPWR _6953_/Q sky130_fd_sc_hd__dfrtp_2
X_6884_ _7156_/CLK _6884_/D fanout884/X VGND VGND VPWR VPWR _6884_/Q sky130_fd_sc_hd__dfrtp_2
X_5904_ _6709_/Q wire680/X wire664/X _6615_/Q VGND VGND VPWR VPWR _5904_/X sky130_fd_sc_hd__a22o_1
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5835_ wire489/X _5685_/X _5689_/X _6907_/Q VGND VGND VPWR VPWR _5835_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length708 _5921_/A2 VGND VGND VPWR VPWR _5974_/A2 sky130_fd_sc_hd__buf_6
X_5766_ _7178_/Q _6110_/S _5764_/X _5765_/X VGND VGND VPWR VPWR _7178_/D sky130_fd_sc_hd__o22a_1
XFILLER_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4717_ _5164_/B _4717_/B VGND VGND VPWR VPWR _5022_/C sky130_fd_sc_hd__nor2_1
X_5697_ _5864_/B _5702_/B _5703_/B VGND VGND VPWR VPWR _5697_/X sky130_fd_sc_hd__and3_4
XFILLER_108_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4648_ _4671_/A _4648_/B VGND VGND VPWR VPWR _4708_/B sky130_fd_sc_hd__nor2_1
XFILLER_108_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold730 _7141_/Q VGND VGND VPWR VPWR hold730/X sky130_fd_sc_hd__bufbuf_16
XFILLER_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4579_ _4818_/C _4965_/B VGND VGND VPWR VPWR _4874_/B sky130_fd_sc_hd__or2_2
Xhold741 _6768_/Q VGND VGND VPWR VPWR hold741/X sky130_fd_sc_hd__bufbuf_16
Xhold763 _7034_/Q VGND VGND VPWR VPWR hold763/X sky130_fd_sc_hd__bufbuf_16
Xhold752 _6800_/Q VGND VGND VPWR VPWR hold752/X sky130_fd_sc_hd__bufbuf_16
Xhold774 _6599_/Q VGND VGND VPWR VPWR hold774/X sky130_fd_sc_hd__bufbuf_16
Xhold785 _6540_/Q VGND VGND VPWR VPWR hold785/X sky130_fd_sc_hd__bufbuf_16
XFILLER_116_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold796 _6619_/Q VGND VGND VPWR VPWR hold796/X sky130_fd_sc_hd__bufbuf_16
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6318_ _6731_/Q wire603/X _6340_/B1 _6597_/Q _6317_/X VGND VGND VPWR VPWR _6321_/C
+ sky130_fd_sc_hd__a221o_1
X_6249_ _6733_/Q _6020_/B wire634/X _6599_/Q VGND VGND VPWR VPWR _6249_/X sky130_fd_sc_hd__a22o_4
XFILLER_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_61_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7095_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_76_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6642_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_187_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_14_csclk _6708_/CLK VGND VGND VPWR VPWR _6623_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_67_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_29_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _6969_/CLK sky130_fd_sc_hd__clkbuf_8
Xhold90 hold90/A VGND VGND VPWR VPWR hold90/X sky130_fd_sc_hd__bufbuf_16
XFILLER_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3950_ _6511_/Q wire837/X _6836_/Q VGND VGND VPWR VPWR _3950_/X sky130_fd_sc_hd__mux2_8
XFILLER_90_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3881_ _6471_/Q _6456_/Q _6666_/Q _3843_/B VGND VGND VPWR VPWR _6456_/D sky130_fd_sc_hd__o211a_1
XFILLER_188_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5620_ _6677_/Q _6679_/Q VGND VGND VPWR VPWR _5620_/Y sky130_fd_sc_hd__nor2_2
XFILLER_157_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5551_ _7110_/Q hold38/X _5557_/S VGND VGND VPWR VPWR hold98/A sky130_fd_sc_hd__mux2_1
X_4502_ _4502_/A _4812_/A VGND VGND VPWR VPWR _5087_/A sky130_fd_sc_hd__nor2_4
XFILLER_145_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5482_ hold529/X _5572_/A0 _5485_/S VGND VGND VPWR VPWR _7049_/D sky130_fd_sc_hd__mux2_1
X_7221_ _7223_/CLK _7221_/D fanout850/X VGND VGND VPWR VPWR _7221_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_144_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4433_ _4818_/A _4672_/A VGND VGND VPWR VPWR _4663_/B sky130_fd_sc_hd__or2_4
X_7152_ _7152_/CLK _7152_/D fanout886/X VGND VGND VPWR VPWR _7152_/Q sky130_fd_sc_hd__dfrtp_2
X_4364_ _4364_/A _4364_/B VGND VGND VPWR VPWR _4478_/C sky130_fd_sc_hd__or2_4
XFILLER_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4295_ _5498_/A0 _6745_/Q _4297_/S VGND VGND VPWR VPWR _6745_/D sky130_fd_sc_hd__mux2_1
X_6103_ _6871_/Q wire593/X wire591/X _6895_/Q _6102_/X VGND VGND VPWR VPWR _6106_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_140_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3315_ hold96/X _3551_/A VGND VGND VPWR VPWR _5261_/A sky130_fd_sc_hd__nor2_8
X_7083_ _7139_/CLK _7083_/D fanout868/X VGND VGND VPWR VPWR _7083_/Q sky130_fd_sc_hd__dfrtp_2
X_3246_ _4958_/A VGND VGND VPWR VPWR _4654_/B sky130_fd_sc_hd__inv_6
XFILLER_112_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6034_ _6036_/A _6034_/B VGND VGND VPWR VPWR _6034_/Y sky130_fd_sc_hd__nor2_8
XFILLER_132_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6936_ _6980_/CLK _6936_/D fanout880/X VGND VGND VPWR VPWR _6936_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6867_ _7147_/CLK _6867_/D fanout886/X VGND VGND VPWR VPWR _6867_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire907 wire907/A VGND VGND VPWR VPWR wire907/X sky130_fd_sc_hd__buf_6
X_5818_ _6946_/Q wire657/X wire651/X _7026_/Q _5817_/X VGND VGND VPWR VPWR _5827_/C
+ sky130_fd_sc_hd__a221o_1
X_6798_ _6824_/CLK _6798_/D _6435_/A VGND VGND VPWR VPWR _6798_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5749_ _6935_/Q wire659/X wire653/A _7055_/Q VGND VGND VPWR VPWR _5749_/X sky130_fd_sc_hd__a22o_1
XFILLER_6_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold560 _6748_/Q VGND VGND VPWR VPWR hold560/X sky130_fd_sc_hd__bufbuf_16
Xhold571 _6847_/Q VGND VGND VPWR VPWR hold571/X sky130_fd_sc_hd__bufbuf_16
XFILLER_173_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold582 _6988_/Q VGND VGND VPWR VPWR hold582/X sky130_fd_sc_hd__bufbuf_16
Xhold593 _5246_/X VGND VGND VPWR VPWR _6839_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_103_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4080_ _6561_/Q wire352/X _4081_/S VGND VGND VPWR VPWR _6561_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4982_ _4758_/A _4634_/B _4554_/A _4863_/B _4766_/A VGND VGND VPWR VPWR _5084_/B
+ sky130_fd_sc_hd__a311o_4
XFILLER_17_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3933_ _3205_/Y input82/X _3970_/B VGND VGND VPWR VPWR _3933_/X sky130_fd_sc_hd__mux2_4
X_6721_ _6851_/CLK _6721_/D fanout851/X VGND VGND VPWR VPWR _6721_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_176_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6652_ _6842_/CLK _6652_/D fanout857/X VGND VGND VPWR VPWR _6652_/Q sky130_fd_sc_hd__dfrtp_2
X_3864_ _6468_/Q _3864_/B VGND VGND VPWR VPWR _3865_/B sky130_fd_sc_hd__nor2_1
XFILLER_32_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5603_ _5611_/A _6679_/Q VGND VGND VPWR VPWR _5665_/B sky130_fd_sc_hd__nor2_4
XFILLER_118_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3795_ _3857_/C _3928_/A VGND VGND VPWR VPWR _3795_/Y sky130_fd_sc_hd__nor2_1
X_6583_ _7208_/CLK _6583_/D VGND VGND VPWR VPWR _6583_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_117_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5534_ wire786/X hold259/X _5539_/S VGND VGND VPWR VPWR _5534_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5465_ wire753/X hold763/X _5467_/S VGND VGND VPWR VPWR _7034_/D sky130_fd_sc_hd__mux2_1
X_4416_ _4722_/A _4416_/B VGND VGND VPWR VPWR _4774_/C sky130_fd_sc_hd__xor2_4
XFILLER_133_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7204_ _7208_/CLK _7204_/D VGND VGND VPWR VPWR _7204_/Q sky130_fd_sc_hd__dfxtp_4
X_5396_ _5396_/A _5594_/B VGND VGND VPWR VPWR _5404_/S sky130_fd_sc_hd__and2_4
XFILLER_99_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7135_ _7135_/CLK _7135_/D fanout864/X VGND VGND VPWR VPWR _7135_/Q sky130_fd_sc_hd__dfrtp_2
X_4347_ _4368_/A _4722_/B VGND VGND VPWR VPWR _4467_/B sky130_fd_sc_hd__nor2_4
XFILLER_160_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7066_ _7154_/CLK _7066_/D fanout884/X VGND VGND VPWR VPWR _7066_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_143_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4278_ _5249_/A0 _6731_/Q _4279_/S VGND VGND VPWR VPWR _4278_/X sky130_fd_sc_hd__mux2_1
X_3229_ _6944_/Q VGND VGND VPWR VPWR _3229_/Y sky130_fd_sc_hd__inv_2
X_6017_ _6019_/A _6034_/B VGND VGND VPWR VPWR _6017_/Y sky130_fd_sc_hd__nor2_8
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_wbbd_sck clkbuf_0_wbbd_sck/X VGND VGND VPWR VPWR _3954_/A2 sky130_fd_sc_hd__clkbuf_8
X_6919_ _6981_/CLK _6919_/D fanout878/X VGND VGND VPWR VPWR _6919_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire715 _4577_/Y VGND VGND VPWR VPWR _4748_/A sky130_fd_sc_hd__buf_8
XFILLER_168_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire737 _4581_/A VGND VGND VPWR VPWR _4987_/A sky130_fd_sc_hd__buf_8
XFILLER_167_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length357 _5584_/S VGND VGND VPWR VPWR _5580_/S sky130_fd_sc_hd__buf_6
XFILLER_191_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold390 _6948_/Q VGND VGND VPWR VPWR hold390/X sky130_fd_sc_hd__bufbuf_16
XFILLER_104_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout870 fanout871/X VGND VGND VPWR VPWR fanout870/X sky130_fd_sc_hd__buf_8
Xfanout881 fanout883/X VGND VGND VPWR VPWR fanout881/X sky130_fd_sc_hd__buf_8
XFILLER_77_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_252 _4236_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_230 wire672/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_241 _5259_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_263 wire912/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_285 hold626/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_274 hold465/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_296 _3821_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3580_ _3238_/A _3295_/Y _4055_/A _6543_/Q _3579_/X VGND VGND VPWR VPWR _3587_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_173_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_586 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5250_ _5599_/A0 hold387/X _5251_/S VGND VGND VPWR VPWR _5250_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4201_ _6411_/A0 hold679/X _4201_/S VGND VGND VPWR VPWR _6663_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5181_ _5095_/X _5166_/X _5180_/X _5161_/X VGND VGND VPWR VPWR _5181_/X sky130_fd_sc_hd__o31a_2
X_4132_ _5247_/A0 hold569/X _4135_/S VGND VGND VPWR VPWR _6605_/D sky130_fd_sc_hd__mux2_1
X_4063_ wire794/X hold668/X _4066_/S VGND VGND VPWR VPWR _6546_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4965_ _4965_/A _4965_/B VGND VGND VPWR VPWR _5069_/D sky130_fd_sc_hd__nor2_1
XFILLER_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6704_ _7220_/CLK _6704_/D _6362_/B VGND VGND VPWR VPWR _6704_/Q sky130_fd_sc_hd__dfrtp_2
X_3916_ _3916_/A _3916_/B VGND VGND VPWR VPWR _6698_/D sky130_fd_sc_hd__nand2_1
XFILLER_149_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4896_ _4987_/A _4586_/B _4736_/B _4689_/Y VGND VGND VPWR VPWR _4905_/C sky130_fd_sc_hd__a22o_2
XFILLER_149_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6635_ _6752_/CLK _6635_/D fanout857/X VGND VGND VPWR VPWR _6635_/Q sky130_fd_sc_hd__dfrtp_2
X_3847_ _6485_/Q _3847_/B VGND VGND VPWR VPWR _3848_/S sky130_fd_sc_hd__nor2_1
X_6566_ _6623_/CLK _6566_/D fanout890/X VGND VGND VPWR VPWR _6566_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3778_ _6530_/Q _4043_/A _4304_/A _6753_/Q _3777_/X VGND VGND VPWR VPWR _3785_/A
+ sky130_fd_sc_hd__a221o_2
X_5517_ _5598_/A0 hold575/X _5517_/S VGND VGND VPWR VPWR _7080_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6497_ _6810_/CLK _6497_/D fanout853/X VGND VGND VPWR VPWR _6497_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_154_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5448_ wire746/X hold740/X _5449_/S VGND VGND VPWR VPWR _7019_/D sky130_fd_sc_hd__mux2_1
X_5379_ _5595_/A0 _6957_/Q _5386_/S VGND VGND VPWR VPWR _6957_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7118_ _7118_/CLK hold53/X fanout869/X VGND VGND VPWR VPWR _7118_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_59_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7049_ _7095_/CLK _7049_/D fanout863/X VGND VGND VPWR VPWR _7049_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire501 _7055_/Q VGND VGND VPWR VPWR wire501/X sky130_fd_sc_hd__buf_4
XFILLER_11_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire512 _7027_/Q VGND VGND VPWR VPWR wire512/X sky130_fd_sc_hd__buf_4
XFILLER_156_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire534 _6934_/Q VGND VGND VPWR VPWR wire534/X sky130_fd_sc_hd__buf_6
Xwire567 _6735_/Q VGND VGND VPWR VPWR wire567/X sky130_fd_sc_hd__buf_6
XFILLER_10_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire556 _6858_/Q VGND VGND VPWR VPWR wire556/X sky130_fd_sc_hd__buf_6
XFILLER_155_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire589 _6010_/Y VGND VGND VPWR VPWR wire589/X sky130_fd_sc_hd__buf_8
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4750_ _4965_/B _4832_/B VGND VGND VPWR VPWR _5144_/B sky130_fd_sc_hd__or2_4
XFILLER_187_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4681_ _4697_/A _4886_/B VGND VGND VPWR VPWR _5033_/B sky130_fd_sc_hd__nor2_1
X_3701_ _7046_/Q _5477_/A _4043_/A _6531_/Q _3700_/X VGND VGND VPWR VPWR _3701_/X
+ sky130_fd_sc_hd__a221o_1
X_6420_ _6420_/A _6421_/B VGND VGND VPWR VPWR _6420_/X sky130_fd_sc_hd__and2_1
X_3632_ _6626_/Q _4154_/A _4097_/A _6578_/Q _3612_/X VGND VGND VPWR VPWR _3635_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6351_ _6638_/Q wire712/X wire625/X _6613_/Q VGND VGND VPWR VPWR _6351_/X sky130_fd_sc_hd__a22o_1
X_5302_ hold150/X hold274/X _5305_/S VGND VGND VPWR VPWR _6889_/D sky130_fd_sc_hd__mux2_1
XFILLER_155_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3563_ _6856_/Q _5261_/A _4196_/A _6662_/Q VGND VGND VPWR VPWR _3563_/X sky130_fd_sc_hd__a22o_1
X_3494_ _3508_/A _3543_/B VGND VGND VPWR VPWR _4196_/A sky130_fd_sc_hd__nor2_8
X_6282_ _6356_/A _6282_/B _6282_/C VGND VGND VPWR VPWR _6282_/X sky130_fd_sc_hd__or3_1
XFILLER_170_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5233_ _5578_/A0 hold362/X _5233_/S VGND VGND VPWR VPWR _6831_/D sky130_fd_sc_hd__mux2_1
X_5164_ _5164_/A _5164_/B VGND VGND VPWR VPWR _5165_/C sky130_fd_sc_hd__nand2_1
XFILLER_130_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4115_ _5408_/A1 _6591_/Q _4117_/S VGND VGND VPWR VPWR _6591_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5095_ _5095_/A _5095_/B _5095_/C _5095_/D VGND VGND VPWR VPWR _5095_/X sky130_fd_sc_hd__or4_4
XFILLER_96_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4046_ hold834/X _6409_/A0 _4048_/S VGND VGND VPWR VPWR _6532_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5997_ _6012_/A _6018_/A _6032_/C VGND VGND VPWR VPWR _6025_/A sky130_fd_sc_hd__and3_4
XFILLER_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4948_ _4949_/B _4537_/X _4959_/A _5130_/A VGND VGND VPWR VPWR _5065_/A sky130_fd_sc_hd__a31o_4
XFILLER_12_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4879_ _5005_/C _4832_/B _4633_/X VGND VGND VPWR VPWR _5145_/A sky130_fd_sc_hd__o21ai_2
XFILLER_193_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6618_ _6623_/CLK _6618_/D fanout872/X VGND VGND VPWR VPWR _6618_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6549_ _6623_/CLK _6549_/D fanout872/X VGND VGND VPWR VPWR _6549_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_106_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput270 _6804_/Q VGND VGND VPWR VPWR pll_div[4] sky130_fd_sc_hd__buf_8
XFILLER_181_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput292 _6505_/Q VGND VGND VPWR VPWR pll_trim[25] sky130_fd_sc_hd__buf_8
Xoutput281 _6495_/Q VGND VGND VPWR VPWR pll_trim[15] sky130_fd_sc_hd__buf_8
XFILLER_181_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire364 _5251_/S VGND VGND VPWR VPWR _5249_/S sky130_fd_sc_hd__buf_6
XFILLER_116_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire375 _6232_/A VGND VGND VPWR VPWR _6306_/A sky130_fd_sc_hd__buf_6
Xwire353 _3379_/X VGND VGND VPWR VPWR wire353/X sky130_fd_sc_hd__buf_8
XFILLER_137_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire397 _3369_/Y VGND VGND VPWR VPWR _5396_/A sky130_fd_sc_hd__buf_8
Xwire386 _5429_/S VGND VGND VPWR VPWR _5431_/S sky130_fd_sc_hd__buf_8
XFILLER_152_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_559 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5920_ _6578_/Q wire684/X wire672/X _6565_/Q _5919_/X VGND VGND VPWR VPWR _5927_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5851_ _5611_/A _7181_/Q wire381/A VGND VGND VPWR VPWR _5851_/X sky130_fd_sc_hd__a21o_1
X_5782_ _3221_/A _5678_/X wire678/X _3213_/A VGND VGND VPWR VPWR _5782_/X sky130_fd_sc_hd__a22o_1
X_4802_ _4802_/A _4802_/B _4802_/C _4802_/D VGND VGND VPWR VPWR _4805_/B sky130_fd_sc_hd__or4_1
X_4733_ _4672_/A _4566_/A _4648_/B _4732_/X VGND VGND VPWR VPWR _4733_/X sky130_fd_sc_hd__o31a_2
XFILLER_175_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6403_ _4236_/A _6371_/B _6402_/X VGND VGND VPWR VPWR _6403_/X sky130_fd_sc_hd__a21o_1
XFILLER_174_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4664_ _5164_/B _4832_/B _4724_/B _4832_/A VGND VGND VPWR VPWR _4664_/X sky130_fd_sc_hd__o22a_1
XFILLER_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4595_ _4949_/C _4595_/B VGND VGND VPWR VPWR _4612_/C sky130_fd_sc_hd__nand2_2
XFILLER_162_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3615_ _6935_/Q _5351_/A _4142_/A _6616_/Q VGND VGND VPWR VPWR _3615_/X sky130_fd_sc_hd__a22o_1
XFILLER_190_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3546_ _3546_/A _3546_/B _3546_/C _3546_/D VGND VGND VPWR VPWR _3547_/D sky130_fd_sc_hd__or4_2
X_6334_ _7200_/Q _6309_/S _6333_/X VGND VGND VPWR VPWR _7200_/D sky130_fd_sc_hd__o21a_1
XFILLER_143_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6265_ _6729_/Q wire603/X _6340_/B1 _6595_/Q VGND VGND VPWR VPWR _6265_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3477_ _3973_/B _3310_/Y _3726_/A _3476_/Y VGND VGND VPWR VPWR _3477_/X sky130_fd_sc_hd__a211o_1
X_5216_ _5216_/A _5576_/B VGND VGND VPWR VPWR _5217_/S sky130_fd_sc_hd__nand2_1
X_6196_ _6891_/Q wire602/X wire581/X wire470/X _6195_/X VGND VGND VPWR VPWR _6196_/X
+ sky130_fd_sc_hd__a221o_4
X_5147_ _5147_/A _5147_/B _5147_/C VGND VGND VPWR VPWR _5148_/B sky130_fd_sc_hd__nor3_1
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5078_ _5078_/A _5078_/B _5078_/C VGND VGND VPWR VPWR _5079_/C sky130_fd_sc_hd__or3_1
XFILLER_56_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4029_ _5598_/A0 hold617/X _4033_/S VGND VGND VPWR VPWR _6517_/D sky130_fd_sc_hd__mux2_1
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_22 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold208 _6746_/Q VGND VGND VPWR VPWR hold208/X sky130_fd_sc_hd__bufbuf_16
XFILLER_172_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4380_ _4740_/A _4395_/D VGND VGND VPWR VPWR _4818_/B sky130_fd_sc_hd__nand2_8
XFILLER_172_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold219 _6617_/Q VGND VGND VPWR VPWR hold219/X sky130_fd_sc_hd__bufbuf_16
X_3400_ _7067_/Q _5495_/A _5207_/A _6817_/Q _3389_/X VGND VGND VPWR VPWR _3400_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_7_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3331_ _3331_/A _3331_/B _3331_/C _3331_/D VGND VGND VPWR VPWR _3379_/B sky130_fd_sc_hd__or4_1
XFILLER_140_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6050_ _7133_/Q _6020_/B wire640/X _6973_/Q _6049_/X VGND VGND VPWR VPWR _6057_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ hold41/X hold99/X _3953_/A VGND VGND VPWR VPWR _3262_/X sky130_fd_sc_hd__mux2_8
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5001_ _5135_/B _5001_/B _5001_/C _5001_/D VGND VGND VPWR VPWR _5001_/X sky130_fd_sc_hd__or4_1
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3193_ _6698_/Q VGND VGND VPWR VPWR _6360_/A sky130_fd_sc_hd__inv_2
XFILLER_78_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6952_ _6971_/CLK _6952_/D fanout879/X VGND VGND VPWR VPWR _6952_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_93_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6883_ _7154_/CLK _6883_/D fanout884/X VGND VGND VPWR VPWR _6883_/Q sky130_fd_sc_hd__dfrtp_2
X_5903_ _6774_/Q wire694/X wire660/X _6605_/Q _5902_/X VGND VGND VPWR VPWR _5910_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_179_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5834_ _6955_/Q _5701_/X _5707_/X wire512/X _5833_/X VGND VGND VPWR VPWR _5839_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5765_ _5663_/A _7177_/Q wire381/A VGND VGND VPWR VPWR _5765_/X sky130_fd_sc_hd__a21o_1
XFILLER_22_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4716_ _4754_/B _4724_/B VGND VGND VPWR VPWR _4797_/C sky130_fd_sc_hd__nor2_1
Xmax_length709 _5669_/X VGND VGND VPWR VPWR _5921_/A2 sky130_fd_sc_hd__buf_6
X_5696_ _5702_/B _5703_/B VGND VGND VPWR VPWR _5698_/B sky130_fd_sc_hd__and2_4
X_4647_ _4654_/B _4422_/Y _4707_/A _4236_/A VGND VGND VPWR VPWR _4917_/B sky130_fd_sc_hd__o31a_4
Xhold720 _5390_/X VGND VGND VPWR VPWR _6967_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_162_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4578_ _4818_/B _4740_/B VGND VGND VPWR VPWR _5062_/A sky130_fd_sc_hd__or2_4
Xhold753 _6616_/Q VGND VGND VPWR VPWR hold753/X sky130_fd_sc_hd__bufbuf_16
XFILLER_89_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold742 _6744_/Q VGND VGND VPWR VPWR hold742/X sky130_fd_sc_hd__bufbuf_16
X_6317_ _6756_/Q _6339_/A2 _6339_/B1 _6771_/Q VGND VGND VPWR VPWR _6317_/X sky130_fd_sc_hd__a22o_1
Xhold764 _6719_/Q VGND VGND VPWR VPWR hold764/X sky130_fd_sc_hd__bufbuf_16
Xhold731 _6647_/Q VGND VGND VPWR VPWR hold731/X sky130_fd_sc_hd__bufbuf_16
Xhold775 _7053_/Q VGND VGND VPWR VPWR hold775/X sky130_fd_sc_hd__bufbuf_16
Xhold797 _6509_/Q VGND VGND VPWR VPWR hold797/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold786 _6589_/Q VGND VGND VPWR VPWR hold786/X sky130_fd_sc_hd__bufbuf_16
X_3529_ _3543_/A hold45/X VGND VGND VPWR VPWR _4112_/A sky130_fd_sc_hd__nor2_8
XFILLER_103_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6248_ _6248_/A _6248_/B _6248_/C VGND VGND VPWR VPWR _6248_/X sky130_fd_sc_hd__or3_4
X_6179_ _6866_/Q _6179_/A2 _6029_/X wire504/X _6178_/X VGND VGND VPWR VPWR _6181_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold80 hold80/A VGND VGND VPWR VPWR hold80/X sky130_fd_sc_hd__bufbuf_16
Xhold91 hold91/A VGND VGND VPWR VPWR hold91/X sky130_fd_sc_hd__bufbuf_16
XFILLER_90_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3880_ _3875_/B _3848_/S _3879_/X _6457_/Q VGND VGND VPWR VPWR _6457_/D sky130_fd_sc_hd__a22o_1
XFILLER_188_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5550_ _7109_/Q _5595_/A0 _5557_/S VGND VGND VPWR VPWR _7109_/D sky130_fd_sc_hd__mux2_1
XFILLER_157_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4501_ _4501_/A _4812_/A VGND VGND VPWR VPWR _4672_/B sky130_fd_sc_hd__nor2_2
XFILLER_145_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5481_ hold601/X wire769/X _5485_/S VGND VGND VPWR VPWR _7048_/D sky130_fd_sc_hd__mux2_1
X_4432_ _4735_/A _4672_/A VGND VGND VPWR VPWR _4470_/B sky130_fd_sc_hd__nor2_8
XFILLER_117_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7220_ _7220_/CLK _7220_/D _6362_/B VGND VGND VPWR VPWR hold68/A sky130_fd_sc_hd__dfrtp_1
XFILLER_144_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4363_ _5050_/A _4413_/C VGND VGND VPWR VPWR _4364_/B sky130_fd_sc_hd__and2_2
X_7151_ _7151_/CLK _7151_/D fanout881/X VGND VGND VPWR VPWR _7151_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_113_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6102_ _6959_/Q wire624/X wire613/X _7055_/Q VGND VGND VPWR VPWR _6102_/X sky130_fd_sc_hd__a22o_1
XFILLER_98_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4294_ wire790/X hold742/X _4297_/S VGND VGND VPWR VPWR _6744_/D sky130_fd_sc_hd__mux2_1
X_3314_ _3314_/A _3314_/B VGND VGND VPWR VPWR _3551_/A sky130_fd_sc_hd__or2_4
X_7082_ _7082_/CLK _7082_/D fanout868/X VGND VGND VPWR VPWR _7082_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_140_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3245_ _4395_/D VGND VGND VPWR VPWR _4819_/A sky130_fd_sc_hd__inv_4
XFILLER_112_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6033_ _6037_/B _6037_/C _6033_/C VGND VGND VPWR VPWR _6033_/X sky130_fd_sc_hd__and3_4
XFILLER_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6935_ _7128_/CLK _6935_/D _6421_/A VGND VGND VPWR VPWR _6935_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6866_ _7154_/CLK _6866_/D fanout886/X VGND VGND VPWR VPWR _6866_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_167_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5817_ _7010_/Q wire701/X wire679/X _7074_/Q VGND VGND VPWR VPWR _5817_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6797_ _3545_/A1 _6797_/D _6455_/X VGND VGND VPWR VPWR _6797_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_50_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire908 wire908/A VGND VGND VPWR VPWR wire908/X sky130_fd_sc_hd__buf_4
X_5748_ _7015_/Q wire697/X wire691/X _7087_/Q _5747_/X VGND VGND VPWR VPWR _5753_/B
+ sky130_fd_sc_hd__a221o_4
XFILLER_10_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length517 _7010_/Q VGND VGND VPWR VPWR _6173_/B2 sky130_fd_sc_hd__buf_6
XFILLER_136_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5679_ _7164_/Q _7163_/Q VGND VGND VPWR VPWR _5707_/C sky130_fd_sc_hd__and2b_4
XFILLER_151_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold561 _6928_/Q VGND VGND VPWR VPWR hold561/X sky130_fd_sc_hd__bufbuf_16
XFILLER_135_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold572 _5255_/X VGND VGND VPWR VPWR _6847_/D sky130_fd_sc_hd__bufbuf_16
Xhold550 _6846_/Q VGND VGND VPWR VPWR hold550/X sky130_fd_sc_hd__bufbuf_16
XFILLER_173_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold583 _5413_/X VGND VGND VPWR VPWR _6988_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold594 _6718_/Q VGND VGND VPWR VPWR hold594/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput170 wb_we_i VGND VGND VPWR VPWR _6372_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_48_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4981_ _5003_/A _5102_/D VGND VGND VPWR VPWR _5121_/B sky130_fd_sc_hd__nand2_2
XFILLER_63_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3932_ _3204_/Y input90/X _3932_/S VGND VGND VPWR VPWR _3932_/X sky130_fd_sc_hd__mux2_8
X_6720_ _6720_/CLK _6720_/D fanout874/X VGND VGND VPWR VPWR _6720_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6651_ _6842_/CLK _6651_/D fanout857/X VGND VGND VPWR VPWR _6651_/Q sky130_fd_sc_hd__dfstp_4
X_3863_ _6469_/Q _3864_/B _3862_/Y _6468_/Q VGND VGND VPWR VPWR _6469_/D sky130_fd_sc_hd__o22a_1
X_5602_ _5602_/A0 hold354/X hold66/X VGND VGND VPWR VPWR _5602_/X sky130_fd_sc_hd__mux2_1
X_6582_ _7208_/CLK _6582_/D VGND VGND VPWR VPWR _6582_/Q sky130_fd_sc_hd__dfxtp_2
X_3794_ _3794_/A _3794_/B _3794_/C _3794_/D VGND VGND VPWR VPWR _3794_/X sky130_fd_sc_hd__or4_1
X_5533_ _5578_/A0 _7094_/Q _5539_/S VGND VGND VPWR VPWR _7094_/D sky130_fd_sc_hd__mux2_1
XFILLER_191_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5464_ hold156/X hold403/X _5467_/S VGND VGND VPWR VPWR _7033_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_60_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7132_/CLK sky130_fd_sc_hd__clkbuf_8
X_4415_ _4529_/A _4529_/B _4414_/B _4533_/A VGND VGND VPWR VPWR _4415_/X sky130_fd_sc_hd__a31o_2
X_5395_ _5602_/A0 hold368/X _5395_/S VGND VGND VPWR VPWR _6972_/D sky130_fd_sc_hd__mux2_1
XFILLER_105_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7203_ _7210_/CLK _7203_/D VGND VGND VPWR VPWR _7203_/Q sky130_fd_sc_hd__dfxtp_4
X_4346_ _4722_/B _4345_/Y _4346_/S VGND VGND VPWR VPWR _4533_/A sky130_fd_sc_hd__mux2_8
XFILLER_132_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7134_ _7134_/CLK _7134_/D fanout864/X VGND VGND VPWR VPWR _7134_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_101_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7065_ _7153_/CLK _7065_/D fanout882/X VGND VGND VPWR VPWR _7065_/Q sky130_fd_sc_hd__dfrtp_2
Xclkbuf_leaf_75_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6771_/CLK sky130_fd_sc_hd__clkbuf_8
X_4277_ _6409_/A0 _6730_/Q _4279_/S VGND VGND VPWR VPWR _6730_/D sky130_fd_sc_hd__mux2_1
X_3228_ _6952_/Q VGND VGND VPWR VPWR _3228_/Y sky130_fd_sc_hd__inv_2
X_6016_ _6032_/A _6035_/A _6018_/A VGND VGND VPWR VPWR _6022_/C sky130_fd_sc_hd__and3_4
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6918_ _6981_/CLK _6918_/D fanout878/X VGND VGND VPWR VPWR _6918_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_168_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_13_csclk _6708_/CLK VGND VGND VPWR VPWR _6621_/CLK sky130_fd_sc_hd__clkbuf_8
X_6849_ _6994_/CLK _6849_/D fanout870/X VGND VGND VPWR VPWR _6849_/Q sky130_fd_sc_hd__dfrtp_1
Xwire716 _4592_/B VGND VGND VPWR VPWR _4947_/B sky130_fd_sc_hd__buf_8
XFILLER_168_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire749 hold57/X VGND VGND VPWR VPWR wire749/X sky130_fd_sc_hd__buf_8
XFILLER_6_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_28_csclk _6987_/CLK VGND VGND VPWR VPWR _6980_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_184_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold380 _6860_/Q VGND VGND VPWR VPWR hold380/X sky130_fd_sc_hd__bufbuf_16
XFILLER_104_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold391 _7078_/Q VGND VGND VPWR VPWR hold391/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout882 fanout883/X VGND VGND VPWR VPWR fanout882/X sky130_fd_sc_hd__buf_8
Xfanout871 fanout871/A VGND VGND VPWR VPWR fanout871/X sky130_fd_sc_hd__buf_8
XFILLER_133_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_242 hold199/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_231 wire672/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_220 wire570/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_286 _6672_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_275 hold465/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_253 _3938_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_264 _3938_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_297 _3876_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length892 fanout871/A VGND VGND VPWR VPWR fanout868/A sky130_fd_sc_hd__buf_8
XFILLER_181_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4200_ _5249_/A0 hold441/X _4201_/S VGND VGND VPWR VPWR _6662_/D sky130_fd_sc_hd__mux2_1
X_5180_ _5180_/A _5180_/B _5180_/C _5179_/X VGND VGND VPWR VPWR _5180_/X sky130_fd_sc_hd__or4b_1
X_4131_ _5487_/A0 hold772/X _4135_/S VGND VGND VPWR VPWR _6604_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4062_ _5487_/A0 hold795/X _4066_/S VGND VGND VPWR VPWR _6545_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4964_ _4536_/B _4959_/X _4906_/C VGND VGND VPWR VPWR _5174_/D sky130_fd_sc_hd__a21o_1
XFILLER_91_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6703_ _7220_/CLK _6703_/D _6362_/B VGND VGND VPWR VPWR _6703_/Q sky130_fd_sc_hd__dfrtp_2
X_3915_ _6360_/A _3915_/B VGND VGND VPWR VPWR _3916_/B sky130_fd_sc_hd__or2_1
XFILLER_20_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4895_ _4987_/A _4409_/Y _4736_/B _4748_/B VGND VGND VPWR VPWR _5129_/A sky130_fd_sc_hd__a22o_1
XFILLER_149_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6634_ _6752_/CLK _6634_/D fanout857/X VGND VGND VPWR VPWR _6634_/Q sky130_fd_sc_hd__dfrtp_2
X_3846_ _3196_/Y _6665_/Q _3201_/Y _3859_/B _6475_/Q VGND VGND VPWR VPWR _6475_/D
+ sky130_fd_sc_hd__a41o_1
XFILLER_164_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6565_ _6720_/CLK _6565_/D fanout873/X VGND VGND VPWR VPWR _6565_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_138_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3777_ _7077_/Q _5513_/A _4178_/A _6644_/Q VGND VGND VPWR VPWR _3777_/X sky130_fd_sc_hd__a22o_1
X_5516_ wire786/X hold384/X _5521_/S VGND VGND VPWR VPWR _7079_/D sky130_fd_sc_hd__mux2_1
X_6496_ _6810_/CLK _6496_/D fanout853/X VGND VGND VPWR VPWR _6496_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_145_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5447_ _5519_/A0 hold833/X _5449_/S VGND VGND VPWR VPWR _7018_/D sky130_fd_sc_hd__mux2_1
XFILLER_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5378_ _5378_/A _5378_/B VGND VGND VPWR VPWR _5386_/S sky130_fd_sc_hd__nand2_8
XFILLER_160_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7117_ _7133_/CLK _7117_/D fanout883/X VGND VGND VPWR VPWR _7117_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_120_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4329_ _6407_/A0 hold747/X _4333_/S VGND VGND VPWR VPWR _6773_/D sky130_fd_sc_hd__mux2_1
XFILLER_170_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7048_ _7132_/CLK _7048_/D fanout863/X VGND VGND VPWR VPWR _7048_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_86_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire502 _7054_/Q VGND VGND VPWR VPWR wire502/X sky130_fd_sc_hd__buf_6
Xwire513 wire513/A VGND VGND VPWR VPWR _3219_/A sky130_fd_sc_hd__buf_6
Xwire524 _6992_/Q VGND VGND VPWR VPWR _3223_/A sky130_fd_sc_hd__buf_8
Xwire546 _6878_/Q VGND VGND VPWR VPWR wire546/X sky130_fd_sc_hd__buf_6
XFILLER_156_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire535 _6930_/Q VGND VGND VPWR VPWR wire535/X sky130_fd_sc_hd__buf_6
Xwire557 _6823_/Q VGND VGND VPWR VPWR wire557/X sky130_fd_sc_hd__buf_6
XFILLER_170_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire579 _6030_/Y VGND VGND VPWR VPWR wire579/X sky130_fd_sc_hd__buf_8
XFILLER_6_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire568 _6661_/Q VGND VGND VPWR VPWR wire568/X sky130_fd_sc_hd__clkbuf_8
XFILLER_124_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3700_ _6551_/Q _3473_/Y _4196_/A _6660_/Q VGND VGND VPWR VPWR _3700_/X sky130_fd_sc_hd__a22o_1
X_4680_ _5099_/A _5024_/A _4680_/C _4670_/X VGND VGND VPWR VPWR _4708_/D sky130_fd_sc_hd__or4b_1
X_3631_ _6903_/Q _5315_/A _5279_/A _6871_/Q _3611_/X VGND VGND VPWR VPWR _3635_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6350_ _6544_/Q wire592/X wire590/X _6567_/Q _6349_/X VGND VGND VPWR VPWR _6355_/B
+ sky130_fd_sc_hd__a221o_1
X_3562_ _6652_/Q _4184_/A _4286_/A _6741_/Q VGND VGND VPWR VPWR _3562_/X sky130_fd_sc_hd__a22o_4
X_5301_ wire773/A hold347/X _5305_/S VGND VGND VPWR VPWR _5301_/X sky130_fd_sc_hd__mux2_1
X_6281_ _6281_/A _6281_/B _6281_/C _6281_/D VGND VGND VPWR VPWR _6282_/C sky130_fd_sc_hd__or4_4
X_3493_ _3514_/A _3493_/B VGND VGND VPWR VPWR _4274_/A sky130_fd_sc_hd__nor2_8
XFILLER_142_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_579 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5232_ wire746/X hold732/X _5233_/S VGND VGND VPWR VPWR _5232_/X sky130_fd_sc_hd__mux2_1
X_5163_ _5163_/A _5163_/B _5163_/C VGND VGND VPWR VPWR _5163_/X sky130_fd_sc_hd__or3_1
XFILLER_130_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4114_ _5247_/A0 hold510/X _4117_/S VGND VGND VPWR VPWR _6590_/D sky130_fd_sc_hd__mux2_1
X_5094_ _4395_/D _4987_/B _4586_/B _5116_/A _4797_/C VGND VGND VPWR VPWR _5095_/D
+ sky130_fd_sc_hd__a311o_1
XFILLER_84_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4045_ hold701/X _6408_/A0 _4048_/S VGND VGND VPWR VPWR _6531_/D sky130_fd_sc_hd__mux2_1
XFILLER_49_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5996_ _6012_/A _6037_/C _6032_/C VGND VGND VPWR VPWR _5996_/X sky130_fd_sc_hd__and3_4
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4947_ _4986_/C _4947_/B VGND VGND VPWR VPWR _4959_/A sky130_fd_sc_hd__nand2_8
XFILLER_24_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4878_ _4878_/A VGND VGND VPWR VPWR _5130_/A sky130_fd_sc_hd__inv_2
XFILLER_32_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6617_ _6712_/CLK _6617_/D fanout872/X VGND VGND VPWR VPWR _6617_/Q sky130_fd_sc_hd__dfrtp_2
X_3829_ _3828_/X _6481_/Q _3840_/S VGND VGND VPWR VPWR _6481_/D sky130_fd_sc_hd__mux2_1
XFILLER_106_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6548_ _6623_/CLK _6548_/D fanout872/X VGND VGND VPWR VPWR _6548_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_4_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6479_ _3957_/A1 _6479_/D _6434_/X VGND VGND VPWR VPWR hold40/A sky130_fd_sc_hd__dfrtp_2
XFILLER_121_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput260 _3962_/A VGND VGND VPWR VPWR pad_flash_io1_oeb sky130_fd_sc_hd__buf_8
Xoutput271 _6798_/Q VGND VGND VPWR VPWR pll_ena sky130_fd_sc_hd__buf_8
XFILLER_99_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput293 _6498_/Q VGND VGND VPWR VPWR pll_trim[2] sky130_fd_sc_hd__buf_8
Xoutput282 _6811_/Q VGND VGND VPWR VPWR pll_trim[16] sky130_fd_sc_hd__buf_8
XFILLER_101_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire365 _5248_/S VGND VGND VPWR VPWR _5251_/S sky130_fd_sc_hd__buf_8
Xwire354 _3351_/X VGND VGND VPWR VPWR _3378_/C sky130_fd_sc_hd__buf_4
XFILLER_11_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire376 _5814_/X VGND VGND VPWR VPWR _5827_/A sky130_fd_sc_hd__buf_4
XFILLER_139_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire387 _3944_/X VGND VGND VPWR VPWR wire387/X sky130_fd_sc_hd__buf_6
XFILLER_171_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5850_ _6859_/Q _5698_/Y _5839_/X _5849_/X _3921_/A VGND VGND VPWR VPWR _5850_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_61_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5781_ _7096_/Q _5856_/A2 _5693_/X _7080_/Q _5780_/X VGND VGND VPWR VPWR _5784_/B
+ sky130_fd_sc_hd__a221o_1
X_4801_ _4758_/C _4719_/X _4789_/X _4800_/X _5078_/A VGND VGND VPWR VPWR _4802_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_34_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4732_ _4562_/B _4812_/C _4723_/X _4727_/Y _4731_/X VGND VGND VPWR VPWR _4732_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4663_ _4663_/A _4663_/B VGND VGND VPWR VPWR _4724_/B sky130_fd_sc_hd__or2_4
X_6402_ _4236_/C _6402_/A2 _6372_/B _4236_/B VGND VGND VPWR VPWR _6402_/X sky130_fd_sc_hd__a22o_1
X_3614_ _7151_/Q hold64/A wire388/X wire558/X VGND VGND VPWR VPWR _3614_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4594_ _4871_/A _4592_/B _4812_/A VGND VGND VPWR VPWR _4595_/B sky130_fd_sc_hd__a21oi_4
XFILLER_115_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3545_ _3545_/A1 _3361_/Y _4055_/A _6544_/Q _3544_/X VGND VGND VPWR VPWR _3546_/D
+ sky130_fd_sc_hd__a221o_2
X_6333_ wire824/X _7199_/Q wire381/X _6332_/X VGND VGND VPWR VPWR _6333_/X sky130_fd_sc_hd__a211o_1
XFILLER_135_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3476_ _5225_/A _3520_/B VGND VGND VPWR VPWR _3476_/Y sky130_fd_sc_hd__nor2_4
X_6264_ _6749_/Q wire575/X _6335_/B _6774_/Q _6261_/X VGND VGND VPWR VPWR _6269_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_142_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5215_ _6818_/Q wire739/X _5215_/S VGND VGND VPWR VPWR _6818_/D sky130_fd_sc_hd__mux2_1
X_6195_ _7115_/Q wire650/X _6021_/B _7155_/Q VGND VGND VPWR VPWR _6195_/X sky130_fd_sc_hd__a22o_1
XFILLER_69_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5146_ _5146_/A _5146_/B VGND VGND VPWR VPWR _5146_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5077_ _5121_/A _5121_/B VGND VGND VPWR VPWR _5077_/Y sky130_fd_sc_hd__nor2_1
XFILLER_178_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4028_ _5248_/A0 hold217/X _4033_/S VGND VGND VPWR VPWR _6516_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5979_ _6752_/Q _5979_/A2 wire662/X _6544_/Q VGND VGND VPWR VPWR _5979_/X sky130_fd_sc_hd__a22o_1
XFILLER_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold209 _4296_/X VGND VGND VPWR VPWR _6746_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_144_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3330_ _6972_/Q _5387_/A _3736_/A2 input51/X _3326_/X VGND VGND VPWR VPWR _3331_/D
+ sky130_fd_sc_hd__a221o_4
XFILLER_125_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5000_ _5121_/B _5081_/C _5000_/C _5136_/D VGND VGND VPWR VPWR _5001_/D sky130_fd_sc_hd__or4_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ hold40/X hold59/X _3845_/A VGND VGND VPWR VPWR hold41/A sky130_fd_sc_hd__mux2_1
XFILLER_66_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3192_ _6459_/Q VGND VGND VPWR VPWR _3192_/Y sky130_fd_sc_hd__inv_2
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6951_ _6951_/CLK _6951_/D _6421_/A VGND VGND VPWR VPWR _6951_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_93_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6882_ _6979_/CLK _6882_/D fanout884/X VGND VGND VPWR VPWR _6882_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_62_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5902_ _6729_/Q wire710/X wire689/X _6640_/Q VGND VGND VPWR VPWR _5902_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5833_ _6915_/Q wire699/X wire666/X wire553/X VGND VGND VPWR VPWR _5833_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5764_ _6855_/Q _5698_/Y _5753_/X _5763_/X _6109_/S VGND VGND VPWR VPWR _5764_/X
+ sky130_fd_sc_hd__o221a_4
X_4715_ _4453_/Y _4692_/C _4695_/X _5166_/A VGND VGND VPWR VPWR _4797_/B sky130_fd_sc_hd__a31o_1
X_5695_ _7077_/Q _5693_/X wire672/X _6893_/Q VGND VGND VPWR VPWR _5695_/X sky130_fd_sc_hd__a22o_1
XFILLER_175_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4646_ _4774_/A _4774_/C VGND VGND VPWR VPWR _4707_/A sky130_fd_sc_hd__or2_2
XFILLER_162_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4577_ _4818_/B _4740_/B VGND VGND VPWR VPWR _4577_/Y sky130_fd_sc_hd__nor2_1
Xhold721 _6895_/Q VGND VGND VPWR VPWR hold721/X sky130_fd_sc_hd__bufbuf_16
XFILLER_146_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold710 _7043_/Q VGND VGND VPWR VPWR hold710/X sky130_fd_sc_hd__bufbuf_16
XFILLER_150_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold732 _6830_/Q VGND VGND VPWR VPWR hold732/X sky130_fd_sc_hd__bufbuf_16
Xhold743 _6535_/Q VGND VGND VPWR VPWR hold743/X sky130_fd_sc_hd__bufbuf_16
Xhold754 _6805_/Q VGND VGND VPWR VPWR hold754/X sky130_fd_sc_hd__bufbuf_16
X_6316_ _6751_/Q wire575/X _6335_/B _6776_/Q _6311_/X VGND VGND VPWR VPWR _6321_/B
+ sky130_fd_sc_hd__a221o_1
X_3528_ _5252_/A _3528_/B VGND VGND VPWR VPWR _4160_/A sky130_fd_sc_hd__nor2_8
Xhold787 _6811_/Q VGND VGND VPWR VPWR hold787/X sky130_fd_sc_hd__bufbuf_16
XFILLER_1_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold765 _4264_/X VGND VGND VPWR VPWR _6719_/D sky130_fd_sc_hd__bufbuf_16
Xhold776 _6644_/Q VGND VGND VPWR VPWR hold776/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold798 _6833_/Q VGND VGND VPWR VPWR hold798/X sky130_fd_sc_hd__bufbuf_16
XFILLER_130_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6247_ _6247_/A _6247_/B _6247_/C _6247_/D VGND VGND VPWR VPWR _6248_/C sky130_fd_sc_hd__or4_1
XFILLER_103_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3459_ _3508_/A _5252_/B VGND VGND VPWR VPWR _4316_/A sky130_fd_sc_hd__nor2_8
XFILLER_39_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6178_ _7106_/Q wire712/X wire625/X _6946_/Q VGND VGND VPWR VPWR _6178_/X sky130_fd_sc_hd__a22o_4
X_5129_ _5129_/A _5129_/B _5123_/C _5123_/B VGND VGND VPWR VPWR _5130_/C sky130_fd_sc_hd__or4bb_1
XFILLER_69_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold92 hold92/A VGND VGND VPWR VPWR hold92/X sky130_fd_sc_hd__bufbuf_16
Xhold81 hold81/A VGND VGND VPWR VPWR hold81/X sky130_fd_sc_hd__bufbuf_16
XFILLER_152_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold70 hold70/A VGND VGND VPWR VPWR hold70/X sky130_fd_sc_hd__bufbuf_16
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4500_ _4500_/A _4586_/B VGND VGND VPWR VPWR _5116_/A sky130_fd_sc_hd__and2_2
X_5480_ wire507/X wire780/X _5485_/S VGND VGND VPWR VPWR _7047_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4431_ _4992_/A _4851_/B _4499_/C _4507_/A VGND VGND VPWR VPWR _4539_/D sky130_fd_sc_hd__o211a_4
XFILLER_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1 _6413_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4362_ _5050_/A _4413_/C VGND VGND VPWR VPWR _4364_/A sky130_fd_sc_hd__nor2_2
X_7150_ _7151_/CLK hold67/X fanout880/X VGND VGND VPWR VPWR _7150_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_125_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4293_ _5487_/A0 hold789/X _4297_/S VGND VGND VPWR VPWR _6743_/D sky130_fd_sc_hd__mux2_1
X_6101_ _6903_/Q wire600/X wire645/X _6935_/Q _6100_/X VGND VGND VPWR VPWR _6106_/B
+ sky130_fd_sc_hd__a221o_1
X_3313_ _6964_/Q _5378_/A _5342_/A _6932_/Q _3312_/X VGND VGND VPWR VPWR _3313_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7081_ _7081_/CLK _7081_/D fanout871/X VGND VGND VPWR VPWR _7081_/Q sky130_fd_sc_hd__dfrtp_2
X_3244_ _4469_/A VGND VGND VPWR VPWR _4740_/A sky130_fd_sc_hd__clkinv_16
XFILLER_140_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6032_ _6032_/A _6037_/C _6032_/C VGND VGND VPWR VPWR _6032_/X sky130_fd_sc_hd__and3_4
XFILLER_100_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6934_ _7128_/CLK _6934_/D _6421_/A VGND VGND VPWR VPWR _6934_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_54_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6865_ _7096_/CLK _6865_/D fanout883/X VGND VGND VPWR VPWR _6865_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_179_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6796_ _3545_/A1 _6796_/D _6454_/X VGND VGND VPWR VPWR _6796_/Q sky130_fd_sc_hd__dfrtn_1
X_5816_ _7098_/Q _5856_/A2 wire677/X _7082_/Q _5815_/X VGND VGND VPWR VPWR _5827_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire909 wire909/A VGND VGND VPWR VPWR _3973_/B sky130_fd_sc_hd__buf_8
X_5747_ _6991_/Q wire692/X wire678/X _7071_/Q VGND VGND VPWR VPWR _5747_/X sky130_fd_sc_hd__a22o_1
XFILLER_157_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5678_ _7165_/Q _5705_/B _5703_/B VGND VGND VPWR VPWR _5678_/X sky130_fd_sc_hd__and3_4
X_4629_ _4996_/A _4749_/C VGND VGND VPWR VPWR _5079_/B sky130_fd_sc_hd__nor2_4
XFILLER_190_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold562 _6525_/Q VGND VGND VPWR VPWR hold562/X sky130_fd_sc_hd__bufbuf_16
Xhold540 _6919_/Q VGND VGND VPWR VPWR hold540/X sky130_fd_sc_hd__bufbuf_16
Xhold551 _5254_/X VGND VGND VPWR VPWR _6846_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_131_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold584 _6685_/Q VGND VGND VPWR VPWR hold584/X sky130_fd_sc_hd__bufbuf_16
Xhold595 _6827_/Q VGND VGND VPWR VPWR hold595/X sky130_fd_sc_hd__bufbuf_16
XFILLER_1_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold573 _7036_/Q VGND VGND VPWR VPWR hold573/X sky130_fd_sc_hd__bufbuf_16
XFILLER_106_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput160 wb_dat_i[6] VGND VGND VPWR VPWR _6396_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_110_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4980_ _4980_/A _4980_/B _4980_/C _4367_/X VGND VGND VPWR VPWR _5121_/A sky130_fd_sc_hd__or4b_4
XFILLER_91_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3931_ _3203_/Y input92/X _3932_/S VGND VGND VPWR VPWR _3931_/X sky130_fd_sc_hd__mux2_8
XFILLER_177_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6650_ _6650_/CLK _6650_/D fanout858/X VGND VGND VPWR VPWR _6650_/Q sky130_fd_sc_hd__dfrtp_2
X_3862_ _6469_/Q _3866_/B _3864_/B VGND VGND VPWR VPWR _3862_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_177_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5601_ _5601_/A0 hold292/X hold66/X VGND VGND VPWR VPWR _5601_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6581_ _7208_/CLK _6581_/D VGND VGND VPWR VPWR _6581_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_192_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5532_ _5532_/A0 hold716/X _5539_/S VGND VGND VPWR VPWR _7093_/D sky130_fd_sc_hd__mux2_1
X_3793_ _3793_/A _3793_/B _3793_/C _3793_/D VGND VGND VPWR VPWR _3794_/D sky130_fd_sc_hd__or4_4
XFILLER_157_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_9_csclk _6708_/CLK VGND VGND VPWR VPWR _6632_/CLK sky130_fd_sc_hd__clkbuf_8
X_5463_ wire769/X hold609/X _5467_/S VGND VGND VPWR VPWR _7032_/D sky130_fd_sc_hd__mux2_1
X_4414_ _4529_/B _4414_/B VGND VGND VPWR VPWR _4416_/B sky130_fd_sc_hd__nand2_8
X_5394_ hold57/X hold270/X _5395_/S VGND VGND VPWR VPWR _6971_/D sky130_fd_sc_hd__mux2_1
X_7202_ _7220_/CLK _7202_/D _6362_/B VGND VGND VPWR VPWR _7202_/Q sky130_fd_sc_hd__dfrtp_2
X_4345_ _4345_/A _4345_/B VGND VGND VPWR VPWR _4345_/Y sky130_fd_sc_hd__nand2_1
X_7133_ _7133_/CLK _7133_/D fanout883/X VGND VGND VPWR VPWR _7133_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_99_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7064_ _7145_/CLK _7064_/D _6421_/A VGND VGND VPWR VPWR _7064_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_140_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4276_ wire790/X hold462/X _4279_/S VGND VGND VPWR VPWR _6729_/D sky130_fd_sc_hd__mux2_1
X_3227_ _6960_/Q VGND VGND VPWR VPWR _3227_/Y sky130_fd_sc_hd__inv_2
X_6015_ _6037_/B _6018_/A _6032_/C VGND VGND VPWR VPWR _6022_/B sky130_fd_sc_hd__and3_4
XFILLER_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6917_ _6981_/CLK _6917_/D fanout878/X VGND VGND VPWR VPWR _6917_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_54_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6848_ _6992_/CLK _6848_/D fanout868/X VGND VGND VPWR VPWR _6848_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_52_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire706 _5674_/X VGND VGND VPWR VPWR wire706/X sky130_fd_sc_hd__buf_8
XFILLER_10_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire717 _4617_/B VGND VGND VPWR VPWR _4989_/A sky130_fd_sc_hd__buf_8
X_6779_ _7218_/CLK _6779_/D _6362_/B VGND VGND VPWR VPWR _6779_/Q sky130_fd_sc_hd__dfrtp_2
Xwire728 _5459_/B VGND VGND VPWR VPWR _5585_/B sky130_fd_sc_hd__buf_8
Xwire739 wire739/A VGND VGND VPWR VPWR wire739/X sky130_fd_sc_hd__buf_8
XFILLER_182_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length359 _5538_/S VGND VGND VPWR VPWR _5539_/S sky130_fd_sc_hd__buf_8
XFILLER_136_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold370 _7068_/Q VGND VGND VPWR VPWR hold370/X sky130_fd_sc_hd__bufbuf_16
XFILLER_117_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold381 _5269_/X VGND VGND VPWR VPWR _6860_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_117_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold392 _7124_/Q VGND VGND VPWR VPWR hold392/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout861 fanout871/A VGND VGND VPWR VPWR fanout861/X sky130_fd_sc_hd__buf_8
Xfanout850 _6447_/A VGND VGND VPWR VPWR fanout850/X sky130_fd_sc_hd__buf_8
Xfanout883 fanout889/X VGND VGND VPWR VPWR fanout883/X sky130_fd_sc_hd__buf_8
Xfanout872 fanout873/X VGND VGND VPWR VPWR fanout872/X sky130_fd_sc_hd__buf_8
XFILLER_46_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_243 hold57/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_232 wire672/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_210 _3220_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_221 wire571/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_276 hold465/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_265 hold38/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_254 wire835/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_287 hold808/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_298 _4235_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length893 fanout891/X VGND VGND VPWR VPWR fanout871/A sky130_fd_sc_hd__buf_8
X_4130_ _4130_/A _4154_/B VGND VGND VPWR VPWR _4135_/S sky130_fd_sc_hd__nand2_8
XFILLER_122_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4061_ _4061_/A _4154_/B VGND VGND VPWR VPWR _4066_/S sky130_fd_sc_hd__nand2_4
XFILLER_37_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4963_ _4971_/B VGND VGND VPWR VPWR _4963_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6702_ _7210_/CLK _6702_/D _6362_/B VGND VGND VPWR VPWR _6702_/Q sky130_fd_sc_hd__dfrtp_2
X_3914_ _6706_/Q _3883_/X _6701_/Q VGND VGND VPWR VPWR _6706_/D sky130_fd_sc_hd__a21o_1
XFILLER_149_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4894_ _4956_/C _4689_/Y _4617_/Y VGND VGND VPWR VPWR _4906_/C sky130_fd_sc_hd__a21o_1
X_6633_ _6633_/CLK _6633_/D fanout858/X VGND VGND VPWR VPWR _6633_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_60_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3845_ _3845_/A _6664_/Q VGND VGND VPWR VPWR _3859_/B sky130_fd_sc_hd__nor2_8
XFILLER_138_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6564_ _6650_/CLK _6564_/D fanout890/X VGND VGND VPWR VPWR _6564_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3776_ _6800_/Q _5194_/A _3771_/X _3773_/X _3775_/X VGND VGND VPWR VPWR _3793_/B
+ sky130_fd_sc_hd__a2111o_2
X_6495_ _6815_/CLK _6495_/D fanout855/X VGND VGND VPWR VPWR _6495_/Q sky130_fd_sc_hd__dfstp_4
X_5515_ _5578_/A0 hold391/X _5521_/S VGND VGND VPWR VPWR _7078_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5446_ _5572_/A0 hold518/X _5449_/S VGND VGND VPWR VPWR _7017_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5377_ hold21/X _6956_/Q _5377_/S VGND VGND VPWR VPWR hold22/A sky130_fd_sc_hd__mux2_1
X_7116_ _7156_/CLK _7116_/D fanout884/X VGND VGND VPWR VPWR _7116_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_113_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4328_ _4328_/A _6406_/B VGND VGND VPWR VPWR _4333_/S sky130_fd_sc_hd__nand2_4
X_4259_ _6715_/Q _5498_/A0 _4261_/S VGND VGND VPWR VPWR _6715_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7047_ _7134_/CLK _7047_/D fanout864/X VGND VGND VPWR VPWR _7047_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire503 _7053_/Q VGND VGND VPWR VPWR wire503/X sky130_fd_sc_hd__buf_8
XFILLER_168_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire536 _6914_/Q VGND VGND VPWR VPWR wire536/X sky130_fd_sc_hd__buf_4
Xwire525 _6980_/Q VGND VGND VPWR VPWR wire525/X sky130_fd_sc_hd__buf_6
Xwire547 _6874_/Q VGND VGND VPWR VPWR wire547/X sky130_fd_sc_hd__buf_6
Xwire558 _6822_/Q VGND VGND VPWR VPWR wire558/X sky130_fd_sc_hd__buf_6
XFILLER_109_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire569 _6658_/Q VGND VGND VPWR VPWR wire569/X sky130_fd_sc_hd__buf_6
XFILLER_124_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_74_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6815_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_159_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3630_ _6927_/Q _5342_/A _4136_/A _6611_/Q _3618_/X VGND VGND VPWR VPWR _3635_/A
+ sky130_fd_sc_hd__a221o_1
X_3561_ _6992_/Q _5414_/A _5468_/A _7040_/Q VGND VGND VPWR VPWR _3561_/X sky130_fd_sc_hd__a22o_2
X_5300_ _5597_/A0 hold285/X _5305_/S VGND VGND VPWR VPWR _6887_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3492_ _6889_/Q _5297_/A wire391/X _6789_/Q _3490_/X VGND VGND VPWR VPWR _3504_/A
+ sky130_fd_sc_hd__a221o_4
X_6280_ _6714_/Q wire640/X wire638/X _6546_/Q _6279_/X VGND VGND VPWR VPWR _6281_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_142_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5231_ wire753/X hold828/X _5233_/S VGND VGND VPWR VPWR _5231_/X sky130_fd_sc_hd__mux2_1
X_5162_ _5164_/A _4636_/A _4664_/X VGND VGND VPWR VPWR _5163_/C sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_12_csclk _6708_/CLK VGND VGND VPWR VPWR _6591_/CLK sky130_fd_sc_hd__clkbuf_8
X_4113_ _5487_/A0 hold786/X _4117_/S VGND VGND VPWR VPWR _6589_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5093_ _5061_/Y _5076_/X _5092_/X _5059_/X VGND VGND VPWR VPWR _6781_/D sky130_fd_sc_hd__a211o_1
XFILLER_111_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4044_ hold748/X _6407_/A0 _4048_/S VGND VGND VPWR VPWR _6530_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_27_csclk _6708_/CLK VGND VGND VPWR VPWR _6981_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5995_ _7168_/Q _7169_/Q VGND VGND VPWR VPWR _6032_/C sky130_fd_sc_hd__and2b_4
XFILLER_178_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4946_ _4946_/A _4946_/B VGND VGND VPWR VPWR _4946_/X sky130_fd_sc_hd__or2_4
XFILLER_52_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4877_ _5147_/A _4877_/B VGND VGND VPWR VPWR _4878_/A sky130_fd_sc_hd__or2_2
XFILLER_20_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6616_ _6626_/CLK _6616_/D fanout874/X VGND VGND VPWR VPWR _6616_/Q sky130_fd_sc_hd__dfstp_2
X_3828_ _3250_/X _3249_/Y _3828_/S VGND VGND VPWR VPWR _3828_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6547_ _6591_/CLK _6547_/D fanout873/X VGND VGND VPWR VPWR _6547_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3759_ _3759_/A _3759_/B _3759_/C _3759_/D VGND VGND VPWR VPWR _3794_/B sky130_fd_sc_hd__or4_2
XFILLER_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6478_ _3957_/A1 _6478_/D _6433_/X VGND VGND VPWR VPWR hold59/A sky130_fd_sc_hd__dfrtp_2
XFILLER_3_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput250 _3938_/X VGND VGND VPWR VPWR mgmt_gpio_out[9] sky130_fd_sc_hd__clkbuf_4
X_5429_ _5519_/A0 hold727/X _5429_/S VGND VGND VPWR VPWR _7002_/D sky130_fd_sc_hd__mux2_1
Xoutput261 _6808_/Q VGND VGND VPWR VPWR pll90_sel[0] sky130_fd_sc_hd__buf_8
XFILLER_121_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput294 _6499_/Q VGND VGND VPWR VPWR pll_trim[3] sky130_fd_sc_hd__buf_8
Xoutput272 _6805_/Q VGND VGND VPWR VPWR pll_sel[0] sky130_fd_sc_hd__buf_8
Xoutput283 _6812_/Q VGND VGND VPWR VPWR pll_trim[17] sky130_fd_sc_hd__buf_8
XFILLER_87_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire355 _3313_/X VGND VGND VPWR VPWR _3331_/B sky130_fd_sc_hd__buf_4
XFILLER_139_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire366 _3711_/X VGND VGND VPWR VPWR wire366/X sky130_fd_sc_hd__buf_6
XFILLER_7_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire377 _5736_/X VGND VGND VPWR VPWR _5741_/A sky130_fd_sc_hd__buf_6
XFILLER_99_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire388 _5218_/A VGND VGND VPWR VPWR wire388/X sky130_fd_sc_hd__buf_8
Xwire399 _3365_/Y VGND VGND VPWR VPWR _5576_/A sky130_fd_sc_hd__buf_8
XFILLER_152_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_1_wb_clk_i clkbuf_1_1_1_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_98_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4800_ _4800_/A _4800_/B _4800_/C _4800_/D VGND VGND VPWR VPWR _4800_/X sky130_fd_sc_hd__or4_1
XFILLER_22_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5780_ _3220_/A _5682_/X _5794_/B1 wire550/X VGND VGND VPWR VPWR _5780_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4731_ _4898_/B _4756_/B _4728_/X _4592_/B _4730_/X VGND VGND VPWR VPWR _4731_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4662_ _4663_/A _4663_/B VGND VGND VPWR VPWR _4758_/C sky130_fd_sc_hd__nor2_8
XFILLER_147_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3613_ wire904/X _3361_/Y wire446/A _7119_/Q VGND VGND VPWR VPWR _3613_/X sky130_fd_sc_hd__a22o_2
X_6401_ _6401_/A1 _4237_/X _5156_/A _3916_/A VGND VGND VPWR VPWR _7219_/D sky130_fd_sc_hd__o211a_2
X_4593_ _4593_/A _4693_/B _5087_/C VGND VGND VPWR VPWR _4593_/Y sky130_fd_sc_hd__nand3_2
XFILLER_162_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3544_ _6492_/Q _3544_/A2 hold64/A _7153_/Q VGND VGND VPWR VPWR _3544_/X sky130_fd_sc_hd__a22o_1
X_6332_ _6533_/Q _6357_/A2 _6321_/X _6331_/X _6308_/S VGND VGND VPWR VPWR _6332_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_142_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3475_ _6881_/Q wire406/X _3739_/B1 _6985_/Q _3474_/X VGND VGND VPWR VPWR _3488_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6263_ _6759_/Q wire589/X _6337_/B1 _6645_/Q _6262_/X VGND VGND VPWR VPWR _6269_/A
+ sky130_fd_sc_hd__a221o_1
X_5214_ _6817_/Q _5547_/A0 _5215_/S VGND VGND VPWR VPWR _6817_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6194_ _6194_/A _6194_/B _6194_/C _6194_/D VGND VGND VPWR VPWR _6207_/B sky130_fd_sc_hd__or4_1
XFILLER_111_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5145_ _5145_/A _5145_/B _5145_/C _5145_/D VGND VGND VPWR VPWR _5146_/B sky130_fd_sc_hd__or4_2
XFILLER_29_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5076_ _5142_/B _5076_/B _5076_/C _5076_/D VGND VGND VPWR VPWR _5076_/X sky130_fd_sc_hd__or4_1
X_4027_ hold38/X hold850/X _4033_/S VGND VGND VPWR VPWR _4027_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5978_ _6580_/Q wire684/X _5967_/X _5977_/X VGND VGND VPWR VPWR _5981_/C sky130_fd_sc_hd__a211o_1
XFILLER_12_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4929_ _4500_/A _4758_/A _4711_/C _4682_/Y VGND VGND VPWR VPWR _4932_/B sky130_fd_sc_hd__a31o_1
XFILLER_165_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _3260_/A _3293_/B _3309_/B VGND VGND VPWR VPWR _3505_/A sky130_fd_sc_hd__or3_4
XFILLER_66_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3191_ _6477_/Q VGND VGND VPWR VPWR _3191_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6950_ _6950_/CLK _6950_/D fanout875/X VGND VGND VPWR VPWR _6950_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5901_ _6564_/Q wire673/X wire653/X _6650_/Q VGND VGND VPWR VPWR _5901_/X sky130_fd_sc_hd__a22o_1
XFILLER_19_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6881_ _7096_/CLK _6881_/D fanout882/X VGND VGND VPWR VPWR _6881_/Q sky130_fd_sc_hd__dfrtp_2
X_5832_ _7083_/Q wire677/X _5694_/X wire542/X _5831_/X VGND VGND VPWR VPWR _5839_/A
+ sky130_fd_sc_hd__a221o_4
XFILLER_62_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5763_ _5763_/A _5763_/B _5763_/C _5763_/D VGND VGND VPWR VPWR _5763_/X sky130_fd_sc_hd__or4_2
X_4714_ _5062_/B _4714_/B VGND VGND VPWR VPWR _5050_/B sky130_fd_sc_hd__or2_2
XFILLER_175_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5694_ _5864_/B _5707_/B _5707_/C VGND VGND VPWR VPWR _5694_/X sky130_fd_sc_hd__and3_4
XFILLER_163_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4645_ _4887_/B _4787_/B _4642_/X _4644_/Y _4567_/X VGND VGND VPWR VPWR _4645_/X
+ sky130_fd_sc_hd__o41a_2
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4576_ _4871_/A _4953_/A VGND VGND VPWR VPWR _4708_/A sky130_fd_sc_hd__nor2_1
XFILLER_146_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold700 _6621_/Q VGND VGND VPWR VPWR hold700/X sky130_fd_sc_hd__bufbuf_16
Xhold711 _6754_/Q VGND VGND VPWR VPWR hold711/X sky130_fd_sc_hd__bufbuf_16
Xhold744 _6927_/Q VGND VGND VPWR VPWR hold744/X sky130_fd_sc_hd__bufbuf_16
Xhold722 _6903_/Q VGND VGND VPWR VPWR hold722/X sky130_fd_sc_hd__bufbuf_16
X_3527_ input48/X _3736_/A2 _5585_/A _7145_/Q wire368/X VGND VGND VPWR VPWR _3533_/B
+ sky130_fd_sc_hd__a221o_4
Xhold755 _6578_/Q VGND VGND VPWR VPWR hold755/X sky130_fd_sc_hd__bufbuf_16
Xhold733 _5232_/X VGND VGND VPWR VPWR _6830_/D sky130_fd_sc_hd__bufbuf_16
X_6315_ _6761_/Q wire589/X _6337_/B1 _6647_/Q _6312_/X VGND VGND VPWR VPWR _6321_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold788 _6995_/Q VGND VGND VPWR VPWR hold788/X sky130_fd_sc_hd__bufbuf_16
Xhold777 _7075_/Q VGND VGND VPWR VPWR hold777/X sky130_fd_sc_hd__bufbuf_16
Xhold766 _7221_/Q VGND VGND VPWR VPWR hold766/X sky130_fd_sc_hd__bufbuf_16
XFILLER_162_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold799 _6723_/Q VGND VGND VPWR VPWR hold799/X sky130_fd_sc_hd__bufbuf_16
X_6246_ _6545_/Q wire638/X wire616/X _6644_/Q _6245_/X VGND VGND VPWR VPWR _6247_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3458_ _7001_/Q wire450/X _4154_/A _6628_/Q _3456_/X VGND VGND VPWR VPWR _3472_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_190_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6177_ _6874_/Q wire593/X wire591/X _6898_/Q _6176_/X VGND VGND VPWR VPWR _6181_/B
+ sky130_fd_sc_hd__a221o_1
X_3389_ input32/X _3283_/Y _5477_/A _7051_/Q VGND VGND VPWR VPWR _3389_/X sky130_fd_sc_hd__a22o_1
X_5128_ _5128_/A _5128_/B _5128_/C _5128_/D VGND VGND VPWR VPWR _5143_/A sky130_fd_sc_hd__or4_4
XFILLER_69_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5059_ _4935_/D _5102_/C _5102_/D _5036_/X _5058_/X VGND VGND VPWR VPWR _5059_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_84_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold82 hold82/A VGND VGND VPWR VPWR hold82/X sky130_fd_sc_hd__bufbuf_16
XFILLER_63_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold71 hold71/A VGND VGND VPWR VPWR hold71/X sky130_fd_sc_hd__bufbuf_16
Xhold60 hold60/A VGND VGND VPWR VPWR hold60/X sky130_fd_sc_hd__bufbuf_16
XFILLER_63_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold93 hold93/A VGND VGND VPWR VPWR hold93/X sky130_fd_sc_hd__bufbuf_16
XFILLER_189_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4430_ _4507_/A _4500_/A _4851_/B _4499_/C VGND VGND VPWR VPWR _5140_/B sky130_fd_sc_hd__and4_2
XANTENNA_2 _6414_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4361_ _4566_/A _4558_/B VGND VGND VPWR VPWR _4502_/A sky130_fd_sc_hd__or2_4
X_6100_ _6951_/Q wire637/X wire635/X _6927_/Q VGND VGND VPWR VPWR _6100_/X sky130_fd_sc_hd__a22o_1
X_7080_ _7152_/CLK _7080_/D fanout883/X VGND VGND VPWR VPWR _7080_/Q sky130_fd_sc_hd__dfrtp_2
X_3312_ input42/X _4023_/S _5549_/A _7116_/Q VGND VGND VPWR VPWR _3312_/X sky130_fd_sc_hd__a22o_1
X_4292_ _4292_/A _5378_/B VGND VGND VPWR VPWR _4297_/S sky130_fd_sc_hd__nand2_8
XFILLER_113_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3243_ _4672_/A VGND VGND VPWR VPWR _4735_/B sky130_fd_sc_hd__inv_4
X_6031_ _6032_/A _6035_/A _6037_/C VGND VGND VPWR VPWR _6031_/X sky130_fd_sc_hd__and3_1
XFILLER_140_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6933_ _7151_/CLK _6933_/D fanout880/X VGND VGND VPWR VPWR _6933_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_82_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6864_ _7096_/CLK _6864_/D fanout883/X VGND VGND VPWR VPWR _6864_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_179_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5815_ _7018_/Q wire697/X wire662/X wire547/X VGND VGND VPWR VPWR _5815_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6795_ _3545_/A1 _6795_/D _6453_/X VGND VGND VPWR VPWR _6795_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_50_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5746_ wire482/X _5675_/X wire664/X _6951_/Q _5745_/X VGND VGND VPWR VPWR _5753_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_50_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5677_ wire483/X _5675_/X wire702/X _6973_/Q VGND VGND VPWR VPWR _5677_/X sky130_fd_sc_hd__a22o_1
XFILLER_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4628_ _4995_/A _4989_/A VGND VGND VPWR VPWR _4628_/Y sky130_fd_sc_hd__nor2_1
Xhold530 _6836_/Q VGND VGND VPWR VPWR hold530/X sky130_fd_sc_hd__bufbuf_16
XFILLER_123_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold563 _4038_/X VGND VGND VPWR VPWR _6525_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_151_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4559_ _4808_/A _5013_/A _4559_/C _4558_/X VGND VGND VPWR VPWR _4559_/X sky130_fd_sc_hd__or4b_1
Xhold541 _6838_/Q VGND VGND VPWR VPWR hold541/X sky130_fd_sc_hd__bufbuf_16
Xhold552 _7037_/Q VGND VGND VPWR VPWR hold552/X sky130_fd_sc_hd__bufbuf_16
Xhold574 _7144_/Q VGND VGND VPWR VPWR hold574/X sky130_fd_sc_hd__bufbuf_16
XFILLER_104_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold585 _4229_/X VGND VGND VPWR VPWR _6685_/D sky130_fd_sc_hd__bufbuf_16
Xhold596 _6823_/Q VGND VGND VPWR VPWR hold596/X sky130_fd_sc_hd__bufbuf_16
X_6229_ _7068_/Q wire648/X wire633/X _6916_/Q VGND VGND VPWR VPWR _6229_/X sky130_fd_sc_hd__a22o_1
XFILLER_58_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput161 wb_dat_i[7] VGND VGND VPWR VPWR _6399_/B1 sky130_fd_sc_hd__clkbuf_4
Xinput150 wb_dat_i[26] VGND VGND VPWR VPWR _6384_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3930_ _6843_/Q input89/X _3932_/S VGND VGND VPWR VPWR _3930_/X sky130_fd_sc_hd__mux2_8
XFILLER_17_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3861_ _6467_/Q _3861_/B VGND VGND VPWR VPWR _3866_/B sky130_fd_sc_hd__nor2_2
XFILLER_176_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5600_ _5600_/A0 hold449/X hold66/X VGND VGND VPWR VPWR _5600_/X sky130_fd_sc_hd__mux2_1
X_6580_ _6650_/CLK _6580_/D fanout858/X VGND VGND VPWR VPWR _6580_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3792_ _3792_/A _3792_/B _3792_/C _3792_/D VGND VGND VPWR VPWR _3793_/D sky130_fd_sc_hd__or4_1
XFILLER_31_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5531_ _5531_/A _5576_/B VGND VGND VPWR VPWR _5538_/S sky130_fd_sc_hd__nand2_4
XFILLER_117_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5462_ wire786/X hold359/X _5467_/S VGND VGND VPWR VPWR _7031_/D sky130_fd_sc_hd__mux2_1
X_7201_ _7220_/CLK _7201_/D fanout853/X VGND VGND VPWR VPWR _7201_/Q sky130_fd_sc_hd__dfrtp_2
X_4413_ _4672_/A _4696_/A _4413_/C _4436_/B VGND VGND VPWR VPWR _4414_/B sky130_fd_sc_hd__and4_4
X_5393_ wire758/X hold282/X _5395_/S VGND VGND VPWR VPWR _6970_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4344_ _4408_/B _4408_/A VGND VGND VPWR VPWR _4553_/A sky130_fd_sc_hd__nand2b_4
XFILLER_113_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7132_ _7132_/CLK _7132_/D fanout868/X VGND VGND VPWR VPWR _7132_/Q sky130_fd_sc_hd__dfrtp_2
X_7063_ _7145_/CLK _7063_/D fanout883/X VGND VGND VPWR VPWR _7063_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_140_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6014_ _6014_/A _6034_/B VGND VGND VPWR VPWR _6014_/Y sky130_fd_sc_hd__nor2_8
X_4275_ _6407_/A0 hold778/X _4279_/S VGND VGND VPWR VPWR _6728_/D sky130_fd_sc_hd__mux2_1
X_3226_ _6968_/Q VGND VGND VPWR VPWR _3226_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6916_ _6980_/CLK _6916_/D fanout880/X VGND VGND VPWR VPWR _6916_/Q sky130_fd_sc_hd__dfrtp_2
X_6847_ _6992_/CLK _6847_/D fanout868/X VGND VGND VPWR VPWR _6847_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire707 _5673_/X VGND VGND VPWR VPWR wire707/X sky130_fd_sc_hd__buf_8
X_6778_ _7190_/CLK _6778_/D _6362_/B VGND VGND VPWR VPWR hold93/A sky130_fd_sc_hd__dfrtp_2
XFILLER_22_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire718 _6376_/A VGND VGND VPWR VPWR _5156_/A sky130_fd_sc_hd__buf_8
XFILLER_167_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5729_ _6958_/Q wire707/X _5681_/X _6918_/Q _5728_/X VGND VGND VPWR VPWR _5734_/B
+ sky130_fd_sc_hd__a221o_4
Xwire729 wire729/A VGND VGND VPWR VPWR wire729/X sky130_fd_sc_hd__buf_8
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold371 _6980_/Q VGND VGND VPWR VPWR hold371/X sky130_fd_sc_hd__bufbuf_16
XFILLER_123_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold360 _7071_/Q VGND VGND VPWR VPWR hold360/X sky130_fd_sc_hd__bufbuf_16
Xhold382 _6924_/Q VGND VGND VPWR VPWR hold382/X sky130_fd_sc_hd__bufbuf_16
Xhold393 _5566_/X VGND VGND VPWR VPWR _7124_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_131_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout851 _6447_/A VGND VGND VPWR VPWR fanout851/X sky130_fd_sc_hd__buf_8
Xfanout884 fanout889/X VGND VGND VPWR VPWR fanout884/X sky130_fd_sc_hd__buf_8
Xfanout873 fanout890/X VGND VGND VPWR VPWR fanout873/X sky130_fd_sc_hd__buf_8
XFILLER_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout862 fanout868/A VGND VGND VPWR VPWR fanout862/X sky130_fd_sc_hd__buf_8
XFILLER_100_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_200 wire485/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_222 wire591/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_233 wire672/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_211 wire519/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_244 _5600_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_277 hold465/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_266 hold150/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_255 _3969_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_299 _5685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_288 hold808/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4060_ _4303_/A0 hold405/X _4060_/S VGND VGND VPWR VPWR _6544_/D sky130_fd_sc_hd__mux2_1
XFILLER_49_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4962_ _4962_/A _4962_/B VGND VGND VPWR VPWR _4971_/B sky130_fd_sc_hd__or2_2
XFILLER_91_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4893_ _4893_/A _4893_/B VGND VGND VPWR VPWR _4906_/B sky130_fd_sc_hd__nand2_1
X_3913_ _6705_/Q _3883_/X _6700_/Q VGND VGND VPWR VPWR _6705_/D sky130_fd_sc_hd__a21o_1
X_6701_ _7208_/CLK _6701_/D _6362_/B VGND VGND VPWR VPWR _6701_/Q sky130_fd_sc_hd__dfrtp_2
X_6632_ _6632_/CLK _6632_/D fanout872/X VGND VGND VPWR VPWR _6632_/Q sky130_fd_sc_hd__dfstp_2
X_3844_ _6457_/Q _6476_/Q _3924_/C VGND VGND VPWR VPWR _6476_/D sky130_fd_sc_hd__mux2_1
XFILLER_177_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6563_ _6591_/CLK _6563_/D fanout873/X VGND VGND VPWR VPWR _6563_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_118_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3775_ _7069_/Q _5504_/A _4190_/A _6654_/Q _3774_/X VGND VGND VPWR VPWR _3775_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_157_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6494_ _6815_/CLK _6494_/D fanout855/X VGND VGND VPWR VPWR _6494_/Q sky130_fd_sc_hd__dfstp_4
X_5514_ wire802/X _7077_/Q _5521_/S VGND VGND VPWR VPWR _7077_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5445_ wire769/X hold600/X _5449_/S VGND VGND VPWR VPWR _7016_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7115_ _7155_/CLK _7115_/D fanout884/X VGND VGND VPWR VPWR _7115_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_154_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5376_ hold57/X hold273/X _5377_/S VGND VGND VPWR VPWR _6955_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4327_ _6411_/A0 hold650/X _4327_/S VGND VGND VPWR VPWR _6772_/D sky130_fd_sc_hd__mux2_1
X_4258_ hold440/X wire794/A _4261_/S VGND VGND VPWR VPWR _6714_/D sky130_fd_sc_hd__mux2_1
X_7046_ _7134_/CLK _7046_/D fanout864/X VGND VGND VPWR VPWR _7046_/Q sky130_fd_sc_hd__dfstp_4
X_3209_ _3209_/A VGND VGND VPWR VPWR _3209_/Y sky130_fd_sc_hd__inv_2
X_4189_ hold398/X _4303_/A0 _4189_/S VGND VGND VPWR VPWR _6653_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire504 _7050_/Q VGND VGND VPWR VPWR wire504/X sky130_fd_sc_hd__buf_6
Xwire515 _7023_/Q VGND VGND VPWR VPWR wire515/X sky130_fd_sc_hd__buf_6
Xwire548 _6873_/Q VGND VGND VPWR VPWR wire548/X sky130_fd_sc_hd__buf_6
XFILLER_155_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire526 _6979_/Q VGND VGND VPWR VPWR wire526/X sky130_fd_sc_hd__buf_6
Xwire537 _6912_/Q VGND VGND VPWR VPWR _3233_/A sky130_fd_sc_hd__buf_6
XFILLER_11_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire559 wire559/A VGND VGND VPWR VPWR wire559/X sky130_fd_sc_hd__clkbuf_8
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold190 hold333/X VGND VGND VPWR VPWR _3293_/B sky130_fd_sc_hd__bufbuf_16
XFILLER_65_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_8_csclk _6744_/CLK VGND VGND VPWR VPWR _6633_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_61_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3560_ _7008_/Q _5432_/A _3368_/Y input14/X VGND VGND VPWR VPWR _3560_/X sky130_fd_sc_hd__a22o_4
XFILLER_155_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3491_ _3508_/A _3732_/B VGND VGND VPWR VPWR _5185_/A sky130_fd_sc_hd__nor2_8
X_5230_ _5255_/A0 hold769/X _5233_/S VGND VGND VPWR VPWR _6828_/D sky130_fd_sc_hd__mux2_1
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5161_ _4940_/B _5101_/C _5161_/C _5161_/D VGND VGND VPWR VPWR _5161_/X sky130_fd_sc_hd__and4bb_1
XFILLER_96_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4112_ _4112_/A _5236_/B VGND VGND VPWR VPWR _4117_/S sky130_fd_sc_hd__nand2_8
X_5092_ _5083_/X _5091_/X _5077_/Y VGND VGND VPWR VPWR _5092_/X sky130_fd_sc_hd__o21a_1
XFILLER_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4043_ _4043_/A _6406_/B VGND VGND VPWR VPWR _4048_/S sky130_fd_sc_hd__and2_4
XFILLER_83_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5994_ _6030_/A _6014_/A VGND VGND VPWR VPWR _6021_/A sky130_fd_sc_hd__nor2_8
XFILLER_64_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4945_ _5095_/B _5022_/D _5180_/B _4945_/D VGND VGND VPWR VPWR _4946_/B sky130_fd_sc_hd__or4_1
XFILLER_52_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4876_ _4617_/B _4970_/B _4898_/B _5147_/B VGND VGND VPWR VPWR _4877_/B sky130_fd_sc_hd__o22a_1
XFILLER_178_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6615_ _6712_/CLK _6615_/D fanout872/X VGND VGND VPWR VPWR _6615_/Q sky130_fd_sc_hd__dfrtp_2
X_3827_ _3845_/A _3830_/B VGND VGND VPWR VPWR _3827_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3758_ _6957_/Q _5378_/A _4256_/A _6713_/Q _3740_/X VGND VGND VPWR VPWR _3759_/D
+ sky130_fd_sc_hd__a221o_4
XFILLER_137_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6546_ _6591_/CLK _6546_/D fanout873/X VGND VGND VPWR VPWR _6546_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_118_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3689_ _6625_/Q _4154_/A _4250_/A _6709_/Q VGND VGND VPWR VPWR _3689_/X sky130_fd_sc_hd__a22o_4
X_6477_ _6668_/CLK _6477_/D _6432_/X VGND VGND VPWR VPWR _6477_/Q sky130_fd_sc_hd__dfrtp_2
Xoutput240 _6841_/Q VGND VGND VPWR VPWR mgmt_gpio_out[34] sky130_fd_sc_hd__buf_8
XFILLER_133_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5428_ wire763/X hold423/X _5431_/S VGND VGND VPWR VPWR _7001_/D sky130_fd_sc_hd__mux2_1
Xoutput262 _6809_/Q VGND VGND VPWR VPWR pll90_sel[1] sky130_fd_sc_hd__buf_8
Xoutput251 _3957_/X VGND VGND VPWR VPWR pad_flash_clk sky130_fd_sc_hd__clkbuf_4
X_5359_ _5602_/A0 hold363/X _5359_/S VGND VGND VPWR VPWR _5359_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput273 _6806_/Q VGND VGND VPWR VPWR pll_sel[1] sky130_fd_sc_hd__buf_8
Xoutput284 _6813_/Q VGND VGND VPWR VPWR pll_trim[18] sky130_fd_sc_hd__buf_8
Xoutput295 _6500_/Q VGND VGND VPWR VPWR pll_trim[4] sky130_fd_sc_hd__buf_8
XFILLER_181_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7029_ _7105_/CLK _7029_/D fanout862/X VGND VGND VPWR VPWR _7029_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_55_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire356 _5580_/S VGND VGND VPWR VPWR _5581_/S sky130_fd_sc_hd__buf_6
XFILLER_183_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire367 _3674_/X VGND VGND VPWR VPWR wire367/X sky130_fd_sc_hd__buf_6
Xwire389 _3543_/Y VGND VGND VPWR VPWR _4055_/A sky130_fd_sc_hd__buf_8
XFILLER_124_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4730_ _4740_/B _5017_/A _4729_/X VGND VGND VPWR VPWR _4730_/X sky130_fd_sc_hd__o21ba_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4661_ _4745_/A _4697_/A VGND VGND VPWR VPWR _4933_/B sky130_fd_sc_hd__nand2_2
XFILLER_9_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6400_ _6399_/X _7218_/Q _6400_/S VGND VGND VPWR VPWR _7218_/D sky130_fd_sc_hd__mux2_1
X_3612_ _6552_/Q _3473_/Y _4055_/A _6542_/Q VGND VGND VPWR VPWR _3612_/X sky130_fd_sc_hd__a22o_1
XFILLER_128_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4592_ _4812_/A _4592_/B VGND VGND VPWR VPWR _5087_/C sky130_fd_sc_hd__nor2_4
XFILLER_128_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6331_ _6356_/A _6331_/B _6331_/C _6331_/D VGND VGND VPWR VPWR _6331_/X sky130_fd_sc_hd__or4_1
XFILLER_143_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3543_ _3543_/A _3543_/B VGND VGND VPWR VPWR _3543_/Y sky130_fd_sc_hd__nor2_4
XFILLER_142_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3474_ _6921_/Q _3582_/A2 _3473_/Y _6554_/Q VGND VGND VPWR VPWR _3474_/X sky130_fd_sc_hd__a22o_1
X_6262_ _6734_/Q wire642/X wire630/X wire561/X VGND VGND VPWR VPWR _6262_/X sky130_fd_sc_hd__a22o_1
X_6193_ _6987_/Q _6028_/X _6034_/Y _6995_/Q _6192_/X VGND VGND VPWR VPWR _6194_/D
+ sky130_fd_sc_hd__a221o_4
X_5213_ _6816_/Q wire753/X _5215_/S VGND VGND VPWR VPWR _6816_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5144_ _5144_/A _5144_/B VGND VGND VPWR VPWR _5145_/D sky130_fd_sc_hd__nand2_1
XFILLER_111_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5075_ _5075_/A _5075_/B _5075_/C _5075_/D VGND VGND VPWR VPWR _5076_/D sky130_fd_sc_hd__or4_1
X_4026_ _5595_/A0 hold749/X _4033_/S VGND VGND VPWR VPWR _6514_/D sky130_fd_sc_hd__mux2_1
XFILLER_65_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5977_ _6593_/Q _5977_/A2 wire667/X _6539_/Q _5964_/X VGND VGND VPWR VPWR _5977_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_52_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4928_ _4932_/A VGND VGND VPWR VPWR _4928_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4859_ _4624_/B _4845_/B _4858_/X _5114_/A _5114_/B VGND VGND VPWR VPWR _4859_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_60_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6529_ _7152_/CLK _6529_/D fanout882/X VGND VGND VPWR VPWR _6529_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_73_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6646_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_28_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_26_csclk _6708_/CLK VGND VGND VPWR VPWR _6833_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_124_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5900_ _6739_/Q wire700/X wire679/X _7222_/Q _5898_/X VGND VGND VPWR VPWR _5915_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_179_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6880_ _6980_/CLK _6880_/D fanout880/X VGND VGND VPWR VPWR _6880_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_81_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5831_ _7107_/Q _5857_/A2 wire689/X _7051_/Q VGND VGND VPWR VPWR _5831_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5762_ _6911_/Q _5680_/X _5687_/X wire507/X _5761_/X VGND VGND VPWR VPWR _5763_/D
+ sky130_fd_sc_hd__a221o_1
X_4713_ _4713_/A _4713_/B _4713_/C _4713_/D VGND VGND VPWR VPWR _4713_/X sky130_fd_sc_hd__or4_1
XFILLER_148_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5693_ _7165_/Q _5702_/B _5701_/C VGND VGND VPWR VPWR _5693_/X sky130_fd_sc_hd__and3_4
XFILLER_163_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4644_ _4917_/A _4897_/B VGND VGND VPWR VPWR _4644_/Y sky130_fd_sc_hd__nand2_1
X_4575_ _4987_/A _4575_/B VGND VGND VPWR VPWR _4575_/Y sky130_fd_sc_hd__nand2_2
Xhold712 _6764_/Q VGND VGND VPWR VPWR hold712/X sky130_fd_sc_hd__bufbuf_16
Xhold701 _6531_/Q VGND VGND VPWR VPWR hold701/X sky130_fd_sc_hd__bufbuf_16
Xhold723 _6552_/Q VGND VGND VPWR VPWR hold723/X sky130_fd_sc_hd__bufbuf_16
XFILLER_116_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6314_ _6716_/Q wire640/X wire632/X _6592_/Q VGND VGND VPWR VPWR _6330_/B sky130_fd_sc_hd__a22o_1
X_3526_ _6815_/Q _5207_/A _3995_/A _6500_/Q VGND VGND VPWR VPWR _3526_/X sky130_fd_sc_hd__a22o_4
Xhold734 _6681_/Q VGND VGND VPWR VPWR hold734/X sky130_fd_sc_hd__bufbuf_16
Xhold745 _6640_/Q VGND VGND VPWR VPWR hold745/X sky130_fd_sc_hd__bufbuf_16
Xhold767 _6609_/Q VGND VGND VPWR VPWR hold767/X sky130_fd_sc_hd__bufbuf_16
XFILLER_143_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold778 _6728_/Q VGND VGND VPWR VPWR hold778/X sky130_fd_sc_hd__bufbuf_16
Xhold756 _6683_/Q VGND VGND VPWR VPWR hold756/X sky130_fd_sc_hd__bufbuf_16
X_6245_ _6763_/Q wire649/X _6335_/B _6773_/Q VGND VGND VPWR VPWR _6245_/X sky130_fd_sc_hd__a22o_4
Xhold789 _6743_/Q VGND VGND VPWR VPWR hold789/X sky130_fd_sc_hd__bufbuf_16
XFILLER_115_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3457_ _3540_/A _5252_/B VGND VGND VPWR VPWR _4154_/A sky130_fd_sc_hd__nor2_8
X_6176_ _6962_/Q wire624/X wire613/X _7058_/Q VGND VGND VPWR VPWR _6176_/X sky130_fd_sc_hd__a22o_1
XFILLER_162_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3388_ wire470/X _3714_/A2 _4234_/S input69/X VGND VGND VPWR VPWR _3388_/X sky130_fd_sc_hd__a22o_1
X_5127_ _5127_/A VGND VGND VPWR VPWR _5146_/A sky130_fd_sc_hd__inv_2
XFILLER_84_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5058_ _6781_/Q _5156_/A _5038_/Y _5057_/X VGND VGND VPWR VPWR _5058_/X sky130_fd_sc_hd__a22o_1
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4009_ hold665/X _5595_/A0 _4021_/S VGND VGND VPWR VPWR _4009_/X sky130_fd_sc_hd__mux2_1
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold50 hold50/A VGND VGND VPWR VPWR hold50/X sky130_fd_sc_hd__bufbuf_16
XFILLER_121_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold83 hold83/A VGND VGND VPWR VPWR hold83/X sky130_fd_sc_hd__bufbuf_16
XFILLER_152_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold72 hold72/A VGND VGND VPWR VPWR hold72/X sky130_fd_sc_hd__bufbuf_16
Xhold61 hold61/A VGND VGND VPWR VPWR hold61/X sky130_fd_sc_hd__bufbuf_16
Xhold94 hold94/A VGND VGND VPWR VPWR hold94/X sky130_fd_sc_hd__bufbuf_16
XFILLER_90_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_2_0_mgmt_gpio_in[4] clkbuf_2_3_0_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR _3545_/A1
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_3 _6424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4360_ _4566_/A _4558_/B VGND VGND VPWR VPWR _4581_/A sky130_fd_sc_hd__nor2_8
X_3311_ _3508_/A hold96/X VGND VGND VPWR VPWR hold97/A sky130_fd_sc_hd__nor2_8
XFILLER_140_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4291_ _6411_/A0 hold555/X _4291_/S VGND VGND VPWR VPWR _4291_/X sky130_fd_sc_hd__mux2_1
X_3242_ _4735_/A VGND VGND VPWR VPWR _4564_/A sky130_fd_sc_hd__clkinv_4
X_6030_ _6030_/A _6036_/A VGND VGND VPWR VPWR _6030_/Y sky130_fd_sc_hd__nor2_8
XFILLER_39_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6932_ _7155_/CLK _6932_/D fanout884/X VGND VGND VPWR VPWR _6932_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_82_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6863_ _7145_/CLK _6863_/D fanout881/X VGND VGND VPWR VPWR _6863_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5814_ _6906_/Q _5814_/A2 _5812_/X _5813_/X VGND VGND VPWR VPWR _5814_/X sky130_fd_sc_hd__a211o_1
XFILLER_22_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6794_ _3545_/A1 _6794_/D _6452_/X VGND VGND VPWR VPWR _6794_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_50_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5745_ _6975_/Q wire702/X _5931_/A2 _6871_/Q VGND VGND VPWR VPWR _5745_/X sky130_fd_sc_hd__a22o_1
XFILLER_163_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5676_ _5864_/B _5705_/B _5701_/C VGND VGND VPWR VPWR _5676_/X sky130_fd_sc_hd__and3_4
XFILLER_135_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4627_ _4986_/C _4990_/A _4623_/X _4624_/Y _4626_/Y VGND VGND VPWR VPWR _4627_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_151_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold520 _7025_/Q VGND VGND VPWR VPWR hold520/X sky130_fd_sc_hd__bufbuf_16
XFILLER_190_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4558_ _4819_/A _4558_/B _4844_/B VGND VGND VPWR VPWR _4558_/X sky130_fd_sc_hd__or3_2
XFILLER_104_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold542 _5244_/X VGND VGND VPWR VPWR _6838_/D sky130_fd_sc_hd__bufbuf_16
Xhold553 _6780_/Q VGND VGND VPWR VPWR hold99/A sky130_fd_sc_hd__bufbuf_16
Xhold531 _6994_/Q VGND VGND VPWR VPWR hold531/X sky130_fd_sc_hd__bufbuf_16
Xhold575 _7080_/Q VGND VGND VPWR VPWR hold575/X sky130_fd_sc_hd__bufbuf_16
Xhold564 _6872_/Q VGND VGND VPWR VPWR hold564/X sky130_fd_sc_hd__bufbuf_16
X_4489_ _4651_/B _4746_/A VGND VGND VPWR VPWR _4659_/A sky130_fd_sc_hd__nor2_8
XFILLER_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold586 _6649_/Q VGND VGND VPWR VPWR hold586/X sky130_fd_sc_hd__bufbuf_16
Xhold597 _6658_/Q VGND VGND VPWR VPWR hold597/X sky130_fd_sc_hd__bufbuf_16
X_3509_ _6826_/Q _3384_/Y _4304_/A _6757_/Q _3507_/X VGND VGND VPWR VPWR _3522_/A
+ sky130_fd_sc_hd__a221o_4
XFILLER_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6228_ wire552/X _6014_/Y wire618/A _7052_/Q _6227_/X VGND VGND VPWR VPWR _6231_/C
+ sky130_fd_sc_hd__a221o_4
XFILLER_66_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ _5611_/A _7192_/Q _5664_/X _6158_/X VGND VGND VPWR VPWR _6159_/X sky130_fd_sc_hd__a211o_2
XFILLER_66_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput140 wb_dat_i[17] VGND VGND VPWR VPWR _6381_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput162 wb_dat_i[8] VGND VGND VPWR VPWR _6377_/B1 sky130_fd_sc_hd__clkbuf_4
Xinput151 wb_dat_i[27] VGND VGND VPWR VPWR _6386_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_95_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3860_ _3898_/A _3810_/B _3859_/Y _3858_/Y VGND VGND VPWR VPWR _3861_/B sky130_fd_sc_hd__o31a_2
XFILLER_176_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3791_ _7021_/Q _3301_/Y _3735_/Y _6825_/Q _3743_/X VGND VGND VPWR VPWR _3792_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5530_ wire739/X hold689/X _5530_/S VGND VGND VPWR VPWR _7092_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5461_ _5578_/A0 _7030_/Q _5467_/S VGND VGND VPWR VPWR _7030_/D sky130_fd_sc_hd__mux2_1
XFILLER_184_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4412_ _4671_/A _4997_/A VGND VGND VPWR VPWR _4412_/Y sky130_fd_sc_hd__nor2_2
XFILLER_117_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7200_ _7220_/CLK _7200_/D fanout854/X VGND VGND VPWR VPWR _7200_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_172_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5392_ hold150/X hold272/X _5395_/S VGND VGND VPWR VPWR _6969_/D sky130_fd_sc_hd__mux2_1
X_7131_ _7147_/CLK _7131_/D fanout888/X VGND VGND VPWR VPWR _7131_/Q sky130_fd_sc_hd__dfrtp_2
X_4343_ _4340_/B _4690_/A _4341_/X VGND VGND VPWR VPWR _4408_/B sky130_fd_sc_hd__o21ai_4
XFILLER_125_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7062_ _7111_/CLK _7062_/D fanout881/X VGND VGND VPWR VPWR _7062_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_113_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4274_ _4274_/A _5242_/B VGND VGND VPWR VPWR _4279_/S sky130_fd_sc_hd__nand2_4
X_3225_ _6976_/Q VGND VGND VPWR VPWR _3225_/Y sky130_fd_sc_hd__inv_2
X_6013_ _6032_/A _6033_/C VGND VGND VPWR VPWR _6034_/B sky130_fd_sc_hd__nand2_8
XFILLER_100_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6915_ _6930_/CLK _6915_/D fanout885/X VGND VGND VPWR VPWR _6915_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_82_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6846_ _7223_/CLK _6846_/D _6455_/A VGND VGND VPWR VPWR _6846_/Q sky130_fd_sc_hd__dfrtp_1
X_6777_ _7225_/CLK _6777_/D fanout850/X VGND VGND VPWR VPWR _6777_/Q sky130_fd_sc_hd__dfrtp_2
X_3989_ hold1/X hold23/X _3991_/S VGND VGND VPWR VPWR hold24/A sky130_fd_sc_hd__mux2_2
XFILLER_176_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5728_ wire529/X wire680/X wire665/X _6950_/Q VGND VGND VPWR VPWR _5728_/X sky130_fd_sc_hd__a22o_2
Xwire719 hold71/X VGND VGND VPWR VPWR hold72/A sky130_fd_sc_hd__buf_6
XFILLER_10_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5659_ _7159_/Q _7160_/Q _5659_/C _7157_/Q VGND VGND VPWR VPWR _5659_/X sky130_fd_sc_hd__or4b_1
XFILLER_184_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold350 _6507_/Q VGND VGND VPWR VPWR hold350/X sky130_fd_sc_hd__bufbuf_16
XFILLER_123_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold361 _6821_/Q VGND VGND VPWR VPWR hold361/X sky130_fd_sc_hd__bufbuf_16
Xhold372 _5404_/X VGND VGND VPWR VPWR _6980_/D sky130_fd_sc_hd__bufbuf_16
Xhold383 _5341_/X VGND VGND VPWR VPWR _6924_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_77_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold394 _7126_/Q VGND VGND VPWR VPWR hold394/X sky130_fd_sc_hd__bufbuf_16
XFILLER_131_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout830 _3877_/Y VGND VGND VPWR VPWR _5252_/C sky130_fd_sc_hd__buf_8
Xfanout852 wire860/A VGND VGND VPWR VPWR _6447_/A sky130_fd_sc_hd__buf_8
Xfanout885 fanout889/X VGND VGND VPWR VPWR fanout885/X sky130_fd_sc_hd__buf_8
Xfanout874 fanout875/X VGND VGND VPWR VPWR fanout874/X sky130_fd_sc_hd__buf_8
XFILLER_58_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout863 fanout864/X VGND VGND VPWR VPWR fanout863/X sky130_fd_sc_hd__buf_8
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_234 wire674/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_223 wire593/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_201 wire492/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_212 wire522/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_256 _7229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_267 hold214/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_245 _4303_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_289 hold848/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_278 hold465/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__1132_ clkbuf_0__1132_/X VGND VGND VPWR VPWR _4108_/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_5_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4961_ _4749_/C _5005_/C _4875_/A VGND VGND VPWR VPWR _4962_/B sky130_fd_sc_hd__a21oi_1
X_4892_ _5005_/C _4756_/B _4623_/D VGND VGND VPWR VPWR _5071_/C sky130_fd_sc_hd__o21ai_2
X_6700_ _7208_/CLK _6700_/D _6362_/B VGND VGND VPWR VPWR _6700_/Q sky130_fd_sc_hd__dfrtp_2
X_3912_ _3905_/X _3909_/Y _3918_/B _6680_/Q VGND VGND VPWR VPWR _6680_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_51_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6631_ _6833_/CLK _6631_/D fanout872/X VGND VGND VPWR VPWR _6631_/Q sky130_fd_sc_hd__dfrtp_2
X_3843_ _6664_/Q _3843_/B VGND VGND VPWR VPWR _3924_/C sky130_fd_sc_hd__nand2_1
XFILLER_32_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6562_ _7210_/CLK _6562_/D VGND VGND VPWR VPWR _6562_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_9_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3774_ _6535_/Q _4049_/A _3551_/Y wire833/X VGND VGND VPWR VPWR _3774_/X sky130_fd_sc_hd__a22o_1
XFILLER_192_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6493_ _6815_/CLK _6493_/D fanout855/X VGND VGND VPWR VPWR _6493_/Q sky130_fd_sc_hd__dfstp_4
X_5513_ _5513_/A _5576_/B VGND VGND VPWR VPWR _5521_/S sky130_fd_sc_hd__nand2_8
XFILLER_160_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5444_ wire780/X hold661/X _5449_/S VGND VGND VPWR VPWR _7015_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7114_ _7155_/CLK _7114_/D fanout884/X VGND VGND VPWR VPWR _7114_/Q sky130_fd_sc_hd__dfrtp_2
X_5375_ _5600_/A0 hold509/X _5377_/S VGND VGND VPWR VPWR _6954_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4326_ _6410_/A0 hold688/X _4327_/S VGND VGND VPWR VPWR _6771_/D sky130_fd_sc_hd__mux2_1
X_4257_ hold770/X _5487_/A0 _4261_/S VGND VGND VPWR VPWR _6713_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7045_ _7134_/CLK _7045_/D fanout861/X VGND VGND VPWR VPWR _7045_/Q sky130_fd_sc_hd__dfstp_4
X_3208_ _7112_/Q VGND VGND VPWR VPWR _3208_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4188_ hold473/X _5249_/A0 _4189_/S VGND VGND VPWR VPWR _6652_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6829_ _7107_/CLK _6829_/D fanout866/X VGND VGND VPWR VPWR _6829_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire505 _7049_/Q VGND VGND VPWR VPWR wire505/X sky130_fd_sc_hd__buf_6
XFILLER_183_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire527 _6978_/Q VGND VGND VPWR VPWR wire527/X sky130_fd_sc_hd__buf_6
XFILLER_149_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire549 _6872_/Q VGND VGND VPWR VPWR _3237_/A sky130_fd_sc_hd__buf_6
Xwire538 _6906_/Q VGND VGND VPWR VPWR wire538/X sky130_fd_sc_hd__buf_6
Xwire516 _7016_/Q VGND VGND VPWR VPWR _3220_/A sky130_fd_sc_hd__buf_8
XFILLER_183_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold180 _5536_/X VGND VGND VPWR VPWR _7097_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold191 _3278_/X VGND VGND VPWR VPWR _3314_/B sky130_fd_sc_hd__bufbuf_16
XFILLER_120_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3490_ _7228_/A _5245_/A _4136_/A _6613_/Q VGND VGND VPWR VPWR _3490_/X sky130_fd_sc_hd__a22o_4
XFILLER_115_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length681 _5690_/X VGND VGND VPWR VPWR _5926_/A2 sky130_fd_sc_hd__buf_6
X_5160_ _4414_/B _4711_/C _4802_/A _5159_/X VGND VGND VPWR VPWR _5161_/D sky130_fd_sc_hd__a211oi_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5091_ _5135_/B _5119_/B _5091_/C VGND VGND VPWR VPWR _5091_/X sky130_fd_sc_hd__or3_1
X_4111_ _6588_/Q wire353/X _4111_/S VGND VGND VPWR VPWR _6588_/D sky130_fd_sc_hd__mux2_1
X_4042_ _5602_/A0 hold278/X hold73/X VGND VGND VPWR VPWR _4042_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5993_ _6019_/A _6033_/C _6035_/C VGND VGND VPWR VPWR _6027_/B sky130_fd_sc_hd__and3b_4
XFILLER_64_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4944_ _4772_/A _4624_/B _5114_/A _4943_/Y VGND VGND VPWR VPWR _4945_/D sky130_fd_sc_hd__a211o_1
X_4875_ _4875_/A _4899_/B VGND VGND VPWR VPWR _4936_/C sky130_fd_sc_hd__nor2_8
XFILLER_60_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6614_ _6626_/CLK _6614_/D fanout874/X VGND VGND VPWR VPWR _6614_/Q sky130_fd_sc_hd__dfrtp_2
X_3826_ _3826_/A _3826_/B VGND VGND VPWR VPWR _6482_/D sky130_fd_sc_hd__xor2_1
XFILLER_165_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3757_ _6733_/Q _4280_/A _5236_/A _6833_/Q _3742_/X VGND VGND VPWR VPWR _3759_/C
+ sky130_fd_sc_hd__a221o_1
X_6545_ _6621_/CLK _6545_/D fanout872/X VGND VGND VPWR VPWR _6545_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3688_ _6942_/Q wire401/X _4268_/A _6724_/Q _3670_/X VGND VGND VPWR VPWR _3693_/A
+ sky130_fd_sc_hd__a221o_1
X_6476_ _3957_/A1 _6476_/D _6431_/X VGND VGND VPWR VPWR _6476_/Q sky130_fd_sc_hd__dfrtp_2
Xoutput230 _6515_/Q VGND VGND VPWR VPWR mgmt_gpio_out[25] sky130_fd_sc_hd__buf_8
Xoutput241 wire460/X VGND VGND VPWR VPWR mgmt_gpio_out[35] sky130_fd_sc_hd__buf_8
X_5427_ _5598_/A0 wire522/A _5431_/S VGND VGND VPWR VPWR _7000_/D sky130_fd_sc_hd__mux2_1
Xoutput252 _3958_/Y VGND VGND VPWR VPWR pad_flash_clk_oeb sky130_fd_sc_hd__buf_8
XFILLER_160_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5358_ _5601_/A0 hold203/X _5359_/S VGND VGND VPWR VPWR _5358_/X sky130_fd_sc_hd__mux2_1
Xoutput263 _6810_/Q VGND VGND VPWR VPWR pll90_sel[2] sky130_fd_sc_hd__buf_8
Xoutput285 _6814_/Q VGND VGND VPWR VPWR pll_trim[19] sky130_fd_sc_hd__buf_8
Xoutput274 _6807_/Q VGND VGND VPWR VPWR pll_sel[2] sky130_fd_sc_hd__buf_8
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput296 _6501_/Q VGND VGND VPWR VPWR pll_trim[5] sky130_fd_sc_hd__buf_8
X_4309_ hold670/X _6411_/A0 _4309_/S VGND VGND VPWR VPWR _6757_/D sky130_fd_sc_hd__mux2_1
X_5289_ _5595_/A0 _6877_/Q _5296_/S VGND VGND VPWR VPWR _6877_/D sky130_fd_sc_hd__mux2_1
XFILLER_75_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7028_ _7095_/CLK _7028_/D fanout865/X VGND VGND VPWR VPWR _7028_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_74_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire379 _6110_/S VGND VGND VPWR VPWR _6309_/S sky130_fd_sc_hd__buf_8
Xwire368 _3526_/X VGND VGND VPWR VPWR wire368/X sky130_fd_sc_hd__buf_6
XFILLER_136_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4660_ _4745_/A _4697_/A VGND VGND VPWR VPWR _4660_/X sky130_fd_sc_hd__and2_4
XFILLER_30_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3611_ input37/X _3310_/Y _4118_/A wire571/X VGND VGND VPWR VPWR _3611_/X sky130_fd_sc_hd__a22o_2
XFILLER_155_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6330_ _6330_/A _6330_/B _6330_/C _6330_/D VGND VGND VPWR VPWR _6331_/D sky130_fd_sc_hd__or4_4
X_4591_ _4898_/B _4591_/B VGND VGND VPWR VPWR _4591_/X sky130_fd_sc_hd__or2_1
X_3542_ _7025_/Q _3301_/Y _3325_/Y _6913_/Q _3541_/X VGND VGND VPWR VPWR _3546_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3473_ _3543_/A _3528_/B VGND VGND VPWR VPWR _3473_/Y sky130_fd_sc_hd__nor2_8
X_6261_ _6655_/Q _6311_/B VGND VGND VPWR VPWR _6261_/X sky130_fd_sc_hd__and2_1
XFILLER_143_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6192_ _7075_/Q _6009_/X _6012_/X _6971_/Q VGND VGND VPWR VPWR _6192_/X sky130_fd_sc_hd__a22o_1
X_5212_ hold659/X _6411_/A0 _5215_/S VGND VGND VPWR VPWR _6815_/D sky130_fd_sc_hd__mux2_1
XFILLER_123_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5143_ _5143_/A _5143_/B _5143_/C VGND VGND VPWR VPWR _5143_/Y sky130_fd_sc_hd__nor3_2
XFILLER_111_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5074_ _5074_/A _5126_/A _5175_/A _5145_/C VGND VGND VPWR VPWR _5075_/D sky130_fd_sc_hd__or4_1
X_4025_ _4025_/A _5378_/B VGND VGND VPWR VPWR _4025_/Y sky130_fd_sc_hd__nand2_8
XFILLER_56_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5976_ _5976_/A _5976_/B _5976_/C _5976_/D VGND VGND VPWR VPWR _5976_/X sky130_fd_sc_hd__or4_2
XFILLER_52_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4927_ _5023_/A _4927_/B VGND VGND VPWR VPWR _4932_/A sky130_fd_sc_hd__nor2_2
X_4858_ _4399_/Y _4845_/B _5171_/A _4856_/X _4857_/X VGND VGND VPWR VPWR _4858_/X
+ sky130_fd_sc_hd__a2111o_4
XFILLER_60_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3809_ _6469_/Q _6468_/Q VGND VGND VPWR VPWR _3810_/B sky130_fd_sc_hd__nor2_1
XFILLER_193_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4789_ _4772_/A _4575_/B _4453_/Y _4719_/X VGND VGND VPWR VPWR _4789_/X sky130_fd_sc_hd__a22o_1
X_6528_ _6931_/CLK _6528_/D fanout885/X VGND VGND VPWR VPWR _6528_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_7_csclk _6744_/CLK VGND VGND VPWR VPWR _6554_/CLK sky130_fd_sc_hd__clkbuf_8
X_6459_ _3957_/A1 _6459_/D _6414_/X VGND VGND VPWR VPWR _6459_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_133_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5830_ _7181_/Q _6110_/S _5828_/X _5829_/X VGND VGND VPWR VPWR _7181_/D sky130_fd_sc_hd__o22a_1
X_5761_ _7063_/Q _5974_/A2 _5926_/A2 wire486/X VGND VGND VPWR VPWR _5761_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4712_ _4922_/A _4712_/B _5069_/B _4936_/A VGND VGND VPWR VPWR _4713_/D sky130_fd_sc_hd__or4_4
XFILLER_187_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5692_ _7165_/Q _5705_/B _5706_/B VGND VGND VPWR VPWR _5692_/X sky130_fd_sc_hd__and3_4
XFILLER_175_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4643_ _4812_/A _4819_/B _5062_/A VGND VGND VPWR VPWR _4897_/B sky130_fd_sc_hd__or3_4
X_4574_ _5128_/A VGND VGND VPWR VPWR _4574_/Y sky130_fd_sc_hd__inv_2
Xhold702 _6820_/Q VGND VGND VPWR VPWR wire559/A sky130_fd_sc_hd__bufbuf_16
Xhold724 _6975_/Q VGND VGND VPWR VPWR hold724/X sky130_fd_sc_hd__bufbuf_16
XFILLER_143_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6313_ _6662_/Q wire647/X wire638/X _6548_/Q VGND VGND VPWR VPWR _6330_/A sky130_fd_sc_hd__a22o_1
X_3525_ _7033_/Q _5459_/A _4292_/A wire564/X _3523_/X VGND VGND VPWR VPWR _3533_/A
+ sky130_fd_sc_hd__a221o_2
Xhold746 _6488_/Q VGND VGND VPWR VPWR hold746/X sky130_fd_sc_hd__bufbuf_16
Xhold713 _6756_/Q VGND VGND VPWR VPWR hold713/X sky130_fd_sc_hd__bufbuf_16
Xhold735 _4221_/X VGND VGND VPWR VPWR _6681_/D sky130_fd_sc_hd__bufbuf_16
XFILLER_143_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6244_ _6540_/Q wire592/X wire612/X _6649_/Q _6243_/X VGND VGND VPWR VPWR _6247_/C
+ sky130_fd_sc_hd__a221o_1
Xhold768 _6822_/Q VGND VGND VPWR VPWR hold768/X sky130_fd_sc_hd__bufbuf_16
Xhold779 _6758_/Q VGND VGND VPWR VPWR hold779/X sky130_fd_sc_hd__bufbuf_16
Xhold757 _4225_/X VGND VGND VPWR VPWR _6683_/D sky130_fd_sc_hd__bufbuf_16
X_3456_ input16/X _3368_/Y _4130_/A _6608_/Q VGND VGND VPWR VPWR _3456_/X sky130_fd_sc_hd__a22o_2
X_3387_ input41/X _4023_/S _5324_/A _6915_/Q VGND VGND VPWR VPWR _3387_/X sky130_fd_sc_hd__a22o_1
X_6175_ _6906_/Q _6021_/A wire646/X wire533/X _6174_/X VGND VGND VPWR VPWR _6181_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_97_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5126_ _5126_/A _5126_/B VGND VGND VPWR VPWR _5127_/A sky130_fd_sc_hd__nor2_1
X_5057_ _5057_/A _5057_/B VGND VGND VPWR VPWR _5057_/X sky130_fd_sc_hd__or2_4
XFILLER_111_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4008_ _4034_/A _6421_/B _4007_/X _4023_/S _5594_/B VGND VGND VPWR VPWR _4024_/S
+ sky130_fd_sc_hd__o221a_4
XFILLER_72_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5959_ _5959_/A _5959_/B _5959_/C _5959_/D VGND VGND VPWR VPWR _5959_/X sky130_fd_sc_hd__or4_1
XFILLER_53_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold40 hold40/A VGND VGND VPWR VPWR hold40/X sky130_fd_sc_hd__bufbuf_16
XFILLER_0_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold51 hold51/A VGND VGND VPWR VPWR hold51/X sky130_fd_sc_hd__bufbuf_16
Xhold73 hold73/A VGND VGND VPWR VPWR hold73/X sky130_fd_sc_hd__bufbuf_16
XFILLER_152_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold62 hold62/A VGND VGND VPWR VPWR hold62/X sky130_fd_sc_hd__bufbuf_16
XFILLER_36_609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold84 hold84/A VGND VGND VPWR VPWR hold84/X sky130_fd_sc_hd__bufbuf_16
XFILLER_152_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold95 hold95/A VGND VGND VPWR VPWR hold95/X sky130_fd_sc_hd__bufbuf_16
XFILLER_189_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_4 _6429_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3310_ _4034_/A _4241_/A VGND VGND VPWR VPWR _3310_/Y sky130_fd_sc_hd__nor2_8
XFILLER_140_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4290_ _6410_/A0 hold566/X _4291_/S VGND VGND VPWR VPWR _4290_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3241_ _7165_/Q VGND VGND VPWR VPWR _3241_/Y sky130_fd_sc_hd__inv_6
XFILLER_113_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6931_ _6931_/CLK _6931_/D fanout885/X VGND VGND VPWR VPWR _6931_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6862_ _7145_/CLK _6862_/D _6421_/A VGND VGND VPWR VPWR _6862_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_179_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5813_ _6914_/Q wire699/X wire666/X _6866_/Q _5811_/X VGND VGND VPWR VPWR _5813_/X
+ sky130_fd_sc_hd__a221o_1
X_6793_ _3545_/A1 _6793_/D _6451_/X VGND VGND VPWR VPWR _6793_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_50_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5744_ _7177_/Q _6110_/S _5742_/X _5743_/X VGND VGND VPWR VPWR _7177_/D sky130_fd_sc_hd__o22a_1
X_5675_ _7165_/Q _5705_/B _5701_/C VGND VGND VPWR VPWR _5675_/X sky130_fd_sc_hd__and3_4
Xclkbuf_leaf_72_csclk _6744_/CLK VGND VGND VPWR VPWR _6736_/CLK sky130_fd_sc_hd__clkbuf_8
X_4626_ _5114_/B VGND VGND VPWR VPWR _4626_/Y sky130_fd_sc_hd__inv_2
XFILLER_163_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold510 _6590_/Q VGND VGND VPWR VPWR hold510/X sky130_fd_sc_hd__bufbuf_16
X_4557_ _4883_/A _5119_/A _4557_/C _4557_/D VGND VGND VPWR VPWR _4559_/C sky130_fd_sc_hd__or4_1
Xhold532 _6650_/Q VGND VGND VPWR VPWR hold532/X sky130_fd_sc_hd__bufbuf_16
Xhold521 _7105_/Q VGND VGND VPWR VPWR hold521/X sky130_fd_sc_hd__bufbuf_16
Xhold554 _4287_/X VGND VGND VPWR VPWR _6738_/D sky130_fd_sc_hd__bufbuf_16
Xhold543 _6845_/Q VGND VGND VPWR VPWR hold543/X sky130_fd_sc_hd__bufbuf_16
Xhold587 _7152_/Q VGND VGND VPWR VPWR hold587/X sky130_fd_sc_hd__bufbuf_16
X_4488_ _4655_/A _4651_/B VGND VGND VPWR VPWR _4488_/X sky130_fd_sc_hd__or2_1
Xhold576 _6614_/Q VGND VGND VPWR VPWR hold576/X sky130_fd_sc_hd__bufbuf_16
XFILLER_104_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3508_ _3508_/A _3733_/B VGND VGND VPWR VPWR _4304_/A sky130_fd_sc_hd__nor2_8
Xhold565 _6659_/Q VGND VGND VPWR VPWR hold565/X sky130_fd_sc_hd__bufbuf_16
XFILLER_104_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6227_ _7108_/Q wire712/X wire625/X _6948_/Q VGND VGND VPWR VPWR _6227_/X sky130_fd_sc_hd__a22o_1
X_3439_ _6882_/Q _3353_/Y _5405_/A _6986_/Q VGND VGND VPWR VPWR _3439_/X sky130_fd_sc_hd__a22o_1
XFILLER_58_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold598 _4195_/X VGND VGND VPWR VPWR _6658_/D sky130_fd_sc_hd__bufbuf_16
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ _6857_/Q _6060_/B _6144_/X _6157_/X _6109_/S VGND VGND VPWR VPWR _6158_/X
+ sky130_fd_sc_hd__o221a_1
X_5109_ _4748_/B _5041_/X _5056_/B _5104_/Y VGND VGND VPWR VPWR _5178_/B sky130_fd_sc_hd__a211o_4
Xclkbuf_leaf_10_csclk _6708_/CLK VGND VGND VPWR VPWR _6712_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6089_ _6975_/Q wire641/X wire639/X _6879_/Q _6087_/X VGND VGND VPWR VPWR _6106_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_73_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_csclk _6708_/CLK VGND VGND VPWR VPWR _6626_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_26_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput141 wb_dat_i[18] VGND VGND VPWR VPWR _6383_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput130 wb_adr_i[9] VGND VGND VPWR VPWR _4351_/A sky130_fd_sc_hd__clkbuf_4
Xinput163 wb_dat_i[9] VGND VGND VPWR VPWR _6380_/B1 sky130_fd_sc_hd__clkbuf_4
Xinput152 wb_dat_i[28] VGND VGND VPWR VPWR _6390_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3790_ _6997_/Q _5423_/A _4310_/A _6758_/Q _3789_/X VGND VGND VPWR VPWR _3792_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5460_ _5532_/A0 hold725/X _5467_/S VGND VGND VPWR VPWR _7029_/D sky130_fd_sc_hd__mux2_1
X_4411_ _4871_/A _4997_/A VGND VGND VPWR VPWR _4411_/Y sky130_fd_sc_hd__nor2_2
XFILLER_145_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5391_ wire773/X hold630/X _5395_/S VGND VGND VPWR VPWR _6968_/D sky130_fd_sc_hd__mux2_1
X_7130_ _7147_/CLK _7130_/D fanout886/X VGND VGND VPWR VPWR _7130_/Q sky130_fd_sc_hd__dfrtp_2
X_4342_ _4654_/A _4654_/B VGND VGND VPWR VPWR _4690_/A sky130_fd_sc_hd__nand2_8
XFILLER_153_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4273_ hold454/X _4303_/A0 _4273_/S VGND VGND VPWR VPWR _4273_/X sky130_fd_sc_hd__mux2_1
X_7061_ _7105_/CLK _7061_/D fanout862/X VGND VGND VPWR VPWR _7061_/Q sky130_fd_sc_hd__dfstp_4
X_3224_ _6984_/Q VGND VGND VPWR VPWR _3224_/Y sky130_fd_sc_hd__inv_2
X_6012_ _6012_/A _6035_/A _6018_/A VGND VGND VPWR VPWR _6012_/X sky130_fd_sc_hd__and3_4
XFILLER_101_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
.ends

