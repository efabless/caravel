* NGSPICE file created from housekeeping.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtn_1 abstract view
.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_1 abstract view
.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_2 abstract view
.subckt sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt housekeeping VGND VPWR debug_in debug_mode debug_oeb debug_out irq[0] irq[1]
+ irq[2] mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13]
+ mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18]
+ mask_rev_in[19] mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23]
+ mask_rev_in[24] mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4]
+ mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14]
+ mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19]
+ mgmt_gpio_in[1] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23]
+ mgmt_gpio_in[24] mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28]
+ mgmt_gpio_in[29] mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32]
+ mgmt_gpio_in[33] mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37]
+ mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7]
+ mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16]
+ mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20]
+ mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2]
+ mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[35] mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4]
+ mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18]
+ mgmt_gpio_out[19] mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22]
+ mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27]
+ mgmt_gpio_out[28] mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31]
+ mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36]
+ mgmt_gpio_out[37] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oeb
+ pad_flash_csb pad_flash_csb_oeb pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ieb
+ pad_flash_io0_oeb pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ieb pad_flash_io1_oeb
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1]
+ pll_div[2] pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0]
+ pll_trim[10] pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16]
+ pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22]
+ pll_trim[23] pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5]
+ pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out[0] pwr_ctrl_out[1]
+ pwr_ctrl_out[2] pwr_ctrl_out[3] qspi_enabled reset ser_rx ser_tx serial_clock serial_data_1
+ serial_data_2 serial_load serial_resetn spi_csb spi_enabled spi_sck spi_sdi spi_sdo
+ spi_sdoenb spimemio_flash_clk spimemio_flash_csb spimemio_flash_io0_di spimemio_flash_io0_do
+ spimemio_flash_io0_oeb spimemio_flash_io1_di spimemio_flash_io1_do spimemio_flash_io1_oeb
+ spimemio_flash_io2_di spimemio_flash_io2_do spimemio_flash_io2_oeb spimemio_flash_io3_di
+ spimemio_flash_io3_do spimemio_flash_io3_oeb trap uart_enabled user_clock usr1_vcc_pwrgood
+ usr1_vdd_pwrgood usr2_vcc_pwrgood usr2_vdd_pwrgood wb_ack_o wb_adr_i[0] wb_adr_i[10]
+ wb_adr_i[11] wb_adr_i[12] wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17]
+ wb_adr_i[18] wb_adr_i[19] wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23]
+ wb_adr_i[24] wb_adr_i[25] wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2]
+ wb_adr_i[30] wb_adr_i[31] wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7]
+ wb_adr_i[8] wb_adr_i[9] wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11]
+ wb_dat_i[12] wb_dat_i[13] wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18]
+ wb_dat_i[19] wb_dat_i[1] wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24]
+ wb_dat_i[25] wb_dat_i[26] wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30]
+ wb_dat_i[31] wb_dat_i[3] wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8]
+ wb_dat_i[9] wb_dat_o[0] wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14]
+ wb_dat_o[15] wb_dat_o[16] wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20]
+ wb_dat_o[21] wb_dat_o[22] wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27]
+ wb_dat_o[28] wb_dat_o[29] wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4]
+ wb_dat_o[5] wb_dat_o[6] wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0]
+ wb_sel_i[1] wb_sel_i[2] wb_sel_i[3] wb_stb_i wb_we_i
XFILLER_79_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6914_ _6963_/CLK _6914_/D _7042_/SET_B VGND VGND VPWR VPWR _6914_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6845_ _7141_/CLK _6845_/D wire3980/X VGND VGND VPWR VPWR _6845_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6776_ _7204_/CLK _6776_/D wire4261/X VGND VGND VPWR VPWR _6776_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3988_ hold700/X _4311_/A0 _3988_/S VGND VGND VPWR VPWR _6486_/D sky130_fd_sc_hd__mux2_1
Xwire709 _5249_/S VGND VGND VPWR VPWR _5248_/S sky130_fd_sc_hd__buf_2
XFILLER_167_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5727_ _6055_/A1 _5727_/A2 _5727_/B1 _6053_/B2 _5726_/X VGND VGND VPWR VPWR _5728_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_109_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5658_ _7151_/Q _7150_/Q VGND VGND VPWR VPWR _5706_/C sky130_fd_sc_hd__and2_2
X_4609_ _4609_/A _4609_/B _4794_/A VGND VGND VPWR VPWR _4644_/C sky130_fd_sc_hd__nor3_1
XFILLER_163_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5589_ _6562_/Q _5648_/C _7143_/Q VGND VGND VPWR VPWR _5589_/X sky130_fd_sc_hd__a21o_1
Xwire4016 wire4016/A VGND VGND VPWR VPWR wire4016/X sky130_fd_sc_hd__clkbuf_1
Xhold340 _6890_/Q VGND VGND VPWR VPWR hold340/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3304 _4610_/X VGND VGND VPWR VPWR _4652_/B sky130_fd_sc_hd__clkbuf_1
Xhold351 _6751_/Q VGND VGND VPWR VPWR hold351/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 _6753_/Q VGND VGND VPWR VPWR hold362/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire4049 wire4049/A VGND VGND VPWR VPWR wire4049/X sky130_fd_sc_hd__clkbuf_2
XFILLER_132_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold373 _7207_/Q VGND VGND VPWR VPWR hold373/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3315 _4673_/A VGND VGND VPWR VPWR _4694_/B sky130_fd_sc_hd__clkbuf_2
Xwire3326 _4562_/X VGND VGND VPWR VPWR _4569_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold384 _7209_/Q VGND VGND VPWR VPWR hold384/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3337 _4638_/B VGND VGND VPWR VPWR _4614_/A sky130_fd_sc_hd__clkbuf_1
Xhold395 _6843_/Q VGND VGND VPWR VPWR hold395/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2603 _4669_/X VGND VGND VPWR VPWR wire2603/X sky130_fd_sc_hd__clkbuf_1
Xwire2614 wire2614/A VGND VGND VPWR VPWR _6262_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_132_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2625 _6307_/A2 VGND VGND VPWR VPWR _6272_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2636 _6329_/B1 VGND VGND VPWR VPWR _6264_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire2647 _6273_/B1 VGND VGND VPWR VPWR _6326_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1902 _6943_/Q VGND VGND VPWR VPWR _5801_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2658 _6033_/X VGND VGND VPWR VPWR _6188_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire1913 _3746_/A1 VGND VGND VPWR VPWR wire1913/X sky130_fd_sc_hd__clkbuf_1
Xwire1924 wire1925/X VGND VGND VPWR VPWR _5993_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire1935 _3389_/A1 VGND VGND VPWR VPWR wire1935/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1946 wire1947/X VGND VGND VPWR VPWR _3611_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_100_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1957 _5811_/A1 VGND VGND VPWR VPWR wire1957/X sky130_fd_sc_hd__clkbuf_1
Xwire1968 wire1969/X VGND VGND VPWR VPWR _6129_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire1979 _5721_/A1 VGND VGND VPWR VPWR _6054_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3860 wire3861/X VGND VGND VPWR VPWR wire3860/X sky130_fd_sc_hd__clkbuf_1
Xwire3871 wire3872/X VGND VGND VPWR VPWR wire3871/X sky130_fd_sc_hd__clkbuf_1
Xwire3882 wire3883/X VGND VGND VPWR VPWR _3785_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_96_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3893 wire3894/X VGND VGND VPWR VPWR wire3893/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4960_ _4960_/A _4960_/B _4959_/X VGND VGND VPWR VPWR _4961_/B sky130_fd_sc_hd__or3b_1
X_3911_ _6346_/A _3888_/B _3191_/Y VGND VGND VPWR VPWR _6691_/D sky130_fd_sc_hd__o21ai_1
XFILLER_44_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4891_ _4516_/B _4871_/Y _4880_/X _4890_/X VGND VGND VPWR VPWR _4891_/X sky130_fd_sc_hd__a211o_1
X_6630_ _7206_/CLK _6630_/D VGND VGND VPWR VPWR _6630_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3842_ _6456_/Q _3794_/B _6458_/Q VGND VGND VPWR VPWR _3842_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6561_ _7110_/CLK _6561_/D wire3999/X VGND VGND VPWR VPWR _6561_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_158_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3773_ _7066_/Q _3292_/Y _4028_/A _6521_/Q VGND VGND VPWR VPWR _3773_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5512_ _5536_/A1 hold707/X _5514_/S VGND VGND VPWR VPWR _7074_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6492_ _6825_/CLK _6492_/D _6495_/SET_B VGND VGND VPWR VPWR _6492_/Q sky130_fd_sc_hd__dfstp_1
X_5443_ _5575_/A0 hold199/X _5444_/S VGND VGND VPWR VPWR _7013_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5374_ _5374_/A0 hold300/X _5375_/S VGND VGND VPWR VPWR _6952_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7113_ _7129_/CLK _7113_/D wire4061/A VGND VGND VPWR VPWR _7113_/Q sky130_fd_sc_hd__dfrtp_1
X_4325_ hold548/X _4325_/A1 _4328_/S VGND VGND VPWR VPWR _6766_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7044_ _7084_/CLK _7044_/D _7035_/SET_B VGND VGND VPWR VPWR _7044_/Q sky130_fd_sc_hd__dfrtp_1
X_4256_ hold399/X _4256_/A1 _4257_/S VGND VGND VPWR VPWR _6709_/D sky130_fd_sc_hd__mux2_1
Xwire1209 wire1210/X VGND VGND VPWR VPWR _5439_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_47_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3207_ _7061_/Q VGND VGND VPWR VPWR _3207_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4187_ _6645_/Q wire374/X _4188_/S VGND VGND VPWR VPWR _6645_/D sky130_fd_sc_hd__mux2_1
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6828_ _7130_/CLK _6828_/D wire4058/X VGND VGND VPWR VPWR _6828_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire506 _5282_/S VGND VGND VPWR VPWR _5281_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire517 _5267_/S VGND VGND VPWR VPWR _5264_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_6759_ _6761_/CLK _6759_/D wire4019/X VGND VGND VPWR VPWR _6759_/Q sky130_fd_sc_hd__dfrtp_1
Xwire528 wire529/X VGND VGND VPWR VPWR _4108_/S sky130_fd_sc_hd__clkbuf_2
Xwire539 wire540/X VGND VGND VPWR VPWR wire539/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3101 _5951_/A2 VGND VGND VPWR VPWR _5944_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3112 wire3112/A VGND VGND VPWR VPWR _5922_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3123 wire3123/A VGND VGND VPWR VPWR _5748_/A2 sky130_fd_sc_hd__clkbuf_2
Xhold170 _6499_/Q VGND VGND VPWR VPWR hold170/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 _7051_/Q VGND VGND VPWR VPWR hold181/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold192 _7138_/Q VGND VGND VPWR VPWR hold192/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3134 _5761_/A2 VGND VGND VPWR VPWR _5749_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_120_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2400 _5908_/A1 VGND VGND VPWR VPWR _6274_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire3145 _5758_/A2 VGND VGND VPWR VPWR _5739_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2411 _6508_/Q VGND VGND VPWR VPWR _6276_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3156 _5995_/A2 VGND VGND VPWR VPWR wire3156/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3167 _4668_/X VGND VGND VPWR VPWR _5072_/A3 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2422 wire2423/X VGND VGND VPWR VPWR _3559_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2433 wire2434/X VGND VGND VPWR VPWR _3345_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2444 wire2444/A VGND VGND VPWR VPWR _3384_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_144_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2455 _6206_/B1 VGND VGND VPWR VPWR _6155_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1710 _5763_/A1 VGND VGND VPWR VPWR _6113_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1721 wire1722/X VGND VGND VPWR VPWR wire1721/X sky130_fd_sc_hd__clkbuf_1
Xwire2466 _6330_/B1 VGND VGND VPWR VPWR _6313_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2477 _6282_/A2 VGND VGND VPWR VPWR _6309_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1732 _7030_/Q VGND VGND VPWR VPWR _5778_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2488 wire2489/X VGND VGND VPWR VPWR _6337_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1743 _5701_/B2 VGND VGND VPWR VPWR wire1743/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1754 _6107_/B2 VGND VGND VPWR VPWR _5767_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire2499 _6181_/A2 VGND VGND VPWR VPWR _6339_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1765 wire1766/X VGND VGND VPWR VPWR wire1765/X sky130_fd_sc_hd__clkbuf_1
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1776 wire1777/X VGND VGND VPWR VPWR _6108_/A1 sky130_fd_sc_hd__clkbuf_1
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1787 _7010_/Q VGND VGND VPWR VPWR wire1787/X sky130_fd_sc_hd__clkbuf_1
Xwire1798 _7005_/Q VGND VGND VPWR VPWR _3553_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout3562 hold21/X VGND VGND VPWR VPWR hold22/A sky130_fd_sc_hd__buf_6
X_4110_ _4110_/A0 hold187/X _4110_/S VGND VGND VPWR VPWR _6579_/D sky130_fd_sc_hd__mux2_1
XFILLER_111_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5090_ _5090_/A _5090_/B _5089_/X VGND VGND VPWR VPWR _5170_/B sky130_fd_sc_hd__or3b_1
XFILLER_110_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3690 _3235_/Y VGND VGND VPWR VPWR _5705_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4041_ _6393_/A0 hold443/X _4045_/S VGND VGND VPWR VPWR _6531_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5992_ _6033_/A _6020_/C _6040_/C VGND VGND VPWR VPWR _5992_/X sky130_fd_sc_hd__and3_1
XFILLER_52_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4943_ _4395_/Y _5060_/B _4833_/Y VGND VGND VPWR VPWR _5053_/B sky130_fd_sc_hd__a21o_1
XFILLER_178_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4874_ _5001_/A _4931_/B _5001_/C VGND VGND VPWR VPWR _4897_/C sky130_fd_sc_hd__and3_1
X_6613_ _6702_/CLK _6613_/D _6440_/A VGND VGND VPWR VPWR _6613_/Q sky130_fd_sc_hd__dfrtp_1
Xmax_length3109 _5663_/X VGND VGND VPWR VPWR _5819_/B1 sky130_fd_sc_hd__clkbuf_1
X_3825_ _3824_/X hold24/A _3828_/S VGND VGND VPWR VPWR _6466_/D sky130_fd_sc_hd__mux2_1
XFILLER_193_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6544_ _3945_/A1 _6544_/D _6432_/X VGND VGND VPWR VPWR _6544_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3756_ _6011_/B2 wire866/X wire851/X _3756_/B2 _3739_/X VGND VGND VPWR VPWR _3760_/A
+ sky130_fd_sc_hd__a221o_1
Xclkbuf_3_5_0_csclk clkbuf_3_5_0_csclk/A VGND VGND VPWR VPWR _6579_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_180_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6475_ _6824_/CLK _6475_/D _6483_/SET_B VGND VGND VPWR VPWR _6475_/Q sky130_fd_sc_hd__dfstp_1
X_3687_ _6995_/Q _3762_/A2 _3687_/B1 _3687_/B2 _3686_/X VGND VGND VPWR VPWR _3687_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5426_ _5462_/A0 hold482/X _5429_/S VGND VGND VPWR VPWR _6998_/D sky130_fd_sc_hd__mux2_1
Xoutput220 _6546_/Q VGND VGND VPWR VPWR mgmt_gpio_out[16] sky130_fd_sc_hd__buf_12
XFILLER_161_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput231 _6828_/Q VGND VGND VPWR VPWR mgmt_gpio_out[26] sky130_fd_sc_hd__buf_12
Xoutput242 wire1488/X VGND VGND VPWR VPWR mgmt_gpio_out[36] sky130_fd_sc_hd__buf_12
Xoutput253 wire3675/X VGND VGND VPWR VPWR pad_flash_csb sky130_fd_sc_hd__buf_12
Xoutput264 _6806_/Q VGND VGND VPWR VPWR pll_bypass sky130_fd_sc_hd__buf_12
X_5357_ _5588_/A0 hold651/X _5357_/S VGND VGND VPWR VPWR _6937_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput275 _6490_/Q VGND VGND VPWR VPWR pll_trim[0] sky130_fd_sc_hd__buf_12
Xoutput286 _6491_/Q VGND VGND VPWR VPWR pll_trim[1] sky130_fd_sc_hd__buf_12
XFILLER_114_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput297 _6496_/Q VGND VGND VPWR VPWR pll_trim[6] sky130_fd_sc_hd__buf_12
X_4308_ _4308_/A0 hold352/X _4311_/S VGND VGND VPWR VPWR _6752_/D sky130_fd_sc_hd__mux2_1
X_5288_ _5477_/A0 hold93/X _5291_/S VGND VGND VPWR VPWR _6875_/D sky130_fd_sc_hd__mux2_1
Xwire1006 _5860_/S VGND VGND VPWR VPWR _5838_/S sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1017 _4642_/X VGND VGND VPWR VPWR _4643_/B1 sky130_fd_sc_hd__clkbuf_1
X_7027_ _7027_/CLK _7027_/D fanout3976/X VGND VGND VPWR VPWR _7027_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1028 _3720_/B1 VGND VGND VPWR VPWR _3539_/B1 sky130_fd_sc_hd__clkbuf_1
X_4239_ _5534_/A1 hold336/X _4239_/S VGND VGND VPWR VPWR _6685_/D sky130_fd_sc_hd__mux2_1
XFILLER_75_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1039 _4046_/A VGND VGND VPWR VPWR _3767_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_74_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire358 wire359/X VGND VGND VPWR VPWR wire358/X sky130_fd_sc_hd__clkbuf_2
XFILLER_139_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire369 wire370/X VGND VGND VPWR VPWR wire369/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length2953 _5842_/A2 VGND VGND VPWR VPWR wire2949/A sky130_fd_sc_hd__clkbuf_1
XFILLER_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length2975 _5685_/X VGND VGND VPWR VPWR wire2967/A sky130_fd_sc_hd__clkbuf_1
XFILLER_136_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2230 _6711_/Q VGND VGND VPWR VPWR wire2230/X sky130_fd_sc_hd__clkbuf_1
Xwire2241 _6704_/Q VGND VGND VPWR VPWR _6305_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2252 _6262_/A1 VGND VGND VPWR VPWR _5890_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2274 wire2275/X VGND VGND VPWR VPWR _6236_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire1540 _7131_/Q VGND VGND VPWR VPWR _6123_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2285 _6662_/Q VGND VGND VPWR VPWR _6277_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2296 _6638_/Q VGND VGND VPWR VPWR _6337_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire1551 hold604/X VGND VGND VPWR VPWR _6198_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1562 _7115_/Q VGND VGND VPWR VPWR wire1562/X sky130_fd_sc_hd__clkbuf_1
Xwire1573 _5548_/A1 VGND VGND VPWR VPWR _6099_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire1584 _6117_/B2 VGND VGND VPWR VPWR wire1584/X sky130_fd_sc_hd__clkbuf_1
Xwire1595 _7092_/Q VGND VGND VPWR VPWR _3648_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3610_ _5906_/B2 _4153_/A _3519_/Y _6286_/A1 VGND VGND VPWR VPWR _3610_/X sky130_fd_sc_hd__a22o_1
X_4590_ _4590_/A _4694_/B VGND VGND VPWR VPWR _4598_/B sky130_fd_sc_hd__nor2_1
X_3541_ _3541_/A _3541_/B _3541_/C _3541_/D VGND VGND VPWR VPWR _3542_/D sky130_fd_sc_hd__or4_1
Xwire870 wire871/X VGND VGND VPWR VPWR wire870/X sky130_fd_sc_hd__clkbuf_2
Xwire881 wire881/A VGND VGND VPWR VPWR wire881/X sky130_fd_sc_hd__clkbuf_1
Xwire892 _3336_/Y VGND VGND VPWR VPWR wire892/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6260_ _6666_/Q _6283_/A2 _6325_/B1 _6682_/Q VGND VGND VPWR VPWR _6260_/X sky130_fd_sc_hd__a22o_1
X_3472_ _3472_/A _3472_/B VGND VGND VPWR VPWR _3472_/Y sky130_fd_sc_hd__nor2_1
Xfanout4060 wire4066/A VGND VGND VPWR VPWR fanout4060/X sky130_fd_sc_hd__buf_6
XFILLER_115_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5211_ _5211_/A0 hold526/X _5211_/S VGND VGND VPWR VPWR _6811_/D sky130_fd_sc_hd__mux2_1
X_6191_ _6191_/A1 _5994_/X _6191_/B1 _6191_/B2 _6191_/C1 VGND VGND VPWR VPWR _6192_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_142_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5142_ _5142_/A _5142_/B _5141_/X VGND VGND VPWR VPWR _5172_/C sky130_fd_sc_hd__or3b_1
Xfanout3392 _5410_/A0 VGND VGND VPWR VPWR _5587_/A0 sky130_fd_sc_hd__buf_6
XFILLER_69_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5073_ _5095_/A _5073_/B _5072_/X VGND VGND VPWR VPWR _5073_/X sky130_fd_sc_hd__or3b_1
XFILLER_84_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4024_ _4024_/A0 _4122_/A0 _4027_/S VGND VGND VPWR VPWR _4024_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5975_ _7157_/Q _7158_/Q VGND VGND VPWR VPWR _6021_/A sky130_fd_sc_hd__or2_2
XFILLER_52_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4926_ _4926_/A _4992_/B VGND VGND VPWR VPWR _5031_/C sky130_fd_sc_hd__nand2_1
XFILLER_138_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4857_ _4857_/A _4857_/B _4857_/C _4857_/D VGND VGND VPWR VPWR _4857_/X sky130_fd_sc_hd__and4_1
XFILLER_193_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3808_ hold24/A _3823_/B VGND VGND VPWR VPWR _3821_/S sky130_fd_sc_hd__and2_1
XFILLER_176_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4788_ _4743_/B _4805_/B2 _4799_/B1 _4679_/B VGND VGND VPWR VPWR _4985_/C sky130_fd_sc_hd__o22ai_1
X_6527_ _6799_/CLK _6527_/D _6743_/SET_B VGND VGND VPWR VPWR _6527_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3739_ _5657_/A1 wire956/X wire895/X _5986_/A1 VGND VGND VPWR VPWR _3739_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6458_ _6545_/CLK _6458_/D _6413_/X VGND VGND VPWR VPWR _6458_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5409_ _5586_/A0 hold599/X _5409_/S VGND VGND VPWR VPWR _6983_/D sky130_fd_sc_hd__mux2_1
X_6389_ _4228_/A _6389_/A2 _6388_/X VGND VGND VPWR VPWR _6389_/X sky130_fd_sc_hd__a21o_1
XFILLER_125_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length4163 input58/X VGND VGND VPWR VPWR wire4162/A sky130_fd_sc_hd__clkbuf_1
XFILLER_156_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length3462 _5540_/A1 VGND VGND VPWR VPWR _4329_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_184_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length3495 _6396_/A0 VGND VGND VPWR VPWR _4316_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_109_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length2772 _6150_/A2 VGND VGND VPWR VPWR _6052_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_125_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2060 _6864_/Q VGND VGND VPWR VPWR _6185_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire2071 wire2072/X VGND VGND VPWR VPWR _6215_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire2082 wire2083/X VGND VGND VPWR VPWR _3575_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_94_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2093 _6847_/Q VGND VGND VPWR VPWR _6169_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1370 hold70/X VGND VGND VPWR VPWR _3489_/B sky130_fd_sc_hd__clkbuf_1
Xwire1381 _3512_/B VGND VGND VPWR VPWR _3711_/A sky130_fd_sc_hd__buf_2
XFILLER_47_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5760_ _7069_/Q _5760_/A2 _5760_/B1 _5760_/B2 _5759_/X VGND VGND VPWR VPWR _5771_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4711_ _4638_/A _4603_/B _4839_/B _4689_/X wire357/X VGND VGND VPWR VPWR _4713_/C
+ sky130_fd_sc_hd__o311a_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5691_ _5693_/A _5691_/B VGND VGND VPWR VPWR _5691_/Y sky130_fd_sc_hd__nand2_1
XFILLER_147_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4642_ _4642_/A _4642_/B _4642_/C _4642_/D VGND VGND VPWR VPWR _4642_/X sky130_fd_sc_hd__and4_1
XFILLER_163_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4573_ _4484_/B _4573_/B VGND VGND VPWR VPWR _4981_/C sky130_fd_sc_hd__nand2b_1
XFILLER_190_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold703 _6984_/Q VGND VGND VPWR VPWR hold703/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold714 _6474_/Q VGND VGND VPWR VPWR hold714/X sky130_fd_sc_hd__dlygate4sd3_1
X_6312_ _6689_/Q _6337_/A2 _6312_/B1 _6312_/B2 VGND VGND VPWR VPWR _6312_/X sky130_fd_sc_hd__a22o_1
X_3524_ _3524_/A _3524_/B _3524_/C _3524_/D VGND VGND VPWR VPWR _3524_/X sky130_fd_sc_hd__or4_1
Xhold725 _7197_/Q VGND VGND VPWR VPWR hold725/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6243_ _6243_/A1 wire977/X _6232_/X _6242_/X _6293_/C1 VGND VGND VPWR VPWR _6243_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_170_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3455_ _3462_/A _3510_/A VGND VGND VPWR VPWR _4040_/A sky130_fd_sc_hd__nor2_2
XFILLER_130_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6174_ _6904_/Q _6174_/A2 _6174_/B1 _6174_/B2 VGND VGND VPWR VPWR _6174_/X sky130_fd_sc_hd__a22o_1
X_3386_ _6190_/A1 _3386_/A2 _5562_/A _7125_/Q _3381_/X VGND VGND VPWR VPWR _3392_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5125_ _5125_/A _5125_/B VGND VGND VPWR VPWR _5128_/C sky130_fd_sc_hd__nor2_1
XFILLER_111_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5056_ _5023_/A _4673_/A _4950_/B _4887_/C VGND VGND VPWR VPWR _5056_/X sky130_fd_sc_hd__o211a_1
XFILLER_38_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4007_ _5481_/A0 hold633/X _4007_/S VGND VGND VPWR VPWR _6503_/D sky130_fd_sc_hd__mux2_1
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_1_wb_clk_i clkbuf_1_0_1_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_25_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5958_ _6328_/B2 _5958_/A2 _5958_/B1 _7094_/Q VGND VGND VPWR VPWR _5958_/X sky130_fd_sc_hd__a22o_1
XFILLER_52_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4909_ _4915_/C VGND VGND VPWR VPWR _4909_/Y sky130_fd_sc_hd__inv_2
X_5889_ _6256_/B2 _5889_/A2 _5958_/B1 _7091_/Q VGND VGND VPWR VPWR _5889_/X sky130_fd_sc_hd__a22o_1
XFILLER_138_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length2068 _6861_/Q VGND VGND VPWR VPWR wire2065/A sky130_fd_sc_hd__clkbuf_1
XFILLER_107_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_2_0_csclk clkbuf_2_3_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_5_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_134_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold30 hold30/A VGND VGND VPWR VPWR hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A VGND VGND VPWR VPWR hold41/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold52 hold52/A VGND VGND VPWR VPWR hold52/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold63 hold63/A VGND VGND VPWR VPWR hold63/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 hold74/A VGND VGND VPWR VPWR hold74/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 hold85/A VGND VGND VPWR VPWR hold85/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 hold96/A VGND VGND VPWR VPWR hold96/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length3281 _5223_/B VGND VGND VPWR VPWR _4270_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_144_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_5 mgmt_gpio_in[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3240_ _4565_/A VGND VGND VPWR VPWR _4610_/A sky130_fd_sc_hd__clkinv_2
XFILLER_112_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6930_ _7131_/CLK _6930_/D wire4055/X VGND VGND VPWR VPWR _6930_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6861_ _7110_/CLK _6861_/D wire3999/X VGND VGND VPWR VPWR _6861_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_6_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _6683_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_62_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5812_ _6160_/B2 _5812_/A2 _5812_/B1 _6162_/A1 _5811_/X VGND VGND VPWR VPWR _5813_/D
+ sky130_fd_sc_hd__a221o_1
X_6792_ _6811_/CLK _6792_/D wire3935/A VGND VGND VPWR VPWR _6792_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR clkbuf_2_1_0_mgmt_gpio_in[4]/A
+ sky130_fd_sc_hd__clkbuf_8
X_5743_ _5743_/A _5743_/B VGND VGND VPWR VPWR _5743_/X sky130_fd_sc_hd__or2_1
XFILLER_188_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5674_ _5674_/A1 _5717_/A2 _5673_/X VGND VGND VPWR VPWR _5681_/C sky130_fd_sc_hd__a21o_1
XFILLER_148_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4625_ _4635_/B _4679_/B VGND VGND VPWR VPWR _5177_/A sky130_fd_sc_hd__nor2_1
XFILLER_148_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold500 _6864_/Q VGND VGND VPWR VPWR hold500/X sky130_fd_sc_hd__dlygate4sd3_1
X_4556_ _4556_/A VGND VGND VPWR VPWR _4783_/A sky130_fd_sc_hd__inv_2
XFILLER_116_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold511 _6823_/Q VGND VGND VPWR VPWR hold511/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 _6818_/Q VGND VGND VPWR VPWR hold522/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire4209 wire4210/X VGND VGND VPWR VPWR wire4209/X sky130_fd_sc_hd__clkbuf_1
Xhold533 _7079_/Q VGND VGND VPWR VPWR hold533/X sky130_fd_sc_hd__dlygate4sd3_1
X_3507_ _3536_/B _3507_/B VGND VGND VPWR VPWR _3507_/Y sky130_fd_sc_hd__nor2_1
Xhold544 _7084_/Q VGND VGND VPWR VPWR hold544/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 _6509_/Q VGND VGND VPWR VPWR hold555/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3508 _5308_/A0 VGND VGND VPWR VPWR _5416_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4487_ _4488_/A _4487_/B VGND VGND VPWR VPWR _4530_/B sky130_fd_sc_hd__nand2_1
Xhold566 _7028_/Q VGND VGND VPWR VPWR hold566/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 _6490_/Q VGND VGND VPWR VPWR hold577/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold588 _6995_/Q VGND VGND VPWR VPWR hold588/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6226_ _6521_/Q _6301_/A2 _6301_/B1 _6761_/Q _6223_/X VGND VGND VPWR VPWR _6232_/A
+ sky130_fd_sc_hd__a221o_1
Xwire2807 _5988_/X VGND VGND VPWR VPWR wire2807/X sky130_fd_sc_hd__clkbuf_1
X_3438_ _3438_/A1 wire954/X _3550_/A2 _3438_/B2 wire842/X VGND VGND VPWR VPWR _3446_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold599 _6983_/Q VGND VGND VPWR VPWR hold599/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire2818 _6334_/A2 VGND VGND VPWR VPWR _6274_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_106_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2829 _5822_/A2 VGND VGND VPWR VPWR _5707_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6157_ _7140_/Q _6157_/A2 _6157_/B1 _6157_/B2 _6147_/X VGND VGND VPWR VPWR _6157_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3369_ _6213_/B2 wire922/X _3548_/B1 _6210_/B2 VGND VGND VPWR VPWR _3369_/X sky130_fd_sc_hd__a22o_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5108_ _5108_/A _5108_/B VGND VGND VPWR VPWR _5109_/D sky130_fd_sc_hd__nor2_1
XFILLER_57_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6088_ _6088_/A1 _6088_/A2 _6132_/B1 _6088_/B2 VGND VGND VPWR VPWR _6088_/X sky130_fd_sc_hd__a22o_1
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5039_ _5039_/A _5039_/B _5038_/X VGND VGND VPWR VPWR _5039_/X sky130_fd_sc_hd__or3b_1
XFILLER_73_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length1120 _3777_/B1 VGND VGND VPWR VPWR _3636_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_119_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout3947 wire4022/A VGND VGND VPWR VPWR wire3948/A sky130_fd_sc_hd__buf_2
Xmax_length1175 _3324_/Y VGND VGND VPWR VPWR _3470_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_162_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length1186 _3581_/A2 VGND VGND VPWR VPWR wire1185/A sky130_fd_sc_hd__clkbuf_1
XFILLER_150_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput120 wb_adr_i[29] VGND VGND VPWR VPWR input120/X sky130_fd_sc_hd__clkbuf_1
Xinput131 wb_cyc_i VGND VGND VPWR VPWR wire4278/A sky130_fd_sc_hd__clkbuf_1
Xinput142 wb_dat_i[19] VGND VGND VPWR VPWR _6372_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput153 wb_dat_i[29] VGND VGND VPWR VPWR _6379_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput164 wb_rstn_i VGND VGND VPWR VPWR wire4269/A sky130_fd_sc_hd__clkbuf_1
XFILLER_36_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4410_ _4433_/C _4436_/B VGND VGND VPWR VPWR _5001_/A sky130_fd_sc_hd__and2b_1
XFILLER_126_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5390_ _5489_/A0 hold527/X _5391_/S VGND VGND VPWR VPWR _6966_/D sky130_fd_sc_hd__mux2_1
X_4341_ _4342_/B _4342_/C VGND VGND VPWR VPWR _4341_/X sky130_fd_sc_hd__and2_1
XFILLER_125_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7060_ _7129_/CLK _7060_/D wire4056/A VGND VGND VPWR VPWR _7060_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4272_ hold475/X _5555_/A0 _4275_/S VGND VGND VPWR VPWR _6722_/D sky130_fd_sc_hd__mux2_1
XFILLER_98_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6011_ _6011_/A1 _6073_/A2 _6055_/B1 _6011_/B2 _6010_/X VGND VGND VPWR VPWR _6012_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_97_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3223_ _6933_/Q VGND VGND VPWR VPWR _3223_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6913_ _7064_/CLK _6913_/D wire4045/X VGND VGND VPWR VPWR _6913_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6844_ _6956_/CLK _6844_/D _7137_/RESET_B VGND VGND VPWR VPWR _6844_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6775_ _6775_/CLK _6775_/D fanout3973/X VGND VGND VPWR VPWR _6775_/Q sky130_fd_sc_hd__dfrtp_1
X_3987_ hold718/X _4286_/A0 _3988_/S VGND VGND VPWR VPWR _6485_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5726_ _6063_/A1 _5735_/B1 _5734_/B1 _6064_/A1 VGND VGND VPWR VPWR _5726_/X sky130_fd_sc_hd__a22o_1
XFILLER_109_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5657_ _5657_/A1 _5724_/A2 _5725_/A2 _6031_/B2 VGND VGND VPWR VPWR _5657_/X sky130_fd_sc_hd__a22o_1
XFILLER_163_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4608_ _4792_/A _4797_/A _4607_/X VGND VGND VPWR VPWR _4644_/B sky130_fd_sc_hd__a21o_1
XFILLER_184_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5588_ _5588_/A0 hold650/X _5588_/S VGND VGND VPWR VPWR _7142_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold330 _6834_/Q VGND VGND VPWR VPWR hold330/X sky130_fd_sc_hd__dlygate4sd3_1
X_4539_ _4819_/C _4819_/D VGND VGND VPWR VPWR _4553_/B sky130_fd_sc_hd__and2_1
Xhold341 _6580_/Q VGND VGND VPWR VPWR hold341/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold352 _6752_/Q VGND VGND VPWR VPWR hold352/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire4039 wire4040/X VGND VGND VPWR VPWR wire4039/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3305 wire3306/X VGND VGND VPWR VPWR _4653_/C sky130_fd_sc_hd__clkbuf_1
Xhold363 _6771_/Q VGND VGND VPWR VPWR hold363/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3316 _4585_/X VGND VGND VPWR VPWR _5018_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xhold374 _7124_/Q VGND VGND VPWR VPWR hold374/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3327 _4561_/Y VGND VGND VPWR VPWR _4563_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold385 _7063_/Q VGND VGND VPWR VPWR hold385/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold396 _6523_/Q VGND VGND VPWR VPWR hold396/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3338 _4958_/B1 VGND VGND VPWR VPWR _4694_/A sky130_fd_sc_hd__clkbuf_2
Xwire3349 _4389_/Y VGND VGND VPWR VPWR _4662_/B sky130_fd_sc_hd__clkbuf_2
Xwire2604 _4631_/B VGND VGND VPWR VPWR _5144_/C1 sky130_fd_sc_hd__clkbuf_1
XFILLER_131_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2626 wire2627/X VGND VGND VPWR VPWR _6307_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire2637 _6329_/B1 VGND VGND VPWR VPWR _6314_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_104_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6209_ _6209_/A1 _6209_/A2 _6209_/B1 _6209_/B2 _6208_/X VGND VGND VPWR VPWR _6217_/B
+ sky130_fd_sc_hd__a221o_1
Xwire1903 wire1904/X VGND VGND VPWR VPWR _3535_/A1 sky130_fd_sc_hd__clkbuf_1
X_7189_ _7193_/CLK _7189_/D VGND VGND VPWR VPWR _7189_/Q sky130_fd_sc_hd__dfxtp_1
Xwire2648 wire2649/X VGND VGND VPWR VPWR _6273_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire2659 _6282_/B1 VGND VGND VPWR VPWR _6309_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1914 _6035_/A1 VGND VGND VPWR VPWR _3746_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire1925 wire1926/X VGND VGND VPWR VPWR wire1925/X sky130_fd_sc_hd__clkbuf_1
Xwire1936 hold99/A VGND VGND VPWR VPWR _3389_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1947 _6074_/B2 VGND VGND VPWR VPWR wire1947/X sky130_fd_sc_hd__clkbuf_1
XFILLER_133_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1958 _6919_/Q VGND VGND VPWR VPWR _5811_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_73_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1969 _5779_/B2 VGND VGND VPWR VPWR wire1969/X sky130_fd_sc_hd__clkbuf_1
XFILLER_46_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length853 _3415_/Y VGND VGND VPWR VPWR wire849/A sky130_fd_sc_hd__clkbuf_1
XFILLER_181_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length897 _3335_/Y VGND VGND VPWR VPWR _3597_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_142_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3850 _4436_/A VGND VGND VPWR VPWR _4621_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_122_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3861 wire3862/X VGND VGND VPWR VPWR wire3861/X sky130_fd_sc_hd__clkbuf_1
Xwire3872 input96/X VGND VGND VPWR VPWR wire3872/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3883 input93/X VGND VGND VPWR VPWR wire3883/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3894 wire3895/X VGND VGND VPWR VPWR wire3894/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_71_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7115_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_36_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3910_ _3906_/X _3908_/Y _6565_/Q _3896_/B VGND VGND VPWR VPWR _6565_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4890_ _5174_/A _4890_/B _4890_/C _4890_/D VGND VGND VPWR VPWR _4890_/X sky130_fd_sc_hd__or4_1
XFILLER_44_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3841_ _6545_/Q _3795_/Y _6459_/Q VGND VGND VPWR VPWR _6459_/D sky130_fd_sc_hd__a21o_1
XFILLER_149_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3772_ _3772_/A1 _3526_/Y _3767_/X _3769_/X _3771_/X VGND VGND VPWR VPWR _3789_/B
+ sky130_fd_sc_hd__a2111o_1
X_6560_ _6811_/CLK _6560_/D _6430_/A VGND VGND VPWR VPWR _6560_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5511_ _5511_/A _5511_/B VGND VGND VPWR VPWR _5519_/S sky130_fd_sc_hd__nand2_1
XFILLER_145_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6491_ _6825_/CLK _6491_/D _6495_/SET_B VGND VGND VPWR VPWR _6491_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_172_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5442_ _5442_/A0 hold182/X _5442_/S VGND VGND VPWR VPWR _7012_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5373_ _5586_/A0 hold603/X _5375_/S VGND VGND VPWR VPWR _6951_/D sky130_fd_sc_hd__mux2_1
XFILLER_126_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_24_csclk _6579_/CLK VGND VGND VPWR VPWR _7111_/CLK sky130_fd_sc_hd__clkbuf_16
X_4324_ _4324_/A _4324_/B VGND VGND VPWR VPWR _4328_/S sky130_fd_sc_hd__and2_1
XFILLER_114_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7112_ _7112_/CLK _7112_/D _7112_/SET_B VGND VGND VPWR VPWR _7112_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_99_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7043_ _7135_/CLK _7043_/D wire4090/X VGND VGND VPWR VPWR hold94/A sky130_fd_sc_hd__dfstp_1
XFILLER_87_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4255_ hold146/X _4255_/A1 _4257_/S VGND VGND VPWR VPWR _6708_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3206_ _3206_/A VGND VGND VPWR VPWR _3206_/Y sky130_fd_sc_hd__inv_2
X_4186_ _6644_/Q wire370/X _4188_/S VGND VGND VPWR VPWR _6644_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_39_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7132_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_67_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_1_0_csclk clkbuf_3_1_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_1_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_94_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6827_ _7130_/CLK hold39/X wire4058/X VGND VGND VPWR VPWR _6827_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire507 _5285_/S VGND VGND VPWR VPWR _5282_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_6758_ _6775_/CLK _6758_/D wire3978/X VGND VGND VPWR VPWR _6758_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_149_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire518 _5232_/Y VGND VGND VPWR VPWR _5240_/S sky130_fd_sc_hd__clkbuf_4
Xwire529 wire530/X VGND VGND VPWR VPWR wire529/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5709_ _6842_/Q _5709_/A2 _5708_/X wire997/X _6047_/A1 VGND VGND VPWR VPWR _5709_/X
+ sky130_fd_sc_hd__o221a_1
X_6689_ _7093_/CLK _6689_/D wire3959/A VGND VGND VPWR VPWR _6689_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_136_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3102 wire3102/A VGND VGND VPWR VPWR _5951_/A2 sky130_fd_sc_hd__clkbuf_1
Xhold160 _4177_/X VGND VGND VPWR VPWR _6636_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 _6915_/Q VGND VGND VPWR VPWR hold171/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3113 _5775_/A2 VGND VGND VPWR VPWR _5735_/A2 sky130_fd_sc_hd__clkbuf_2
Xhold182 _7012_/Q VGND VGND VPWR VPWR hold182/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3124 _5780_/A2 VGND VGND VPWR VPWR _5712_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3135 _5790_/A2 VGND VGND VPWR VPWR _5725_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold193 _6885_/Q VGND VGND VPWR VPWR hold193/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire2401 _6513_/Q VGND VGND VPWR VPWR _5908_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3146 _5855_/A2 VGND VGND VPWR VPWR _5758_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2412 _5900_/B2 VGND VGND VPWR VPWR _6252_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2423 wire2424/X VGND VGND VPWR VPWR wire2423/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3168 _4676_/A2 VGND VGND VPWR VPWR _4683_/B sky130_fd_sc_hd__clkbuf_2
Xwire2434 _6497_/Q VGND VGND VPWR VPWR wire2434/X sky130_fd_sc_hd__clkbuf_1
Xwire3179 _4655_/B VGND VGND VPWR VPWR _4659_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1700 _7040_/Q VGND VGND VPWR VPWR _3394_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2445 _6488_/Q VGND VGND VPWR VPWR wire2445/X sky130_fd_sc_hd__clkbuf_2
XFILLER_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1711 _3210_/A VGND VGND VPWR VPWR _5763_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2456 wire2457/X VGND VGND VPWR VPWR _6206_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_144_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1722 _3769_/B2 VGND VGND VPWR VPWR wire1722/X sky130_fd_sc_hd__clkbuf_1
XFILLER_93_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2467 _6330_/B1 VGND VGND VPWR VPWR _6286_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1733 hold92/A VGND VGND VPWR VPWR _6108_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire2478 wire2478/A VGND VGND VPWR VPWR _6322_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire2489 _6023_/D VGND VGND VPWR VPWR wire2489/X sky130_fd_sc_hd__clkbuf_1
Xwire1744 _7026_/Q VGND VGND VPWR VPWR _5701_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1755 wire1756/X VGND VGND VPWR VPWR _6107_/B2 sky130_fd_sc_hd__clkbuf_1
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1766 _3736_/B2 VGND VGND VPWR VPWR wire1766/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1777 _7013_/Q VGND VGND VPWR VPWR wire1777/X sky130_fd_sc_hd__clkbuf_1
XFILLER_73_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1788 wire1789/X VGND VGND VPWR VPWR _6202_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire1799 wire1800/X VGND VGND VPWR VPWR _3214_/A sky130_fd_sc_hd__clkbuf_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_671 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout4297 wire4302/A VGND VGND VPWR VPWR _4570_/D sky130_fd_sc_hd__buf_6
XFILLER_111_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3680 wire3681/X VGND VGND VPWR VPWR _5872_/B sky130_fd_sc_hd__clkbuf_1
X_4040_ _4040_/A _6392_/B VGND VGND VPWR VPWR _4045_/S sky130_fd_sc_hd__nand2_2
XFILLER_110_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2990 _5760_/B1 VGND VGND VPWR VPWR _5748_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_77_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5991_ _6019_/A _6039_/C _6030_/C VGND VGND VPWR VPWR _6029_/B sky130_fd_sc_hd__and3b_1
XFILLER_52_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4942_ _4942_/A _4942_/B VGND VGND VPWR VPWR _5060_/B sky130_fd_sc_hd__nand2_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4873_ _5050_/A _5050_/B VGND VGND VPWR VPWR _4873_/Y sky130_fd_sc_hd__nand2_1
XFILLER_178_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6612_ _6702_/CLK _6612_/D _6440_/A VGND VGND VPWR VPWR _6612_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3824_ hold66/A _3820_/A _3816_/Y _3823_/X VGND VGND VPWR VPWR _3824_/X sky130_fd_sc_hd__a22o_1
XFILLER_32_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length2409 _6302_/A1 VGND VGND VPWR VPWR _5931_/B2 sky130_fd_sc_hd__clkbuf_1
X_6543_ _3945_/A1 _6543_/D _6431_/X VGND VGND VPWR VPWR _6543_/Q sky130_fd_sc_hd__dfrtp_2
X_3755_ _3755_/A _3755_/B _3755_/C _3755_/D VGND VGND VPWR VPWR _3790_/B sky130_fd_sc_hd__or4_1
XFILLER_9_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3686_ _5432_/A1 _3763_/B1 _3686_/B1 _3686_/B2 VGND VGND VPWR VPWR _3686_/X sky130_fd_sc_hd__a22o_1
X_6474_ _6824_/CLK _6474_/D _6483_/SET_B VGND VGND VPWR VPWR _6474_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_133_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5425_ _5539_/A1 hold509/X _5429_/S VGND VGND VPWR VPWR _6997_/D sky130_fd_sc_hd__mux2_1
Xoutput210 _3227_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[7] sky130_fd_sc_hd__buf_12
Xoutput221 _6547_/Q VGND VGND VPWR VPWR mgmt_gpio_out[17] sky130_fd_sc_hd__buf_12
XFILLER_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput232 _6829_/Q VGND VGND VPWR VPWR mgmt_gpio_out[27] sky130_fd_sc_hd__buf_12
XFILLER_161_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput243 wire1490/X VGND VGND VPWR VPWR mgmt_gpio_out[37] sky130_fd_sc_hd__buf_12
XFILLER_161_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput254 _3944_/Y VGND VGND VPWR VPWR pad_flash_csb_oeb sky130_fd_sc_hd__buf_12
X_5356_ _5356_/A0 hold684/X _5356_/S VGND VGND VPWR VPWR _6936_/D sky130_fd_sc_hd__mux2_1
Xoutput265 _6792_/Q VGND VGND VPWR VPWR pll_dco_ena sky130_fd_sc_hd__buf_12
Xoutput276 _6484_/Q VGND VGND VPWR VPWR pll_trim[10] sky130_fd_sc_hd__buf_12
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput287 _6478_/Q VGND VGND VPWR VPWR pll_trim[20] sky130_fd_sc_hd__buf_12
Xoutput298 _6497_/Q VGND VGND VPWR VPWR pll_trim[7] sky130_fd_sc_hd__buf_12
X_4307_ _5212_/C hold351/X _4311_/S VGND VGND VPWR VPWR _6751_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5287_ _5581_/A0 hold318/X _5291_/S VGND VGND VPWR VPWR _6874_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1007 wire1008/X VGND VGND VPWR VPWR _5948_/S sky130_fd_sc_hd__clkbuf_2
Xwire1018 wire1019/X VGND VGND VPWR VPWR wire1018/X sky130_fd_sc_hd__clkbuf_2
X_7026_ _7027_/CLK _7026_/D fanout3976/X VGND VGND VPWR VPWR _7026_/Q sky130_fd_sc_hd__dfstp_1
X_4238_ _4250_/A0 hold334/X _4239_/S VGND VGND VPWR VPWR _6684_/D sky130_fd_sc_hd__mux2_1
Xwire1029 _4222_/A VGND VGND VPWR VPWR _3720_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4169_ _6629_/Q wire366/X _4173_/S VGND VGND VPWR VPWR _6629_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3600 _5477_/A0 VGND VGND VPWR VPWR _5522_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_128_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length3633 _4235_/A0 VGND VGND VPWR VPWR _4211_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_139_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length3644 _5554_/A0 VGND VGND VPWR VPWR _5440_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_183_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire359 _3790_/X VGND VGND VPWR VPWR wire359/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2220 _6717_/Q VGND VGND VPWR VPWR _6258_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire2231 _6710_/Q VGND VGND VPWR VPWR _6327_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire2242 _6704_/Q VGND VGND VPWR VPWR _3574_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire2253 _6687_/Q VGND VGND VPWR VPWR _6262_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2264 _4225_/A1 VGND VGND VPWR VPWR _6287_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1530 _7209_/Q VGND VGND VPWR VPWR _6273_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2275 _6670_/Q VGND VGND VPWR VPWR wire2275/X sky130_fd_sc_hd__clkbuf_1
Xwire1541 wire1542/X VGND VGND VPWR VPWR _3597_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_93_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1552 wire1553/X VGND VGND VPWR VPWR _3199_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2297 wire2298/X VGND VGND VPWR VPWR _3576_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire1563 wire1564/X VGND VGND VPWR VPWR _3578_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_171_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1585 wire1586/X VGND VGND VPWR VPWR _6117_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_46_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7159__4309 VGND VGND VPWR VPWR _7159_/D _7159__4309/LO sky130_fd_sc_hd__conb_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3540_ _3540_/A1 _3540_/A2 wire902/X _3540_/B2 wire561/X VGND VGND VPWR VPWR _3541_/D
+ sky130_fd_sc_hd__a221o_1
Xwire860 _3343_/Y VGND VGND VPWR VPWR wire860/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire871 wire872/X VGND VGND VPWR VPWR wire871/X sky130_fd_sc_hd__dlymetal6s2s_1
Xwire882 wire886/X VGND VGND VPWR VPWR wire882/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_142_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3471_ _3507_/B _3528_/B VGND VGND VPWR VPWR _4318_/A sky130_fd_sc_hd__nor2_1
XFILLER_115_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout4050 wire4066/A VGND VGND VPWR VPWR wire4052/A sky130_fd_sc_hd__buf_6
XFILLER_170_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5210_ _5210_/A _5210_/B VGND VGND VPWR VPWR _5211_/S sky130_fd_sc_hd__nand2_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6190_ _6190_/A1 _6212_/A2 _6190_/B1 _6976_/Q VGND VGND VPWR VPWR _6190_/X sky130_fd_sc_hd__a22o_1
XFILLER_97_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout3371 wire3387/A VGND VGND VPWR VPWR _5561_/A0 sky130_fd_sc_hd__buf_6
X_5141_ _4872_/A _4728_/Y _4916_/A _4618_/C VGND VGND VPWR VPWR _5141_/X sky130_fd_sc_hd__o211a_1
XFILLER_69_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5072_ _4645_/X _4665_/B _5072_/A3 _4611_/A VGND VGND VPWR VPWR _5072_/X sky130_fd_sc_hd__a31o_1
XFILLER_56_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4023_ hold313/X _5530_/A1 _4027_/S VGND VGND VPWR VPWR _4023_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5974_ _7157_/Q _7158_/Q VGND VGND VPWR VPWR _6020_/C sky130_fd_sc_hd__nor2_2
XFILLER_80_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4925_ _5095_/A _4925_/B _4924_/Y VGND VGND VPWR VPWR _4925_/X sky130_fd_sc_hd__or3b_1
XFILLER_80_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4856_ _4759_/A _4395_/Y _4502_/A _4833_/Y VGND VGND VPWR VPWR _4857_/D sky130_fd_sc_hd__a211oi_1
XFILLER_193_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3807_ hold66/A _3807_/B hold81/A VGND VGND VPWR VPWR _3823_/B sky130_fd_sc_hd__and3_1
XFILLER_20_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4787_ _4718_/B _4689_/B _4770_/C VGND VGND VPWR VPWR _4982_/B sky130_fd_sc_hd__o21bai_1
XFILLER_119_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6526_ _7090_/CLK _6526_/D wire3935/X VGND VGND VPWR VPWR _6526_/Q sky130_fd_sc_hd__dfrtp_1
X_3738_ _6858_/Q wire936/X _3738_/B1 _6004_/B2 VGND VGND VPWR VPWR _3738_/X sky130_fd_sc_hd__a22o_1
XFILLER_109_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6457_ _6545_/CLK _6457_/D _6412_/X VGND VGND VPWR VPWR _6457_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3669_ _3669_/A _3669_/B _3669_/C _3669_/D VGND VGND VPWR VPWR _3723_/A sky130_fd_sc_hd__or4_1
XFILLER_118_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5408_ _5540_/A1 hold558/X _5408_/S VGND VGND VPWR VPWR _6982_/D sky130_fd_sc_hd__mux2_1
XFILLER_192_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6388_ _4228_/C _6357_/A _6358_/B _4228_/B VGND VGND VPWR VPWR _6388_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5339_ _5339_/A0 hold539/X _5339_/S VGND VGND VPWR VPWR _6921_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7009_ _7080_/CLK _7009_/D wire3992/X VGND VGND VPWR VPWR _7009_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_75_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2050 _3571_/A1 VGND VGND VPWR VPWR wire2050/X sky130_fd_sc_hd__clkbuf_1
XFILLER_182_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2061 _6863_/Q VGND VGND VPWR VPWR _6162_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire2072 _6857_/Q VGND VGND VPWR VPWR wire2072/X sky130_fd_sc_hd__clkbuf_1
XFILLER_66_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2083 _5263_/A1 VGND VGND VPWR VPWR wire2083/X sky130_fd_sc_hd__clkbuf_1
Xwire2094 wire2095/X VGND VGND VPWR VPWR _3233_/A sky130_fd_sc_hd__clkbuf_2
Xwire1360 wire1361/X VGND VGND VPWR VPWR wire1360/X sky130_fd_sc_hd__clkbuf_1
Xwire1371 _3510_/B VGND VGND VPWR VPWR _3482_/B sky130_fd_sc_hd__clkbuf_1
Xwire1382 hold168/X VGND VGND VPWR VPWR _3512_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1393 _3285_/Y VGND VGND VPWR VPWR _3322_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4710_ _4848_/A1 _4677_/B _4710_/B1 _4710_/B2 _4709_/X VGND VGND VPWR VPWR _4710_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5690_ _5705_/A _5705_/B _5703_/B VGND VGND VPWR VPWR _5690_/X sky130_fd_sc_hd__and3_1
X_4641_ _4639_/A _4624_/B _4710_/B1 _4799_/B1 _4640_/X VGND VGND VPWR VPWR _4642_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_30_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4572_ _4981_/A _4981_/B _4571_/X VGND VGND VPWR VPWR _4572_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_128_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold704 _7095_/Q VGND VGND VPWR VPWR hold704/X sky130_fd_sc_hd__dlygate4sd3_1
X_6311_ _6311_/A1 _6340_/A2 _6337_/B1 _6311_/B2 _6310_/X VGND VGND VPWR VPWR _6315_/B
+ sky130_fd_sc_hd__a221o_1
Xhold715 _6475_/Q VGND VGND VPWR VPWR hold715/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire690 _5357_/S VGND VGND VPWR VPWR _5356_/S sky130_fd_sc_hd__clkbuf_1
X_3523_ _3523_/A1 _3698_/A2 wire920/A _5775_/A1 _3522_/X VGND VGND VPWR VPWR _3524_/D
+ sky130_fd_sc_hd__a221o_1
Xhold726 _3967_/X VGND VGND VPWR VPWR hold726/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6242_ _6316_/A _6242_/B _6242_/C _6242_/D VGND VGND VPWR VPWR _6242_/X sky130_fd_sc_hd__or4_1
X_3454_ _3528_/B _3454_/B VGND VGND VPWR VPWR _3454_/Y sky130_fd_sc_hd__nor2_1
XFILLER_143_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3385_ _3385_/A1 _5511_/A _5430_/A _7008_/Q VGND VGND VPWR VPWR _3385_/X sky130_fd_sc_hd__a22o_1
X_6173_ _6968_/Q _6173_/A2 _6173_/B1 _6173_/B2 _6172_/X VGND VGND VPWR VPWR _6173_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_97_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout3190 _4718_/B VGND VGND VPWR VPWR _4976_/A1 sky130_fd_sc_hd__buf_6
X_5124_ _5124_/A _5124_/B _5124_/C _4708_/B VGND VGND VPWR VPWR _5125_/B sky130_fd_sc_hd__or4b_1
XFILLER_57_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5055_ _5126_/B _5162_/B _5126_/C _5162_/C VGND VGND VPWR VPWR _5067_/B sky130_fd_sc_hd__or4_1
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4006_ _5585_/A0 hold259/X _4007_/S VGND VGND VPWR VPWR _6502_/D sky130_fd_sc_hd__mux2_1
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5957_ _5957_/A _5957_/B _5957_/C _5957_/D VGND VGND VPWR VPWR _5957_/X sky130_fd_sc_hd__or4_1
XFILLER_111_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4908_ _4958_/B1 _4913_/B1 _4630_/A _5152_/A1 VGND VGND VPWR VPWR _4915_/C sky130_fd_sc_hd__o22ai_1
X_5888_ _6264_/B2 _5888_/A2 _5887_/X VGND VGND VPWR VPWR _5891_/C sky130_fd_sc_hd__a21o_1
XFILLER_139_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4839_ _4839_/A _4839_/B VGND VGND VPWR VPWR _5127_/B sky130_fd_sc_hd__nor2_1
XFILLER_193_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length2003 _5758_/A1 VGND VGND VPWR VPWR _6114_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_193_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6509_ _6701_/CLK _6509_/D _6429_/A VGND VGND VPWR VPWR _6509_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold20 hold20/A VGND VGND VPWR VPWR hold20/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold31 hold31/A VGND VGND VPWR VPWR hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A VGND VGND VPWR VPWR hold42/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold53 hold53/A VGND VGND VPWR VPWR hold53/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold64 hold64/A VGND VGND VPWR VPWR hold64/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A VGND VGND VPWR VPWR hold75/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 hold86/A VGND VGND VPWR VPWR hold86/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold97 hold97/A VGND VGND VPWR VPWR hold97/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_6 mgmt_gpio_in[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1190 wire1191/X VGND VGND VPWR VPWR _3684_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_35_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6860_ _7129_/CLK _6860_/D wire4056/X VGND VGND VPWR VPWR _6860_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5811_ _5811_/A1 _5811_/A2 _5811_/B1 _7079_/Q VGND VGND VPWR VPWR _5811_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6791_ _6811_/CLK _6791_/D wire3935/A VGND VGND VPWR VPWR _6791_/Q sky130_fd_sc_hd__dfrtp_1
X_5742_ _7012_/Q _5762_/B1 _5742_/B1 _5742_/B2 _5742_/C1 VGND VGND VPWR VPWR _5750_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_188_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5673_ _5673_/A1 _5715_/A2 _5745_/A2 _5673_/B2 VGND VGND VPWR VPWR _5673_/X sky130_fd_sc_hd__a22o_1
XFILLER_163_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4624_ _4661_/B _4624_/B VGND VGND VPWR VPWR _4679_/B sky130_fd_sc_hd__or2_4
XFILLER_148_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold501 _6706_/Q VGND VGND VPWR VPWR hold501/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4555_ _4802_/B _4802_/C VGND VGND VPWR VPWR _4556_/A sky130_fd_sc_hd__nor2_1
Xhold512 _6593_/Q VGND VGND VPWR VPWR hold512/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 _6816_/Q VGND VGND VPWR VPWR hold523/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 _6977_/Q VGND VGND VPWR VPWR hold534/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 _6508_/Q VGND VGND VPWR VPWR hold545/X sky130_fd_sc_hd__dlygate4sd3_1
X_3506_ _3506_/A1 wire937/X _3502_/Y _6320_/B2 wire564/X VGND VGND VPWR VPWR _3506_/X
+ sky130_fd_sc_hd__a221o_1
Xhold556 _7092_/Q VGND VGND VPWR VPWR hold556/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3509 _5506_/A0 VGND VGND VPWR VPWR _5308_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
X_4486_ _4486_/A _4942_/A VGND VGND VPWR VPWR _5065_/A sky130_fd_sc_hd__nor2_1
Xhold567 _7101_/Q VGND VGND VPWR VPWR hold567/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold578 _6901_/Q VGND VGND VPWR VPWR hold578/X sky130_fd_sc_hd__dlygate4sd3_1
X_6225_ _6225_/A1 _6225_/A2 _6225_/B1 _6225_/B2 VGND VGND VPWR VPWR _6241_/B sky130_fd_sc_hd__a22o_1
Xhold589 _6590_/Q VGND VGND VPWR VPWR hold589/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3437_ _3437_/A1 _3437_/A2 wire885/X _3437_/B2 wire571/X VGND VGND VPWR VPWR _3446_/A
+ sky130_fd_sc_hd__a221o_1
Xwire2808 _6337_/A2 VGND VGND VPWR VPWR _6262_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire2819 wire2819/A VGND VGND VPWR VPWR _6334_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_106_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3368_ _6205_/B2 _3368_/A2 wire878/X _6215_/A1 _3346_/X VGND VGND VPWR VPWR _3371_/C
+ sky130_fd_sc_hd__a221o_1
X_6156_ _6156_/A _6156_/B _6156_/C _6156_/D VGND VGND VPWR VPWR _6156_/X sky130_fd_sc_hd__or4_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5107_ _5107_/A _5107_/B _5107_/C _4676_/X VGND VGND VPWR VPWR _5178_/B sky130_fd_sc_hd__or4b_1
X_3299_ _3303_/A hold84/X VGND VGND VPWR VPWR hold85/A sky130_fd_sc_hd__nand2_2
XFILLER_85_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6087_ _6087_/A1 _6087_/A2 _6087_/B1 _6956_/Q _6086_/X VGND VGND VPWR VPWR _6094_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_111_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5038_ _4396_/X _4668_/X _4836_/Y _4453_/A VGND VGND VPWR VPWR _5038_/X sky130_fd_sc_hd__a31o_1
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6989_ _6989_/CLK _6989_/D wire3995/X VGND VGND VPWR VPWR _6989_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length1132 _3332_/Y VGND VGND VPWR VPWR wire1130/A sky130_fd_sc_hd__clkbuf_1
XFILLER_162_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout3937 wire3948/A VGND VGND VPWR VPWR _3946_/B sky130_fd_sc_hd__buf_6
XFILLER_150_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput110 wb_adr_i[1] VGND VGND VPWR VPWR _4570_/A sky130_fd_sc_hd__clkbuf_2
Xinput121 wb_adr_i[2] VGND VGND VPWR VPWR wire4302/A sky130_fd_sc_hd__clkbuf_1
Xinput132 wb_dat_i[0] VGND VGND VPWR VPWR _6363_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput143 wb_dat_i[1] VGND VGND VPWR VPWR _6367_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput154 wb_dat_i[2] VGND VGND VPWR VPWR _6370_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput165 wb_sel_i[0] VGND VGND VPWR VPWR _6360_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_17_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4340_ _4348_/A _4348_/B _4348_/C VGND VGND VPWR VPWR _4404_/B sky130_fd_sc_hd__and3_1
XFILLER_126_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4271_ hold372/X _5224_/A0 _4275_/S VGND VGND VPWR VPWR _6721_/D sky130_fd_sc_hd__mux2_1
X_3222_ _3222_/A VGND VGND VPWR VPWR _3222_/Y sky130_fd_sc_hd__inv_2
X_6010_ _6010_/A1 _6067_/A2 _6057_/A2 _6010_/B2 VGND VGND VPWR VPWR _6010_/X sky130_fd_sc_hd__a22o_1
XFILLER_140_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_588 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6912_ _7064_/CLK _6912_/D wire4045/X VGND VGND VPWR VPWR _6912_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_82_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6843_ _6956_/CLK _6843_/D wire4039/X VGND VGND VPWR VPWR _6843_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_90_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6774_ _7036_/CLK _6774_/D fanout3973/X VGND VGND VPWR VPWR _6774_/Q sky130_fd_sc_hd__dfrtp_1
X_3986_ hold717/X _4333_/A0 _3988_/S VGND VGND VPWR VPWR _6484_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5725_ _6060_/B2 _5725_/A2 _5735_/A2 _6064_/B2 _5724_/X VGND VGND VPWR VPWR _5728_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5656_ _7152_/Q _5706_/B _5703_/B VGND VGND VPWR VPWR _5656_/X sky130_fd_sc_hd__and3_1
XFILLER_175_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4607_ _4981_/C _4607_/B _4778_/A _4607_/D VGND VGND VPWR VPWR _4607_/X sky130_fd_sc_hd__and4b_1
X_5587_ _5587_/A0 hold649/X _5587_/S VGND VGND VPWR VPWR _7141_/D sky130_fd_sc_hd__mux2_1
Xwire4007 wire4007/A VGND VGND VPWR VPWR wire4007/X sky130_fd_sc_hd__clkbuf_2
Xhold320 _6978_/Q VGND VGND VPWR VPWR hold320/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4018 wire4018/A VGND VGND VPWR VPWR wire4018/X sky130_fd_sc_hd__clkbuf_1
Xhold331 _6670_/Q VGND VGND VPWR VPWR hold331/X sky130_fd_sc_hd__dlygate4sd3_1
X_4538_ _4538_/A _4538_/B VGND VGND VPWR VPWR _4538_/Y sky130_fd_sc_hd__nand2_1
Xwire4029 wire4029/A VGND VGND VPWR VPWR wire4029/X sky130_fd_sc_hd__clkbuf_2
XFILLER_132_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold342 _6922_/Q VGND VGND VPWR VPWR hold342/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 _6754_/Q VGND VGND VPWR VPWR hold353/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3306 _4645_/B VGND VGND VPWR VPWR wire3306/X sky130_fd_sc_hd__clkbuf_1
Xhold364 _6772_/Q VGND VGND VPWR VPWR hold364/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold375 _6820_/Q VGND VGND VPWR VPWR hold375/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3317 _4623_/A VGND VGND VPWR VPWR _4784_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3328 _5169_/A1 VGND VGND VPWR VPWR _4683_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold386 _6572_/Q VGND VGND VPWR VPWR hold386/X sky130_fd_sc_hd__dlygate4sd3_1
X_4469_ _4474_/A _4832_/B VGND VGND VPWR VPWR _4839_/A sky130_fd_sc_hd__or2_1
XFILLER_77_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3339 _4958_/B1 VGND VGND VPWR VPWR _4848_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold397 _6763_/Q VGND VGND VPWR VPWR hold397/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire2605 _4639_/A VGND VGND VPWR VPWR _4633_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_104_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2616 _6339_/B1 VGND VGND VPWR VPWR _6312_/B1 sky130_fd_sc_hd__clkbuf_2
X_6208_ _7142_/Q _6208_/A2 _6208_/B1 _6208_/B2 _6208_/C1 VGND VGND VPWR VPWR _6208_/X
+ sky130_fd_sc_hd__a221o_1
Xwire2627 _6039_/X VGND VGND VPWR VPWR wire2627/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2638 wire2639/X VGND VGND VPWR VPWR _6329_/B1 sky130_fd_sc_hd__clkbuf_2
X_7188_ _7206_/CLK _7188_/D _4189_/B VGND VGND VPWR VPWR _7188_/Q sky130_fd_sc_hd__dfrtp_1
Xwire2649 _6033_/X VGND VGND VPWR VPWR wire2649/X sky130_fd_sc_hd__clkbuf_1
Xwire1904 _5780_/B2 VGND VGND VPWR VPWR wire1904/X sky130_fd_sc_hd__clkbuf_1
Xwire1915 _6938_/Q VGND VGND VPWR VPWR _6035_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_133_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1926 wire1927/X VGND VGND VPWR VPWR wire1926/X sky130_fd_sc_hd__clkbuf_1
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6139_ _6139_/A1 _6139_/A2 _6139_/B1 _6886_/Q _6138_/X VGND VGND VPWR VPWR _6142_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1937 _6927_/Q VGND VGND VPWR VPWR _5801_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_46_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1948 wire1949/X VGND VGND VPWR VPWR _6074_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire1959 _6918_/Q VGND VGND VPWR VPWR _5776_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_85_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length821 hold30/X VGND VGND VPWR VPWR wire820/A sky130_fd_sc_hd__clkbuf_1
XFILLER_158_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_5_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _6702_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_174_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3840 _4070_/A2 VGND VGND VPWR VPWR wire3840/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3862 input98/X VGND VGND VPWR VPWR wire3862/X sky130_fd_sc_hd__clkbuf_1
Xwire3873 wire3874/X VGND VGND VPWR VPWR _3585_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire3884 wire3885/X VGND VGND VPWR VPWR _3920_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire3895 wire3896/X VGND VGND VPWR VPWR wire3895/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3840_ _6460_/Q _6445_/Q _3840_/S VGND VGND VPWR VPWR _6460_/D sky130_fd_sc_hd__mux2_1
XFILLER_189_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3771_ _3771_/A1 _3771_/A2 _3771_/B1 _6222_/A _3770_/X VGND VGND VPWR VPWR _3771_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5510_ _5552_/A0 hold559/X _5510_/S VGND VGND VPWR VPWR _7073_/D sky130_fd_sc_hd__mux2_1
XFILLER_157_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6490_ _6803_/CLK _6490_/D _6495_/SET_B VGND VGND VPWR VPWR _6490_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_9_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5441_ _5573_/A0 hold183/X _5441_/S VGND VGND VPWR VPWR _7011_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5372_ _5489_/A0 hold453/X _5372_/S VGND VGND VPWR VPWR _6950_/D sky130_fd_sc_hd__mux2_1
X_7111_ _7111_/CLK _7111_/D _6401_/A VGND VGND VPWR VPWR _7111_/Q sky130_fd_sc_hd__dfstp_1
X_4323_ hold390/X _4323_/A1 _4323_/S VGND VGND VPWR VPWR _6765_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7042_ _7135_/CLK _7042_/D _7042_/SET_B VGND VGND VPWR VPWR _7042_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_99_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4254_ hold674/X _5531_/A1 _4257_/S VGND VGND VPWR VPWR _6707_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3205_ _3205_/A VGND VGND VPWR VPWR _3205_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4185_ _6643_/Q _6353_/A1 _4188_/S VGND VGND VPWR VPWR _6643_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6826_ _7130_/CLK _6826_/D wire4058/X VGND VGND VPWR VPWR _6826_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6757_ _6761_/CLK _6757_/D wire4019/X VGND VGND VPWR VPWR _6757_/Q sky130_fd_sc_hd__dfrtp_1
Xwire508 wire508/A VGND VGND VPWR VPWR _5274_/S sky130_fd_sc_hd__clkbuf_1
X_3969_ hold35/X hold729/X _3979_/S VGND VGND VPWR VPWR hold36/A sky130_fd_sc_hd__mux2_1
Xwire519 _5145_/X VGND VGND VPWR VPWR _5170_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3837 _6437_/B VGND VGND VPWR VPWR _6431_/B sky130_fd_sc_hd__clkbuf_2
X_5708_ _5708_/A _5708_/B _5708_/C _5708_/D VGND VGND VPWR VPWR _5708_/X sky130_fd_sc_hd__or4_1
XFILLER_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6688_ _6705_/CLK _6688_/D wire3959/A VGND VGND VPWR VPWR _6688_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_176_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5639_ _5634_/Y _5638_/Y _5643_/B VGND VGND VPWR VPWR _7157_/D sky130_fd_sc_hd__a21oi_1
XFILLER_136_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold150 _5528_/X VGND VGND VPWR VPWR _7089_/D sky130_fd_sc_hd__dlygate4sd3_1
Xwire3103 _5739_/B1 VGND VGND VPWR VPWR _5887_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_105_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3114 wire3119/X VGND VGND VPWR VPWR _5775_/A2 sky130_fd_sc_hd__clkbuf_1
Xhold161 _6972_/Q VGND VGND VPWR VPWR hold161/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 _6701_/Q VGND VGND VPWR VPWR hold172/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 _7011_/Q VGND VGND VPWR VPWR hold183/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3125 _5802_/A2 VGND VGND VPWR VPWR _5780_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire3136 _5761_/A2 VGND VGND VPWR VPWR _5790_/A2 sky130_fd_sc_hd__clkbuf_1
Xhold194 _6914_/Q VGND VGND VPWR VPWR hold194/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire2402 wire2403/X VGND VGND VPWR VPWR _6250_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire3147 _5812_/A2 VGND VGND VPWR VPWR _5724_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_144_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3158 _5642_/X VGND VGND VPWR VPWR _5995_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire2413 _6507_/Q VGND VGND VPWR VPWR _5900_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire2424 _6115_/A1 VGND VGND VPWR VPWR wire2424/X sky130_fd_sc_hd__clkbuf_1
Xwire3169 _4662_/Y VGND VGND VPWR VPWR _4676_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire2435 wire2436/X VGND VGND VPWR VPWR _3398_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire1701 _7039_/Q VGND VGND VPWR VPWR _5800_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1712 hold189/X VGND VGND VPWR VPWR _3210_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2457 _6038_/Y VGND VGND VPWR VPWR wire2457/X sky130_fd_sc_hd__clkbuf_1
Xwire1723 _7034_/Q VGND VGND VPWR VPWR _3769_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire2468 wire2469/X VGND VGND VPWR VPWR _6330_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire1734 wire1735/X VGND VGND VPWR VPWR _6093_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire1745 _7024_/Q VGND VGND VPWR VPWR _6176_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_86_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1756 wire1757/X VGND VGND VPWR VPWR wire1756/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1767 _7018_/Q VGND VGND VPWR VPWR _3736_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1778 wire1779/X VGND VGND VPWR VPWR _3640_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_58_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1789 _7009_/Q VGND VGND VPWR VPWR wire1789/X sky130_fd_sc_hd__clkbuf_1
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length673 _5404_/S VGND VGND VPWR VPWR _5406_/S sky130_fd_sc_hd__clkbuf_1
XFILLER_127_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length695 _5353_/S VGND VGND VPWR VPWR wire694/A sky130_fd_sc_hd__clkbuf_1
XFILLER_185_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout3542 wire3555/A VGND VGND VPWR VPWR _4162_/A1 sky130_fd_sc_hd__buf_6
XFILLER_69_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout3597 hold38/A VGND VGND VPWR VPWR _5477_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_150_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3670 wire3671/X VGND VGND VPWR VPWR wire3670/X sky130_fd_sc_hd__clkbuf_2
Xwire3681 _5683_/A VGND VGND VPWR VPWR wire3681/X sky130_fd_sc_hd__clkbuf_1
Xwire3692 _6342_/C1 VGND VGND VPWR VPWR _6268_/C1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2980 _5781_/B1 VGND VGND VPWR VPWR _5737_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2991 _5714_/A2 VGND VGND VPWR VPWR _5684_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5990_ _5990_/A1 _5990_/A2 _5990_/B1 _5990_/B2 VGND VGND VPWR VPWR _5990_/X sky130_fd_sc_hd__a22o_1
XFILLER_91_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4941_ _4459_/B _4446_/Y _4843_/B _4940_/Y VGND VGND VPWR VPWR _5126_/C sky130_fd_sc_hd__a211o_1
XFILLER_33_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4872_ _4872_/A _4872_/B VGND VGND VPWR VPWR _4894_/C sky130_fd_sc_hd__nor2_1
XFILLER_33_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6611_ _6705_/CLK _6611_/D wire3959/X VGND VGND VPWR VPWR _6611_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_178_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3823_ hold24/A _3823_/B VGND VGND VPWR VPWR _3823_/X sky130_fd_sc_hd__or2_1
XFILLER_60_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6542_ _6545_/CLK _6542_/D _6430_/X VGND VGND VPWR VPWR _6542_/Q sky130_fd_sc_hd__dfrtp_1
X_3754_ _3754_/A1 _3310_/Y _3754_/B1 _3754_/B2 _3738_/X VGND VGND VPWR VPWR _3755_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_192_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6473_ _6545_/CLK _6473_/D _6428_/X VGND VGND VPWR VPWR _6473_/Q sky130_fd_sc_hd__dfrtp_2
X_3685_ _3685_/A1 _3685_/A2 _3502_/Y _6246_/B2 wire763/X VGND VGND VPWR VPWR _3688_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_106_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5424_ _5469_/A1 hold585/X _5424_/S VGND VGND VPWR VPWR _6996_/D sky130_fd_sc_hd__mux2_1
Xoutput200 _3202_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[32] sky130_fd_sc_hd__buf_12
Xoutput211 _3226_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[8] sky130_fd_sc_hd__buf_12
XFILLER_133_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput222 _6548_/Q VGND VGND VPWR VPWR mgmt_gpio_out[18] sky130_fd_sc_hd__buf_12
Xoutput233 hold33/A VGND VGND VPWR VPWR mgmt_gpio_out[28] sky130_fd_sc_hd__buf_12
Xoutput244 _6557_/Q VGND VGND VPWR VPWR mgmt_gpio_out[3] sky130_fd_sc_hd__buf_12
XFILLER_114_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5355_ _5481_/A0 hold629/X _5355_/S VGND VGND VPWR VPWR _6935_/D sky130_fd_sc_hd__mux2_1
Xoutput255 _3951_/X VGND VGND VPWR VPWR pad_flash_io0_do sky130_fd_sc_hd__buf_12
Xoutput266 _6793_/Q VGND VGND VPWR VPWR pll_div[0] sky130_fd_sc_hd__buf_12
Xoutput277 _6485_/Q VGND VGND VPWR VPWR pll_trim[11] sky130_fd_sc_hd__buf_12
XFILLER_99_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput288 _6479_/Q VGND VGND VPWR VPWR pll_trim[21] sky130_fd_sc_hd__buf_12
X_4306_ _4306_/A _5229_/B VGND VGND VPWR VPWR _4311_/S sky130_fd_sc_hd__nand2_2
Xoutput299 _6482_/Q VGND VGND VPWR VPWR pll_trim[8] sky130_fd_sc_hd__buf_12
XFILLER_102_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5286_ _5286_/A _5286_/B VGND VGND VPWR VPWR _5291_/S sky130_fd_sc_hd__nand2_2
XFILLER_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1008 wire1009/X VGND VGND VPWR VPWR wire1008/X sky130_fd_sc_hd__clkbuf_1
X_7025_ _7109_/CLK _7025_/D wire4004/X VGND VGND VPWR VPWR _7025_/Q sky130_fd_sc_hd__dfrtp_1
Xwire1019 wire1020/X VGND VGND VPWR VPWR wire1019/X sky130_fd_sc_hd__clkbuf_1
X_4237_ _4237_/A0 hold349/X _4239_/S VGND VGND VPWR VPWR _6683_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4168_ _6628_/Q wire363/X _4170_/S VGND VGND VPWR VPWR _6628_/D sky130_fd_sc_hd__mux2_1
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4099_ hold184/X _4098_/X _4103_/S VGND VGND VPWR VPWR _6571_/D sky130_fd_sc_hd__mux2_1
XFILLER_82_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6809_ _7081_/CLK _6809_/D _7159_/RESET_B VGND VGND VPWR VPWR _6809_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length3601 _5477_/A0 VGND VGND VPWR VPWR _5573_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length3612 _5459_/A0 VGND VGND VPWR VPWR _5432_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_156_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_70_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7076_/CLK sky130_fd_sc_hd__clkbuf_16
Xmax_length2944 _5691_/B VGND VGND VPWR VPWR wire2937/A sky130_fd_sc_hd__clkbuf_1
Xmax_length2955 _5688_/X VGND VGND VPWR VPWR _5820_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_191_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2210 _6724_/Q VGND VGND VPWR VPWR wire2210/X sky130_fd_sc_hd__clkbuf_1
Xwire2221 _4263_/A0 VGND VGND VPWR VPWR _5960_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2232 _6709_/Q VGND VGND VPWR VPWR _6297_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire2243 _6273_/A1 VGND VGND VPWR VPWR _5906_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_120_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2254 _6685_/Q VGND VGND VPWR VPWR _6325_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1520 _3307_/Y VGND VGND VPWR VPWR _3607_/B sky130_fd_sc_hd__clkbuf_2
Xwire1531 _7138_/Q VGND VGND VPWR VPWR _6117_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2276 _6669_/Q VGND VGND VPWR VPWR _6333_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2287 _4206_/A0 VGND VGND VPWR VPWR _5899_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire1542 wire1543/X VGND VGND VPWR VPWR wire1542/X sky130_fd_sc_hd__clkbuf_1
Xwire1553 wire1554/X VGND VGND VPWR VPWR wire1553/X sky130_fd_sc_hd__clkbuf_1
Xwire2298 _6637_/Q VGND VGND VPWR VPWR wire2298/X sky130_fd_sc_hd__clkbuf_1
Xwire1564 _6102_/A1 VGND VGND VPWR VPWR wire1564/X sky130_fd_sc_hd__clkbuf_1
Xwire1575 _6079_/B2 VGND VGND VPWR VPWR _3616_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_74_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1586 wire1587/X VGND VGND VPWR VPWR wire1586/X sky130_fd_sc_hd__clkbuf_1
Xwire1597 _3363_/A1 VGND VGND VPWR VPWR _6198_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_23_csclk _6579_/CLK VGND VGND VPWR VPWR _7083_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_38_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7133_/CLK sky130_fd_sc_hd__clkbuf_16
Xwire850 wire851/X VGND VGND VPWR VPWR _4104_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire861 wire862/X VGND VGND VPWR VPWR _5322_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xwire872 _3339_/Y VGND VGND VPWR VPWR wire872/X sky130_fd_sc_hd__clkbuf_1
Xwire883 _4085_/S VGND VGND VPWR VPWR _4079_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_6_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire894 wire895/X VGND VGND VPWR VPWR wire894/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3470_ _5778_/A1 _3470_/A2 wire864/X _6129_/B2 _3469_/X VGND VGND VPWR VPWR _3484_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_182_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout4073 wire4082/X VGND VGND VPWR VPWR fanout4073/X sky130_fd_sc_hd__buf_6
XFILLER_170_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5140_ _5140_/A _5140_/B _5119_/Y VGND VGND VPWR VPWR _5140_/X sky130_fd_sc_hd__or3b_1
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire4190 input48/X VGND VGND VPWR VPWR wire4190/X sky130_fd_sc_hd__clkbuf_1
XFILLER_123_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5071_ _5071_/A _5112_/C _5071_/C VGND VGND VPWR VPWR _5156_/A sky130_fd_sc_hd__or3_1
X_4022_ _4022_/A _4135_/B VGND VGND VPWR VPWR _4027_/S sky130_fd_sc_hd__and2_2
XFILLER_65_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5973_ _6019_/A _6006_/B VGND VGND VPWR VPWR _6023_/A sky130_fd_sc_hd__nor2_1
XFILLER_80_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4924_ _4924_/A _4924_/B VGND VGND VPWR VPWR _4924_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4855_ _4461_/B _4613_/B _4910_/B1 _4784_/A _4837_/X VGND VGND VPWR VPWR _4857_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_178_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3806_ _6541_/Q _3806_/B VGND VGND VPWR VPWR _3833_/S sky130_fd_sc_hd__nand2b_1
X_4786_ _4425_/B _4798_/B2 _4598_/B VGND VGND VPWR VPWR _4786_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_193_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6525_ _7067_/CLK _6525_/D wire3968/A VGND VGND VPWR VPWR _6525_/Q sky130_fd_sc_hd__dfrtp_1
X_3737_ _6665_/Q _4210_/A _4159_/A _6621_/Q VGND VGND VPWR VPWR _3737_/X sky130_fd_sc_hd__a22o_1
X_6456_ _6545_/CLK _6456_/D _6411_/X VGND VGND VPWR VPWR _6456_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3668_ _7136_/Q wire950/X _3668_/B1 _3668_/B2 _3667_/X VGND VGND VPWR VPWR _3669_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5407_ _5584_/A0 hold188/X _5409_/S VGND VGND VPWR VPWR _6981_/D sky130_fd_sc_hd__mux2_1
XFILLER_134_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6387_ _6387_/A1 _4230_/X _4231_/Y _3191_/Y VGND VGND VPWR VPWR _7205_/D sky130_fd_sc_hd__o211a_2
X_3599_ _3599_/A1 _3599_/A2 _3617_/B1 _3599_/B2 _3598_/X VGND VGND VPWR VPWR _3600_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5338_ _5356_/A0 hold663/X _5338_/S VGND VGND VPWR VPWR _6920_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5269_ _5269_/A0 hold515/X _5269_/S VGND VGND VPWR VPWR _6858_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7008_ _7080_/CLK _7008_/D wire3992/A VGND VGND VPWR VPWR _7008_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length2785 _5992_/X VGND VGND VPWR VPWR _6024_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_124_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2040 _6873_/Q VGND VGND VPWR VPWR _6199_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire2051 _3872_/B VGND VGND VPWR VPWR _3571_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire2062 _5788_/B2 VGND VGND VPWR VPWR _3506_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2073 _3388_/B2 VGND VGND VPWR VPWR _6185_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2084 _6105_/A1 VGND VGND VPWR VPWR _5754_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire2095 wire2096/X VGND VGND VPWR VPWR wire2095/X sky130_fd_sc_hd__clkbuf_1
Xwire1350 wire1351/X VGND VGND VPWR VPWR wire1350/X sky130_fd_sc_hd__clkbuf_2
XFILLER_47_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1361 wire1362/X VGND VGND VPWR VPWR wire1361/X sky130_fd_sc_hd__clkbuf_1
Xwire1372 wire1372/A VGND VGND VPWR VPWR _3510_/B sky130_fd_sc_hd__buf_2
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1394 wire1394/A VGND VGND VPWR VPWR _3525_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_46_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4640_ _5152_/A1 _4620_/A _4799_/B1 VGND VGND VPWR VPWR _4640_/X sky130_fd_sc_hd__a21o_1
XFILLER_175_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4571_ _4562_/X _4565_/X _4568_/X _4484_/A VGND VGND VPWR VPWR _4571_/X sky130_fd_sc_hd__o211a_1
XFILLER_156_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6310_ _6310_/A1 _6310_/A2 _6310_/B1 _6684_/Q VGND VGND VPWR VPWR _6310_/X sky130_fd_sc_hd__a22o_1
XFILLER_128_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold705 _6489_/Q VGND VGND VPWR VPWR hold705/X sky130_fd_sc_hd__dlygate4sd3_1
X_3522_ _6125_/A1 _3522_/A2 _3522_/B1 _7062_/Q VGND VGND VPWR VPWR _3522_/X sky130_fd_sc_hd__a22o_1
Xwire680 _5381_/S VGND VGND VPWR VPWR _5378_/S sky130_fd_sc_hd__clkbuf_2
Xwire691 wire694/A VGND VGND VPWR VPWR _5357_/S sky130_fd_sc_hd__clkbuf_2
Xhold716 _7002_/Q VGND VGND VPWR VPWR hold716/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold727 _6468_/Q VGND VGND VPWR VPWR _3244_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6241_ _6241_/A _6241_/B _6241_/C _6241_/D VGND VGND VPWR VPWR _6242_/D sky130_fd_sc_hd__or4_1
XFILLER_116_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3453_ _3453_/A1 _3317_/Y _3453_/B1 _6323_/A1 _3452_/X VGND VGND VPWR VPWR _3468_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6172_ _6172_/A1 _6172_/A2 _6172_/B1 _6172_/B2 VGND VGND VPWR VPWR _6172_/X sky130_fd_sc_hd__a22o_1
X_3384_ _6984_/Q _3384_/A2 _3384_/B1 _3384_/B2 VGND VGND VPWR VPWR _3384_/X sky130_fd_sc_hd__a22o_1
XFILLER_97_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5123_ _5123_/A _5123_/B _5123_/C VGND VGND VPWR VPWR _5123_/X sky130_fd_sc_hd__and3_1
XFILLER_85_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5054_ _5054_/A _5054_/B VGND VGND VPWR VPWR _5162_/C sky130_fd_sc_hd__nand2_1
XFILLER_85_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4005_ _5575_/A0 hold209/X _4007_/S VGND VGND VPWR VPWR _6501_/D sky130_fd_sc_hd__mux2_1
XFILLER_65_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5956_ _6322_/A1 _5956_/A2 _5956_/B1 _6327_/A1 _5955_/X VGND VGND VPWR VPWR _5957_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4907_ _4984_/A _4983_/A _4986_/A _5079_/A VGND VGND VPWR VPWR _4915_/B sky130_fd_sc_hd__or4_1
X_5887_ _5887_/A1 _5887_/A2 _5927_/A2 _6617_/Q VGND VGND VPWR VPWR _5887_/X sky130_fd_sc_hd__a22o_1
XFILLER_178_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4838_ _4951_/B _4846_/D VGND VGND VPWR VPWR _4868_/A sky130_fd_sc_hd__and2_1
XFILLER_5_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4769_ _4446_/Y _4870_/B _4741_/X _5134_/A _4768_/X VGND VGND VPWR VPWR _4770_/B
+ sky130_fd_sc_hd__a2111o_1
X_6508_ _6701_/CLK _6508_/D _6429_/A VGND VGND VPWR VPWR _6508_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_119_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6439_ _6440_/A _6440_/B VGND VGND VPWR VPWR _6439_/X sky130_fd_sc_hd__and2_1
XFILLER_122_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold10 hold10/A VGND VGND VPWR VPWR hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A VGND VGND VPWR VPWR hold21/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold32 hold32/A VGND VGND VPWR VPWR hold32/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A VGND VGND VPWR VPWR hold43/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold54 hold54/A VGND VGND VPWR VPWR hold54/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold65 hold65/A VGND VGND VPWR VPWR hold65/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_188_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold76 hold76/A VGND VGND VPWR VPWR hold76/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold87 hold87/A VGND VGND VPWR VPWR hold87/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold98 hold98/A VGND VGND VPWR VPWR hold98/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_7 mgmt_gpio_in[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1180 _3323_/Y VGND VGND VPWR VPWR _3537_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1191 wire1192/X VGND VGND VPWR VPWR wire1191/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5810_ _6903_/Q _5817_/A2 _5810_/B1 _6164_/A1 _5809_/X VGND VGND VPWR VPWR _5813_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_35_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6790_ _6545_/CLK _6790_/D _6441_/X VGND VGND VPWR VPWR _6790_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_62_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5741_ hold91/A _5741_/A2 _5741_/B1 hold89/A VGND VGND VPWR VPWR _5741_/X sky130_fd_sc_hd__a22o_1
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5672_ _5688_/A _5699_/B _5699_/C VGND VGND VPWR VPWR _5672_/X sky130_fd_sc_hd__and3_1
XFILLER_175_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4623_ _4623_/A _4639_/B VGND VGND VPWR VPWR _4627_/C sky130_fd_sc_hd__nor2_1
XFILLER_163_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4554_ _4792_/A _4792_/C _4792_/B VGND VGND VPWR VPWR _4802_/C sky130_fd_sc_hd__o21bai_1
XFILLER_144_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold502 _6762_/Q VGND VGND VPWR VPWR hold502/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 _6813_/Q VGND VGND VPWR VPWR hold513/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 _6660_/Q VGND VGND VPWR VPWR hold524/X sky130_fd_sc_hd__dlygate4sd3_1
X_3505_ _6659_/Q _4198_/A _3504_/Y _5959_/B2 VGND VGND VPWR VPWR _3505_/X sky130_fd_sc_hd__a22o_1
Xhold535 _6975_/Q VGND VGND VPWR VPWR hold535/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4485_ _4485_/A _4485_/B VGND VGND VPWR VPWR _4887_/C sky130_fd_sc_hd__nand2_1
Xhold546 _6821_/Q VGND VGND VPWR VPWR hold546/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 _7099_/Q VGND VGND VPWR VPWR hold557/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold568 _7098_/Q VGND VGND VPWR VPWR hold568/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6224_ _6224_/A1 _6335_/A2 _6300_/B1 _6224_/B2 VGND VGND VPWR VPWR _6241_/A sky130_fd_sc_hd__a22o_1
Xhold579 _6720_/Q VGND VGND VPWR VPWR hold579/X sky130_fd_sc_hd__dlygate4sd3_1
X_3436_ _5801_/B2 _3436_/A2 wire894/X _6147_/A1 VGND VGND VPWR VPWR _3436_/X sky130_fd_sc_hd__a22o_1
XFILLER_103_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2809 _6237_/A2 VGND VGND VPWR VPWR _6337_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6155_ _6975_/Q _6190_/B1 _6155_/B1 _6155_/B2 _6154_/X VGND VGND VPWR VPWR _6156_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ _7001_/Q _5421_/A _5466_/A _7041_/Q _3345_/X VGND VGND VPWR VPWR _3367_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_106_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5106_ _5106_/A _5106_/B _5106_/C _5105_/X VGND VGND VPWR VPWR _5156_/C sky130_fd_sc_hd__or4b_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6086_ _6086_/A1 _6086_/A2 _6086_/B1 _6086_/B2 VGND VGND VPWR VPWR _6086_/X sky130_fd_sc_hd__a22o_1
X_3298_ _3526_/A _3476_/A VGND VGND VPWR VPWR _3298_/Y sky130_fd_sc_hd__nor2_1
X_5037_ _4485_/A _5035_/Y _5036_/Y _4418_/B VGND VGND VPWR VPWR _5136_/A sky130_fd_sc_hd__a22o_1
XFILLER_38_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6988_ _7076_/CLK _6988_/D wire3978/X VGND VGND VPWR VPWR _6988_/Q sky130_fd_sc_hd__dfrtp_1
X_5939_ _6310_/A1 _5950_/A2 _5961_/B2 _5938_/X VGND VGND VPWR VPWR _5939_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_22 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout3949 wire3956/A VGND VGND VPWR VPWR wire3950/A sky130_fd_sc_hd__buf_6
XFILLER_1_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput100 wb_adr_i[10] VGND VGND VPWR VPWR _4339_/D sky130_fd_sc_hd__clkbuf_1
Xinput111 wb_adr_i[20] VGND VGND VPWR VPWR _4654_/A sky130_fd_sc_hd__clkbuf_2
Xinput122 wb_adr_i[30] VGND VGND VPWR VPWR _3884_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_49_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput133 wb_dat_i[10] VGND VGND VPWR VPWR _6369_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput144 wb_dat_i[20] VGND VGND VPWR VPWR _6375_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput155 wb_dat_i[30] VGND VGND VPWR VPWR _6381_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput166 wb_sel_i[1] VGND VGND VPWR VPWR _6389_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4270_ _4270_/A _4270_/B VGND VGND VPWR VPWR _4275_/S sky130_fd_sc_hd__and2_2
XFILLER_180_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3221_ _3221_/A VGND VGND VPWR VPWR _3221_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6911_ _7031_/CLK _6911_/D wire4044/X VGND VGND VPWR VPWR _6911_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_63_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6842_ _7115_/CLK _6842_/D wire3980/X VGND VGND VPWR VPWR _6842_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_50_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6773_ _6824_/CLK _6773_/D fanout3973/X VGND VGND VPWR VPWR _6773_/Q sky130_fd_sc_hd__dfstp_1
X_3985_ hold720/X _5231_/A0 _3988_/S VGND VGND VPWR VPWR _6483_/D sky130_fd_sc_hd__mux2_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5724_ _6062_/B2 _5724_/A2 _5724_/B1 hold93/A VGND VGND VPWR VPWR _5724_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5655_ _5688_/A _5700_/C _5699_/B VGND VGND VPWR VPWR _5655_/X sky130_fd_sc_hd__and3_1
XFILLER_176_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4606_ _4802_/C _4606_/B _4606_/C _4793_/B VGND VGND VPWR VPWR _4607_/D sky130_fd_sc_hd__and4b_1
XFILLER_136_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5586_ _5586_/A0 hold594/X _5586_/S VGND VGND VPWR VPWR _7140_/D sky130_fd_sc_hd__mux2_1
Xhold310 _6888_/Q VGND VGND VPWR VPWR hold310/X sky130_fd_sc_hd__dlygate4sd3_1
X_4537_ _4570_/A _4570_/B _4570_/C _4570_/D VGND VGND VPWR VPWR _4971_/B sky130_fd_sc_hd__and4_1
Xhold321 _6850_/Q VGND VGND VPWR VPWR hold321/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire4019 wire4019/A VGND VGND VPWR VPWR wire4019/X sky130_fd_sc_hd__clkbuf_2
Xhold332 _6671_/Q VGND VGND VPWR VPWR hold332/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold343 _6953_/Q VGND VGND VPWR VPWR hold343/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold354 _6620_/Q VGND VGND VPWR VPWR hold354/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 _6773_/Q VGND VGND VPWR VPWR hold365/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3318 _4581_/X VGND VGND VPWR VPWR _4582_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4468_ _4489_/A _4484_/B _4352_/B VGND VGND VPWR VPWR _4468_/X sky130_fd_sc_hd__or3b_1
Xhold376 _6735_/Q VGND VGND VPWR VPWR hold376/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 _6826_/Q VGND VGND VPWR VPWR hold387/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3329 _4545_/X VGND VGND VPWR VPWR _5169_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold398 _6844_/Q VGND VGND VPWR VPWR hold398/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2606 _4823_/A VGND VGND VPWR VPWR _5127_/A sky130_fd_sc_hd__clkbuf_2
X_6207_ _7073_/Q _6207_/A2 _6202_/X _6204_/X _6206_/X VGND VGND VPWR VPWR _6207_/X
+ sky130_fd_sc_hd__a2111o_1
Xwire2617 wire2617/A VGND VGND VPWR VPWR _6339_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3419_ _6162_/A1 wire934/X _3419_/B1 _5801_/A1 VGND VGND VPWR VPWR _3419_/X sky130_fd_sc_hd__a22o_1
X_7187_ _7187_/CLK _7187_/D wire3984/X VGND VGND VPWR VPWR _7187_/Q sky130_fd_sc_hd__dfrtp_1
Xwire2628 _6090_/B1 VGND VGND VPWR VPWR _6248_/B sky130_fd_sc_hd__clkbuf_1
X_4399_ _4420_/A _4596_/A VGND VGND VPWR VPWR _4400_/B sky130_fd_sc_hd__or2_1
Xwire2639 _6181_/B1 VGND VGND VPWR VPWR wire2639/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1905 _6942_/Q VGND VGND VPWR VPWR _5780_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1916 _6935_/Q VGND VGND VPWR VPWR _6163_/B2 sky130_fd_sc_hd__clkbuf_2
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6138_ _6950_/Q _6138_/A2 _6138_/B1 _6138_/B2 VGND VGND VPWR VPWR _6138_/X sky130_fd_sc_hd__a22o_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1927 wire1927/A VGND VGND VPWR VPWR wire1927/X sky130_fd_sc_hd__clkbuf_1
Xwire1938 wire1939/X VGND VGND VPWR VPWR _5778_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire1949 _6924_/Q VGND VGND VPWR VPWR wire1949/X sky130_fd_sc_hd__clkbuf_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6069_ _6069_/A _6069_/B _6069_/C _6069_/D VGND VGND VPWR VPWR _6069_/X sky130_fd_sc_hd__or4_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length888 _3337_/Y VGND VGND VPWR VPWR wire881/A sky130_fd_sc_hd__clkbuf_1
Xmax_length899 _3335_/Y VGND VGND VPWR VPWR _3509_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_107_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3830 _4341_/X VGND VGND VPWR VPWR _4412_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_174_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3841 _6440_/B VGND VGND VPWR VPWR _6435_/B sky130_fd_sc_hd__clkbuf_2
Xwire3852 _4533_/A VGND VGND VPWR VPWR _4607_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire3863 wire3864/X VGND VGND VPWR VPWR _3649_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_89_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3874 wire3875/X VGND VGND VPWR VPWR wire3874/X sky130_fd_sc_hd__clkbuf_1
Xwire3885 input92/X VGND VGND VPWR VPWR wire3885/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3896 input88/X VGND VGND VPWR VPWR wire3896/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3770_ _5864_/B2 _3770_/A2 _3547_/Y _3770_/B2 VGND VGND VPWR VPWR _3770_/X sky130_fd_sc_hd__a22o_1
XFILLER_32_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5440_ _5440_/A0 hold412/X _5440_/S VGND VGND VPWR VPWR _7010_/D sky130_fd_sc_hd__mux2_1
XFILLER_157_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5371_ _5389_/A0 hold227/X _5375_/S VGND VGND VPWR VPWR _6949_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7110_ _7110_/CLK _7110_/D _7110_/RESET_B VGND VGND VPWR VPWR _7110_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_114_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4322_ hold391/X _4322_/A1 _4323_/S VGND VGND VPWR VPWR _6764_/D sky130_fd_sc_hd__mux2_1
XFILLER_153_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7041_ _7080_/CLK _7041_/D wire3991/X VGND VGND VPWR VPWR _7041_/Q sky130_fd_sc_hd__dfrtp_1
X_4253_ hold501/X _4259_/A1 _4257_/S VGND VGND VPWR VPWR _6706_/D sky130_fd_sc_hd__mux2_1
X_3204_ _3204_/A VGND VGND VPWR VPWR _3204_/Y sky130_fd_sc_hd__inv_2
X_4184_ _6642_/Q wire366/X _4188_/S VGND VGND VPWR VPWR _6642_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A VGND VGND VPWR VPWR _7204_/CLK sky130_fd_sc_hd__clkbuf_8
X_6825_ _6825_/CLK _6825_/D wire3954/X VGND VGND VPWR VPWR _6825_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6756_ _6761_/CLK _6756_/D wire4019/X VGND VGND VPWR VPWR _6756_/Q sky130_fd_sc_hd__dfrtp_1
X_3968_ hold714/X _3984_/A1 _3976_/S VGND VGND VPWR VPWR _6474_/D sky130_fd_sc_hd__mux2_1
XFILLER_148_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3816 _4693_/A VGND VGND VPWR VPWR _4661_/B sky130_fd_sc_hd__clkbuf_2
Xmax_length3827 _4657_/B VGND VGND VPWR VPWR _4667_/B sky130_fd_sc_hd__clkbuf_2
X_5707_ _5707_/A1 _5707_/A2 _5707_/B1 _6498_/Q _5707_/C1 VGND VGND VPWR VPWR _5708_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6687_ _7093_/CLK _6687_/D wire3961/X VGND VGND VPWR VPWR _6687_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_148_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3899_ _5592_/B _3899_/B _7146_/Q _7147_/Q VGND VGND VPWR VPWR _3908_/B sky130_fd_sc_hd__and4b_1
XFILLER_164_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5638_ _7157_/Q _5643_/A VGND VGND VPWR VPWR _5638_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5569_ _5569_/A0 hold510/X _5569_/S VGND VGND VPWR VPWR _7125_/D sky130_fd_sc_hd__mux2_1
XFILLER_163_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold140 _6779_/Q VGND VGND VPWR VPWR hold140/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 _6907_/Q VGND VGND VPWR VPWR hold151/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold162 _6859_/Q VGND VGND VPWR VPWR hold162/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3104 _5727_/A2 VGND VGND VPWR VPWR _5805_/A2 sky130_fd_sc_hd__clkbuf_2
Xhold173 _6956_/Q VGND VGND VPWR VPWR hold173/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3126 _5841_/A2 VGND VGND VPWR VPWR _5802_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold184 _6571_/Q VGND VGND VPWR VPWR hold184/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3137 _5853_/A2 VGND VGND VPWR VPWR _5804_/A2 sky130_fd_sc_hd__clkbuf_1
Xhold195 _6906_/Q VGND VGND VPWR VPWR hold195/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire2403 wire2403/A VGND VGND VPWR VPWR wire2403/X sky130_fd_sc_hd__clkbuf_1
Xwire3148 _5855_/A2 VGND VGND VPWR VPWR _5812_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire2414 _6506_/Q VGND VGND VPWR VPWR _6227_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3159 _6163_/A2 VGND VGND VPWR VPWR _6140_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire2425 _5755_/B2 VGND VGND VPWR VPWR _6115_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2436 _6496_/Q VGND VGND VPWR VPWR wire2436/X sky130_fd_sc_hd__clkbuf_1
Xwire2447 wire2448/X VGND VGND VPWR VPWR _3361_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire1702 wire1703/X VGND VGND VPWR VPWR _6141_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_58_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1713 _5742_/B2 VGND VGND VPWR VPWR _6076_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire2458 _6057_/B1 VGND VGND VPWR VPWR _6042_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_58_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2469 _6182_/B1 VGND VGND VPWR VPWR wire2469/X sky130_fd_sc_hd__clkbuf_1
Xwire1735 _7028_/Q VGND VGND VPWR VPWR wire1735/X sky130_fd_sc_hd__clkbuf_1
Xwire1746 wire1747/X VGND VGND VPWR VPWR _6152_/A1 sky130_fd_sc_hd__clkbuf_2
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1757 wire1757/A VGND VGND VPWR VPWR wire1757/X sky130_fd_sc_hd__clkbuf_1
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1768 _3351_/B2 VGND VGND VPWR VPWR _6201_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_18_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1779 _6089_/A1 VGND VGND VPWR VPWR wire1779/X sky130_fd_sc_hd__clkbuf_1
XFILLER_170_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3660 _5545_/A0 VGND VGND VPWR VPWR _5350_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3671 wire3672/X VGND VGND VPWR VPWR wire3671/X sky130_fd_sc_hd__clkbuf_1
Xwire3682 _5693_/A VGND VGND VPWR VPWR _5683_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3693 _5946_/C1 VGND VGND VPWR VPWR _6342_/C1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2970 _5779_/B1 VGND VGND VPWR VPWR _5721_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2992 _5789_/B1 VGND VGND VPWR VPWR _5714_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_92_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4940_ _4940_/A _4940_/B VGND VGND VPWR VPWR _4940_/Y sky130_fd_sc_hd__nor2_1
XFILLER_92_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4871_ _4871_/A _4871_/B VGND VGND VPWR VPWR _4871_/Y sky130_fd_sc_hd__nand2_1
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3822_ _3821_/X _6467_/Q _3828_/S VGND VGND VPWR VPWR _6467_/D sky130_fd_sc_hd__mux2_1
X_6610_ _7208_/CLK _6610_/D wire4026/A VGND VGND VPWR VPWR _6610_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_177_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6541_ _3945_/A1 _6541_/D _6429_/X VGND VGND VPWR VPWR _6541_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_193_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3753_ _3753_/A1 wire830/X _5223_/A _6820_/Q wire541/X VGND VGND VPWR VPWR _3755_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6472_ _3945_/A1 _6472_/D _6427_/X VGND VGND VPWR VPWR _6472_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_146_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3684_ _7075_/Q _3684_/A2 _3684_/B1 _5711_/A1 VGND VGND VPWR VPWR _3684_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5423_ _5537_/A1 hold588/X _5424_/S VGND VGND VPWR VPWR _6995_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput201 _3201_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[33] sky130_fd_sc_hd__buf_12
Xoutput212 _3225_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[9] sky130_fd_sc_hd__buf_12
Xoutput223 _6549_/Q VGND VGND VPWR VPWR mgmt_gpio_out[19] sky130_fd_sc_hd__buf_12
Xoutput234 _6831_/Q VGND VGND VPWR VPWR mgmt_gpio_out[29] sky130_fd_sc_hd__buf_12
X_5354_ _5576_/A0 hold133/X _5354_/S VGND VGND VPWR VPWR _6934_/D sky130_fd_sc_hd__mux2_1
Xoutput245 _6558_/Q VGND VGND VPWR VPWR mgmt_gpio_out[4] sky130_fd_sc_hd__buf_12
Xoutput256 _3948_/A VGND VGND VPWR VPWR pad_flash_io0_ieb sky130_fd_sc_hd__buf_12
XFILLER_114_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput267 _6794_/Q VGND VGND VPWR VPWR pll_div[1] sky130_fd_sc_hd__buf_12
X_4305_ _4305_/A0 hold236/X hold31/X VGND VGND VPWR VPWR _6750_/D sky130_fd_sc_hd__mux2_1
Xoutput278 _6486_/Q VGND VGND VPWR VPWR pll_trim[12] sky130_fd_sc_hd__buf_12
X_5285_ _5348_/A0 _6873_/Q _5285_/S VGND VGND VPWR VPWR hold86/A sky130_fd_sc_hd__mux2_1
Xoutput289 _6480_/Q VGND VGND VPWR VPWR pll_trim[22] sky130_fd_sc_hd__buf_12
XFILLER_59_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7024_ _7080_/CLK _7024_/D _6562_/SET_B VGND VGND VPWR VPWR _7024_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4236_ _4248_/A0 hold347/X _4239_/S VGND VGND VPWR VPWR _6682_/D sky130_fd_sc_hd__mux2_1
Xwire1009 _5651_/Y VGND VGND VPWR VPWR wire1009/X sky130_fd_sc_hd__clkbuf_1
X_4167_ _6627_/Q wire361/X _4173_/S VGND VGND VPWR VPWR _6627_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4098_ hold121/X _5247_/A0 _4102_/S VGND VGND VPWR VPWR _4098_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_4_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _6705_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_51_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4303 _4396_/A VGND VGND VPWR VPWR _4419_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_11_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6808_ _7081_/CLK _6808_/D _7159_/RESET_B VGND VGND VPWR VPWR _6808_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_168_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3602 _5477_/A0 VGND VGND VPWR VPWR _5342_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6739_ _6979_/CLK _6739_/D fanout4027/X VGND VGND VPWR VPWR _6739_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length3635 _5536_/A1 VGND VGND VPWR VPWR _5467_/A1 sky130_fd_sc_hd__clkbuf_1
Xmax_length3657 wire3656/A VGND VGND VPWR VPWR _5233_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_109_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2200 _3753_/A1 VGND VGND VPWR VPWR wire2200/X sky130_fd_sc_hd__clkbuf_1
Xwire2211 _3621_/B2 VGND VGND VPWR VPWR _6279_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2233 _5927_/B2 VGND VGND VPWR VPWR _3558_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire2244 _6703_/Q VGND VGND VPWR VPWR _6273_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1510 _3378_/Y VGND VGND VPWR VPWR _3460_/B sky130_fd_sc_hd__clkbuf_1
Xwire2255 _6683_/Q VGND VGND VPWR VPWR _5921_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1521 _3305_/Y VGND VGND VPWR VPWR _3318_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2266 _6676_/Q VGND VGND VPWR VPWR _3720_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire1532 _7134_/Q VGND VGND VPWR VPWR _6197_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_171_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2277 _6668_/Q VGND VGND VPWR VPWR _6310_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_120_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1543 wire1544/X VGND VGND VPWR VPWR wire1543/X sky130_fd_sc_hd__clkbuf_1
Xwire2299 _6637_/Q VGND VGND VPWR VPWR _6311_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1554 wire1555/X VGND VGND VPWR VPWR wire1554/X sky130_fd_sc_hd__clkbuf_1
Xwire1565 _7114_/Q VGND VGND VPWR VPWR _6102_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1576 _7105_/Q VGND VGND VPWR VPWR _6079_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1587 _7098_/Q VGND VGND VPWR VPWR wire1587/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1598 _7089_/Q VGND VGND VPWR VPWR _3363_/A1 sky130_fd_sc_hd__clkbuf_1
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire840 _3439_/X VGND VGND VPWR VPWR wire840/X sky130_fd_sc_hd__clkbuf_1
XFILLER_127_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire851 wire852/X VGND VGND VPWR VPWR wire851/X sky130_fd_sc_hd__dlymetal6s2s_1
Xwire862 wire863/X VGND VGND VPWR VPWR wire862/X sky130_fd_sc_hd__clkbuf_1
XFILLER_182_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire884 wire885/X VGND VGND VPWR VPWR _4085_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_127_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire895 wire896/X VGND VGND VPWR VPWR wire895/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_127_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4180 input51/X VGND VGND VPWR VPWR wire4180/X sky130_fd_sc_hd__clkbuf_1
XFILLER_123_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4191 wire4192/X VGND VGND VPWR VPWR _3709_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5070_ _5071_/A _5112_/C _5071_/C VGND VGND VPWR VPWR _5070_/Y sky130_fd_sc_hd__nor3_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3490 _6396_/A0 VGND VGND VPWR VPWR _4208_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4021_ _4045_/A0 hold299/X _4021_/S VGND VGND VPWR VPWR _6515_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5972_ _6000_/A _6039_/C VGND VGND VPWR VPWR _6006_/B sky130_fd_sc_hd__nand2_1
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4923_ _5153_/A _5109_/A _4923_/C _4923_/D VGND VGND VPWR VPWR _4924_/B sky130_fd_sc_hd__or4_1
XFILLER_178_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4854_ _4932_/A _4942_/B _4675_/A _4503_/C VGND VGND VPWR VPWR _4857_/B sky130_fd_sc_hd__o31a_1
XFILLER_60_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3805_ _6543_/Q _3834_/B _3890_/B _3850_/A VGND VGND VPWR VPWR _3806_/B sky130_fd_sc_hd__a31o_1
X_4785_ _4735_/A _4425_/B _5015_/B VGND VGND VPWR VPWR _4785_/X sky130_fd_sc_hd__a21o_1
XFILLER_165_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3736_ _5995_/B2 _3736_/A2 _3736_/B1 _3736_/B2 VGND VGND VPWR VPWR _3736_/X sky130_fd_sc_hd__a22o_1
X_6524_ _7066_/CLK _6524_/D wire3970/X VGND VGND VPWR VPWR _6524_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6455_ _6545_/CLK _6455_/D _6410_/X VGND VGND VPWR VPWR _6455_/Q sky130_fd_sc_hd__dfrtp_1
X_3667_ _3667_/A1 _3667_/A2 _3667_/B1 _6252_/A1 VGND VGND VPWR VPWR _3667_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5406_ _5406_/A0 hold89/X _5406_/S VGND VGND VPWR VPWR hold90/A sky130_fd_sc_hd__mux2_1
X_6386_ _6385_/X _7204_/Q _6386_/S VGND VGND VPWR VPWR _7204_/D sky130_fd_sc_hd__mux2_1
X_3598_ _3598_/A1 wire882/X _4264_/A _6308_/A1 _3597_/X VGND VGND VPWR VPWR _3598_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5337_ _5526_/A0 hold661/X _5337_/S VGND VGND VPWR VPWR _6919_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5268_ _5268_/A _5268_/B VGND VGND VPWR VPWR _5268_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7007_ _7027_/CLK _7007_/D wire3992/A VGND VGND VPWR VPWR _7007_/Q sky130_fd_sc_hd__dfrtp_1
X_4219_ _4237_/A0 hold339/X _4221_/S VGND VGND VPWR VPWR _6672_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5199_ _5199_/A0 hold450/X _5199_/S VGND VGND VPWR VPWR _6803_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length3421 _5481_/A0 VGND VGND VPWR VPWR _5364_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_137_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3487 hold15/X VGND VGND VPWR VPWR wire3486/A sky130_fd_sc_hd__clkbuf_1
XFILLER_164_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2030 _6879_/Q VGND VGND VPWR VPWR _6147_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2041 _5833_/A1 VGND VGND VPWR VPWR _3396_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_93_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2052 _5281_/A1 VGND VGND VPWR VPWR _3872_/B sky130_fd_sc_hd__clkbuf_2
Xwire2063 _6139_/A1 VGND VGND VPWR VPWR _5788_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2074 wire2075/X VGND VGND VPWR VPWR _3388_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire2085 wire2086/X VGND VGND VPWR VPWR _6105_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1340 _4965_/B VGND VGND VPWR VPWR _4894_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1351 wire1352/X VGND VGND VPWR VPWR wire1351/X sky130_fd_sc_hd__clkbuf_1
Xwire2096 _3555_/A1 VGND VGND VPWR VPWR wire2096/X sky130_fd_sc_hd__clkbuf_1
XFILLER_59_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1362 wire1363/X VGND VGND VPWR VPWR wire1362/X sky130_fd_sc_hd__clkbuf_1
XFILLER_46_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1384 _3482_/A VGND VGND VPWR VPWR _3534_/A sky130_fd_sc_hd__buf_2
Xwire1395 _3331_/A VGND VGND VPWR VPWR _3510_/A sky130_fd_sc_hd__buf_2
XFILLER_46_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4570_ _4570_/A _4570_/B _4570_/C _4570_/D VGND VGND VPWR VPWR _4664_/B sky130_fd_sc_hd__or4_2
XFILLER_162_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3521_ _5776_/A1 _5331_/A _3566_/B1 _7123_/Q VGND VGND VPWR VPWR _3524_/C sky130_fd_sc_hd__a22o_1
Xwire670 _5409_/S VGND VGND VPWR VPWR wire670/X sky130_fd_sc_hd__clkbuf_1
XFILLER_156_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold706 _6488_/Q VGND VGND VPWR VPWR hold706/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire692 _5355_/S VGND VGND VPWR VPWR _5354_/S sky130_fd_sc_hd__clkbuf_2
Xhold717 _6484_/Q VGND VGND VPWR VPWR hold717/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold728 _6692_/Q VGND VGND VPWR VPWR _6697_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6240_ _6601_/Q _6314_/A2 _6314_/B1 _6516_/Q _6239_/X VGND VGND VPWR VPWR _6241_/D
+ sky130_fd_sc_hd__a221o_1
X_3452_ _5778_/B2 _3452_/A2 wire833/X _3452_/B2 VGND VGND VPWR VPWR _3452_/X sky130_fd_sc_hd__a22o_1
XFILLER_171_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6171_ _7180_/Q _6170_/X _6171_/S VGND VGND VPWR VPWR _7180_/D sky130_fd_sc_hd__mux2_1
XFILLER_143_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3383_ _6182_/A1 _3383_/A2 _3383_/B1 _7016_/Q VGND VGND VPWR VPWR _3383_/X sky130_fd_sc_hd__a22o_1
XFILLER_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5122_ _4582_/B _5164_/A3 _4504_/A _4504_/B VGND VGND VPWR VPWR _5123_/C sky130_fd_sc_hd__o211a_1
XFILLER_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5053_ _5053_/A _5053_/B _5052_/X VGND VGND VPWR VPWR _5067_/A sky130_fd_sc_hd__or3b_1
X_4004_ _5514_/A0 hold569/X _4004_/S VGND VGND VPWR VPWR _6500_/D sky130_fd_sc_hd__mux2_1
XFILLER_1_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5955_ _6674_/Q _5955_/A2 _5955_/B1 _6325_/B2 VGND VGND VPWR VPWR _5955_/X sky130_fd_sc_hd__a22o_1
XFILLER_111_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4906_ _5021_/A _5023_/C _5021_/C VGND VGND VPWR VPWR _5079_/A sky130_fd_sc_hd__nor3_1
XFILLER_33_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5886_ _6622_/Q _5922_/A2 _5886_/B1 _5886_/B2 _5885_/X VGND VGND VPWR VPWR _5891_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_139_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_84_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6811_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_139_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4837_ _4652_/X _4836_/Y _4932_/A VGND VGND VPWR VPWR _4837_/X sky130_fd_sc_hd__a21o_1
XFILLER_193_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4768_ _4993_/A _4524_/B _4818_/B _4894_/A _4767_/X VGND VGND VPWR VPWR _4768_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_147_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6507_ _6702_/CLK _6507_/D _6440_/A VGND VGND VPWR VPWR _6507_/Q sky130_fd_sc_hd__dfrtp_1
X_3719_ _6052_/B2 _3719_/A2 _3719_/B1 _6762_/Q VGND VGND VPWR VPWR _3719_/X sky130_fd_sc_hd__a22o_1
X_4699_ _4699_/A _4699_/B _4860_/B _4699_/D VGND VGND VPWR VPWR _4699_/X sky130_fd_sc_hd__and4_1
Xmax_length1348 _4486_/A VGND VGND VPWR VPWR _4996_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_162_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6438_ _6438_/A _6440_/B VGND VGND VPWR VPWR _6438_/X sky130_fd_sc_hd__and2_1
XFILLER_20_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6369_ _4228_/B _6369_/A2 _6369_/B1 _4228_/A VGND VGND VPWR VPWR _6369_/X sky130_fd_sc_hd__a22o_1
XFILLER_96_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_22_csclk _6579_/CLK VGND VGND VPWR VPWR _7046_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_88_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold11 hold11/A VGND VGND VPWR VPWR hold11/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold22 hold22/A VGND VGND VPWR VPWR hold22/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 hold33/A VGND VGND VPWR VPWR hold33/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold44 hold44/A VGND VGND VPWR VPWR hold44/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold55 hold55/A VGND VGND VPWR VPWR hold55/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A VGND VGND VPWR VPWR hold66/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 hold77/A VGND VGND VPWR VPWR hold77/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 hold88/A VGND VGND VPWR VPWR hold88/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 hold99/A VGND VGND VPWR VPWR hold99/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_37_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7116_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_44_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_mgmt_gpio_in[4] mgmt_gpio_in[4] VGND VGND VPWR VPWR clkbuf_0_mgmt_gpio_in[4]/X
+ sky130_fd_sc_hd__clkbuf_16
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3251 _5529_/B VGND VGND VPWR VPWR _6392_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_172_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3273 _5553_/B VGND VGND VPWR VPWR _5520_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA_8 mgmt_gpio_in[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1170 _3325_/Y VGND VGND VPWR VPWR _3612_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1181 _3322_/Y VGND VGND VPWR VPWR _3747_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1192 _3321_/Y VGND VGND VPWR VPWR wire1192/X sky130_fd_sc_hd__clkbuf_1
XFILLER_62_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5740_ _5740_/A _5740_/B _5740_/C _5740_/D VGND VGND VPWR VPWR _5740_/X sky130_fd_sc_hd__or4_1
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5671_ _7152_/Q _5706_/B _5699_/C VGND VGND VPWR VPWR _5671_/X sky130_fd_sc_hd__and3_1
XFILLER_30_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4622_ _4639_/B VGND VGND VPWR VPWR _4622_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4553_ _4553_/A _4553_/B VGND VGND VPWR VPWR _4792_/C sky130_fd_sc_hd__nor2_1
XFILLER_175_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold503 _7067_/Q VGND VGND VPWR VPWR hold503/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold514 _6817_/Q VGND VGND VPWR VPWR hold514/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold525 _6717_/Q VGND VGND VPWR VPWR hold525/X sky130_fd_sc_hd__dlygate4sd3_1
X_3504_ _3504_/A _3538_/B VGND VGND VPWR VPWR _3504_/Y sky130_fd_sc_hd__nor2_1
XFILLER_116_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4484_ _4484_/A _4484_/B _4352_/B VGND VGND VPWR VPWR _4484_/X sky130_fd_sc_hd__or3b_1
Xhold536 _7071_/Q VGND VGND VPWR VPWR hold536/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 _6861_/Q VGND VGND VPWR VPWR hold547/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold558 _6982_/Q VGND VGND VPWR VPWR hold558/X sky130_fd_sc_hd__dlygate4sd3_1
X_6223_ _6223_/A1 _6334_/A2 _6299_/B1 _6223_/B2 VGND VGND VPWR VPWR _6223_/X sky130_fd_sc_hd__a22o_1
Xhold569 _6500_/Q VGND VGND VPWR VPWR hold569/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3435_ _6975_/Q _3570_/A2 wire910/X _6166_/A1 _3434_/X VGND VGND VPWR VPWR _3447_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6154_ _6959_/Q _6154_/A2 _6154_/B1 _6154_/B2 VGND VGND VPWR VPWR _6154_/X sky130_fd_sc_hd__a22o_1
X_3366_ _5842_/A1 wire933/X _3366_/B1 _3366_/B2 wire854/X VGND VGND VPWR VPWR _3371_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_662 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5105_ _5105_/A1 _5105_/A2 _5023_/C _5105_/B2 _4713_/A VGND VGND VPWR VPWR _5105_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6085_ _6085_/A _6085_/B VGND VGND VPWR VPWR _6085_/X sky130_fd_sc_hd__or2_1
X_3297_ _3297_/A _3301_/C hold26/X VGND VGND VPWR VPWR _3297_/X sky130_fd_sc_hd__or3b_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5036_ _5036_/A _5036_/B VGND VGND VPWR VPWR _5036_/Y sky130_fd_sc_hd__nand2_1
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6987_ _7121_/CLK _6987_/D wire4042/X VGND VGND VPWR VPWR _6987_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5938_ _5938_/A _5960_/B VGND VGND VPWR VPWR _5938_/X sky130_fd_sc_hd__or2_1
XFILLER_179_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5869_ _5869_/A _5869_/B _5869_/C _5869_/D VGND VGND VPWR VPWR _5869_/X sky130_fd_sc_hd__or4_1
XFILLER_178_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length1123 _3709_/A2 VGND VGND VPWR VPWR _3733_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_107_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length1145 _3329_/Y VGND VGND VPWR VPWR _3771_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_134_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput101 wb_adr_i[11] VGND VGND VPWR VPWR _4339_/C sky130_fd_sc_hd__clkbuf_1
Xinput112 wb_adr_i[21] VGND VGND VPWR VPWR _4390_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_88_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput123 wb_adr_i[31] VGND VGND VPWR VPWR _3884_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_102_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput134 wb_dat_i[11] VGND VGND VPWR VPWR _6372_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput145 wb_dat_i[21] VGND VGND VPWR VPWR _6378_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput156 wb_dat_i[31] VGND VGND VPWR VPWR _6384_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput167 wb_sel_i[2] VGND VGND VPWR VPWR _6358_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_102_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_646 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3220_ _6957_/Q VGND VGND VPWR VPWR _3220_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6910_ _7140_/CLK _6910_/D fanout4057/X VGND VGND VPWR VPWR _6910_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_82_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6841_ _7131_/CLK hold9/X fanout4057/X VGND VGND VPWR VPWR _6841_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6772_ _6824_/CLK _6772_/D _6483_/SET_B VGND VGND VPWR VPWR _6772_/Q sky130_fd_sc_hd__dfrtp_1
X_3984_ hold719/X _3984_/A1 _3988_/S VGND VGND VPWR VPWR _6482_/D sky130_fd_sc_hd__mux2_1
X_5723_ _5723_/A1 _5723_/A2 _5746_/B1 _6065_/A1 _5722_/X VGND VGND VPWR VPWR _5728_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_31_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5654_ _7148_/Q _7149_/Q VGND VGND VPWR VPWR _5699_/B sky130_fd_sc_hd__and2b_1
X_4605_ _4605_/A _4610_/A _4609_/A VGND VGND VPWR VPWR _4606_/C sky130_fd_sc_hd__or3_1
XFILLER_176_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5585_ _5585_/A0 hold282/X _5586_/S VGND VGND VPWR VPWR _7139_/D sky130_fd_sc_hd__mux2_1
XFILLER_163_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold300 _6952_/Q VGND VGND VPWR VPWR hold300/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 _6614_/Q VGND VGND VPWR VPWR hold311/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_191_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4536_ _4926_/A _4493_/X _4531_/X _4824_/A _4930_/A VGND VGND VPWR VPWR _4536_/Y
+ sky130_fd_sc_hd__a41oi_1
XFILLER_144_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold322 _6519_/Q VGND VGND VPWR VPWR hold322/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold333 _6569_/Q VGND VGND VPWR VPWR hold333/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold344 _6825_/Q VGND VGND VPWR VPWR hold344/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 _6679_/Q VGND VGND VPWR VPWR hold355/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold366 _6736_/Q VGND VGND VPWR VPWR hold366/X sky130_fd_sc_hd__dlygate4sd3_1
X_4467_ _4467_/A _4654_/B _4467_/C VGND VGND VPWR VPWR _4484_/B sky130_fd_sc_hd__or3_2
Xwire3319 _4684_/B VGND VGND VPWR VPWR _4800_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold377 _6731_/Q VGND VGND VPWR VPWR hold377/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold388 _6549_/Q VGND VGND VPWR VPWR hold388/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6206_ _6206_/A1 _6206_/A2 _6206_/B1 _6985_/Q _6205_/X VGND VGND VPWR VPWR _6206_/X
+ sky130_fd_sc_hd__a221o_1
Xhold399 _6709_/Q VGND VGND VPWR VPWR hold399/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire2607 _4823_/A VGND VGND VPWR VPWR _5148_/A sky130_fd_sc_hd__clkbuf_2
X_3418_ _6951_/Q _3418_/A2 wire921/X _6887_/Q VGND VGND VPWR VPWR _3418_/X sky130_fd_sc_hd__a22o_1
X_4398_ _4846_/A _4846_/B _4398_/C VGND VGND VPWR VPWR _4538_/B sky130_fd_sc_hd__and3_4
X_7186_ _7187_/CLK _7186_/D wire3984/X VGND VGND VPWR VPWR _7186_/Q sky130_fd_sc_hd__dfrtp_1
Xwire2618 _6138_/B1 VGND VGND VPWR VPWR _6063_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2629 _6207_/A2 VGND VGND VPWR VPWR _6090_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_58_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1906 _3222_/A VGND VGND VPWR VPWR _6113_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire1917 _6934_/Q VGND VGND VPWR VPWR _6140_/B2 sky130_fd_sc_hd__clkbuf_2
X_3349_ _6505_/Q _4001_/A _3394_/A2 _3349_/B2 VGND VGND VPWR VPWR _3349_/X sky130_fd_sc_hd__a22o_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6137_ _6137_/A1 _6160_/A2 _6137_/B1 _6137_/B2 _6136_/X VGND VGND VPWR VPWR _6142_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1928 wire1929/X VGND VGND VPWR VPWR _5674_/A1 sky130_fd_sc_hd__clkbuf_2
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1939 _6137_/A1 VGND VGND VPWR VPWR wire1939/X sky130_fd_sc_hd__clkbuf_1
XFILLER_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6068_ _6068_/A _6068_/B _6068_/C _6068_/D VGND VGND VPWR VPWR _6068_/X sky130_fd_sc_hd__or4_1
XFILLER_45_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5019_ _5019_/A _5019_/B _5083_/C _5106_/B VGND VGND VPWR VPWR _5030_/A sky130_fd_sc_hd__or4_1
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout3758 hold243/X VGND VGND VPWR VPWR _3963_/B sky130_fd_sc_hd__buf_4
XFILLER_150_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3831 _4547_/A VGND VGND VPWR VPWR _4378_/B sky130_fd_sc_hd__clkbuf_2
Xfanout3769 wire3778/X VGND VGND VPWR VPWR _5593_/B sky130_fd_sc_hd__buf_6
Xwire3842 _4120_/C VGND VGND VPWR VPWR _6440_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_89_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3853 _4533_/A VGND VGND VPWR VPWR _4846_/C sky130_fd_sc_hd__clkbuf_2
Xwire3864 wire3865/X VGND VGND VPWR VPWR wire3864/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3875 wire3876/X VGND VGND VPWR VPWR wire3875/X sky130_fd_sc_hd__clkbuf_1
Xwire3886 input91/X VGND VGND VPWR VPWR _3918_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3897 wire3898/X VGND VGND VPWR VPWR _7213_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_76_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5370_ _5547_/A0 _5735_/B2 _5372_/S VGND VGND VPWR VPWR _6948_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4321_ hold397/X _4321_/A1 _4321_/S VGND VGND VPWR VPWR _6763_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7040_ _7056_/CLK _7040_/D wire3992/X VGND VGND VPWR VPWR _7040_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4252_ _4252_/A _5223_/B VGND VGND VPWR VPWR _4257_/S sky130_fd_sc_hd__and2_2
XFILLER_101_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3203_ _3203_/A VGND VGND VPWR VPWR _3203_/Y sky130_fd_sc_hd__inv_2
X_4183_ _6641_/Q wire363/X _4188_/S VGND VGND VPWR VPWR _6641_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6824_ _6824_/CLK _6824_/D wire3954/X VGND VGND VPWR VPWR _6824_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6755_ _6755_/CLK _6755_/D wire3950/X VGND VGND VPWR VPWR _6755_/Q sky130_fd_sc_hd__dfrtp_1
X_3967_ _3967_/A0 hold152/X _3981_/S VGND VGND VPWR VPWR _3967_/X sky130_fd_sc_hd__mux2_1
X_5706_ _7152_/Q _5706_/B _5706_/C VGND VGND VPWR VPWR _5706_/X sky130_fd_sc_hd__and3_1
XFILLER_50_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6686_ _6705_/CLK _6686_/D wire3959/A VGND VGND VPWR VPWR _6686_/Q sky130_fd_sc_hd__dfrtp_1
X_3898_ _7144_/Q _7145_/Q VGND VGND VPWR VPWR _3899_/B sky130_fd_sc_hd__nor2_1
XFILLER_148_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5637_ _7157_/Q _5637_/B _6039_/A VGND VGND VPWR VPWR _5643_/B sky130_fd_sc_hd__and3_1
XFILLER_148_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5568_ _5568_/A0 hold374/X _5569_/S VGND VGND VPWR VPWR _7124_/D sky130_fd_sc_hd__mux2_1
Xhold130 _6926_/Q VGND VGND VPWR VPWR hold130/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold141 _3258_/X VGND VGND VPWR VPWR hold141/X sky130_fd_sc_hd__dlygate4sd3_1
X_4519_ _4871_/A _4994_/A _4515_/X _4850_/A _4518_/Y VGND VGND VPWR VPWR _4519_/X
+ sky130_fd_sc_hd__o2111a_1
Xhold152 hold725/X VGND VGND VPWR VPWR hold152/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3105 _5739_/B1 VGND VGND VPWR VPWR _5727_/A2 sky130_fd_sc_hd__clkbuf_2
Xhold163 _6547_/Q VGND VGND VPWR VPWR hold163/X sky130_fd_sc_hd__dlygate4sd3_1
X_5499_ _5577_/A0 hold385/X _5499_/S VGND VGND VPWR VPWR _7063_/D sky130_fd_sc_hd__mux2_1
Xhold174 _6551_/Q VGND VGND VPWR VPWR hold174/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3116 _5846_/A2 VGND VGND VPWR VPWR _5831_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold185 _7061_/Q VGND VGND VPWR VPWR hold185/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold196 _7130_/Q VGND VGND VPWR VPWR hold196/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3149 _5824_/A2 VGND VGND VPWR VPWR _5855_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire2415 wire2416/X VGND VGND VPWR VPWR _6214_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_144_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2426 _6501_/Q VGND VGND VPWR VPWR _5755_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire2437 wire2437/A VGND VGND VPWR VPWR _3425_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire2448 wire2448/A VGND VGND VPWR VPWR wire2448/X sky130_fd_sc_hd__clkbuf_1
X_7169_ _7180_/CLK _7169_/D wire3996/X VGND VGND VPWR VPWR _7169_/Q sky130_fd_sc_hd__dfrtp_1
Xwire1703 wire1703/A VGND VGND VPWR VPWR wire1703/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1714 wire1715/X VGND VGND VPWR VPWR _5742_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire2459 _6256_/B1 VGND VGND VPWR VPWR _6057_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire1725 wire1726/X VGND VGND VPWR VPWR _6202_/A1 sky130_fd_sc_hd__clkbuf_2
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1747 wire1748/X VGND VGND VPWR VPWR wire1747/X sky130_fd_sc_hd__clkbuf_1
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1769 _5447_/A1 VGND VGND VPWR VPWR _3351_/B2 sky130_fd_sc_hd__clkbuf_2
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length653 _5440_/S VGND VGND VPWR VPWR _5441_/S sky130_fd_sc_hd__clkbuf_1
XFILLER_154_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout4256 wire4264/A VGND VGND VPWR VPWR _4189_/B sky130_fd_sc_hd__buf_6
XFILLER_38_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout3577 _4242_/A1 VGND VGND VPWR VPWR _4206_/A1 sky130_fd_sc_hd__buf_6
XFILLER_96_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3650 _5224_/A0 VGND VGND VPWR VPWR _4259_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire3661 wire3661/A VGND VGND VPWR VPWR _5545_/A0 sky130_fd_sc_hd__clkbuf_1
Xwire3672 wire3673/X VGND VGND VPWR VPWR wire3672/X sky130_fd_sc_hd__clkbuf_1
Xwire3694 _6293_/C1 VGND VGND VPWR VPWR _5946_/C1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2960 _5791_/B1 VGND VGND VPWR VPWR _5723_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_77_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2971 _5802_/B1 VGND VGND VPWR VPWR _5779_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire2982 wire2983/X VGND VGND VPWR VPWR _5781_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_76_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2993 _5760_/B1 VGND VGND VPWR VPWR _5789_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_92_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4870_ _4931_/B _4870_/B VGND VGND VPWR VPWR _4872_/B sky130_fd_sc_hd__nor2_1
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3821_ hold25/A _3248_/Y _3821_/S VGND VGND VPWR VPWR _3821_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6540_ _7090_/CLK _6540_/D wire3948/X VGND VGND VPWR VPWR _6540_/Q sky130_fd_sc_hd__dfrtp_1
X_3752_ _3752_/A1 _3503_/Y _3733_/X VGND VGND VPWR VPWR _3755_/B sky130_fd_sc_hd__a21o_1
XFILLER_192_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6471_ _6545_/CLK _6471_/D _6426_/X VGND VGND VPWR VPWR _6471_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_185_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3683_ _3683_/A1 wire834/X _5187_/A _6794_/Q wire764/X VGND VGND VPWR VPWR _3683_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_145_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5422_ _5422_/A0 hold587/X _5424_/S VGND VGND VPWR VPWR _6994_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput202 _3200_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[34] sky130_fd_sc_hd__buf_12
Xoutput213 wire1453/X VGND VGND VPWR VPWR mgmt_gpio_out[0] sky130_fd_sc_hd__buf_12
XFILLER_145_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput224 wire1018/X VGND VGND VPWR VPWR mgmt_gpio_out[1] sky130_fd_sc_hd__buf_12
XFILLER_114_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput235 _6556_/Q VGND VGND VPWR VPWR mgmt_gpio_out[2] sky130_fd_sc_hd__buf_12
X_5353_ _5353_/A0 hold576/X _5353_/S VGND VGND VPWR VPWR _6933_/D sky130_fd_sc_hd__mux2_1
XFILLER_126_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput246 _6559_/Q VGND VGND VPWR VPWR mgmt_gpio_out[5] sky130_fd_sc_hd__buf_12
Xoutput257 _3948_/Y VGND VGND VPWR VPWR pad_flash_io0_oeb sky130_fd_sc_hd__buf_12
Xoutput268 _6795_/Q VGND VGND VPWR VPWR pll_div[2] sky130_fd_sc_hd__buf_12
X_4304_ _4304_/A0 hold139/X hold31/X VGND VGND VPWR VPWR _6749_/D sky130_fd_sc_hd__mux2_1
Xoutput279 _6487_/Q VGND VGND VPWR VPWR pll_trim[13] sky130_fd_sc_hd__buf_12
XFILLER_87_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5284_ _5365_/A0 hold100/X _5285_/S VGND VGND VPWR VPWR _6872_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7023_ _7056_/CLK _7023_/D wire3992/X VGND VGND VPWR VPWR _7023_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4235_ _4235_/A0 hold346/X _4239_/S VGND VGND VPWR VPWR _6681_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4166_ _6626_/Q wire359/X _4173_/S VGND VGND VPWR VPWR _6626_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4097_ hold231/X _4096_/X _4097_/S VGND VGND VPWR VPWR _6570_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6807_ _7081_/CLK _6807_/D _7159_/RESET_B VGND VGND VPWR VPWR _6807_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4999_ _4999_/A _4999_/B VGND VGND VPWR VPWR _4999_/Y sky130_fd_sc_hd__nand2_1
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6738_ _6740_/CLK hold23/X fanout4027/X VGND VGND VPWR VPWR _6738_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6669_ _6702_/CLK _6669_/D wire3959/X VGND VGND VPWR VPWR _6669_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2946 _5929_/B1 VGND VGND VPWR VPWR _5950_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_152_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_587 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2201 _6736_/Q VGND VGND VPWR VPWR _3753_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2212 _6723_/Q VGND VGND VPWR VPWR _3621_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2223 wire2223/A VGND VGND VPWR VPWR _3579_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire2234 _6709_/Q VGND VGND VPWR VPWR _5927_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire1500 wire1501/X VGND VGND VPWR VPWR _3729_/B sky130_fd_sc_hd__clkbuf_2
Xwire1511 _3379_/B VGND VGND VPWR VPWR _3485_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2256 _6682_/Q VGND VGND VPWR VPWR _5899_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1522 _3305_/Y VGND VGND VPWR VPWR _3674_/B sky130_fd_sc_hd__clkbuf_2
Xwire2267 wire2268/X VGND VGND VPWR VPWR _6239_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2278 _6667_/Q VGND VGND VPWR VPWR _3623_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_93_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1533 wire1534/X VGND VGND VPWR VPWR _6183_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire2289 _6660_/Q VGND VGND VPWR VPWR _6228_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1544 _6100_/A1 VGND VGND VPWR VPWR wire1544/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1555 wire1555/A VGND VGND VPWR VPWR wire1555/X sky130_fd_sc_hd__clkbuf_1
XFILLER_171_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1566 _7113_/Q VGND VGND VPWR VPWR _6083_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_86_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1577 _7103_/Q VGND VGND VPWR VPWR _6011_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_46_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1588 _7097_/Q VGND VGND VPWR VPWR _6092_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire1599 wire1600/X VGND VGND VPWR VPWR _6189_/A1 sky130_fd_sc_hd__clkbuf_2
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire830 _3460_/Y VGND VGND VPWR VPWR wire830/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_167_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire841 _3426_/X VGND VGND VPWR VPWR wire841/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire852 _3415_/Y VGND VGND VPWR VPWR wire852/X sky130_fd_sc_hd__clkbuf_1
Xwire863 wire864/X VGND VGND VPWR VPWR wire863/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire874 wire875/X VGND VGND VPWR VPWR wire874/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire885 wire886/X VGND VGND VPWR VPWR wire885/X sky130_fd_sc_hd__clkbuf_2
XFILLER_182_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire896 _3335_/Y VGND VGND VPWR VPWR wire896/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout4031 wire4090/X VGND VGND VPWR VPWR _6404_/A sky130_fd_sc_hd__buf_6
XFILLER_155_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout4064 wire4083/X VGND VGND VPWR VPWR wire4066/A sky130_fd_sc_hd__clkbuf_2
XFILLER_170_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire4170 wire4171/X VGND VGND VPWR VPWR wire4170/X sky130_fd_sc_hd__clkbuf_1
Xwire4181 wire4182/X VGND VGND VPWR VPWR _3402_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_69_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4192 wire4193/X VGND VGND VPWR VPWR wire4192/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3480 hold16/X VGND VGND VPWR VPWR _5291_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
X_4020_ _4208_/A1 hold267/X _4021_/S VGND VGND VPWR VPWR _6514_/D sky130_fd_sc_hd__mux2_1
Xwire2790 _6308_/B1 VGND VGND VPWR VPWR _6338_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5971_ _7154_/Q _7153_/Q VGND VGND VPWR VPWR _6039_/C sky130_fd_sc_hd__nor2_2
XFILLER_64_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4922_ _5177_/A _4922_/B _5177_/B _4920_/X VGND VGND VPWR VPWR _4923_/D sky130_fd_sc_hd__or4b_1
XFILLER_33_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4853_ _4683_/A _4707_/B _4447_/Y VGND VGND VPWR VPWR _4860_/C sky130_fd_sc_hd__o21a_1
XFILLER_193_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3804_ _6455_/Q _6454_/Q _6453_/Q VGND VGND VPWR VPWR _3890_/B sky130_fd_sc_hd__or3b_1
XFILLER_159_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4784_ _4784_/A _4784_/B VGND VGND VPWR VPWR _5015_/B sky130_fd_sc_hd__nor2_1
XFILLER_159_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_opt_2_0_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR clkbuf_opt_2_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_16
X_6523_ _7067_/CLK _6523_/D wire3968/X VGND VGND VPWR VPWR _6523_/Q sky130_fd_sc_hd__dfstp_1
X_3735_ _6482_/Q _3735_/A2 _3735_/B1 _3731_/Y VGND VGND VPWR VPWR _3735_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length1508 _3380_/X VGND VGND VPWR VPWR wire1507/A sky130_fd_sc_hd__clkbuf_1
X_6454_ _3945_/A1 _6454_/D _6409_/X VGND VGND VPWR VPWR _6454_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length1519 _3607_/B VGND VGND VPWR VPWR _3731_/B sky130_fd_sc_hd__clkbuf_1
X_3666_ _6063_/A1 _3666_/A2 _3666_/B1 _6061_/B2 wire770/X VGND VGND VPWR VPWR _3669_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_133_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5405_ _5495_/A0 hold301/X _5405_/S VGND VGND VPWR VPWR _6979_/D sky130_fd_sc_hd__mux2_1
X_6385_ _4228_/B _6385_/A2 _6385_/B1 _4228_/Y _6384_/X VGND VGND VPWR VPWR _6385_/X
+ sky130_fd_sc_hd__a221o_1
X_3597_ _3597_/A1 _3597_/A2 wire800/X _3597_/B2 VGND VGND VPWR VPWR _3597_/X sky130_fd_sc_hd__a22o_1
X_5336_ _5585_/A0 hold281/X _5336_/S VGND VGND VPWR VPWR _6918_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5267_ _5561_/A0 hold124/X _5267_/S VGND VGND VPWR VPWR _6857_/D sky130_fd_sc_hd__mux2_1
X_7006_ _7027_/CLK _7006_/D fanout3976/X VGND VGND VPWR VPWR _7006_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_75_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4218_ _5531_/A1 hold332/X _4221_/S VGND VGND VPWR VPWR _6671_/D sky130_fd_sc_hd__mux2_1
X_5198_ _5198_/A0 hold455/X _5199_/S VGND VGND VPWR VPWR _6802_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4149_ _4248_/A0 hold294/X _4152_/S VGND VGND VPWR VPWR _6612_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length3444 hold107/X VGND VGND VPWR VPWR hold108/A sky130_fd_sc_hd__clkbuf_1
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length3455 _5534_/A1 VGND VGND VPWR VPWR _4251_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_164_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2020 _6885_/Q VGND VGND VPWR VPWR wire2020/X sky130_fd_sc_hd__clkbuf_1
Xwire2031 hold75/A VGND VGND VPWR VPWR _6123_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_94_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2042 _6174_/B2 VGND VGND VPWR VPWR _5833_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2053 _6869_/Q VGND VGND VPWR VPWR _6106_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire2064 hold18/A VGND VGND VPWR VPWR _6139_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_93_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1330 _5784_/X VGND VGND VPWR VPWR wire1330/X sky130_fd_sc_hd__clkbuf_1
Xwire2075 hold98/A VGND VGND VPWR VPWR wire2075/X sky130_fd_sc_hd__clkbuf_1
Xwire1341 _4644_/C VGND VGND VPWR VPWR _5095_/A sky130_fd_sc_hd__clkbuf_1
Xwire2086 hold51/A VGND VGND VPWR VPWR wire2086/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1352 wire1353/X VGND VGND VPWR VPWR wire1352/X sky130_fd_sc_hd__clkbuf_1
Xwire2097 _6845_/Q VGND VGND VPWR VPWR _3555_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1363 _3922_/X VGND VGND VPWR VPWR wire1363/X sky130_fd_sc_hd__clkbuf_1
XFILLER_93_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1374 _3477_/A VGND VGND VPWR VPWR _3538_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1385 _3297_/X VGND VGND VPWR VPWR _3482_/A sky130_fd_sc_hd__clkbuf_2
Xwire1396 _3536_/A VGND VGND VPWR VPWR _3331_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_74_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire660 _5416_/S VGND VGND VPWR VPWR _5418_/S sky130_fd_sc_hd__clkbuf_1
X_3520_ _6730_/Q _4276_/A _3692_/A2 _3520_/B2 VGND VGND VPWR VPWR _3520_/X sky130_fd_sc_hd__a22o_1
XFILLER_116_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire671 _5406_/S VGND VGND VPWR VPWR _5409_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_171_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire682 _5376_/Y VGND VGND VPWR VPWR _5381_/S sky130_fd_sc_hd__dlymetal6s2s_1
Xhold707 _7074_/Q VGND VGND VPWR VPWR hold707/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire693 _5351_/S VGND VGND VPWR VPWR _5355_/S sky130_fd_sc_hd__clkbuf_1
Xhold718 _6485_/Q VGND VGND VPWR VPWR hold718/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold729 _7198_/Q VGND VGND VPWR VPWR hold729/X sky130_fd_sc_hd__dlygate4sd3_1
X_3451_ _3451_/A _3478_/B VGND VGND VPWR VPWR _3451_/Y sky130_fd_sc_hd__nor2_1
XFILLER_170_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3382_ _6480_/Q _3420_/A2 _5484_/A _7056_/Q VGND VGND VPWR VPWR _3382_/X sky130_fd_sc_hd__a22o_1
X_6170_ _6170_/A1 _7179_/Q wire450/X VGND VGND VPWR VPWR _6170_/X sky130_fd_sc_hd__a21o_1
XFILLER_130_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_3_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _7093_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_111_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5121_ _5140_/B _5121_/B VGND VGND VPWR VPWR _5139_/B sky130_fd_sc_hd__and2b_1
XFILLER_111_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5052_ _4461_/B _4613_/B _4652_/B _5161_/A2 VGND VGND VPWR VPWR _5052_/X sky130_fd_sc_hd__o22a_1
XFILLER_111_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4003_ _5513_/A0 hold170/X _4003_/S VGND VGND VPWR VPWR _6499_/D sky130_fd_sc_hd__mux2_1
XFILLER_37_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5954_ _6334_/B2 _5954_/A2 _5953_/X VGND VGND VPWR VPWR _5957_/C sky130_fd_sc_hd__a21o_1
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4905_ _4905_/A _4905_/B VGND VGND VPWR VPWR _4925_/B sky130_fd_sc_hd__nand2_1
X_5885_ _6248_/A _5885_/A2 _5885_/B1 _6250_/A1 VGND VGND VPWR VPWR _5885_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4836_ _4836_/A _5001_/B VGND VGND VPWR VPWR _4836_/Y sky130_fd_sc_hd__nand2_1
XFILLER_138_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4767_ _4993_/A _4454_/Y _5049_/B _4983_/B _4766_/X VGND VGND VPWR VPWR _4767_/X
+ sky130_fd_sc_hd__a2111o_1
X_6506_ _7090_/CLK _6506_/D wire3945/A VGND VGND VPWR VPWR _6506_/Q sky130_fd_sc_hd__dfrtp_1
X_3718_ _7120_/Q wire889/X wire852/X _3718_/B2 wire748/X VGND VGND VPWR VPWR _3721_/C
+ sky130_fd_sc_hd__a221o_1
X_4698_ wire2602/X _4698_/B _4698_/C _4698_/D VGND VGND VPWR VPWR _4699_/D sky130_fd_sc_hd__and4b_1
XFILLER_119_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6437_ _6437_/A _6437_/B VGND VGND VPWR VPWR _6437_/X sky130_fd_sc_hd__and2_1
XFILLER_106_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3649_ _6500_/Q _3287_/Y _3547_/Y _3649_/B2 VGND VGND VPWR VPWR _3649_/X sky130_fd_sc_hd__a22o_1
XFILLER_136_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6368_ _6367_/X _7198_/Q _6386_/S VGND VGND VPWR VPWR _7198_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5319_ _5586_/A0 hold598/X _5319_/S VGND VGND VPWR VPWR _6903_/D sky130_fd_sc_hd__mux2_1
X_6299_ _6299_/A1 _6334_/A2 _6299_/B1 _6299_/B2 VGND VGND VPWR VPWR _6299_/X sky130_fd_sc_hd__a22o_1
Xhold12 hold12/A VGND VGND VPWR VPWR hold12/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold23 hold23/A VGND VGND VPWR VPWR hold23/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold34 hold34/A VGND VGND VPWR VPWR hold34/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold45 hold45/A VGND VGND VPWR VPWR hold45/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A VGND VGND VPWR VPWR hold56/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hold67/A VGND VGND VPWR VPWR hold67/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A VGND VGND VPWR VPWR hold78/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold89 hold89/A VGND VGND VPWR VPWR hold89/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_90_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length3263 _5268_/B VGND VGND VPWR VPWR wire3262/A sky130_fd_sc_hd__clkbuf_1
XFILLER_125_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_9 mgmt_gpio_in[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1160 _3452_/A2 VGND VGND VPWR VPWR _3423_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire1171 _3419_/B1 VGND VGND VPWR VPWR _5340_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1182 _3516_/B1 VGND VGND VPWR VPWR _3613_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_35_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1193 wire1194/X VGND VGND VPWR VPWR _3469_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_47_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5670_ _5683_/A _5706_/B _5699_/C VGND VGND VPWR VPWR _5670_/X sky130_fd_sc_hd__and3_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4621_ _4621_/A _4621_/B _4621_/C VGND VGND VPWR VPWR _4621_/X sky130_fd_sc_hd__or3_1
XFILLER_129_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4552_ _4553_/B _4552_/B VGND VGND VPWR VPWR _4792_/B sky130_fd_sc_hd__nor2_1
XFILLER_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold504 _6522_/Q VGND VGND VPWR VPWR hold504/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3503_ _3504_/A _3511_/A VGND VGND VPWR VPWR _3503_/Y sky130_fd_sc_hd__nor2_1
Xhold515 _6858_/Q VGND VGND VPWR VPWR hold515/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire490 _5322_/X VGND VGND VPWR VPWR _5330_/S sky130_fd_sc_hd__buf_2
XFILLER_183_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4483_ _4483_/A VGND VGND VPWR VPWR _5106_/A sky130_fd_sc_hd__inv_2
Xhold526 _6811_/Q VGND VGND VPWR VPWR hold526/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold537 _6760_/Q VGND VGND VPWR VPWR hold537/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold548 _6766_/Q VGND VGND VPWR VPWR hold548/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6222_ _6222_/A _6272_/B VGND VGND VPWR VPWR _6222_/X sky130_fd_sc_hd__and2_1
Xhold559 _7073_/Q VGND VGND VPWR VPWR hold559/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3434_ _6149_/A1 _5520_/A _5349_/A _6163_/B2 VGND VGND VPWR VPWR _3434_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6153_ _6153_/A1 _6175_/A2 _6153_/B1 _6911_/Q _6152_/X VGND VGND VPWR VPWR _6156_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3365_ _6212_/A1 _3386_/A2 _3419_/B1 _3365_/B2 VGND VGND VPWR VPWR _3365_/X sky130_fd_sc_hd__a22o_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5104_ _5104_/A _5104_/B _5104_/C _5104_/D VGND VGND VPWR VPWR _5104_/X sky130_fd_sc_hd__or4_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6084_ _6084_/A _6084_/B _6084_/C _6084_/D VGND VGND VPWR VPWR _6085_/B sky130_fd_sc_hd__or4_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3296_ _3320_/A _3331_/A VGND VGND VPWR VPWR _3296_/Y sky130_fd_sc_hd__nor2_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5035_ _5035_/A _5035_/B VGND VGND VPWR VPWR _5035_/Y sky130_fd_sc_hd__nand2_1
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6986_ _7027_/CLK _6986_/D fanout3976/X VGND VGND VPWR VPWR _6986_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_80_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5937_ _6311_/B2 _5953_/A2 _5965_/A2 _6300_/B2 _5936_/X VGND VGND VPWR VPWR _5945_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5868_ _6239_/B2 _5868_/A2 _5936_/B1 _6237_/B2 _5867_/X VGND VGND VPWR VPWR _5869_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_139_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4819_ _4544_/X _4981_/C _4819_/C _4819_/D VGND VGND VPWR VPWR _4821_/C sky130_fd_sc_hd__and4bb_1
X_5799_ _6151_/B2 _5799_/A2 _5799_/B1 _6149_/A1 _5798_/X VGND VGND VPWR VPWR _5799_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_154_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput102 wb_adr_i[12] VGND VGND VPWR VPWR _4338_/B sky130_fd_sc_hd__clkbuf_1
Xinput113 wb_adr_i[22] VGND VGND VPWR VPWR _4390_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput124 wb_adr_i[3] VGND VGND VPWR VPWR _4570_/C sky130_fd_sc_hd__buf_6
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput135 wb_dat_i[12] VGND VGND VPWR VPWR _6376_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_193_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput146 wb_dat_i[22] VGND VGND VPWR VPWR _6382_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput157 wb_dat_i[3] VGND VGND VPWR VPWR _6373_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput168 wb_sel_i[3] VGND VGND VPWR VPWR _6357_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_56_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_83_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6799_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_39_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6840_ _6973_/CLK _6840_/D fanout4078/X VGND VGND VPWR VPWR _6840_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_62_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6771_ _6824_/CLK _6771_/D fanout3973/X VGND VGND VPWR VPWR _6771_/Q sky130_fd_sc_hd__dfrtp_1
X_3983_ _3983_/A _5430_/B VGND VGND VPWR VPWR _3991_/S sky130_fd_sc_hd__and2_1
XFILLER_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5722_ _6063_/B2 _5722_/A2 _5744_/B2 _6971_/Q _5722_/C1 VGND VGND VPWR VPWR _5722_/X
+ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_21_csclk _6579_/CLK VGND VGND VPWR VPWR _7135_/CLK sky130_fd_sc_hd__clkbuf_16
X_5653_ _7151_/Q _7150_/Q VGND VGND VPWR VPWR _5700_/C sky130_fd_sc_hd__and2b_1
XFILLER_30_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4604_ _4342_/C _4819_/D _4793_/A VGND VGND VPWR VPWR _4606_/B sky130_fd_sc_hd__a21o_1
XFILLER_148_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5584_ _5584_/A0 hold192/X _5586_/S VGND VGND VPWR VPWR _7138_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_36_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7140_/CLK sky130_fd_sc_hd__clkbuf_16
X_4535_ _4745_/A _4535_/B VGND VGND VPWR VPWR _4824_/A sky130_fd_sc_hd__or2_1
Xhold301 _6979_/Q VGND VGND VPWR VPWR hold301/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 _6892_/Q VGND VGND VPWR VPWR hold312/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 _4026_/X VGND VGND VPWR VPWR _6519_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 _6684_/Q VGND VGND VPWR VPWR hold334/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold345 _6761_/Q VGND VGND VPWR VPWR hold345/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4466_ _4846_/C _4951_/B VGND VGND VPWR VPWR _4493_/B sky130_fd_sc_hd__nand2_1
Xwire3309 _5074_/A2 VGND VGND VPWR VPWR _4686_/B sky130_fd_sc_hd__clkbuf_1
Xhold356 _6715_/Q VGND VGND VPWR VPWR hold356/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 _6726_/Q VGND VGND VPWR VPWR hold367/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 _6734_/Q VGND VGND VPWR VPWR hold378/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold389 _6855_/Q VGND VGND VPWR VPWR hold389/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6205_ _6205_/A1 _6205_/A2 _6205_/B1 _6205_/B2 VGND VGND VPWR VPWR _6205_/X sky130_fd_sc_hd__a22o_1
X_3417_ _3417_/A _3456_/B VGND VGND VPWR VPWR _3417_/Y sky130_fd_sc_hd__nor2_2
Xwire2608 _4462_/Y VGND VGND VPWR VPWR _4955_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
X_7185_ _7185_/CLK _7185_/D _7185_/RESET_B VGND VGND VPWR VPWR _7185_/Q sky130_fd_sc_hd__dfrtp_1
X_4397_ _4397_/A _4667_/B VGND VGND VPWR VPWR _4484_/A sky130_fd_sc_hd__nand2_1
XFILLER_98_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2619 _6173_/B1 VGND VGND VPWR VPWR _6138_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6136_ _6918_/Q _6136_/A2 _6159_/B1 _6942_/Q VGND VGND VPWR VPWR _6136_/X sky130_fd_sc_hd__a22o_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3348_ _6993_/Q _3387_/A2 _3426_/B1 _7057_/Q wire857/X VGND VGND VPWR VPWR _3355_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1907 hold97/A VGND VGND VPWR VPWR _3222_/A sky130_fd_sc_hd__clkbuf_2
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1918 _6933_/Q VGND VGND VPWR VPWR _6104_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1929 _6930_/Q VGND VGND VPWR VPWR wire1929/X sky130_fd_sc_hd__clkbuf_1
XFILLER_97_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6067_ _6867_/Q _6067_/A2 _6078_/A2 _6067_/B2 _6066_/X VGND VGND VPWR VPWR _6068_/D
+ sky130_fd_sc_hd__a221o_1
X_3279_ hold62/X hold27/X VGND VGND VPWR VPWR _3451_/A sky130_fd_sc_hd__or2_1
XFILLER_39_761 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5018_ _5018_/A _5023_/C _5018_/C VGND VGND VPWR VPWR _5106_/B sky130_fd_sc_hd__nor3_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6969_ _7088_/CLK _6969_/D wire4069/A VGND VGND VPWR VPWR _6969_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_41_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length879 _3338_/Y VGND VGND VPWR VPWR wire878/A sky130_fd_sc_hd__clkbuf_1
XFILLER_135_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3810 _5023_/B VGND VGND VPWR VPWR _4660_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3821 wire3822/X VGND VGND VPWR VPWR _4611_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3843 wire3844/X VGND VGND VPWR VPWR _4120_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_110_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3854 _4667_/C VGND VGND VPWR VPWR _4451_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_1_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3865 wire3866/X VGND VGND VPWR VPWR wire3865/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3876 wire3877/X VGND VGND VPWR VPWR wire3876/X sky130_fd_sc_hd__clkbuf_1
XFILLER_150_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3887 wire3888/X VGND VGND VPWR VPWR _3921_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3898 wire3899/X VGND VGND VPWR VPWR wire3898/X sky130_fd_sc_hd__clkbuf_1
XFILLER_67_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4320_ hold502/X _5504_/A0 _4321_/S VGND VGND VPWR VPWR _6762_/D sky130_fd_sc_hd__mux2_1
XFILLER_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4251_ _4251_/A0 hold224/X _4251_/S VGND VGND VPWR VPWR _6705_/D sky130_fd_sc_hd__mux2_1
X_3202_ _3202_/A VGND VGND VPWR VPWR _3202_/Y sky130_fd_sc_hd__inv_2
X_4182_ _6640_/Q wire360/X _4188_/S VGND VGND VPWR VPWR _6640_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6823_ _7075_/CLK _6823_/D wire4041/X VGND VGND VPWR VPWR _6823_/Q sky130_fd_sc_hd__dfrtp_1
X_6754_ _6825_/CLK _6754_/D wire3954/X VGND VGND VPWR VPWR _6754_/Q sky130_fd_sc_hd__dfrtp_1
X_3966_ _3966_/A _5430_/B VGND VGND VPWR VPWR _3982_/S sky130_fd_sc_hd__and2_1
XFILLER_176_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5705_ _5705_/A _5705_/B _5706_/C VGND VGND VPWR VPWR _5705_/X sky130_fd_sc_hd__and3_1
X_6685_ _6702_/CLK _6685_/D _6685_/RESET_B VGND VGND VPWR VPWR _6685_/Q sky130_fd_sc_hd__dfrtp_1
X_3897_ _5615_/A _5590_/A2 _3896_/X VGND VGND VPWR VPWR _6562_/D sky130_fd_sc_hd__o21ai_1
XFILLER_176_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5636_ _7156_/Q _5624_/B _5634_/Y _5635_/X VGND VGND VPWR VPWR _7156_/D sky130_fd_sc_hd__a31o_1
XFILLER_191_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5567_ _5567_/A0 hold250/X _5570_/S VGND VGND VPWR VPWR _7123_/D sky130_fd_sc_hd__mux2_1
XFILLER_163_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold120 _5498_/X VGND VGND VPWR VPWR _7062_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 _6870_/Q VGND VGND VPWR VPWR hold131/X sky130_fd_sc_hd__dlygate4sd3_1
X_4518_ _5124_/A VGND VGND VPWR VPWR _4518_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold142 _3519_/Y VGND VGND VPWR VPWR _4141_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold153 hold726/X VGND VGND VPWR VPWR hold153/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5498_ _5498_/A0 _7062_/Q _5498_/S VGND VGND VPWR VPWR _5498_/X sky130_fd_sc_hd__mux2_1
Xwire3106 _5781_/A2 VGND VGND VPWR VPWR _5739_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_132_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3117 _5756_/A2 VGND VGND VPWR VPWR _5846_/A2 sky130_fd_sc_hd__clkbuf_1
Xhold164 _6838_/Q VGND VGND VPWR VPWR hold164/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 _4065_/X VGND VGND VPWR VPWR _6551_/D sky130_fd_sc_hd__dlygate4sd3_1
Xwire3128 wire3129/X VGND VGND VPWR VPWR _5841_/A2 sky130_fd_sc_hd__clkbuf_2
Xhold186 _6939_/Q VGND VGND VPWR VPWR hold186/X sky130_fd_sc_hd__dlygate4sd3_1
X_4449_ _4932_/A _4742_/A _4836_/A VGND VGND VPWR VPWR _4502_/A sky130_fd_sc_hd__and3b_1
Xhold197 _7202_/Q VGND VGND VPWR VPWR hold197/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3139 _5827_/A2 VGND VGND VPWR VPWR _5853_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire2405 _6511_/Q VGND VGND VPWR VPWR _3766_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire2416 wire2417/X VGND VGND VPWR VPWR wire2416/X sky130_fd_sc_hd__clkbuf_1
X_7168_ _3937_/A1 _7168_/D wire4001/X VGND VGND VPWR VPWR _7168_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_132_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1715 wire1716/X VGND VGND VPWR VPWR wire1715/X sky130_fd_sc_hd__clkbuf_1
Xwire1726 _7033_/Q VGND VGND VPWR VPWR wire1726/X sky130_fd_sc_hd__clkbuf_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6119_ _6119_/A _6119_/B _6119_/C _6119_/D VGND VGND VPWR VPWR _6119_/X sky130_fd_sc_hd__or4_1
XFILLER_100_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1737 _3685_/A1 VGND VGND VPWR VPWR _6049_/A sky130_fd_sc_hd__clkbuf_1
Xwire1748 wire1749/X VGND VGND VPWR VPWR wire1748/X sky130_fd_sc_hd__clkbuf_1
X_7099_ _7137_/CLK _7099_/D wire4007/X VGND VGND VPWR VPWR _7099_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_100_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1759 _5739_/B2 VGND VGND VPWR VPWR _6074_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_73_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length665 _5417_/S VGND VGND VPWR VPWR _5413_/S sky130_fd_sc_hd__clkbuf_1
XFILLER_182_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length687 _5369_/S VGND VGND VPWR VPWR _5372_/S sky130_fd_sc_hd__clkbuf_2
Xfanout3512 wire3523/A VGND VGND VPWR VPWR _5479_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_135_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout3534 _4249_/A0 VGND VGND VPWR VPWR _5532_/A1 sky130_fd_sc_hd__buf_6
XFILLER_135_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout3556 _5343_/A0 VGND VGND VPWR VPWR _5574_/A0 sky130_fd_sc_hd__buf_6
XFILLER_78_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3640 wire3641/X VGND VGND VPWR VPWR _5251_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_150_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3651 _5563_/A0 VGND VGND VPWR VPWR _5224_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3662 wire3663/X VGND VGND VPWR VPWR wire3662/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3673 wire3674/X VGND VGND VPWR VPWR wire3673/X sky130_fd_sc_hd__clkbuf_1
XFILLER_78_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3684 wire3685/X VGND VGND VPWR VPWR _5894_/B sky130_fd_sc_hd__clkbuf_1
Xwire3695 _6318_/S VGND VGND VPWR VPWR _6293_/C1 sky130_fd_sc_hd__clkbuf_2
Xwire2950 _5788_/B1 VGND VGND VPWR VPWR _5734_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2961 _5798_/B1 VGND VGND VPWR VPWR _5791_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2972 _5851_/A2 VGND VGND VPWR VPWR _5802_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2983 _5683_/X VGND VGND VPWR VPWR wire2983/X sky130_fd_sc_hd__clkbuf_1
XFILLER_94_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2994 _5843_/B1 VGND VGND VPWR VPWR _5760_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3820_ _3820_/A _3823_/B VGND VGND VPWR VPWR _3820_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3751_ _3751_/A1 wire901/X wire882/X _3751_/B2 _3750_/X VGND VGND VPWR VPWR _3751_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_9_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6470_ _6545_/CLK _6470_/D _6425_/X VGND VGND VPWR VPWR _6470_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3682_ input12/X _3682_/A2 _3682_/B1 input21/X VGND VGND VPWR VPWR _3682_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5421_ _5421_/A _5535_/B VGND VGND VPWR VPWR _5429_/S sky130_fd_sc_hd__nand2_2
XFILLER_161_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput203 wire1356/X VGND VGND VPWR VPWR mgmt_gpio_oeb[35] sky130_fd_sc_hd__buf_12
X_5352_ _5352_/A0 hold461/X _5354_/S VGND VGND VPWR VPWR _6932_/D sky130_fd_sc_hd__mux2_1
Xoutput214 _3926_/X VGND VGND VPWR VPWR mgmt_gpio_out[10] sky130_fd_sc_hd__buf_12
Xoutput225 _6550_/Q VGND VGND VPWR VPWR mgmt_gpio_out[20] sky130_fd_sc_hd__buf_12
XFILLER_99_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput236 _6832_/Q VGND VGND VPWR VPWR mgmt_gpio_out[30] sky130_fd_sc_hd__buf_12
XFILLER_99_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput247 wire1458/X VGND VGND VPWR VPWR mgmt_gpio_out[6] sky130_fd_sc_hd__buf_12
XFILLER_114_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput258 _7213_/X VGND VGND VPWR VPWR pad_flash_io1_do sky130_fd_sc_hd__buf_12
X_4303_ hold22/X _6748_/Q hold31/X VGND VGND VPWR VPWR hold32/A sky130_fd_sc_hd__mux2_1
XFILLER_153_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5283_ _5481_/A0 hold636/X _5285_/S VGND VGND VPWR VPWR _6871_/D sky130_fd_sc_hd__mux2_1
Xoutput269 _6796_/Q VGND VGND VPWR VPWR pll_div[3] sky130_fd_sc_hd__buf_12
XFILLER_87_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7022_ _7027_/CLK _7022_/D fanout3976/X VGND VGND VPWR VPWR _7022_/Q sky130_fd_sc_hd__dfrtp_1
X_4234_ _4234_/A _4234_/B VGND VGND VPWR VPWR _4239_/S sky130_fd_sc_hd__nand2_2
XFILLER_101_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4165_ _6695_/Q _6348_/B VGND VGND VPWR VPWR _4170_/S sky130_fd_sc_hd__and2_1
XFILLER_95_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4096_ hold164/X _5246_/A0 _4100_/S VGND VGND VPWR VPWR _4096_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6806_ _7036_/CLK _6806_/D wire3974/X VGND VGND VPWR VPWR _6806_/Q sky130_fd_sc_hd__dfstp_1
X_4998_ _4999_/A _4450_/Y _4741_/C _4734_/Y _4894_/C VGND VGND VPWR VPWR _5045_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_168_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3949_ _6459_/Q _3949_/B VGND VGND VPWR VPWR _3950_/A sky130_fd_sc_hd__or2_2
X_6737_ _6979_/CLK _6737_/D fanout4027/X VGND VGND VPWR VPWR _6737_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length3637 _5536_/A1 VGND VGND VPWR VPWR _5485_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_109_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6668_ _6702_/CLK _6668_/D _6685_/RESET_B VGND VGND VPWR VPWR _6668_/Q sky130_fd_sc_hd__dfrtp_1
Xmax_length3659 _5350_/A0 VGND VGND VPWR VPWR wire3656/A sky130_fd_sc_hd__clkbuf_1
XFILLER_176_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5619_ _5622_/B VGND VGND VPWR VPWR _5619_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6599_ _7090_/CLK _6599_/D wire3948/X VGND VGND VPWR VPWR _6599_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_164_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length2969 _5851_/A2 VGND VGND VPWR VPWR wire2968/A sky130_fd_sc_hd__clkbuf_1
XFILLER_152_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2202 _6735_/Q VGND VGND VPWR VPWR _6334_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_105_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2213 _6722_/Q VGND VGND VPWR VPWR _6256_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2224 wire2225/X VGND VGND VPWR VPWR _5938_/A sky130_fd_sc_hd__clkbuf_2
Xwire2235 _6708_/Q VGND VGND VPWR VPWR _3625_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_120_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1501 _3414_/Y VGND VGND VPWR VPWR wire1501/X sky130_fd_sc_hd__clkbuf_1
Xwire2246 _6702_/Q VGND VGND VPWR VPWR _5900_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1512 _3472_/B VGND VGND VPWR VPWR _3379_/B sky130_fd_sc_hd__clkbuf_2
Xwire2257 wire2258/X VGND VGND VPWR VPWR _6235_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire1523 _3303_/Y VGND VGND VPWR VPWR _3528_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2268 _6675_/Q VGND VGND VPWR VPWR wire2268/X sky130_fd_sc_hd__clkbuf_1
Xwire2279 _6665_/Q VGND VGND VPWR VPWR _6235_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1534 wire1535/X VGND VGND VPWR VPWR wire1534/X sky130_fd_sc_hd__clkbuf_1
Xwire1545 _7130_/Q VGND VGND VPWR VPWR _6100_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_74_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1567 _7111_/Q VGND VGND VPWR VPWR _3748_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_171_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1578 _7102_/Q VGND VGND VPWR VPWR _6208_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1589 wire1590/X VGND VGND VPWR VPWR _6050_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_46_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire820 wire820/A VGND VGND VPWR VPWR wire820/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_167_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire831 _3457_/X VGND VGND VPWR VPWR wire831/X sky130_fd_sc_hd__clkbuf_1
Xwire842 wire843/X VGND VGND VPWR VPWR wire842/X sky130_fd_sc_hd__clkbuf_1
XFILLER_127_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire864 _3343_/Y VGND VGND VPWR VPWR wire864/X sky130_fd_sc_hd__clkbuf_2
XFILLER_182_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire875 _3338_/Y VGND VGND VPWR VPWR wire875/X sky130_fd_sc_hd__dlymetal6s2s_1
Xwire886 wire887/X VGND VGND VPWR VPWR wire886/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length473 _5569_/S VGND VGND VPWR VPWR _5570_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_182_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout4043 wire4080/X VGND VGND VPWR VPWR wire4046/A sky130_fd_sc_hd__buf_6
Xmax_length495 _5320_/S VGND VGND VPWR VPWR _5317_/S sky130_fd_sc_hd__clkbuf_2
Xfanout4054 fanout4054/A VGND VGND VPWR VPWR wire4056/A sky130_fd_sc_hd__buf_6
XFILLER_123_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout4087 wire4094/X VGND VGND VPWR VPWR wire4092/A sky130_fd_sc_hd__buf_6
Xwire4160 _3926_/A1 VGND VGND VPWR VPWR wire4160/X sky130_fd_sc_hd__clkbuf_1
Xwire4171 input55/X VGND VGND VPWR VPWR wire4171/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4182 wire4183/X VGND VGND VPWR VPWR wire4182/X sky130_fd_sc_hd__clkbuf_1
Xwire4193 wire4194/X VGND VGND VPWR VPWR wire4193/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3470 _4116_/A0 VGND VGND VPWR VPWR _5576_/A0 sky130_fd_sc_hd__clkbuf_2
Xwire3481 wire3482/X VGND VGND VPWR VPWR _5498_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_84_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2780 _6163_/B1 VGND VGND VPWR VPWR _6081_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire2791 _6029_/B VGND VGND VPWR VPWR _6308_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_92_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5970_ _7174_/Q wire397/X _5970_/S VGND VGND VPWR VPWR _7174_/D sky130_fd_sc_hd__mux2_1
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4921_ _4674_/A _4684_/A _4622_/Y _4635_/Y VGND VGND VPWR VPWR _4922_/B sky130_fd_sc_hd__a31o_1
XFILLER_33_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4852_ _4674_/A _4684_/A _4595_/B _4506_/Y VGND VGND VPWR VPWR _4862_/B sky130_fd_sc_hd__a31o_1
XFILLER_33_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3803_ _6471_/Q _3838_/B VGND VGND VPWR VPWR _3890_/A sky130_fd_sc_hd__nand2_1
X_4783_ _4783_/A _4802_/D VGND VGND VPWR VPWR _4783_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6522_ _7067_/CLK _6522_/D wire3968/X VGND VGND VPWR VPWR _6522_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3734_ _7026_/Q _3326_/Y _5203_/A _6806_/Q VGND VGND VPWR VPWR _3734_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6453_ _3945_/A1 _6453_/D _6408_/X VGND VGND VPWR VPWR _6453_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3665_ _6258_/B2 _3665_/A2 _3665_/B1 _3665_/B2 VGND VGND VPWR VPWR _3665_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5404_ _5554_/A0 hold320/X _5404_/S VGND VGND VPWR VPWR _6978_/D sky130_fd_sc_hd__mux2_1
XFILLER_134_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6384_ _4228_/C _6384_/A2 _6384_/B1 _4228_/A VGND VGND VPWR VPWR _6384_/X sky130_fd_sc_hd__a22o_1
X_3596_ _3596_/A1 _3596_/A2 _3596_/B1 _3596_/B2 wire780/X VGND VGND VPWR VPWR _3600_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5335_ _5353_/A0 hold519/X _5339_/S VGND VGND VPWR VPWR _6917_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5266_ _5365_/A0 hold98/X _5267_/S VGND VGND VPWR VPWR _6856_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7005_ _7027_/CLK _7005_/D fanout3976/X VGND VGND VPWR VPWR _7005_/Q sky130_fd_sc_hd__dfrtp_1
X_4217_ _4223_/A0 hold331/X _4221_/S VGND VGND VPWR VPWR _6670_/D sky130_fd_sc_hd__mux2_1
X_5197_ _5197_/A0 hold451/X _5199_/S VGND VGND VPWR VPWR _6801_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4148_ _4247_/A0 hold306/X _4152_/S VGND VGND VPWR VPWR _6611_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4079_ hold609/X _5309_/A0 _4079_/S VGND VGND VPWR VPWR _4079_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3401 _5374_/A0 VGND VGND VPWR VPWR _5392_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3456 _5534_/A1 VGND VGND VPWR VPWR _4215_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_137_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length2733 _6086_/A2 VGND VGND VPWR VPWR _6132_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_180_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length2766 _6202_/A2 VGND VGND VPWR VPWR wire2765/A sky130_fd_sc_hd__clkbuf_1
XFILLER_166_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2010 _6035_/B2 VGND VGND VPWR VPWR _5657_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2021 _6883_/Q VGND VGND VPWR VPWR _6064_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2032 wire2033/X VGND VGND VPWR VPWR _3230_/A sky130_fd_sc_hd__clkbuf_1
Xwire2043 _6872_/Q VGND VGND VPWR VPWR _6174_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire1320 _5993_/X VGND VGND VPWR VPWR wire1320/X sky130_fd_sc_hd__clkbuf_1
Xwire2065 wire2065/A VGND VGND VPWR VPWR _3231_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_120_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2076 _6855_/Q VGND VGND VPWR VPWR _6164_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1331 wire1332/X VGND VGND VPWR VPWR _5785_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_115_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1342 _4599_/X VGND VGND VPWR VPWR _4600_/C1 sky130_fd_sc_hd__clkbuf_1
XFILLER_47_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1353 _3935_/X VGND VGND VPWR VPWR wire1353/X sky130_fd_sc_hd__clkbuf_1
Xwire2098 _6845_/Q VGND VGND VPWR VPWR _6120_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire1364 wire1365/X VGND VGND VPWR VPWR wire1364/X sky130_fd_sc_hd__clkbuf_2
XFILLER_46_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1375 hold63/X VGND VGND VPWR VPWR _3477_/A sky130_fd_sc_hd__clkbuf_1
Xwire1386 _3507_/B VGND VGND VPWR VPWR _3476_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1397 _3281_/X VGND VGND VPWR VPWR _3536_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_61_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_670 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire650 wire651/X VGND VGND VPWR VPWR _5446_/S sky130_fd_sc_hd__clkbuf_1
XFILLER_128_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire661 wire661/A VGND VGND VPWR VPWR _5416_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_183_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire672 _5404_/S VGND VGND VPWR VPWR _5405_/S sky130_fd_sc_hd__clkbuf_1
Xhold708 _6487_/Q VGND VGND VPWR VPWR hold708/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire683 wire684/X VGND VGND VPWR VPWR _5384_/S sky130_fd_sc_hd__clkbuf_2
Xhold719 _6482_/Q VGND VGND VPWR VPWR hold719/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire694 wire694/A VGND VGND VPWR VPWR _5351_/S sky130_fd_sc_hd__clkbuf_1
XFILLER_183_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3450_ _3510_/A _3607_/B VGND VGND VPWR VPWR _3450_/Y sky130_fd_sc_hd__nor2_1
XFILLER_143_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3381_ _6976_/Q _5394_/A wire870/X _3381_/B2 VGND VGND VPWR VPWR _3381_/X sky130_fd_sc_hd__a22o_1
X_5120_ _5171_/A _5172_/A _5119_/Y VGND VGND VPWR VPWR _5121_/B sky130_fd_sc_hd__or3b_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5051_ _5044_/X _5048_/X wire400/X VGND VGND VPWR VPWR _5104_/A sky130_fd_sc_hd__o21a_1
XFILLER_85_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4002_ _5536_/A1 hold673/X _4004_/S VGND VGND VPWR VPWR _6498_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5953_ _6337_/B2 _5953_/A2 _5953_/B1 _6705_/Q VGND VGND VPWR VPWR _5953_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4904_ _4633_/B _4589_/B _4902_/X _4638_/A _4903_/X VGND VGND VPWR VPWR _4905_/B
+ sky130_fd_sc_hd__o221a_1
X_5884_ _6707_/Q _5927_/B1 _5959_/B1 _6265_/A1 _5883_/X VGND VGND VPWR VPWR _5891_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_60_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4835_ _4932_/A _4835_/B VGND VGND VPWR VPWR _4857_/A sky130_fd_sc_hd__or2_1
XFILLER_178_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4766_ _4993_/A _4516_/B _4815_/A _4987_/B _4765_/X VGND VGND VPWR VPWR _4766_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_193_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6505_ _7056_/CLK _6505_/D wire3992/X VGND VGND VPWR VPWR _6505_/Q sky130_fd_sc_hd__dfrtp_1
X_3717_ _6475_/Q _3782_/A2 _3735_/A2 _6483_/Q VGND VGND VPWR VPWR _3717_/X sky130_fd_sc_hd__a22o_1
XFILLER_147_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4697_ _4693_/C _4683_/B _4696_/X _4653_/X VGND VGND VPWR VPWR _4698_/D sky130_fd_sc_hd__o211a_1
XFILLER_107_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3648_ _3648_/A1 _3450_/Y _3496_/Y _6293_/A1 _3647_/X VGND VGND VPWR VPWR _3651_/C
+ sky130_fd_sc_hd__a221o_1
X_6436_ _6437_/A _6437_/B VGND VGND VPWR VPWR _6436_/X sky130_fd_sc_hd__and2_1
XFILLER_106_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6367_ _4228_/B _6367_/A2 _6367_/B1 _4228_/Y _6366_/X VGND VGND VPWR VPWR _6367_/X
+ sky130_fd_sc_hd__a221o_1
X_3579_ _3579_/A1 wire970/X _3579_/B1 _3579_/B2 _3578_/X VGND VGND VPWR VPWR _3582_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5318_ _5489_/A0 hold456/X _5318_/S VGND VGND VPWR VPWR _6902_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6298_ _7093_/Q _6298_/A2 _6298_/B1 _6298_/B2 VGND VGND VPWR VPWR _6298_/X sky130_fd_sc_hd__a22o_1
XFILLER_114_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold13 hold13/A VGND VGND VPWR VPWR hold13/X sky130_fd_sc_hd__dlygate4sd3_1
X_5249_ hold3/X _6841_/Q _5249_/S VGND VGND VPWR VPWR hold9/A sky130_fd_sc_hd__mux2_1
Xhold24 hold24/A VGND VGND VPWR VPWR hold24/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 hold35/A VGND VGND VPWR VPWR hold35/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold46 hold46/A VGND VGND VPWR VPWR hold46/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold57 hold57/A VGND VGND VPWR VPWR hold57/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 hold68/A VGND VGND VPWR VPWR hold68/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold79 hold79/A VGND VGND VPWR VPWR hold79/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_68_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3264 _5502_/B VGND VGND VPWR VPWR _5268_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_165_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1150 _3328_/Y VGND VGND VPWR VPWR _3561_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1161 _3645_/A2 VGND VGND VPWR VPWR _3452_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire1172 _3738_/B1 VGND VGND VPWR VPWR _3419_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire1183 _3516_/B1 VGND VGND VPWR VPWR _5385_/A sky130_fd_sc_hd__clkbuf_1
Xwire1194 _3736_/A2 VGND VGND VPWR VPWR wire1194/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_721 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4620_ _4620_/A _4635_/B VGND VGND VPWR VPWR _5115_/B sky130_fd_sc_hd__nor2_1
XFILLER_148_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4551_ _4341_/X _4819_/D _4476_/A VGND VGND VPWR VPWR _4552_/B sky130_fd_sc_hd__a21oi_1
XFILLER_156_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3502_ _3518_/A _3502_/B VGND VGND VPWR VPWR _3502_/Y sky130_fd_sc_hd__nor2_1
Xwire480 _5553_/Y VGND VGND VPWR VPWR _5561_/S sky130_fd_sc_hd__clkbuf_2
Xhold505 _7000_/Q VGND VGND VPWR VPWR hold505/X sky130_fd_sc_hd__dlygate4sd3_1
X_4482_ _4596_/A _4482_/B VGND VGND VPWR VPWR _4483_/A sky130_fd_sc_hd__or2_1
Xhold516 _7094_/Q VGND VGND VPWR VPWR hold516/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire491 _5321_/S VGND VGND VPWR VPWR _5314_/S sky130_fd_sc_hd__clkbuf_1
XFILLER_128_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold527 _6966_/Q VGND VGND VPWR VPWR hold527/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold538 _7065_/Q VGND VGND VPWR VPWR hold538/X sky130_fd_sc_hd__dlygate4sd3_1
X_6221_ _6726_/Q _6296_/A2 _6296_/B1 _6221_/B2 VGND VGND VPWR VPWR _6221_/X sky130_fd_sc_hd__a22o_1
Xhold549 _6768_/Q VGND VGND VPWR VPWR hold549/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3433_ _6163_/A1 _3433_/A2 _3557_/B1 _6155_/B2 _3432_/X VGND VGND VPWR VPWR _3447_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_171_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6152_ _6152_/A1 _6152_/A2 _6152_/B1 _6152_/B2 VGND VGND VPWR VPWR _6152_/X sky130_fd_sc_hd__a22o_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ _7025_/Q _3364_/A2 wire868/X _7110_/Q _3363_/X VGND VGND VPWR VPWR _3372_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5103_ _5103_/A _5103_/B VGND VGND VPWR VPWR _5104_/D sky130_fd_sc_hd__nor2_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _6948_/Q _6138_/A2 _6102_/A2 _6083_/B2 _6082_/X VGND VGND VPWR VPWR _6084_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3295_ _3344_/A _3339_/B VGND VGND VPWR VPWR _3295_/Y sky130_fd_sc_hd__nor2_1
XFILLER_97_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _4962_/Y _4991_/Y _5033_/X _5034_/B1 _6778_/Q VGND VGND VPWR VPWR _6778_/D
+ sky130_fd_sc_hd__o32a_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6985_ _7102_/CLK _6985_/D wire4004/A VGND VGND VPWR VPWR _6985_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_41_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5936_ _6624_/Q _5936_/A2 _5936_/B1 _6312_/B2 VGND VGND VPWR VPWR _5936_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5867_ _6225_/B2 _5918_/A2 _5932_/A2 _6228_/A1 VGND VGND VPWR VPWR _5867_/X sky130_fd_sc_hd__a22o_1
XFILLER_33_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4818_ _4818_/A _4818_/B _4618_/C VGND VGND VPWR VPWR _4818_/X sky130_fd_sc_hd__or3b_1
X_5798_ _6148_/A _5798_/A2 _5798_/B1 _6150_/B2 _5797_/X VGND VGND VPWR VPWR _5798_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_193_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4749_ _4638_/B _4749_/B _4749_/C VGND VGND VPWR VPWR _4965_/B sky130_fd_sc_hd__and3b_1
XFILLER_134_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6419_ _6429_/A _6432_/B VGND VGND VPWR VPWR _6419_/X sky130_fd_sc_hd__and2_1
Xmax_length1169 _3612_/A2 VGND VGND VPWR VPWR wire1168/A sky130_fd_sc_hd__clkbuf_1
XFILLER_162_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput103 wb_adr_i[13] VGND VGND VPWR VPWR _4338_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_163_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput114 wb_adr_i[23] VGND VGND VPWR VPWR _4390_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput125 wb_adr_i[4] VGND VGND VPWR VPWR _4342_/C sky130_fd_sc_hd__buf_6
XFILLER_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput136 wb_dat_i[13] VGND VGND VPWR VPWR _6379_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput147 wb_dat_i[23] VGND VGND VPWR VPWR _6385_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput158 wb_dat_i[4] VGND VGND VPWR VPWR _6375_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput169 wb_stb_i VGND VGND VPWR VPWR wire4255/A sky130_fd_sc_hd__clkbuf_1
XFILLER_76_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_2_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7092_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_24_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length2360 _6538_/Q VGND VGND VPWR VPWR wire2357/A sky130_fd_sc_hd__clkbuf_1
XFILLER_4_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3982_ hold630/X _3991_/A1 _3982_/S VGND VGND VPWR VPWR _6481_/D sky130_fd_sc_hd__mux2_1
X_6770_ _6770_/CLK _6770_/D fanout4005/X VGND VGND VPWR VPWR _6770_/Q sky130_fd_sc_hd__dfrtp_1
X_5721_ _5721_/A1 _5721_/A2 _5721_/B1 _5721_/B2 _5720_/X VGND VGND VPWR VPWR _5728_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_188_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5652_ _6171_/S VGND VGND VPWR VPWR _5652_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4603_ _4745_/A _4603_/B VGND VGND VPWR VPWR _5059_/A sky130_fd_sc_hd__nor2_1
XFILLER_175_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5583_ _5583_/A0 hold403/X _5583_/S VGND VGND VPWR VPWR _7137_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4534_ _4745_/A _4802_/A VGND VGND VPWR VPWR _4964_/A sky130_fd_sc_hd__nor2_1
XFILLER_175_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold302 _6744_/Q VGND VGND VPWR VPWR hold302/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold313 _6516_/Q VGND VGND VPWR VPWR hold313/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold324 _6866_/Q VGND VGND VPWR VPWR hold324/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 _6824_/Q VGND VGND VPWR VPWR hold335/X sky130_fd_sc_hd__dlygate4sd3_1
X_4465_ _4846_/C _4951_/B VGND VGND VPWR VPWR _4465_/X sky130_fd_sc_hd__and2_1
Xhold346 _6681_/Q VGND VGND VPWR VPWR hold346/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold357 _6710_/Q VGND VGND VPWR VPWR hold357/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold368 _6727_/Q VGND VGND VPWR VPWR hold368/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold379 _6774_/Q VGND VGND VPWR VPWR hold379/X sky130_fd_sc_hd__dlygate4sd3_1
X_3416_ _3416_/A _3416_/B VGND VGND VPWR VPWR _3416_/Y sky130_fd_sc_hd__nand2_1
X_6204_ _7025_/Q _6204_/A2 _6204_/B1 _7110_/Q _6203_/X VGND VGND VPWR VPWR _6204_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7184_ _7185_/CLK _7184_/D wire3984/X VGND VGND VPWR VPWR _7184_/Q sky130_fd_sc_hd__dfrtp_1
X_4396_ _4396_/A _4596_/A _5021_/A VGND VGND VPWR VPWR _4396_/X sky130_fd_sc_hd__or3_2
Xwire2609 _4444_/Y VGND VGND VPWR VPWR _4724_/B sky130_fd_sc_hd__clkbuf_2
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6135_ _6135_/A1 _6158_/A2 _6158_/B1 _6135_/B2 _6134_/X VGND VGND VPWR VPWR _6143_/B
+ sky130_fd_sc_hd__a221o_1
X_3347_ _3347_/A1 _3407_/A2 _5250_/A _6218_/B2 VGND VGND VPWR VPWR _3347_/X sky130_fd_sc_hd__a22o_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1908 wire1909/X VGND VGND VPWR VPWR _5738_/B2 sky130_fd_sc_hd__clkbuf_2
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1919 _6081_/B2 VGND VGND VPWR VPWR _5736_/A1 sky130_fd_sc_hd__clkbuf_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6066_ _7051_/Q _6124_/A2 _6126_/A2 _6066_/B2 VGND VGND VPWR VPWR _6066_/X sky130_fd_sc_hd__a22o_1
X_3278_ _3546_/A _3324_/A VGND VGND VPWR VPWR _3278_/Y sky130_fd_sc_hd__nor2_1
X_5017_ _5017_/A _5017_/B VGND VGND VPWR VPWR _5083_/C sky130_fd_sc_hd__nor2_1
XFILLER_39_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6968_ _6973_/CLK _6968_/D wire4069/X VGND VGND VPWR VPWR _6968_/Q sky130_fd_sc_hd__dfrtp_1
X_5919_ _6276_/B2 _5930_/A2 _5944_/B1 _6287_/B2 VGND VGND VPWR VPWR _5919_/X sky130_fd_sc_hd__a22o_1
X_6899_ _7046_/CLK _6899_/D wire4052/X VGND VGND VPWR VPWR _6899_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_139_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3800 _4842_/A1 VGND VGND VPWR VPWR _4581_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3811 _4472_/X VGND VGND VPWR VPWR _5023_/B sky130_fd_sc_hd__clkbuf_2
Xwire3822 _4390_/X VGND VGND VPWR VPWR wire3822/X sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3833 _6432_/B VGND VGND VPWR VPWR _6428_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3844 _4070_/A2 VGND VGND VPWR VPWR wire3844/X sky130_fd_sc_hd__clkbuf_1
Xwire3855 _4570_/B VGND VGND VPWR VPWR _4450_/A sky130_fd_sc_hd__buf_2
XFILLER_89_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3866 wire3867/X VGND VGND VPWR VPWR wire3866/X sky130_fd_sc_hd__clkbuf_1
XFILLER_150_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3877 input95/X VGND VGND VPWR VPWR wire3877/X sky130_fd_sc_hd__clkbuf_1
XFILLER_67_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3888 input90/X VGND VGND VPWR VPWR wire3888/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3899 wire3900/X VGND VGND VPWR VPWR wire3899/X sky130_fd_sc_hd__clkbuf_1
XFILLER_67_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4250_ _4250_/A0 hold226/X _4251_/S VGND VGND VPWR VPWR _6704_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3201_ _7106_/Q VGND VGND VPWR VPWR _3201_/Y sky130_fd_sc_hd__inv_2
X_4181_ _6639_/Q wire358/X _4188_/S VGND VGND VPWR VPWR _6639_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6822_ _7139_/CLK _6822_/D _6499_/SET_B VGND VGND VPWR VPWR _6822_/Q sky130_fd_sc_hd__dfrtp_1
X_6753_ _6755_/CLK _6753_/D wire3950/X VGND VGND VPWR VPWR _6753_/Q sky130_fd_sc_hd__dfstp_1
X_3965_ _3965_/A1 _3963_/B hold55/X VGND VGND VPWR VPWR hold7/A sky130_fd_sc_hd__o21ai_1
XFILLER_149_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5704_ _6978_/Q _5741_/B1 _5746_/B1 _5981_/B2 VGND VGND VPWR VPWR _5704_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3896_ _5648_/C _3896_/B VGND VGND VPWR VPWR _3896_/X sky130_fd_sc_hd__or2_1
X_6684_ _6702_/CLK _6684_/D wire3958/X VGND VGND VPWR VPWR _6684_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_31_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5635_ _6564_/Q _6000_/A _6033_/A VGND VGND VPWR VPWR _5635_/X sky130_fd_sc_hd__and3_1
XFILLER_136_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5566_ _5566_/A0 hold605/X _5570_/S VGND VGND VPWR VPWR _7122_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold110 _6550_/Q VGND VGND VPWR VPWR hold110/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 _6839_/Q VGND VGND VPWR VPWR hold121/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold132 _7107_/Q VGND VGND VPWR VPWR hold132/X sky130_fd_sc_hd__dlygate4sd3_1
X_4517_ _4942_/A _4520_/B VGND VGND VPWR VPWR _5124_/A sky130_fd_sc_hd__nor2_1
X_5497_ _5584_/A0 hold185/X _5497_/S VGND VGND VPWR VPWR _7061_/D sky130_fd_sc_hd__mux2_1
Xhold143 _4144_/X VGND VGND VPWR VPWR _6608_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 _5545_/X VGND VGND VPWR VPWR _7103_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 _6467_/Q VGND VGND VPWR VPWR hold165/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 _7042_/Q VGND VGND VPWR VPWR hold176/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3129 _5659_/X VGND VGND VPWR VPWR wire3129/X sky130_fd_sc_hd__clkbuf_1
X_4448_ _4516_/A _4448_/B VGND VGND VPWR VPWR _4510_/A sky130_fd_sc_hd__nand2_1
Xhold187 _6579_/Q VGND VGND VPWR VPWR hold187/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire2406 _6511_/Q VGND VGND VPWR VPWR _6223_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold198 _5256_/X VGND VGND VPWR VPWR _6847_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_120_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2417 _6505_/Q VGND VGND VPWR VPWR wire2417/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4379_ _4379_/A _4402_/A _4379_/C _4407_/A VGND VGND VPWR VPWR _4657_/B sky130_fd_sc_hd__nor4_2
X_7167_ _3937_/A1 _7167_/D wire4001/X VGND VGND VPWR VPWR _7167_/Q sky130_fd_sc_hd__dfrtp_1
Xwire2428 wire2429/X VGND VGND VPWR VPWR _6080_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2439 _6490_/Q VGND VGND VPWR VPWR _3769_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire1705 _7038_/Q VGND VGND VPWR VPWR _5777_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1716 _7036_/Q VGND VGND VPWR VPWR wire1716/X sky130_fd_sc_hd__clkbuf_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1727 wire1728/X VGND VGND VPWR VPWR _6186_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_86_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6118_ _6118_/A1 _6118_/A2 _6115_/X _6117_/X VGND VGND VPWR VPWR _6119_/D sky130_fd_sc_hd__a211o_1
X_7098_ _7101_/CLK _7098_/D wire3996/A VGND VGND VPWR VPWR _7098_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1738 wire1739/X VGND VGND VPWR VPWR _3685_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_100_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1749 _7023_/Q VGND VGND VPWR VPWR wire1749/X sky130_fd_sc_hd__clkbuf_1
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6049_ _6049_/A _6049_/B VGND VGND VPWR VPWR _6049_/X sky130_fd_sc_hd__and2_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_82_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6803_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_10_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length622 _5484_/Y VGND VGND VPWR VPWR _5491_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length655 wire654/A VGND VGND VPWR VPWR wire651/A sky130_fd_sc_hd__clkbuf_1
XFILLER_185_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length666 _5417_/S VGND VGND VPWR VPWR wire661/A sky130_fd_sc_hd__clkbuf_1
XFILLER_5_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout3524 hold48/X VGND VGND VPWR VPWR hold49/A sky130_fd_sc_hd__clkbuf_1
XFILLER_118_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3630 _5503_/A0 VGND VGND VPWR VPWR _4325_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3641 wire3642/X VGND VGND VPWR VPWR wire3641/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3652 wire3652/A VGND VGND VPWR VPWR _5563_/A0 sky130_fd_sc_hd__clkbuf_2
Xwire3663 wire3664/X VGND VGND VPWR VPWR wire3663/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_20_csclk _6579_/CLK VGND VGND VPWR VPWR _7127_/CLK sky130_fd_sc_hd__clkbuf_16
Xwire3674 _3952_/X VGND VGND VPWR VPWR wire3674/X sky130_fd_sc_hd__clkbuf_1
Xwire3685 _5743_/B VGND VGND VPWR VPWR wire3685/X sky130_fd_sc_hd__clkbuf_1
Xwire2940 _5796_/B1 VGND VGND VPWR VPWR _5768_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire3696 _3907_/A VGND VGND VPWR VPWR _6318_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_49_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2951 _5759_/B1 VGND VGND VPWR VPWR _5788_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2962 _5839_/B1 VGND VGND VPWR VPWR _5798_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire2973 wire2974/X VGND VGND VPWR VPWR _5851_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire2984 _5845_/A2 VGND VGND VPWR VPWR _5806_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_134_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2995 _5682_/X VGND VGND VPWR VPWR _5843_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_134_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_35_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7134_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_17_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3750_ _6716_/Q _4264_/A wire800/X _6228_/B2 VGND VGND VPWR VPWR _3750_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3681_ _5714_/A1 _3681_/A2 _3681_/B1 _6522_/Q _3680_/X VGND VGND VPWR VPWR _3688_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5420_ _5552_/A0 hold698/X _5420_/S VGND VGND VPWR VPWR _6993_/D sky130_fd_sc_hd__mux2_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput204 wire1364/X VGND VGND VPWR VPWR mgmt_gpio_oeb[36] sky130_fd_sc_hd__buf_12
X_5351_ _5351_/A0 hold222/X _5351_/S VGND VGND VPWR VPWR _6931_/D sky130_fd_sc_hd__mux2_1
Xoutput215 wire2347/X VGND VGND VPWR VPWR mgmt_gpio_out[11] sky130_fd_sc_hd__buf_12
XFILLER_126_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput226 _6551_/Q VGND VGND VPWR VPWR mgmt_gpio_out[21] sky130_fd_sc_hd__buf_12
XFILLER_154_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput237 hold40/A VGND VGND VPWR VPWR mgmt_gpio_out[31] sky130_fd_sc_hd__buf_12
Xoutput248 _6561_/Q VGND VGND VPWR VPWR mgmt_gpio_out[7] sky130_fd_sc_hd__buf_12
X_4302_ _5387_/A0 hold293/X hold31/X VGND VGND VPWR VPWR _6747_/D sky130_fd_sc_hd__mux2_1
X_5282_ _5576_/A0 hold131/X _5282_/S VGND VGND VPWR VPWR _6870_/D sky130_fd_sc_hd__mux2_1
Xoutput259 _3950_/Y VGND VGND VPWR VPWR pad_flash_io1_ieb sky130_fd_sc_hd__buf_12
X_7021_ _7056_/CLK _7021_/D fanout3976/X VGND VGND VPWR VPWR _7021_/Q sky130_fd_sc_hd__dfrtp_1
X_4233_ _6346_/A _3963_/B _6697_/Q _4230_/X _6391_/A3 VGND VGND VPWR VPWR _6680_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_114_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4164_ hold288/X _4215_/A1 _4164_/S VGND VGND VPWR VPWR _6625_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4095_ hold333/X _4094_/X _4097_/S VGND VGND VPWR VPWR _6569_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6805_ _7036_/CLK _6805_/D wire3974/A VGND VGND VPWR VPWR _6805_/Q sky130_fd_sc_hd__dfstp_1
X_4997_ _4997_/A _5036_/B VGND VGND VPWR VPWR _5009_/A sky130_fd_sc_hd__nor2_1
XFILLER_23_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6736_ _6979_/CLK _6736_/D fanout4027/X VGND VGND VPWR VPWR _6736_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_177_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3948_ _3948_/A VGND VGND VPWR VPWR _3948_/Y sky130_fd_sc_hd__inv_2
Xmax_length3627 _5212_/C VGND VGND VPWR VPWR _3984_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_176_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length3638 _5536_/A1 VGND VGND VPWR VPWR _5422_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_139_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6667_ _6683_/CLK _6667_/D wire3965/A VGND VGND VPWR VPWR _6667_/Q sky130_fd_sc_hd__dfstp_1
X_3879_ _4339_/A _4339_/B _3879_/C VGND VGND VPWR VPWR _3887_/A sky130_fd_sc_hd__or3_1
XFILLER_176_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5618_ _7150_/Q _5618_/B VGND VGND VPWR VPWR _5622_/B sky130_fd_sc_hd__or2_1
X_6598_ _6799_/CLK _6598_/D wire3948/A VGND VGND VPWR VPWR _6598_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5549_ _5576_/A0 hold132/X _5550_/S VGND VGND VPWR VPWR _7107_/D sky130_fd_sc_hd__mux2_1
XFILLER_3_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2203 _6734_/Q VGND VGND VPWR VPWR _6303_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2214 wire2215/X VGND VGND VPWR VPWR _6231_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire2225 _6714_/Q VGND VGND VPWR VPWR wire2225/X sky130_fd_sc_hd__clkbuf_1
Xwire2236 _6290_/B2 VGND VGND VPWR VPWR _5918_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2247 _6701_/Q VGND VGND VPWR VPWR _6230_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_559 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1513 _3378_/Y VGND VGND VPWR VPWR _3472_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2258 _6681_/Q VGND VGND VPWR VPWR wire2258/X sky130_fd_sc_hd__clkbuf_1
XFILLER_171_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1524 _3324_/A VGND VGND VPWR VPWR _3526_/A sky130_fd_sc_hd__clkbuf_2
Xwire2269 _6674_/Q VGND VGND VPWR VPWR _6340_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire1535 wire1536/X VGND VGND VPWR VPWR wire1535/X sky130_fd_sc_hd__clkbuf_1
XFILLER_171_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1557 _3351_/A1 VGND VGND VPWR VPWR _6209_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire1568 _7108_/Q VGND VGND VPWR VPWR _6152_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_58_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1579 wire1580/X VGND VGND VPWR VPWR _6157_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_73_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire810 wire811/X VGND VGND VPWR VPWR wire810/X sky130_fd_sc_hd__clkbuf_1
Xwire832 wire833/X VGND VGND VPWR VPWR wire832/X sky130_fd_sc_hd__clkbuf_1
Xwire843 _3425_/X VGND VGND VPWR VPWR wire843/X sky130_fd_sc_hd__clkbuf_1
Xwire854 _3365_/X VGND VGND VPWR VPWR wire854/X sky130_fd_sc_hd__clkbuf_1
XFILLER_127_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire865 wire866/X VGND VGND VPWR VPWR _5544_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xwire876 wire877/X VGND VGND VPWR VPWR _5259_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_182_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout4011 wire4018/X VGND VGND VPWR VPWR wire4016/A sky130_fd_sc_hd__buf_6
Xwire887 _3337_/Y VGND VGND VPWR VPWR wire887/X sky130_fd_sc_hd__clkbuf_2
Xwire898 _3335_/Y VGND VGND VPWR VPWR wire898/X sky130_fd_sc_hd__clkbuf_1
XFILLER_115_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout4077 wire4081/X VGND VGND VPWR VPWR fanout4077/X sky130_fd_sc_hd__clkbuf_4
Xwire4150 _3859_/A1 VGND VGND VPWR VPWR _3832_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A VGND VGND VPWR VPWR _7196_/CLK sky130_fd_sc_hd__clkbuf_8
Xwire4161 wire4162/X VGND VGND VPWR VPWR _3926_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_97_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire4172 wire4173/X VGND VGND VPWR VPWR _3626_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire4183 wire4184/X VGND VGND VPWR VPWR wire4183/X sky130_fd_sc_hd__clkbuf_1
Xwire4194 wire4195/X VGND VGND VPWR VPWR wire4194/X sky130_fd_sc_hd__clkbuf_1
XFILLER_97_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout3398 hold45/X VGND VGND VPWR VPWR _4118_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_150_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3482 wire3483/X VGND VGND VPWR VPWR wire3482/X sky130_fd_sc_hd__clkbuf_1
Xwire3493 _4286_/A0 VGND VGND VPWR VPWR _4334_/A0 sky130_fd_sc_hd__clkbuf_1
Xwire2770 _5995_/B1 VGND VGND VPWR VPWR _6301_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2781 _6104_/A2 VGND VGND VPWR VPWR _6163_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_37_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2792 _6300_/B1 VGND VGND VPWR VPWR _6325_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4920_ _4655_/B _4635_/B _4920_/B1 _4581_/B _4920_/C1 VGND VGND VPWR VPWR _4920_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_45_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4851_ _4639_/B _4692_/B _4510_/C VGND VGND VPWR VPWR _4862_/A sky130_fd_sc_hd__o21ai_1
XFILLER_60_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3802_ _6473_/Q _6472_/Q _6471_/Q VGND VGND VPWR VPWR _3834_/B sky130_fd_sc_hd__and3_2
X_4782_ _4606_/B _4606_/C _4793_/B VGND VGND VPWR VPWR _4802_/D sky130_fd_sc_hd__a21bo_1
X_6521_ _6761_/CLK _6521_/D wire3970/X VGND VGND VPWR VPWR _6521_/Q sky130_fd_sc_hd__dfrtp_1
X_3733_ _6010_/B2 _3733_/A2 _3733_/B1 _5679_/A1 VGND VGND VPWR VPWR _3733_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6452_ _3927_/A1 _6452_/D _6407_/X VGND VGND VPWR VPWR hold1/A sky130_fd_sc_hd__dfrtp_1
X_3664_ _3664_/A1 wire957/X _3664_/B1 _3664_/B2 VGND VGND VPWR VPWR _3669_/B sky130_fd_sc_hd__a22o_1
XFILLER_146_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5403_ _5403_/A _5403_/B VGND VGND VPWR VPWR _5404_/S sky130_fd_sc_hd__nand2_1
X_6383_ _6382_/X _7203_/Q _6386_/S VGND VGND VPWR VPWR _7203_/D sky130_fd_sc_hd__mux2_1
X_3595_ _3595_/A1 _3595_/A2 _5421_/A _6997_/Q wire783/X VGND VGND VPWR VPWR _3595_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_133_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5334_ _5442_/A0 hold177/X _5334_/S VGND VGND VPWR VPWR _6916_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5265_ _5577_/A0 hold389/X _5267_/S VGND VGND VPWR VPWR _6855_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7004_ _7036_/CLK _7004_/D wire3974/A VGND VGND VPWR VPWR _7004_/Q sky130_fd_sc_hd__dfrtp_1
X_4216_ _4216_/A _4234_/B VGND VGND VPWR VPWR _4221_/S sky130_fd_sc_hd__nand2_2
XFILLER_102_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5196_ _5196_/A0 hold458/X _5199_/S VGND VGND VPWR VPWR _6800_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4147_ _4147_/A _4240_/B VGND VGND VPWR VPWR _4152_/S sky130_fd_sc_hd__nand2_2
XFILLER_18_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4078_ hold694/X _4077_/X _4078_/S VGND VGND VPWR VPWR _6557_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length4125 input66/X VGND VGND VPWR VPWR wire4123/A sky130_fd_sc_hd__clkbuf_1
Xmax_length3402 _5482_/A0 VGND VGND VPWR VPWR _5374_/A0 sky130_fd_sc_hd__clkbuf_2
X_6719_ _7036_/CLK _6719_/D wire3974/X VGND VGND VPWR VPWR _6719_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_137_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3457 _4179_/A0 VGND VGND VPWR VPWR _5534_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_109_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3479 _5291_/A0 VGND VGND VPWR VPWR _5480_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_166_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2000 wire2001/X VGND VGND VPWR VPWR _3529_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_105_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2011 _6890_/Q VGND VGND VPWR VPWR _6035_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_132_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2022 _6882_/Q VGND VGND VPWR VPWR _6032_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2033 wire2034/X VGND VGND VPWR VPWR wire2033/X sky130_fd_sc_hd__clkbuf_1
Xwire2044 _6871_/Q VGND VGND VPWR VPWR _6166_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire1310 wire1311/X VGND VGND VPWR VPWR _6180_/B sky130_fd_sc_hd__clkbuf_1
Xwire2055 wire2056/X VGND VGND VPWR VPWR _6089_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1321 _5922_/X VGND VGND VPWR VPWR _5923_/D sky130_fd_sc_hd__clkbuf_1
Xwire2066 _6112_/B2 VGND VGND VPWR VPWR _3572_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_93_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1332 _5780_/X VGND VGND VPWR VPWR wire1332/X sky130_fd_sc_hd__clkbuf_1
Xwire2077 _6141_/A1 VGND VGND VPWR VPWR _5786_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire2088 _6852_/Q VGND VGND VPWR VPWR _6081_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_115_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1354 wire1355/X VGND VGND VPWR VPWR wire1354/X sky130_fd_sc_hd__clkbuf_2
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2099 _6843_/Q VGND VGND VPWR VPWR _6070_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_101_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1365 _3921_/X VGND VGND VPWR VPWR wire1365/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1376 _3465_/B VGND VGND VPWR VPWR _3511_/B sky130_fd_sc_hd__clkbuf_2
Xwire1387 _3297_/X VGND VGND VPWR VPWR _3507_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire640 _5465_/S VGND VGND VPWR VPWR wire640/X sky130_fd_sc_hd__clkbuf_1
Xwire651 wire651/A VGND VGND VPWR VPWR wire651/X sky130_fd_sc_hd__clkbuf_1
Xwire662 wire663/X VGND VGND VPWR VPWR _5414_/S sky130_fd_sc_hd__clkbuf_1
XFILLER_155_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire684 _5382_/S VGND VGND VPWR VPWR wire684/X sky130_fd_sc_hd__clkbuf_1
Xhold709 _7018_/Q VGND VGND VPWR VPWR hold709/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_109_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3380_ _7187_/Q _6817_/Q _3380_/S VGND VGND VPWR VPWR _3380_/X sky130_fd_sc_hd__mux2_2
XFILLER_97_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5050_ _5050_/A _5050_/B _5050_/C VGND VGND VPWR VPWR _5050_/X sky130_fd_sc_hd__and3_1
XFILLER_69_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4001_ _4001_/A _5535_/B VGND VGND VPWR VPWR _4009_/S sky130_fd_sc_hd__nand2_1
Xwire3290 wire3291/X VGND VGND VPWR VPWR _3866_/S sky130_fd_sc_hd__buf_6
XFILLER_77_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5952_ _5952_/A1 _5952_/A2 _5952_/B1 _6328_/A1 _5951_/X VGND VGND VPWR VPWR _5957_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4903_ _5013_/A _5016_/A _4781_/Y _4477_/X VGND VGND VPWR VPWR _4903_/X sky130_fd_sc_hd__o22a_1
X_5883_ _7208_/Q _5883_/A2 _5883_/B1 _6262_/B2 VGND VGND VPWR VPWR _5883_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4834_ _4947_/A _4933_/A _5035_/B _4652_/A _4784_/A VGND VGND VPWR VPWR _4835_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_178_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4765_ _4993_/A _4512_/B _4746_/Y _4985_/B _4764_/X VGND VGND VPWR VPWR _4765_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_193_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6504_ _7001_/CLK _6504_/D wire3991/X VGND VGND VPWR VPWR _6504_/Q sky130_fd_sc_hd__dfrtp_1
X_3716_ _7059_/Q _3716_/A2 wire875/X _6065_/A1 wire752/X VGND VGND VPWR VPWR _3721_/B
+ sky130_fd_sc_hd__a221o_1
X_4696_ _5076_/A _4694_/B _4651_/X _4696_/B2 VGND VGND VPWR VPWR _4696_/X sky130_fd_sc_hd__o22a_1
XFILLER_119_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6435_ _6437_/A _6435_/B VGND VGND VPWR VPWR _6435_/X sky130_fd_sc_hd__and2_1
X_3647_ _3647_/A1 _3647_/A2 _3607_/Y _3647_/B2 VGND VGND VPWR VPWR _3647_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6366_ _4228_/C _6366_/A2 _6366_/B1 _4228_/A VGND VGND VPWR VPWR _6366_/X sky130_fd_sc_hd__a22o_1
X_3578_ _3578_/A1 wire966/X _4276_/A _6729_/Q VGND VGND VPWR VPWR _3578_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5317_ _5353_/A0 hold578/X _5317_/S VGND VGND VPWR VPWR _6901_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6297_ _6614_/Q _6335_/B1 _6327_/B1 _6297_/B2 VGND VGND VPWR VPWR _6297_/X sky130_fd_sc_hd__a22o_1
XFILLER_114_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold14 hold14/A VGND VGND VPWR VPWR hold14/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5248_ _5248_/A0 hold105/X _5248_/S VGND VGND VPWR VPWR _6840_/D sky130_fd_sc_hd__mux2_1
Xhold25 hold25/A VGND VGND VPWR VPWR hold25/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold36 hold36/A VGND VGND VPWR VPWR hold36/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold47 hold47/A VGND VGND VPWR VPWR hold47/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold58 hold58/A VGND VGND VPWR VPWR hold58/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 hold69/A VGND VGND VPWR VPWR hold69/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5179_ _4659_/A _4679_/B _4679_/X _4510_/A _4510_/B VGND VGND VPWR VPWR _5180_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_29_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length2531 _6185_/B1 VGND VGND VPWR VPWR wire2526/A sky130_fd_sc_hd__clkbuf_1
XFILLER_4_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length1863 _6974_/Q VGND VGND VPWR VPWR wire1862/A sky130_fd_sc_hd__clkbuf_1
XFILLER_193_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1001 wire1011/X VGND VGND VPWR VPWR _5860_/S sky130_fd_sc_hd__buf_6
XFILLER_79_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1151 _3328_/Y VGND VGND VPWR VPWR _5484_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1162 _3326_/Y VGND VGND VPWR VPWR _5457_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_47_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1173 _3667_/A2 VGND VGND VPWR VPWR _3738_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1184 _3581_/A2 VGND VGND VPWR VPWR _3516_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1195 _3736_/A2 VGND VGND VPWR VPWR _5511_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_733 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4550_ _4565_/A _4971_/B VGND VGND VPWR VPWR _4793_/B sky130_fd_sc_hd__xnor2_1
XFILLER_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3501_ _7115_/Q wire961/X _3501_/B1 _3501_/B2 _3500_/X VGND VGND VPWR VPWR _3501_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire470 _5586_/S VGND VGND VPWR VPWR wire470/X sky130_fd_sc_hd__clkbuf_1
Xhold506 _7069_/Q VGND VGND VPWR VPWR hold506/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire481 wire482/X VGND VGND VPWR VPWR _5552_/S sky130_fd_sc_hd__clkbuf_2
Xwire492 _5317_/S VGND VGND VPWR VPWR _5321_/S sky130_fd_sc_hd__clkbuf_1
XFILLER_156_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4481_ _5018_/A _4638_/B VGND VGND VPWR VPWR _4482_/B sky130_fd_sc_hd__or2_1
Xhold517 _6815_/Q VGND VGND VPWR VPWR hold517/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold528 _6911_/Q VGND VGND VPWR VPWR hold528/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6220_ _7182_/Q _6219_/X _6319_/S VGND VGND VPWR VPWR _7182_/D sky130_fd_sc_hd__mux2_1
Xhold539 _6921_/Q VGND VGND VPWR VPWR hold539/X sky130_fd_sc_hd__dlygate4sd3_1
X_3432_ _6154_/B2 _5493_/A _3432_/B1 _3432_/B2 VGND VGND VPWR VPWR _3432_/X sky130_fd_sc_hd__a22o_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3363_ _3363_/A1 _3363_/A2 wire928/X _6905_/Q _3362_/X VGND VGND VPWR VPWR _3363_/X
+ sky130_fd_sc_hd__a221o_1
X_6151_ _6151_/A1 _6151_/A2 _6151_/B1 _6151_/B2 _6148_/X VGND VGND VPWR VPWR _6156_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _5102_/A _5102_/B VGND VGND VPWR VPWR _5103_/B sky130_fd_sc_hd__nor2_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3294_ _3331_/A _3546_/B VGND VGND VPWR VPWR _3294_/Y sky130_fd_sc_hd__nor2_1
XFILLER_58_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6082_ _6082_/A1 _6082_/A2 _6082_/B1 _6884_/Q VGND VGND VPWR VPWR _6082_/X sky130_fd_sc_hd__a22o_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _5033_/A _5033_/B _5033_/C VGND VGND VPWR VPWR _5033_/X sky130_fd_sc_hd__or3_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6984_ _7016_/CLK _6984_/D wire4001/A VGND VGND VPWR VPWR _6984_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5935_ _5935_/A _5935_/B _5935_/C _5935_/D VGND VGND VPWR VPWR _5935_/X sky130_fd_sc_hd__or4_1
XFILLER_80_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5866_ _6660_/Q _5934_/A2 _5865_/X VGND VGND VPWR VPWR _5869_/C sky130_fd_sc_hd__a21o_1
X_4817_ _4983_/C _4817_/B _4817_/C _4816_/X VGND VGND VPWR VPWR _4818_/A sky130_fd_sc_hd__or4b_1
XFILLER_178_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5797_ _6163_/B2 _5797_/A2 _5797_/B1 _6154_/B2 VGND VGND VPWR VPWR _5797_/X sky130_fd_sc_hd__a22o_1
XFILLER_193_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4748_ _4748_/A _4872_/A VGND VGND VPWR VPWR _4818_/B sky130_fd_sc_hd__nor2_1
XFILLER_107_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4679_ _4940_/B _4679_/B VGND VGND VPWR VPWR _4679_/X sky130_fd_sc_hd__or2_1
X_6418_ _6441_/A _6441_/B VGND VGND VPWR VPWR _6418_/X sky130_fd_sc_hd__and2_1
Xmax_length1148 _3654_/B1 VGND VGND VPWR VPWR wire1146/A sky130_fd_sc_hd__clkbuf_1
XFILLER_115_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6349_ _7189_/Q wire359/X _6353_/S VGND VGND VPWR VPWR _7189_/D sky130_fd_sc_hd__mux2_1
XFILLER_163_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput104 wb_adr_i[14] VGND VGND VPWR VPWR _4338_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput115 wb_adr_i[24] VGND VGND VPWR VPWR _3880_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput126 wb_adr_i[5] VGND VGND VPWR VPWR _4605_/A sky130_fd_sc_hd__buf_6
Xinput137 wb_dat_i[14] VGND VGND VPWR VPWR _6381_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput148 wb_dat_i[24] VGND VGND VPWR VPWR _6364_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput159 wb_dat_i[5] VGND VGND VPWR VPWR _6378_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3040 _5955_/A2 VGND VGND VPWR VPWR _5892_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_184_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3981_ hold1/X _7204_/Q _3981_/S VGND VGND VPWR VPWR hold2/A sky130_fd_sc_hd__mux2_1
XFILLER_22_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5720_ _6062_/A1 _5745_/A2 _5745_/B1 _6066_/B2 VGND VGND VPWR VPWR _5720_/X sky130_fd_sc_hd__a22o_1
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5651_ _5651_/A _5651_/B VGND VGND VPWR VPWR _5651_/Y sky130_fd_sc_hd__nor2_1
XFILLER_175_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4602_ _4846_/A _4570_/B _4398_/C _4778_/B _4601_/X VGND VGND VPWR VPWR _4647_/A
+ sky130_fd_sc_hd__a41o_1
XFILLER_175_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5582_ _5582_/A0 hold467/X _5582_/S VGND VGND VPWR VPWR _7136_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4533_ _4533_/A _4778_/A VGND VGND VPWR VPWR _4535_/B sky130_fd_sc_hd__nand2_1
XFILLER_7_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold303 _4298_/X VGND VGND VPWR VPWR _6744_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 _4023_/X VGND VGND VPWR VPWR _6516_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold325 _6938_/Q VGND VGND VPWR VPWR hold325/X sky130_fd_sc_hd__dlygate4sd3_1
X_4464_ _4846_/D VGND VGND VPWR VPWR _4464_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold336 _6685_/Q VGND VGND VPWR VPWR hold336/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 _6682_/Q VGND VGND VPWR VPWR hold347/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 _6656_/Q VGND VGND VPWR VPWR hold358/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 _6622_/Q VGND VGND VPWR VPWR hold369/X sky130_fd_sc_hd__dlygate4sd3_1
X_6203_ _6993_/Q _6203_/A2 _6203_/B1 _6203_/B2 VGND VGND VPWR VPWR _6203_/X sky130_fd_sc_hd__a22o_1
X_3415_ _3518_/B _3415_/B VGND VGND VPWR VPWR _3415_/Y sky130_fd_sc_hd__nor2_1
X_7183_ _7187_/CLK _7183_/D wire3984/X VGND VGND VPWR VPWR _7183_/Q sky130_fd_sc_hd__dfrtp_1
X_4395_ _4461_/B VGND VGND VPWR VPWR _4395_/Y sky130_fd_sc_hd__inv_2
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6134_ _7139_/Q _6157_/A2 _6157_/B1 _6134_/B2 _6123_/X VGND VGND VPWR VPWR _6134_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3346_ _6937_/Q _3346_/A2 _3564_/A2 _6921_/Q VGND VGND VPWR VPWR _3346_/X sky130_fd_sc_hd__a22o_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1909 _6082_/A1 VGND VGND VPWR VPWR wire1909/X sky130_fd_sc_hd__clkbuf_1
XFILLER_85_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065_ _6065_/A1 _6065_/A2 _6065_/B1 hold72/A _6048_/X VGND VGND VPWR VPWR _6068_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3277_ _3293_/A _3416_/B VGND VGND VPWR VPWR _3324_/A sky130_fd_sc_hd__nand2_1
X_5016_ _5016_/A _5016_/B VGND VGND VPWR VPWR _5017_/B sky130_fd_sc_hd__and2_1
XFILLER_100_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6967_ _7116_/CLK _6967_/D wire4071/A VGND VGND VPWR VPWR _6967_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_41_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5918_ _5918_/A1 _5918_/A2 _5931_/B1 _6276_/A1 _5917_/X VGND VGND VPWR VPWR _5923_/B
+ sky130_fd_sc_hd__a221o_1
X_6898_ _6956_/CLK _6898_/D wire4040/X VGND VGND VPWR VPWR _6898_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_179_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5849_ _5849_/A1 _5849_/A2 _5849_/B1 _6202_/A1 _5848_/X VGND VGND VPWR VPWR _5857_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length859 wire860/X VGND VGND VPWR VPWR wire858/A sky130_fd_sc_hd__clkbuf_1
XFILLER_108_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3801 _4646_/A VGND VGND VPWR VPWR _4842_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3812 _4942_/B VGND VGND VPWR VPWR _4940_/B sky130_fd_sc_hd__clkbuf_2
Xwire3823 _4380_/X VGND VGND VPWR VPWR _5021_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_122_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3856 _4570_/B VGND VGND VPWR VPWR _4538_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3867 input97/X VGND VGND VPWR VPWR wire3867/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3878 wire3879/X VGND VGND VPWR VPWR _3938_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_131_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3889 wire3890/X VGND VGND VPWR VPWR _3919_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_103_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3200_ _7114_/Q VGND VGND VPWR VPWR _3200_/Y sky130_fd_sc_hd__inv_2
X_4180_ _6693_/Q _6348_/B VGND VGND VPWR VPWR _4188_/S sky130_fd_sc_hd__and2_2
XFILLER_95_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6821_ _7139_/CLK _6821_/D _6499_/SET_B VGND VGND VPWR VPWR _6821_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_63_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6752_ _6825_/CLK _6752_/D wire3954/X VGND VGND VPWR VPWR _6752_/Q sky130_fd_sc_hd__dfrtp_1
X_3964_ _3965_/A1 _3963_/B hold55/X VGND VGND VPWR VPWR hold56/A sky130_fd_sc_hd__o21a_1
XFILLER_189_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5703_ _5705_/A _5703_/B _5703_/C VGND VGND VPWR VPWR _5703_/X sky130_fd_sc_hd__and3_1
XFILLER_176_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6683_ _6683_/CLK _6683_/D fanout3964/A VGND VGND VPWR VPWR _6683_/Q sky130_fd_sc_hd__dfstp_1
Xmax_length3809 _4971_/B VGND VGND VPWR VPWR _4819_/D sky130_fd_sc_hd__clkbuf_2
X_3895_ _7144_/Q _7146_/Q _7147_/Q _7145_/Q VGND VGND VPWR VPWR _3896_/B sky130_fd_sc_hd__or4b_1
XFILLER_176_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5634_ _5637_/B _6039_/A VGND VGND VPWR VPWR _5634_/Y sky130_fd_sc_hd__nand2_1
XFILLER_148_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5565_ _5565_/A0 _7121_/Q _5565_/S VGND VGND VPWR VPWR hold78/A sky130_fd_sc_hd__mux2_1
XFILLER_191_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold100 _6872_/Q VGND VGND VPWR VPWR hold100/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 _4063_/X VGND VGND VPWR VPWR _6550_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4516_ _4516_/A _4516_/B VGND VGND VPWR VPWR _4850_/A sky130_fd_sc_hd__nand2_1
XFILLER_172_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold122 _6974_/Q VGND VGND VPWR VPWR hold122/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 _6934_/Q VGND VGND VPWR VPWR hold133/X sky130_fd_sc_hd__dlygate4sd3_1
X_5496_ _5574_/A0 hold255/X _5497_/S VGND VGND VPWR VPWR _7060_/D sky130_fd_sc_hd__mux2_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold144 _6867_/Q VGND VGND VPWR VPWR hold144/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold155 _6851_/Q VGND VGND VPWR VPWR hold155/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3108 _5819_/B1 VGND VGND VPWR VPWR _5781_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_104_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold166 _3253_/X VGND VGND VPWR VPWR hold166/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3119 wire3120/X VGND VGND VPWR VPWR wire3119/X sky130_fd_sc_hd__clkbuf_2
X_4447_ _4516_/A _4460_/A VGND VGND VPWR VPWR _4447_/Y sky130_fd_sc_hd__nand2_1
Xhold177 _6916_/Q VGND VGND VPWR VPWR hold177/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 _6981_/Q VGND VGND VPWR VPWR hold188/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 _7013_/Q VGND VGND VPWR VPWR hold199/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2407 _6510_/Q VGND VGND VPWR VPWR _6330_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2418 _6504_/Q VGND VGND VPWR VPWR _6182_/A1 sky130_fd_sc_hd__clkbuf_2
X_7166_ _3937_/A1 _7166_/D wire4001/A VGND VGND VPWR VPWR _7166_/Q sky130_fd_sc_hd__dfrtp_1
X_4378_ _4546_/A _4378_/B VGND VGND VPWR VPWR _4721_/A sky130_fd_sc_hd__or2_1
Xwire2429 _5732_/B2 VGND VGND VPWR VPWR wire2429/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_1_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6701_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1706 wire1707/X VGND VGND VPWR VPWR _3551_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_85_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6117_ _6117_/A1 _6157_/A2 _6157_/B1 _6117_/B2 _6116_/X VGND VGND VPWR VPWR _6117_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3329_ _3331_/A hold85/A VGND VGND VPWR VPWR _3329_/Y sky130_fd_sc_hd__nor2_1
XFILLER_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1717 _5721_/B2 VGND VGND VPWR VPWR _3700_/A1 sky130_fd_sc_hd__clkbuf_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7097_ _7115_/CLK _7097_/D wire3980/X VGND VGND VPWR VPWR _7097_/Q sky130_fd_sc_hd__dfrtp_1
Xwire1728 _5834_/B2 VGND VGND VPWR VPWR wire1728/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1739 wire1740/X VGND VGND VPWR VPWR wire1739/X sky130_fd_sc_hd__clkbuf_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6048_ _6499_/Q _6140_/A2 _6081_/B1 _6048_/B2 VGND VGND VPWR VPWR _6048_/X sky130_fd_sc_hd__a22o_1
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length656 _5439_/Y VGND VGND VPWR VPWR wire654/A sky130_fd_sc_hd__clkbuf_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout3503 wire3530/X VGND VGND VPWR VPWR wire3511/A sky130_fd_sc_hd__clkbuf_1
XFILLER_123_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout4259 wire4265/X VGND VGND VPWR VPWR wire4264/A sky130_fd_sc_hd__clkbuf_1
XFILLER_78_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_0_0_mgmt_gpio_in[4] clkbuf_2_1_0_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR _3945_/A1
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_123_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire3620 hold37/A VGND VGND VPWR VPWR wire3620/X sky130_fd_sc_hd__clkbuf_1
XFILLER_123_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3631 _4247_/A0 VGND VGND VPWR VPWR _5503_/A0 sky130_fd_sc_hd__clkbuf_2
Xwire3642 wire3642/A VGND VGND VPWR VPWR wire3642/X sky130_fd_sc_hd__clkbuf_1
XFILLER_150_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3664 hold153/X VGND VGND VPWR VPWR wire3664/X sky130_fd_sc_hd__clkbuf_1
Xwire2930 wire2931/X VGND VGND VPWR VPWR _5783_/C1 sky130_fd_sc_hd__clkbuf_2
Xwire3675 _3943_/X VGND VGND VPWR VPWR wire3675/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2941 _5851_/B1 VGND VGND VPWR VPWR _5796_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire3686 _5796_/A2 VGND VGND VPWR VPWR _5743_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3697 _5858_/C1 VGND VGND VPWR VPWR _6219_/S sky130_fd_sc_hd__clkbuf_2
Xwire2952 _5842_/A2 VGND VGND VPWR VPWR _5759_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_103_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2974 _5685_/X VGND VGND VPWR VPWR wire2974/X sky130_fd_sc_hd__clkbuf_1
Xwire2985 wire2986/X VGND VGND VPWR VPWR _5845_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_18_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3680_ _6707_/Q _4252_/A wire802/X _5899_/A1 VGND VGND VPWR VPWR _3680_/X sky130_fd_sc_hd__a22o_1
XFILLER_159_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5350_ _5350_/A0 hold213/X _5354_/S VGND VGND VPWR VPWR _6930_/D sky130_fd_sc_hd__mux2_1
Xoutput205 wire1366/X VGND VGND VPWR VPWR mgmt_gpio_oeb[37] sky130_fd_sc_hd__buf_12
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput216 _6570_/Q VGND VGND VPWR VPWR mgmt_gpio_out[12] sky130_fd_sc_hd__buf_12
Xoutput227 hold87/A VGND VGND VPWR VPWR mgmt_gpio_out[22] sky130_fd_sc_hd__buf_12
XFILLER_5_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput238 wire1480/X VGND VGND VPWR VPWR mgmt_gpio_out[32] sky130_fd_sc_hd__buf_12
XFILLER_141_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4301_ _5476_/A0 hold190/X hold31/X VGND VGND VPWR VPWR _6746_/D sky130_fd_sc_hd__mux2_1
Xoutput249 _3928_/X VGND VGND VPWR VPWR mgmt_gpio_out[8] sky130_fd_sc_hd__buf_12
X_5281_ _5281_/A0 _5281_/A1 _5281_/S VGND VGND VPWR VPWR hold50/A sky130_fd_sc_hd__mux2_1
XFILLER_99_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7020_ _7074_/CLK _7020_/D fanout3976/X VGND VGND VPWR VPWR _7020_/Q sky130_fd_sc_hd__dfrtp_1
X_4232_ _6696_/Q _4232_/B VGND VGND VPWR VPWR _4232_/X sky130_fd_sc_hd__or2_1
XFILLER_114_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4163_ hold290/X _4214_/A1 _4164_/S VGND VGND VPWR VPWR _6624_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4094_ hold228/X _5389_/A0 _4100_/S VGND VGND VPWR VPWR _4094_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6804_ _6824_/CLK _6804_/D wire3974/A VGND VGND VPWR VPWR _6804_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_63_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4996_ _4996_/A _5003_/B VGND VGND VPWR VPWR _5008_/B sky130_fd_sc_hd__nor2_1
X_6735_ _6755_/CLK _6735_/D fanout3952/X VGND VGND VPWR VPWR _6735_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_189_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3947_ _6460_/Q _3947_/B VGND VGND VPWR VPWR _3948_/A sky130_fd_sc_hd__nand2b_2
XFILLER_23_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6666_ _6702_/CLK _6666_/D wire3965/A VGND VGND VPWR VPWR _6666_/Q sky130_fd_sc_hd__dfrtp_2
X_3878_ _4339_/C _4339_/D _4338_/A _4338_/B VGND VGND VPWR VPWR _3879_/C sky130_fd_sc_hd__or4_1
XFILLER_164_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length2927 _5693_/X VGND VGND VPWR VPWR wire2920/A sky130_fd_sc_hd__clkbuf_1
X_5617_ _5650_/B _5705_/B _5706_/B _7149_/Q _5610_/X VGND VGND VPWR VPWR _7149_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_137_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6597_ _7090_/CLK _6597_/D wire3948/X VGND VGND VPWR VPWR _6597_/Q sky130_fd_sc_hd__dfrtp_1
X_5548_ _5575_/A0 _5548_/A1 _5550_/S VGND VGND VPWR VPWR _7106_/D sky130_fd_sc_hd__mux2_1
XFILLER_105_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5479_ _5479_/A0 hold95/X _5479_/S VGND VGND VPWR VPWR _7045_/D sky130_fd_sc_hd__mux2_1
Xwire2204 _6733_/Q VGND VGND VPWR VPWR _6277_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2215 wire2216/X VGND VGND VPWR VPWR wire2215/X sky130_fd_sc_hd__clkbuf_1
Xwire2237 _6708_/Q VGND VGND VPWR VPWR _6290_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
X_7149_ _7180_/CLK _7149_/D wire3996/X VGND VGND VPWR VPWR _7149_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_48_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2248 _6690_/Q VGND VGND VPWR VPWR _6337_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1503 wire1504/X VGND VGND VPWR VPWR _3432_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_113_590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1514 _3342_/B VGND VGND VPWR VPWR _3338_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_101_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2259 wire2259/A VGND VGND VPWR VPWR _3539_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire1525 _3320_/A VGND VGND VPWR VPWR _5212_/B sky130_fd_sc_hd__clkbuf_2
Xwire1536 hold52/A VGND VGND VPWR VPWR wire1536/X sky130_fd_sc_hd__clkbuf_1
Xwire1547 _7129_/Q VGND VGND VPWR VPWR _6075_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1558 _7118_/Q VGND VGND VPWR VPWR _3351_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_86_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1569 wire1570/X VGND VGND VPWR VPWR _6130_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire800 wire801/X VGND VGND VPWR VPWR wire800/X sky130_fd_sc_hd__clkbuf_2
Xwire811 wire812/X VGND VGND VPWR VPWR wire811/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire822 _3481_/X VGND VGND VPWR VPWR wire822/X sky130_fd_sc_hd__clkbuf_1
Xwire833 wire833/A VGND VGND VPWR VPWR wire833/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire844 wire845/X VGND VGND VPWR VPWR wire844/X sky130_fd_sc_hd__clkbuf_1
XFILLER_182_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire855 wire856/X VGND VGND VPWR VPWR wire855/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire866 wire867/X VGND VGND VPWR VPWR wire866/X sky130_fd_sc_hd__clkbuf_1
XFILLER_127_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire877 wire878/X VGND VGND VPWR VPWR wire877/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_129_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length486 wire485/A VGND VGND VPWR VPWR wire483/A sky130_fd_sc_hd__clkbuf_1
XFILLER_142_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout4067 wire4071/X VGND VGND VPWR VPWR wire4069/A sky130_fd_sc_hd__buf_6
Xfanout4078 wire4081/X VGND VGND VPWR VPWR fanout4078/X sky130_fd_sc_hd__buf_8
XFILLER_89_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4140 wire4141/X VGND VGND VPWR VPWR wire4140/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire4162 wire4162/A VGND VGND VPWR VPWR wire4162/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire4173 input54/X VGND VGND VPWR VPWR wire4173/X sky130_fd_sc_hd__clkbuf_1
Xfanout3377 _5240_/A0 VGND VGND VPWR VPWR wire3387/A sky130_fd_sc_hd__clkbuf_1
XFILLER_151_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire4184 wire4185/X VGND VGND VPWR VPWR wire4184/X sky130_fd_sc_hd__clkbuf_1
Xwire4195 input47/X VGND VGND VPWR VPWR wire4195/X sky130_fd_sc_hd__clkbuf_1
Xwire3450 _6397_/A0 VGND VGND VPWR VPWR _4209_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3461 _4329_/A1 VGND VGND VPWR VPWR _5558_/A0 sky130_fd_sc_hd__clkbuf_2
Xwire3472 hold16/X VGND VGND VPWR VPWR _5237_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3483 hold15/X VGND VGND VPWR VPWR wire3483/X sky130_fd_sc_hd__clkbuf_1
Xwire3494 _6396_/A0 VGND VGND VPWR VPWR _4286_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2760 wire2761/X VGND VGND VPWR VPWR _6302_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_37_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2771 _5994_/X VGND VGND VPWR VPWR _5995_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2782 _6214_/B1 VGND VGND VPWR VPWR _6104_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2793 _5990_/B1 VGND VGND VPWR VPWR _6300_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4850_ _4850_/A _4850_/B VGND VGND VPWR VPWR _5124_/B sky130_fd_sc_hd__nand2_1
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3801_ _6471_/Q _3801_/B VGND VGND VPWR VPWR _6471_/D sky130_fd_sc_hd__xor2_1
X_4781_ _4781_/A _4781_/B VGND VGND VPWR VPWR _4781_/Y sky130_fd_sc_hd__nand2_1
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6520_ _6701_/CLK _6520_/D wire3945/X VGND VGND VPWR VPWR _6520_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3732_ _3732_/A1 _4052_/B wire946/X _7135_/Q VGND VGND VPWR VPWR _3732_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6451_ _3927_/A1 _6451_/D _6406_/X VGND VGND VPWR VPWR hold42/A sky130_fd_sc_hd__dfrtp_1
X_3663_ _6987_/Q _3663_/A2 _3733_/A2 _6057_/A1 VGND VGND VPWR VPWR _3669_/A sky130_fd_sc_hd__a22o_1
XFILLER_118_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5402_ hold534/X _5501_/A0 _5402_/S VGND VGND VPWR VPWR _6977_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6382_ _4228_/B _6382_/A2 _6382_/B1 _4228_/Y _6381_/X VGND VGND VPWR VPWR _6382_/X
+ sky130_fd_sc_hd__a221o_1
X_3594_ _3594_/A1 _3329_/Y _3594_/B1 _3594_/B2 _3555_/X VGND VGND VPWR VPWR _3600_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5333_ _5333_/A0 hold171/X _5333_/S VGND VGND VPWR VPWR _6915_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5264_ _5576_/A0 hold135/X _5264_/S VGND VGND VPWR VPWR _6854_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7003_ _7036_/CLK _7003_/D wire3974/A VGND VGND VPWR VPWR _7003_/Q sky130_fd_sc_hd__dfstp_1
X_4215_ hold406/X _4215_/A1 _4215_/S VGND VGND VPWR VPWR _6669_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5195_ _5195_/A0 hold446/X _5199_/S VGND VGND VPWR VPWR _6799_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_81_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7210_/CLK sky130_fd_sc_hd__clkbuf_16
X_4146_ _4263_/A1 hold238/X _4146_/S VGND VGND VPWR VPWR _6610_/D sky130_fd_sc_hd__mux2_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4077_ hold590/X _5416_/A0 _4079_/S VGND VGND VPWR VPWR _4077_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4979_ _4979_/A _5114_/B _4979_/C _4979_/D VGND VGND VPWR VPWR _4979_/X sky130_fd_sc_hd__or4_1
Xmax_length3403 _5365_/A0 VGND VGND VPWR VPWR _5482_/A0 sky130_fd_sc_hd__clkbuf_1
X_6718_ _7036_/CLK _6718_/D wire3974/X VGND VGND VPWR VPWR _6718_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6649_ _7206_/CLK _6649_/D VGND VGND VPWR VPWR _6649_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_34_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7130_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_180_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2001 wire2002/X VGND VGND VPWR VPWR wire2001/X sky130_fd_sc_hd__clkbuf_1
XFILLER_59_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2012 _6889_/Q VGND VGND VPWR VPWR _6213_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2023 _3361_/B2 VGND VGND VPWR VPWR _5844_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_182_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2034 _3570_/B2 VGND VGND VPWR VPWR wire2034/X sky130_fd_sc_hd__clkbuf_1
XFILLER_120_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1300 _3475_/A2 VGND VGND VPWR VPWR _3407_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire2045 wire2046/X VGND VGND VPWR VPWR _5781_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire1311 _6175_/X VGND VGND VPWR VPWR wire1311/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_49_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7125_/CLK sky130_fd_sc_hd__clkbuf_16
Xwire2056 _6868_/Q VGND VGND VPWR VPWR wire2056/X sky130_fd_sc_hd__clkbuf_1
Xwire1322 _5910_/X VGND VGND VPWR VPWR _5913_/C sky130_fd_sc_hd__clkbuf_1
Xwire2067 _6861_/Q VGND VGND VPWR VPWR _6112_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire2078 _6854_/Q VGND VGND VPWR VPWR _6141_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1333 _5735_/X VGND VGND VPWR VPWR _5740_/B sky130_fd_sc_hd__clkbuf_1
Xwire2089 _6851_/Q VGND VGND VPWR VPWR _6065_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1355 _3934_/X VGND VGND VPWR VPWR wire1355/X sky130_fd_sc_hd__clkbuf_1
Xwire1366 wire1367/X VGND VGND VPWR VPWR wire1366/X sky130_fd_sc_hd__clkbuf_2
XFILLER_74_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1377 _3454_/B VGND VGND VPWR VPWR _3465_/B sky130_fd_sc_hd__clkbuf_2
Xwire1388 _3316_/A VGND VGND VPWR VPWR _3546_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_62_606 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire630 wire631/X VGND VGND VPWR VPWR wire630/X sky130_fd_sc_hd__clkbuf_1
Xwire641 _5465_/S VGND VGND VPWR VPWR _5462_/S sky130_fd_sc_hd__clkbuf_2
Xwire652 _5440_/S VGND VGND VPWR VPWR _5442_/S sky130_fd_sc_hd__clkbuf_1
XFILLER_10_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire663 _5415_/S VGND VGND VPWR VPWR wire663/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire674 _5399_/S VGND VGND VPWR VPWR _5397_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire685 _5376_/Y VGND VGND VPWR VPWR _5382_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_155_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire696 _5345_/S VGND VGND VPWR VPWR _5343_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_170_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3280 _4270_/B VGND VGND VPWR VPWR wire3280/X sky130_fd_sc_hd__clkbuf_1
X_4000_ hold563/X _4000_/A1 _4000_/S VGND VGND VPWR VPWR _6497_/D sky130_fd_sc_hd__mux2_1
Xwire3291 wire3292/X VGND VGND VPWR VPWR wire3291/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5951_ _6321_/A1 _5951_/A2 _5951_/B1 _7211_/Q VGND VGND VPWR VPWR _5951_/X sky130_fd_sc_hd__a22o_1
XFILLER_18_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4902_ _5023_/B _4589_/B _4900_/X _4912_/A1 _5072_/A3 VGND VGND VPWR VPWR _4902_/X
+ sky130_fd_sc_hd__o221a_1
X_5882_ _7170_/Q _5881_/X _5948_/S VGND VGND VPWR VPWR _7170_/D sky130_fd_sc_hd__mux2_1
XFILLER_61_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4833_ _4461_/B _4652_/A _4484_/X VGND VGND VPWR VPWR _4833_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_21_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4764_ _4764_/A _4986_/B _4764_/C VGND VGND VPWR VPWR _4764_/X sky130_fd_sc_hd__or3_1
XFILLER_147_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6503_ _7133_/CLK _6503_/D _7047_/RESET_B VGND VGND VPWR VPWR _6503_/Q sky130_fd_sc_hd__dfrtp_1
X_3715_ _6732_/Q _4282_/A _5229_/A _6825_/Q VGND VGND VPWR VPWR _3715_/X sky130_fd_sc_hd__a22o_1
X_4695_ _5076_/A _4581_/X _4694_/B _4660_/X _4694_/X VGND VGND VPWR VPWR _4698_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_119_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6434_ _6438_/A _6435_/B VGND VGND VPWR VPWR _6434_/X sky130_fd_sc_hd__and2_1
XFILLER_146_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3646_ _6476_/Q _3646_/A2 _3769_/B1 _7036_/Q _3645_/X VGND VGND VPWR VPWR _3651_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6365_ _6364_/X _7197_/Q _6386_/S VGND VGND VPWR VPWR _7197_/D sky130_fd_sc_hd__mux2_1
X_3577_ _3577_/A1 wire924/X wire863/X _6111_/B2 _3576_/X VGND VGND VPWR VPWR _3582_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_136_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5316_ _5487_/A0 hold445/X _5318_/S VGND VGND VPWR VPWR _6900_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6296_ _6729_/Q _6296_/A2 _6296_/B1 _6296_/B2 VGND VGND VPWR VPWR _6296_/X sky130_fd_sc_hd__a22o_1
X_5247_ _5247_/A0 hold121/X _5249_/S VGND VGND VPWR VPWR _6839_/D sky130_fd_sc_hd__mux2_1
Xhold15 hold15/A VGND VGND VPWR VPWR hold15/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 hold26/A VGND VGND VPWR VPWR hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A VGND VGND VPWR VPWR hold37/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 hold48/A VGND VGND VPWR VPWR hold48/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold59 hold59/A VGND VGND VPWR VPWR hold59/X sky130_fd_sc_hd__dlygate4sd3_1
X_5178_ _5178_/A _5178_/B _5178_/C _5178_/D VGND VGND VPWR VPWR _5178_/X sky130_fd_sc_hd__or4_1
XFILLER_56_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4129_ _4129_/A _5529_/B VGND VGND VPWR VPWR _4134_/S sky130_fd_sc_hd__and2_2
XFILLER_84_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length3222 _4491_/B VGND VGND VPWR VPWR _4745_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_177_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length3266 _4318_/B VGND VGND VPWR VPWR wire3260/A sky130_fd_sc_hd__clkbuf_1
XFILLER_153_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length1842 _6991_/Q VGND VGND VPWR VPWR _3423_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_4_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1130 wire1130/A VGND VGND VPWR VPWR _3553_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1141 _3368_/A2 VGND VGND VPWR VPWR _5493_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1152 _3635_/B1 VGND VGND VPWR VPWR _3698_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_47_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1174 _3324_/Y VGND VGND VPWR VPWR _3667_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1185 wire1185/A VGND VGND VPWR VPWR _3441_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_90_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire460 _5924_/X VGND VGND VPWR VPWR wire460/X sky130_fd_sc_hd__clkbuf_1
X_3500_ _3500_/A1 _3500_/A2 _5421_/A _6998_/Q VGND VGND VPWR VPWR _3500_/X sky130_fd_sc_hd__a22o_1
Xwire471 _5579_/S VGND VGND VPWR VPWR _5576_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_128_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4480_ _4588_/A _4935_/A _4621_/A _4621_/B VGND VGND VPWR VPWR _4638_/B sky130_fd_sc_hd__or4_1
Xhold507 _7001_/Q VGND VGND VPWR VPWR hold507/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire482 _5544_/Y VGND VGND VPWR VPWR wire482/X sky130_fd_sc_hd__clkbuf_1
Xhold518 _6525_/Q VGND VGND VPWR VPWR hold518/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire493 _5319_/S VGND VGND VPWR VPWR _5318_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_183_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold529 _6505_/Q VGND VGND VPWR VPWR hold529/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3431_ _3431_/A _3431_/B _3431_/C _3431_/D VGND VGND VPWR VPWR _3447_/A sky130_fd_sc_hd__or4_1
X_6150_ _7079_/Q _6150_/A2 _6150_/B1 _6150_/B2 _6149_/X VGND VGND VPWR VPWR _6156_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3362_ _6897_/Q wire959/X wire862/X _6203_/B2 VGND VGND VPWR VPWR _3362_/X sky130_fd_sc_hd__a22o_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _5114_/C _5145_/B _5112_/D _5101_/D VGND VGND VPWR VPWR _5102_/B sky130_fd_sc_hd__or4_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6081_ _6081_/A1 _6141_/A2 _6081_/B1 _6081_/B2 _6080_/X VGND VGND VPWR VPWR _6084_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ _3293_/A _3313_/B VGND VGND VPWR VPWR _3316_/A sky130_fd_sc_hd__nand2_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5032_ _5012_/X _5032_/A2 _5031_/X VGND VGND VPWR VPWR _5033_/C sky130_fd_sc_hd__o21ba_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6983_ _7116_/CLK _6983_/D wire4071/A VGND VGND VPWR VPWR _6983_/Q sky130_fd_sc_hd__dfrtp_1
X_5934_ _6303_/B2 _5934_/A2 _5934_/B1 _5934_/B2 _5933_/X VGND VGND VPWR VPWR _5935_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_40_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5865_ _6235_/A1 _5865_/A2 _5934_/B1 _6516_/Q VGND VGND VPWR VPWR _5865_/X sky130_fd_sc_hd__a22o_1
X_4816_ _4997_/A _4816_/A2 _4590_/A _4587_/B VGND VGND VPWR VPWR _4816_/X sky130_fd_sc_hd__o22a_1
X_5796_ _6975_/Q _5796_/A2 _5796_/B1 VGND VGND VPWR VPWR _5796_/X sky130_fd_sc_hd__o21a_1
XFILLER_193_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4747_ _5003_/A _4752_/B VGND VGND VPWR VPWR _4985_/B sky130_fd_sc_hd__nor2_1
XFILLER_119_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length1105 _3473_/C1 VGND VGND VPWR VPWR wire1103/A sky130_fd_sc_hd__clkbuf_1
XFILLER_134_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4678_ _5018_/C _4680_/B VGND VGND VPWR VPWR _4916_/B sky130_fd_sc_hd__or2_1
XFILLER_135_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length1127 _3334_/Y VGND VGND VPWR VPWR _3709_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6417_ _6430_/A _6433_/B VGND VGND VPWR VPWR _6417_/X sky130_fd_sc_hd__and2_1
XFILLER_107_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3629_ _3629_/A1 wire903/X wire799/X _3629_/B2 wire555/X VGND VGND VPWR VPWR _3632_/B
+ sky130_fd_sc_hd__a221o_1
X_6348_ _6692_/Q _6348_/B VGND VGND VPWR VPWR _6353_/S sky130_fd_sc_hd__and2_2
XFILLER_103_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput105 wb_adr_i[15] VGND VGND VPWR VPWR _4338_/C sky130_fd_sc_hd__clkbuf_1
X_6279_ _5916_/A _6333_/A2 _6306_/B1 _6279_/B2 _6273_/X VGND VGND VPWR VPWR _6280_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_102_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput116 wb_adr_i[25] VGND VGND VPWR VPWR input116/X sky130_fd_sc_hd__clkbuf_1
Xinput127 wb_adr_i[6] VGND VGND VPWR VPWR wire4285/A sky130_fd_sc_hd__clkbuf_1
XFILLER_130_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput138 wb_dat_i[15] VGND VGND VPWR VPWR _6384_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput149 wb_dat_i[25] VGND VGND VPWR VPWR _6366_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_69_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3074 _5784_/A2 VGND VGND VPWR VPWR _5724_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_165_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length2395 hold316/X VGND VGND VPWR VPWR _4024_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_98_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length1672 hold647/X VGND VGND VPWR VPWR _5483_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_140_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3980_ hold631/X _5437_/A0 _3982_/S VGND VGND VPWR VPWR _6480_/D sky130_fd_sc_hd__mux2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5650_ _5650_/A _5650_/B VGND VGND VPWR VPWR _5650_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4601_ _4749_/C _4572_/Y _4600_/X _4952_/A _5112_/A VGND VGND VPWR VPWR _4601_/X
+ sky130_fd_sc_hd__a2111o_1
X_5581_ _5581_/A0 hold315/X _5581_/S VGND VGND VPWR VPWR _7135_/D sky130_fd_sc_hd__mux2_1
XFILLER_191_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4532_ _4570_/D _4532_/B VGND VGND VPWR VPWR _4971_/A sky130_fd_sc_hd__nor2_2
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold304 _6511_/Q VGND VGND VPWR VPWR hold304/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold315 _7135_/Q VGND VGND VPWR VPWR hold315/X sky130_fd_sc_hd__dlygate4sd3_1
X_4463_ _4474_/A _4944_/A _4462_/Y VGND VGND VPWR VPWR _4487_/B sky130_fd_sc_hd__nor3b_2
Xhold326 _7082_/Q VGND VGND VPWR VPWR hold326/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 _7111_/Q VGND VGND VPWR VPWR hold337/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 _6945_/Q VGND VGND VPWR VPWR hold348/X sky130_fd_sc_hd__dlygate4sd3_1
X_6202_ _6202_/A1 _6202_/A2 _6202_/B1 _6202_/B2 VGND VGND VPWR VPWR _6202_/X sky130_fd_sc_hd__a22o_1
X_3414_ _3416_/A _3414_/B VGND VGND VPWR VPWR _3414_/Y sky130_fd_sc_hd__nand2_1
Xhold359 _4200_/X VGND VGND VPWR VPWR _6656_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7182_ _7187_/CLK _7182_/D wire4015/X VGND VGND VPWR VPWR _7182_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4394_ _4489_/A _4932_/A VGND VGND VPWR VPWR _4461_/B sky130_fd_sc_hd__or2_2
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6133_ _6133_/A1 _6186_/B1 _6128_/X _6130_/X _6132_/X VGND VGND VPWR VPWR _6133_/X
+ sky130_fd_sc_hd__a2111o_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3345_ _3345_/A1 _3425_/B1 _5511_/A _3345_/B2 VGND VGND VPWR VPWR _3345_/X sky130_fd_sc_hd__a22o_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6064_ _6064_/A1 _6064_/A2 _6082_/B1 _6064_/B2 _6063_/X VGND VGND VPWR VPWR _6068_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3276_ _3282_/A hold68/X VGND VGND VPWR VPWR _3416_/B sky130_fd_sc_hd__nor2_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _5107_/C _5015_/B _5015_/C VGND VGND VPWR VPWR _5019_/B sky130_fd_sc_hd__or3_1
XFILLER_38_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6966_ _7075_/CLK _6966_/D wire4066/X VGND VGND VPWR VPWR _6966_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_41_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5917_ _6278_/A1 _5944_/A2 _5917_/B1 _5916_/X VGND VGND VPWR VPWR _5917_/X sky130_fd_sc_hd__a22o_1
X_6897_ _6921_/CLK _6897_/D wire4045/X VGND VGND VPWR VPWR _6897_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5848_ _6202_/B2 _5848_/A2 _5848_/B1 _5848_/B2 VGND VGND VPWR VPWR _5848_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length827 _3678_/B1 VGND VGND VPWR VPWR _4210_/A sky130_fd_sc_hd__clkbuf_2
X_5779_ _6950_/Q _5805_/B1 _5779_/B1 _5779_/B2 VGND VGND VPWR VPWR _5779_/X sky130_fd_sc_hd__a22o_1
Xmax_length838 _3451_/Y VGND VGND VPWR VPWR wire833/A sky130_fd_sc_hd__clkbuf_1
XFILLER_147_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3802 _4712_/B VGND VGND VPWR VPWR _4814_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3813 _4603_/B VGND VGND VPWR VPWR _4942_/B sky130_fd_sc_hd__clkbuf_2
Xwire3824 _4981_/A VGND VGND VPWR VPWR _4668_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_122_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3835 _6441_/B VGND VGND VPWR VPWR _6432_/B sky130_fd_sc_hd__clkbuf_2
Xwire3846 _5241_/C VGND VGND VPWR VPWR _6407_/B sky130_fd_sc_hd__clkbuf_2
Xwire3857 input99/X VGND VGND VPWR VPWR _4570_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3868 wire3869/X VGND VGND VPWR VPWR _3712_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire3879 wire3880/X VGND VGND VPWR VPWR wire3879/X sky130_fd_sc_hd__clkbuf_1
XFILLER_191_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length2192 _6740_/Q VGND VGND VPWR VPWR _3461_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_114_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6820_ _7112_/CLK _6820_/D _7112_/SET_B VGND VGND VPWR VPWR _6820_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6751_ _6825_/CLK _6751_/D wire3954/X VGND VGND VPWR VPWR _6751_/Q sky130_fd_sc_hd__dfrtp_1
X_3963_ hold54/X _3963_/B VGND VGND VPWR VPWR hold55/A sky130_fd_sc_hd__nand2b_1
X_5702_ _7152_/Q _5703_/B _5703_/C VGND VGND VPWR VPWR _5702_/X sky130_fd_sc_hd__and3_1
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_1_1_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
X_6682_ _6683_/CLK _6682_/D fanout3964/A VGND VGND VPWR VPWR _6682_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3894_ _6700_/Q _3876_/X _6695_/Q VGND VGND VPWR VPWR _6700_/D sky130_fd_sc_hd__a21o_1
X_5633_ _7156_/Q _7155_/Q VGND VGND VPWR VPWR _6039_/A sky130_fd_sc_hd__and2_2
XFILLER_191_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5564_ _5582_/A0 hold468/X _5565_/S VGND VGND VPWR VPWR _7120_/D sky130_fd_sc_hd__mux2_1
XFILLER_191_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold101 _6944_/Q VGND VGND VPWR VPWR hold101/X sky130_fd_sc_hd__dlygate4sd3_1
X_4515_ _4515_/A _4515_/B _4515_/C _4863_/A VGND VGND VPWR VPWR _4515_/X sky130_fd_sc_hd__and4_1
Xhold112 _7017_/Q VGND VGND VPWR VPWR hold112/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5495_ _5495_/A0 hold440/X _5495_/S VGND VGND VPWR VPWR _7059_/D sky130_fd_sc_hd__mux2_1
Xhold123 _5399_/X VGND VGND VPWR VPWR _6974_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold134 _6969_/Q VGND VGND VPWR VPWR hold134/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 _7105_/Q VGND VGND VPWR VPWR hold145/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 _6891_/Q VGND VGND VPWR VPWR hold156/X sky130_fd_sc_hd__dlygate4sd3_1
X_4446_ _4872_/A VGND VGND VPWR VPWR _4446_/Y sky130_fd_sc_hd__inv_2
Xhold167 _3270_/B VGND VGND VPWR VPWR _3301_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 _7031_/Q VGND VGND VPWR VPWR hold178/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 _7037_/Q VGND VGND VPWR VPWR hold189/X sky130_fd_sc_hd__dlygate4sd3_1
X_7165_ _3937_/A1 _7165_/D _7176_/RESET_B VGND VGND VPWR VPWR _7165_/Q sky130_fd_sc_hd__dfrtp_1
X_4377_ _4546_/A _4378_/B VGND VGND VPWR VPWR _4657_/A sky130_fd_sc_hd__nor2_1
Xwire2408 _6302_/A1 VGND VGND VPWR VPWR _3596_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire2419 _6503_/Q VGND VGND VPWR VPWR _6163_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6116_ _6116_/A1 _6190_/B1 _6158_/B1 _6116_/B2 VGND VGND VPWR VPWR _6116_/X sky130_fd_sc_hd__a22o_1
X_3328_ _3526_/A _3510_/A VGND VGND VPWR VPWR _3328_/Y sky130_fd_sc_hd__nor2_1
Xwire1707 wire1708/X VGND VGND VPWR VPWR wire1707/X sky130_fd_sc_hd__clkbuf_1
X_7096_ _7115_/CLK _7096_/D wire3980/X VGND VGND VPWR VPWR _7096_/Q sky130_fd_sc_hd__dfstp_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1718 hold72/A VGND VGND VPWR VPWR _5721_/B2 sky130_fd_sc_hd__clkbuf_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1729 hold616/X VGND VGND VPWR VPWR _5834_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6047_ _6047_/A1 wire456/X _6046_/X _5652_/Y _7175_/Q VGND VGND VPWR VPWR _7175_/D
+ sky130_fd_sc_hd__a32o_1
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3259_ hold66/X _3807_/B _3820_/A VGND VGND VPWR VPWR hold67/A sky130_fd_sc_hd__mux2_1
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6949_ _6973_/CLK _6949_/D _7087_/RESET_B VGND VGND VPWR VPWR _6949_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_41_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4300 _4398_/C VGND VGND VPWR VPWR _4376_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_118_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout3548 wire3571/X VGND VGND VPWR VPWR wire3555/A sky130_fd_sc_hd__buf_6
XFILLER_150_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3632 _4211_/A1 VGND VGND VPWR VPWR _4247_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_78_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold690 _7117_/Q VGND VGND VPWR VPWR hold690/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_110_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2920 wire2920/A VGND VGND VPWR VPWR _5695_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire3665 wire3666/X VGND VGND VPWR VPWR wire3665/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3676 _3917_/A VGND VGND VPWR VPWR _3791_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_77_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2931 wire2932/X VGND VGND VPWR VPWR wire2931/X sky130_fd_sc_hd__clkbuf_1
Xwire2942 _5829_/B1 VGND VGND VPWR VPWR _5851_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire3687 _5850_/B VGND VGND VPWR VPWR _5796_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_134_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3698 _6169_/C1 VGND VGND VPWR VPWR _6070_/C1 sky130_fd_sc_hd__clkbuf_1
Xwire2964 _5686_/X VGND VGND VPWR VPWR _5839_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2986 _5683_/X VGND VGND VPWR VPWR wire2986/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2997 _5949_/A2 VGND VGND VPWR VPWR _5920_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput206 _3189_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[3] sky130_fd_sc_hd__buf_12
Xoutput217 wire1452/X VGND VGND VPWR VPWR mgmt_gpio_out[13] sky130_fd_sc_hd__buf_12
XFILLER_99_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4300_ _4300_/A _4300_/B VGND VGND VPWR VPWR hold31/A sky130_fd_sc_hd__nand2_2
Xoutput228 hold12/A VGND VGND VPWR VPWR mgmt_gpio_out[23] sky130_fd_sc_hd__buf_12
Xoutput239 wire1472/X VGND VGND VPWR VPWR mgmt_gpio_out[33] sky130_fd_sc_hd__buf_12
X_5280_ _5487_/A0 hold425/X _5282_/S VGND VGND VPWR VPWR _6868_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4231_ _6696_/Q _4232_/B VGND VGND VPWR VPWR _4231_/Y sky130_fd_sc_hd__nor2_1
XFILLER_141_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4162_ hold249/X _4162_/A1 _4162_/S VGND VGND VPWR VPWR _6623_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4093_ hold284/X _4092_/X _4097_/S VGND VGND VPWR VPWR _4093_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6803_ _6803_/CLK _6803_/D _6495_/SET_B VGND VGND VPWR VPWR _6803_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4995_ _4995_/A _5003_/B VGND VGND VPWR VPWR _5007_/B sky130_fd_sc_hd__nor2_1
X_6734_ _6755_/CLK _6734_/D wire3950/X VGND VGND VPWR VPWR _6734_/Q sky130_fd_sc_hd__dfrtp_1
X_3946_ _6459_/Q _3946_/B VGND VGND VPWR VPWR _3946_/Y sky130_fd_sc_hd__nor2_1
XFILLER_149_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length3629 _4325_/A1 VGND VGND VPWR VPWR wire3628/A sky130_fd_sc_hd__clkbuf_2
X_6665_ _6702_/CLK _6665_/D wire3958/X VGND VGND VPWR VPWR _6665_/Q sky130_fd_sc_hd__dfrtp_1
X_3877_ _3877_/A1 _3965_/A1 _4120_/C VGND VGND VPWR VPWR _3962_/B sky130_fd_sc_hd__o21ai_1
XFILLER_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5616_ _6562_/Q _5650_/B VGND VGND VPWR VPWR _5624_/B sky130_fd_sc_hd__nand2_2
XFILLER_136_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6596_ _6799_/CLK _6596_/D wire3948/X VGND VGND VPWR VPWR _6596_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_152_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5547_ _5547_/A0 hold145/X _5547_/S VGND VGND VPWR VPWR _7105_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5478_ _5487_/A0 hold444/X _5479_/S VGND VGND VPWR VPWR _7044_/D sky130_fd_sc_hd__mux2_1
X_4429_ _4933_/A _4944_/B VGND VGND VPWR VPWR _4836_/A sky130_fd_sc_hd__nor2_1
Xwire2205 _6253_/A1 VGND VGND VPWR VPWR _5886_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire2216 _6721_/Q VGND VGND VPWR VPWR wire2216/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2227 _3630_/B2 VGND VGND VPWR VPWR _5916_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_120_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7148_ _7180_/CLK _7148_/D wire3996/X VGND VGND VPWR VPWR _7148_/Q sky130_fd_sc_hd__dfrtp_2
Xwire2238 _6706_/Q VGND VGND VPWR VPWR _3754_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_58_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1504 wire1505/X VGND VGND VPWR VPWR wire1504/X sky130_fd_sc_hd__clkbuf_1
Xwire2249 wire2250/X VGND VGND VPWR VPWR _3621_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_86_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1515 _3342_/B VGND VGND VPWR VPWR _3711_/B sky130_fd_sc_hd__clkbuf_1
Xwire1526 hold117/X VGND VGND VPWR VPWR _3462_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_59_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1537 _7132_/Q VGND VGND VPWR VPWR _6147_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_101_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7079_ _7079_/CLK _7079_/D wire4049/X VGND VGND VPWR VPWR _7079_/Q sky130_fd_sc_hd__dfrtp_1
Xwire1548 wire1549/X VGND VGND VPWR VPWR _6059_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire1559 _7116_/Q VGND VGND VPWR VPWR _6158_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_39_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire801 wire802/X VGND VGND VPWR VPWR wire801/X sky130_fd_sc_hd__clkbuf_2
XFILLER_168_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire812 _3508_/X VGND VGND VPWR VPWR wire812/X sky130_fd_sc_hd__clkbuf_1
Xwire823 wire824/X VGND VGND VPWR VPWR wire823/X sky130_fd_sc_hd__clkbuf_1
Xwire834 wire835/X VGND VGND VPWR VPWR wire834/X sky130_fd_sc_hd__clkbuf_1
XFILLER_127_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire845 wire846/X VGND VGND VPWR VPWR wire845/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire856 _3356_/X VGND VGND VPWR VPWR wire856/X sky130_fd_sc_hd__clkbuf_1
XFILLER_129_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire867 _3342_/Y VGND VGND VPWR VPWR wire867/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout4002 wire4013/X VGND VGND VPWR VPWR wire4004/A sky130_fd_sc_hd__clkbuf_2
Xwire878 wire878/A VGND VGND VPWR VPWR wire878/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire889 _3336_/Y VGND VGND VPWR VPWR wire889/X sky130_fd_sc_hd__clkbuf_2
XFILLER_129_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout4024 wire4029/A VGND VGND VPWR VPWR wire4026/A sky130_fd_sc_hd__buf_6
XFILLER_142_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length487 _5544_/Y VGND VGND VPWR VPWR wire485/A sky130_fd_sc_hd__clkbuf_1
Xfanout4035 wire4091/X VGND VGND VPWR VPWR _6401_/A sky130_fd_sc_hd__buf_6
XFILLER_89_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout4057 fanout4060/X VGND VGND VPWR VPWR fanout4057/X sky130_fd_sc_hd__buf_6
XFILLER_108_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4130 input64/X VGND VGND VPWR VPWR wire4130/X sky130_fd_sc_hd__clkbuf_1
XFILLER_151_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout4079 wire4088/X VGND VGND VPWR VPWR wire4086/A sky130_fd_sc_hd__buf_6
Xwire4141 input62/X VGND VGND VPWR VPWR wire4141/X sky130_fd_sc_hd__clkbuf_1
Xwire4152 wire4153/X VGND VGND VPWR VPWR _3859_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_123_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4174 wire4175/X VGND VGND VPWR VPWR _3694_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire4185 input50/X VGND VGND VPWR VPWR wire4185/X sky130_fd_sc_hd__clkbuf_1
XFILLER_123_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3440 wire3441/X VGND VGND VPWR VPWR _5463_/A0 sky130_fd_sc_hd__clkbuf_1
Xwire3451 _4033_/A1 VGND VGND VPWR VPWR _6397_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_151_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4196 wire4197/X VGND VGND VPWR VPWR _3566_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_104_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3473 _4305_/A0 VGND VGND VPWR VPWR _4263_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire3484 wire3485/X VGND VGND VPWR VPWR wire3484/X sky130_fd_sc_hd__clkbuf_1
Xwire2750 _6340_/A2 VGND VGND VPWR VPWR _6284_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2761 _6000_/X VGND VGND VPWR VPWR wire2761/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2783 _6184_/A2 VGND VGND VPWR VPWR _6214_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_92_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2794 _6022_/B VGND VGND VPWR VPWR _5990_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3800_ _3800_/A _3800_/B VGND VGND VPWR VPWR _6472_/D sky130_fd_sc_hd__nor2_1
X_4780_ _4780_/A _4981_/C VGND VGND VPWR VPWR _5119_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3731_ _5212_/A _3731_/B VGND VGND VPWR VPWR _3731_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_0_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7090_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_174_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6450_ _3927_/A1 _6450_/D _6405_/X VGND VGND VPWR VPWR _6450_/Q sky130_fd_sc_hd__dfrtp_1
X_3662_ _3661_/X _6785_/Q _3917_/A VGND VGND VPWR VPWR _6785_/D sky130_fd_sc_hd__mux2_1
XFILLER_158_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5401_ hold580/X _5464_/A0 _5402_/S VGND VGND VPWR VPWR _6976_/D sky130_fd_sc_hd__mux2_1
X_6381_ _4228_/C _6381_/A2 _6381_/B1 _4228_/A VGND VGND VPWR VPWR _6381_/X sky130_fd_sc_hd__a22o_1
X_3593_ _3593_/A _3593_/B _3593_/C _3593_/D VGND VGND VPWR VPWR _3593_/X sky130_fd_sc_hd__or4_1
X_5332_ _5476_/A0 hold194/X _5333_/S VGND VGND VPWR VPWR _6914_/D sky130_fd_sc_hd__mux2_1
XFILLER_126_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5263_ _5281_/A0 _5263_/A1 _5263_/S VGND VGND VPWR VPWR _6853_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_718 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7002_ _7036_/CLK _7002_/D wire3974/A VGND VGND VPWR VPWR _7002_/Q sky130_fd_sc_hd__dfstp_1
X_4214_ hold404/X _4214_/A1 _4215_/S VGND VGND VPWR VPWR _6668_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5194_ _5211_/A0 hold422/X _5199_/S VGND VGND VPWR VPWR _6798_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4145_ _4256_/A1 hold247/X _4146_/S VGND VGND VPWR VPWR _6609_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4076_ hold691/X _4075_/X _4078_/S VGND VGND VPWR VPWR _6556_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4978_ _4494_/Y _4783_/Y _5095_/C _5145_/A VGND VGND VPWR VPWR _4979_/D sky130_fd_sc_hd__a211o_1
X_6717_ _6770_/CLK _6717_/D _6767_/RESET_B VGND VGND VPWR VPWR _6717_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_177_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3929_ _3929_/A0 input77/X _3957_/B VGND VGND VPWR VPWR _3929_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6648_ _7206_/CLK _6648_/D VGND VGND VPWR VPWR _6648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6579_ _6579_/CLK _6579_/D _6405_/A VGND VGND VPWR VPWR _6579_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2002 _6894_/Q VGND VGND VPWR VPWR wire2002/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2013 wire2014/X VGND VGND VPWR VPWR _6182_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire2024 wire2025/X VGND VGND VPWR VPWR _3361_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire2035 _6100_/B2 VGND VGND VPWR VPWR _3570_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire1301 _3647_/A2 VGND VGND VPWR VPWR _3475_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_59_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2046 wire2047/X VGND VGND VPWR VPWR wire2046/X sky130_fd_sc_hd__clkbuf_1
Xwire1312 wire1313/X VGND VGND VPWR VPWR _6180_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_120_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2057 _6867_/Q VGND VGND VPWR VPWR _5714_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1323 _5906_/X VGND VGND VPWR VPWR _5913_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_86_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2079 wire2080/X VGND VGND VPWR VPWR _3232_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_59_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1334 wire1335/X VGND VGND VPWR VPWR _5708_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1345 _4487_/B VGND VGND VPWR VPWR _4846_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_47_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1356 wire1357/X VGND VGND VPWR VPWR wire1356/X sky130_fd_sc_hd__buf_6
XFILLER_86_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1367 _3920_/X VGND VGND VPWR VPWR wire1367/X sky130_fd_sc_hd__clkbuf_1
Xwire1378 hold63/X VGND VGND VPWR VPWR _3454_/B sky130_fd_sc_hd__clkbuf_1
Xwire1389 _3536_/B VGND VGND VPWR VPWR _3726_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire620 wire621/X VGND VGND VPWR VPWR wire620/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire631 _5471_/S VGND VGND VPWR VPWR wire631/X sky130_fd_sc_hd__clkbuf_1
Xwire642 _5455_/S VGND VGND VPWR VPWR _5453_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_183_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire664 _5417_/S VGND VGND VPWR VPWR _5415_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3971 _6685_/RESET_B VGND VGND VPWR VPWR fanout3964/A sky130_fd_sc_hd__buf_2
Xwire675 _5402_/S VGND VGND VPWR VPWR _5399_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire686 _5372_/S VGND VGND VPWR VPWR _5375_/S sky130_fd_sc_hd__clkbuf_2
Xwire697 _5348_/S VGND VGND VPWR VPWR _5345_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3270 _5225_/B VGND VGND VPWR VPWR _5286_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_38_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3292 wire3293/X VGND VGND VPWR VPWR wire3292/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2580 _6183_/A2 VGND VGND VPWR VPWR wire2580/X sky130_fd_sc_hd__clkbuf_1
Xwire2591 _5691_/Y VGND VGND VPWR VPWR _5836_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1890 _6952_/Q VGND VGND VPWR VPWR _6190_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5950_ _6333_/B2 _5950_/A2 _5950_/B1 _6326_/A1 _5949_/X VGND VGND VPWR VPWR _5957_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_46_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4901_ _5027_/A _5152_/A1 _4679_/B _5152_/B2 _4901_/B1 VGND VGND VPWR VPWR _4901_/X
+ sky130_fd_sc_hd__a41o_1
X_5881_ _5969_/A1 _5881_/A2 _5880_/X VGND VGND VPWR VPWR _5881_/X sky130_fd_sc_hd__a21o_1
XFILLER_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4832_ _4932_/A _4832_/B _4839_/B VGND VGND VPWR VPWR _4843_/B sky130_fd_sc_hd__nor3_1
XFILLER_21_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4763_ _4763_/A1 _4448_/B _4753_/Y _4762_/X VGND VGND VPWR VPWR _4764_/C sky130_fd_sc_hd__a211o_1
XFILLER_159_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6502_ _7131_/CLK _6502_/D wire4058/A VGND VGND VPWR VPWR _6502_/Q sky130_fd_sc_hd__dfrtp_1
X_3714_ _3714_/A _3714_/B VGND VGND VPWR VPWR _5229_/A sky130_fd_sc_hd__nor2_1
X_4694_ _4694_/A _4694_/B VGND VGND VPWR VPWR _4694_/X sky130_fd_sc_hd__or2_1
XFILLER_174_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6433_ _6433_/A _6433_/B VGND VGND VPWR VPWR _6433_/X sky130_fd_sc_hd__and2_1
X_3645_ _3645_/A1 _3645_/A2 _3767_/B1 _3645_/B2 VGND VGND VPWR VPWR _3645_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6364_ _4228_/C _6364_/A2 _6364_/B1 _4228_/A _6363_/X VGND VGND VPWR VPWR _6364_/X
+ sky130_fd_sc_hd__a221o_1
X_3576_ _5758_/A1 wire960/X wire832/X _3576_/B2 VGND VGND VPWR VPWR _3576_/X sky130_fd_sc_hd__a22o_1
XFILLER_136_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5315_ _5396_/A1 _6066_/B2 _5318_/S VGND VGND VPWR VPWR _6899_/D sky130_fd_sc_hd__mux2_1
X_6295_ _7185_/Q _6319_/S wire444/X _6294_/X VGND VGND VPWR VPWR _7185_/D sky130_fd_sc_hd__o22a_1
XFILLER_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5246_ _5246_/A0 hold164/X _5248_/S VGND VGND VPWR VPWR _6838_/D sky130_fd_sc_hd__mux2_1
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold16 hold16/A VGND VGND VPWR VPWR hold16/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold27 hold27/A VGND VGND VPWR VPWR hold27/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold38 hold38/A VGND VGND VPWR VPWR hold38/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 hold49/A VGND VGND VPWR VPWR hold49/X sky130_fd_sc_hd__dlygate4sd3_1
X_5177_ _5177_/A _5177_/B _5176_/X VGND VGND VPWR VPWR _5178_/D sky130_fd_sc_hd__or3b_1
X_4128_ _5552_/A0 hold419/X _4128_/S VGND VGND VPWR VPWR _6595_/D sky130_fd_sc_hd__mux2_1
XFILLER_29_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4059_ hold646/X _4058_/X _4061_/S VGND VGND VPWR VPWR _6548_/D sky130_fd_sc_hd__mux2_1
XFILLER_43_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_662 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length3234 _4367_/Y VGND VGND VPWR VPWR _4471_/B sky130_fd_sc_hd__clkbuf_1
Xmax_length2500 _6055_/B1 VGND VGND VPWR VPWR _6079_/B1 sky130_fd_sc_hd__clkbuf_1
Xmax_length3256 _5535_/B VGND VGND VPWR VPWR _5430_/B sky130_fd_sc_hd__clkbuf_2
Xmax_length2533 _6001_/Y VGND VGND VPWR VPWR _6025_/A sky130_fd_sc_hd__clkbuf_1
Xmax_length3278 _5475_/B VGND VGND VPWR VPWR _5493_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_137_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length1854 _6988_/Q VGND VGND VPWR VPWR wire1853/A sky130_fd_sc_hd__clkbuf_1
XFILLER_106_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1131 _3332_/Y VGND VGND VPWR VPWR _3533_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1142 _3401_/A2 VGND VGND VPWR VPWR _3368_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_86_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1153 _3635_/B1 VGND VGND VPWR VPWR _3364_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_19_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1164 _3746_/A2 VGND VGND VPWR VPWR _3666_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_35_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1197 _3615_/B1 VGND VGND VPWR VPWR _3744_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_80_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6755_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_7_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire450 wire451/X VGND VGND VPWR VPWR wire450/X sky130_fd_sc_hd__clkbuf_1
Xwire461 wire462/X VGND VGND VPWR VPWR wire461/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire472 _5570_/S VGND VGND VPWR VPWR _5565_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_183_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire483 wire483/A VGND VGND VPWR VPWR _5546_/S sky130_fd_sc_hd__clkbuf_1
XFILLER_156_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold508 _6999_/Q VGND VGND VPWR VPWR hold508/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire494 _5320_/S VGND VGND VPWR VPWR _5319_/S sky130_fd_sc_hd__clkbuf_1
Xhold519 _6917_/Q VGND VGND VPWR VPWR hold519/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3430_ _3430_/A1 _5232_/A _5580_/A _7140_/Q _3418_/X VGND VGND VPWR VPWR _3431_/D
+ sky130_fd_sc_hd__a221o_1
X_3361_ _3361_/A1 _3361_/A2 _3361_/B1 _3361_/B2 _3360_/X VGND VGND VPWR VPWR _3373_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_124_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5100_ _5100_/A _5140_/A _5142_/B _5100_/D VGND VGND VPWR VPWR _5101_/D sky130_fd_sc_hd__or4_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6080_ _6080_/A1 _6140_/A2 _6124_/A2 _7052_/Q VGND VGND VPWR VPWR _6080_/X sky130_fd_sc_hd__a22o_1
X_3292_ _3536_/A _3339_/B VGND VGND VPWR VPWR _3292_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _5031_/A _5031_/B _5031_/C VGND VGND VPWR VPWR _5031_/X sky130_fd_sc_hd__or3_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6982_ _7068_/CLK _6982_/D wire4007/X VGND VGND VPWR VPWR _6982_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_81_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5933_ _6305_/A1 _5953_/B1 _5961_/A2 _5933_/B2 VGND VGND VPWR VPWR _5933_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_33_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7131_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_15_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5864_ _6231_/B2 _5930_/B1 _5912_/B1 _5864_/B2 _5863_/X VGND VGND VPWR VPWR _5869_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4815_ _4815_/A _4987_/C _4815_/C _4814_/X VGND VGND VPWR VPWR _4817_/C sky130_fd_sc_hd__or4b_1
XFILLER_21_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5795_ _7166_/Q _5794_/X _6171_/S VGND VGND VPWR VPWR _7166_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_48_csclk clkbuf_opt_2_0_csclk/X VGND VGND VPWR VPWR _6921_/CLK sky130_fd_sc_hd__clkbuf_16
X_4746_ _4748_/A _4994_/A VGND VGND VPWR VPWR _4746_/Y sky130_fd_sc_hd__nor2_1
XFILLER_193_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4677_ _4677_/A _4677_/B VGND VGND VPWR VPWR _5054_/B sky130_fd_sc_hd__or2_1
Xmax_length1117 _3652_/A2 VGND VGND VPWR VPWR _3486_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_135_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6416_ _6432_/A _6432_/B VGND VGND VPWR VPWR _6416_/X sky130_fd_sc_hd__and2_1
X_3628_ _5922_/B2 _3747_/B1 wire804/X _5922_/A1 _3609_/X VGND VGND VPWR VPWR _3632_/A
+ sky130_fd_sc_hd__a221o_1
X_6347_ _7188_/Q _3888_/Y _6346_/Y _6345_/X VGND VGND VPWR VPWR _7188_/D sky130_fd_sc_hd__a31o_1
XFILLER_103_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3559_ _3559_/A1 _3287_/Y _4324_/A _6769_/Q VGND VGND VPWR VPWR _3559_/X sky130_fd_sc_hd__a22o_1
XFILLER_103_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6278_ _6278_/A1 _6278_/A2 _6278_/B1 _6758_/Q _6277_/X VGND VGND VPWR VPWR _6280_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput106 wb_adr_i[16] VGND VGND VPWR VPWR _4337_/B sky130_fd_sc_hd__clkbuf_1
Xinput117 wb_adr_i[26] VGND VGND VPWR VPWR input117/X sky130_fd_sc_hd__clkbuf_1
XFILLER_130_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput128 wb_adr_i[7] VGND VGND VPWR VPWR _4553_/A sky130_fd_sc_hd__buf_6
XFILLER_48_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput139 wb_dat_i[16] VGND VGND VPWR VPWR _6363_/A2 sky130_fd_sc_hd__clkbuf_1
X_5229_ _5229_/A _5229_/B VGND VGND VPWR VPWR _5231_/S sky130_fd_sc_hd__nand2_1
XFILLER_29_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_90 _5990_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3097 _5848_/A2 VGND VGND VPWR VPWR wire3092/A sky130_fd_sc_hd__clkbuf_1
XFILLER_153_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_79_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4600_ _4367_/B _5106_/A _4574_/Y _4600_/C1 _5127_/A VGND VGND VPWR VPWR _4600_/X
+ sky130_fd_sc_hd__a2111o_1
X_5580_ _5580_/A _5580_/B VGND VGND VPWR VPWR _5586_/S sky130_fd_sc_hd__nand2_2
XFILLER_191_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4531_ _4846_/C _4369_/B _4464_/Y _5050_/A _4530_/X VGND VGND VPWR VPWR _4531_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_190_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold305 _6882_/Q VGND VGND VPWR VPWR hold305/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold316 _6517_/Q VGND VGND VPWR VPWR hold316/X sky130_fd_sc_hd__dlygate4sd3_1
X_4462_ _4591_/A _4462_/B VGND VGND VPWR VPWR _4462_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold327 _6962_/Q VGND VGND VPWR VPWR hold327/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 _6518_/Q VGND VGND VPWR VPWR hold338/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 _6683_/Q VGND VGND VPWR VPWR hold349/X sky130_fd_sc_hd__dlygate4sd3_1
X_6201_ _6201_/A1 _6201_/A2 _6201_/B1 _6201_/B2 _6198_/X VGND VGND VPWR VPWR _6201_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3413_ _7174_/Q _6816_/Q _6818_/Q VGND VGND VPWR VPWR _3413_/X sky130_fd_sc_hd__mux2_2
XFILLER_144_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4393_ _4351_/A _4351_/B _4391_/Y VGND VGND VPWR VPWR _4393_/X sky130_fd_sc_hd__a21o_1
X_7181_ _3937_/A1 _7181_/D wire4015/X VGND VGND VPWR VPWR _7181_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3344_ _3344_/A _3546_/B VGND VGND VPWR VPWR _3344_/Y sky130_fd_sc_hd__nor2_1
X_6132_ _6132_/A1 _6132_/A2 _6132_/B1 _6982_/Q _6132_/C1 VGND VGND VPWR VPWR _6132_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_98_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3275_ _3546_/A _3320_/A VGND VGND VPWR VPWR _3275_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6063_ _6063_/A1 _6138_/A2 _6063_/B1 _6063_/B2 VGND VGND VPWR VPWR _6063_/X sky130_fd_sc_hd__a22o_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5014_ _4400_/B _5013_/B _5105_/B2 VGND VGND VPWR VPWR _5015_/C sky130_fd_sc_hd__a21oi_1
XFILLER_39_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6965_ _7088_/CLK _6965_/D wire4069/X VGND VGND VPWR VPWR _6965_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5916_ _5916_/A _5960_/B VGND VGND VPWR VPWR _5916_/X sky130_fd_sc_hd__or2_1
XFILLER_179_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6896_ _6989_/CLK _6896_/D wire3995/X VGND VGND VPWR VPWR _6896_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5847_ _5847_/A _5847_/B _5847_/C _5847_/D VGND VGND VPWR VPWR _5847_/X sky130_fd_sc_hd__or4_1
XFILLER_22_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5778_ _5778_/A1 _5778_/A2 _5778_/B1 _5778_/B2 _5777_/X VGND VGND VPWR VPWR _5785_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_166_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length828 _3466_/Y VGND VGND VPWR VPWR _3678_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_154_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4729_ _4753_/A _4871_/B VGND VGND VPWR VPWR _4729_/Y sky130_fd_sc_hd__nand2_1
XFILLER_181_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3803 _4664_/B VGND VGND VPWR VPWR _4712_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3814 _4472_/X VGND VGND VPWR VPWR _4603_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3825 _4380_/X VGND VGND VPWR VPWR _4981_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_107_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3847 wire3847/A VGND VGND VPWR VPWR _5241_/C sky130_fd_sc_hd__clkbuf_2
Xwire3858 wire3859/X VGND VGND VPWR VPWR _3770_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire3869 wire3870/X VGND VGND VPWR VPWR wire3869/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6750_ _6963_/CLK _6750_/D _6401_/A VGND VGND VPWR VPWR _6750_/Q sky130_fd_sc_hd__dfrtp_1
X_3962_ _6700_/Q _3962_/B VGND VGND VPWR VPWR _6692_/D sky130_fd_sc_hd__and2_1
X_5701_ _5990_/A1 _5701_/A2 _5701_/B1 _5701_/B2 _5698_/X VGND VGND VPWR VPWR _5708_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6681_ _6683_/CLK _6681_/D fanout3964/A VGND VGND VPWR VPWR _6681_/Q sky130_fd_sc_hd__dfrtp_1
X_3893_ _6699_/Q _3876_/X _6694_/Q VGND VGND VPWR VPWR _6699_/D sky130_fd_sc_hd__a21o_1
XFILLER_188_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5632_ _7155_/Q _5637_/B _5631_/Y VGND VGND VPWR VPWR _7155_/D sky130_fd_sc_hd__a21oi_1
XFILLER_176_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5563_ _5563_/A0 hold216/X _5565_/S VGND VGND VPWR VPWR _7119_/D sky130_fd_sc_hd__mux2_1
XFILLER_157_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4514_ _4516_/B _4514_/B VGND VGND VPWR VPWR _4863_/A sky130_fd_sc_hd__nand2_1
Xhold102 _6581_/Q VGND VGND VPWR VPWR hold102/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 _6464_/Q VGND VGND VPWR VPWR hold113/X sky130_fd_sc_hd__dlygate4sd3_1
X_5494_ _5554_/A0 hold328/X _5494_/S VGND VGND VPWR VPWR _7058_/D sky130_fd_sc_hd__mux2_1
Xhold124 _6857_/Q VGND VGND VPWR VPWR hold124/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 _6854_/Q VGND VGND VPWR VPWR hold135/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold146 _6708_/Q VGND VGND VPWR VPWR hold146/X sky130_fd_sc_hd__dlygate4sd3_1
X_4445_ _4445_/A _4724_/B VGND VGND VPWR VPWR _4872_/A sky130_fd_sc_hd__or2_4
Xhold157 _6470_/Q VGND VGND VPWR VPWR _3242_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 _3301_/X VGND VGND VPWR VPWR hold168/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold179 _5463_/X VGND VGND VPWR VPWR _7031_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7164_ _3937_/A1 _7164_/D _7176_/RESET_B VGND VGND VPWR VPWR _7164_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_144_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4376_ _4376_/A _4951_/B VGND VGND VPWR VPWR _4492_/A sky130_fd_sc_hd__nand2_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6115_ _6115_/A1 _6214_/A2 _6115_/B1 _6115_/B2 VGND VGND VPWR VPWR _6115_/X sky130_fd_sc_hd__a22o_1
XFILLER_112_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3327_ _5212_/B _3534_/A VGND VGND VPWR VPWR _3327_/Y sky130_fd_sc_hd__nor2_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7095_ _7115_/CLK _7095_/D wire3981/X VGND VGND VPWR VPWR _7095_/Q sky130_fd_sc_hd__dfstp_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1708 wire1709/X VGND VGND VPWR VPWR wire1708/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1719 wire1720/X VGND VGND VPWR VPWR _6037_/B2 sky130_fd_sc_hd__clkbuf_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ _6842_/Q _6046_/B VGND VGND VPWR VPWR _6046_/X sky130_fd_sc_hd__or2_1
X_3258_ _3257_/X _3258_/A1 _3941_/A VGND VGND VPWR VPWR _3258_/X sky130_fd_sc_hd__mux2_1
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3189_ _3189_/A VGND VGND VPWR VPWR _3189_/Y sky130_fd_sc_hd__inv_2
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6948_ _7135_/CLK _6948_/D _7035_/SET_B VGND VGND VPWR VPWR _6948_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_41_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6879_ _7134_/CLK _6879_/D _7134_/RESET_B VGND VGND VPWR VPWR _6879_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_10_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length614 _5501_/S VGND VGND VPWR VPWR wire613/A sky130_fd_sc_hd__clkbuf_1
XFILLER_139_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length647 _5448_/Y VGND VGND VPWR VPWR _5455_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_154_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4301 _4570_/D VGND VGND VPWR VPWR _4398_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_163_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3611 _5459_/A0 VGND VGND VPWR VPWR _5220_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold680 _6927_/Q VGND VGND VPWR VPWR hold680/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3622 _6393_/A0 VGND VGND VPWR VPWR _5530_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_150_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold691 _6556_/Q VGND VGND VPWR VPWR hold691/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire2910 _5820_/B1 VGND VGND VPWR VPWR _5695_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire3655 _5269_/A0 VGND VGND VPWR VPWR _5314_/A0 sky130_fd_sc_hd__clkbuf_1
Xwire3666 wire3667/X VGND VGND VPWR VPWR wire3666/X sky130_fd_sc_hd__clkbuf_1
Xwire2921 _5786_/A2 VGND VGND VPWR VPWR _5745_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3677 _3241_/X VGND VGND VPWR VPWR _3791_/A sky130_fd_sc_hd__clkbuf_4
Xwire2932 wire2933/X VGND VGND VPWR VPWR wire2932/X sky130_fd_sc_hd__clkbuf_1
Xwire2943 _5691_/B VGND VGND VPWR VPWR _5829_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3688 wire3689/X VGND VGND VPWR VPWR _5850_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_49_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2954 _5688_/X VGND VGND VPWR VPWR _5842_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire3699 _5858_/C1 VGND VGND VPWR VPWR _6169_/C1 sky130_fd_sc_hd__clkbuf_2
Xwire2965 _5934_/A2 VGND VGND VPWR VPWR _5964_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_134_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2976 _5931_/A2 VGND VGND VPWR VPWR _5959_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire2987 _5843_/B1 VGND VGND VPWR VPWR _5799_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire2998 wire2999/X VGND VGND VPWR VPWR _5949_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput207 _3230_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[4] sky130_fd_sc_hd__buf_12
XFILLER_126_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput218 _3937_/X VGND VGND VPWR VPWR mgmt_gpio_out[14] sky130_fd_sc_hd__clkbuf_1
Xoutput229 _6826_/Q VGND VGND VPWR VPWR mgmt_gpio_out[24] sky130_fd_sc_hd__buf_12
XFILLER_99_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4230_ _6692_/Q _6693_/Q _6695_/Q _6694_/Q VGND VGND VPWR VPWR _4230_/X sky130_fd_sc_hd__or4_1
XFILLER_99_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4161_ hold369/X _4200_/A1 _4162_/S VGND VGND VPWR VPWR _4161_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4092_ _6836_/Q _4092_/A1 _4100_/S VGND VGND VPWR VPWR _4092_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6802_ _6803_/CLK _6802_/D wire3950/A VGND VGND VPWR VPWR _6802_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_91_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4994_ _4994_/A _5003_/B VGND VGND VPWR VPWR _5008_/A sky130_fd_sc_hd__nor2_1
XFILLER_168_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6733_ _6755_/CLK _6733_/D fanout3952/X VGND VGND VPWR VPWR _6733_/Q sky130_fd_sc_hd__dfstp_1
X_3945_ _3945_/A0 _3945_/A1 _6459_/Q VGND VGND VPWR VPWR _3945_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6664_ _6701_/CLK _6664_/D wire3945/X VGND VGND VPWR VPWR _6664_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3876_ _3877_/A1 _3965_/A1 _4120_/C VGND VGND VPWR VPWR _3876_/X sky130_fd_sc_hd__o21a_1
XFILLER_176_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5615_ _5615_/A _6564_/Q VGND VGND VPWR VPWR _5643_/A sky130_fd_sc_hd__nor2_1
X_6595_ _7110_/CLK _6595_/D wire3999/X VGND VGND VPWR VPWR _6595_/Q sky130_fd_sc_hd__dfrtp_1
Xmax_length2929 _5783_/C1 VGND VGND VPWR VPWR _5768_/C1 sky130_fd_sc_hd__clkbuf_1
XFILLER_136_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5546_ _5582_/A0 hold470/X _5546_/S VGND VGND VPWR VPWR _7104_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5477_ _5477_/A0 hold94/X _5480_/S VGND VGND VPWR VPWR _7043_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4428_ _4591_/A _4428_/B VGND VGND VPWR VPWR _4944_/B sky130_fd_sc_hd__nand2_1
Xwire2206 _6732_/Q VGND VGND VPWR VPWR _6253_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_160_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2217 _6719_/Q VGND VGND VPWR VPWR _6308_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7147_ _7187_/CLK _7147_/D _7161_/RESET_B VGND VGND VPWR VPWR _7147_/Q sky130_fd_sc_hd__dfrtp_1
Xwire2228 _6713_/Q VGND VGND VPWR VPWR _3630_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
X_4359_ _4575_/B _4359_/B VGND VGND VPWR VPWR _4363_/B sky130_fd_sc_hd__xnor2_1
Xwire2239 wire2240/X VGND VGND VPWR VPWR _6225_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_98_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1505 wire1506/X VGND VGND VPWR VPWR wire1505/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1516 wire1517/X VGND VGND VPWR VPWR _4111_/B sky130_fd_sc_hd__clkbuf_2
Xwire1527 hold117/X VGND VGND VPWR VPWR _3518_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7078_ _7142_/CLK _7078_/D wire4039/X VGND VGND VPWR VPWR _7078_/Q sky130_fd_sc_hd__dfrtp_1
Xwire1538 wire1539/X VGND VGND VPWR VPWR _3509_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire1549 _7128_/Q VGND VGND VPWR VPWR wire1549/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6029_ _6040_/B _6029_/B _6029_/C _6029_/D VGND VGND VPWR VPWR _6029_/X sky130_fd_sc_hd__or4_1
XFILLER_73_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire802 _3531_/Y VGND VGND VPWR VPWR wire802/X sky130_fd_sc_hd__dlymetal6s2s_1
Xwire813 _3504_/Y VGND VGND VPWR VPWR wire813/X sky130_fd_sc_hd__clkbuf_2
Xwire824 _3479_/X VGND VGND VPWR VPWR wire824/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire835 _3451_/Y VGND VGND VPWR VPWR wire835/X sky130_fd_sc_hd__clkbuf_1
XFILLER_182_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire846 _3422_/X VGND VGND VPWR VPWR wire846/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire857 _3347_/X VGND VGND VPWR VPWR wire857/X sky130_fd_sc_hd__clkbuf_1
Xwire868 _3342_/Y VGND VGND VPWR VPWR wire868/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout4047 fanout4047/A VGND VGND VPWR VPWR wire4049/A sky130_fd_sc_hd__clkbuf_2
Xwire4120 wire4121/X VGND VGND VPWR VPWR _7215_/A sky130_fd_sc_hd__clkbuf_1
Xwire4131 wire4132/X VGND VGND VPWR VPWR _3958_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_151_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4142 wire4143/X VGND VGND VPWR VPWR _3756_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire4153 wire4154/X VGND VGND VPWR VPWR wire4153/X sky130_fd_sc_hd__clkbuf_1
Xwire4164 input57/X VGND VGND VPWR VPWR _3430_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_145_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3430 _5427_/A0 VGND VGND VPWR VPWR _5454_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire4175 wire4176/X VGND VGND VPWR VPWR wire4175/X sky130_fd_sc_hd__clkbuf_1
Xwire3441 wire3442/X VGND VGND VPWR VPWR wire3441/X sky130_fd_sc_hd__clkbuf_1
Xwire4186 wire4187/X VGND VGND VPWR VPWR _3444_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire3452 _4323_/A1 VGND VGND VPWR VPWR _4335_/A0 sky130_fd_sc_hd__clkbuf_1
Xwire4197 wire4198/X VGND VGND VPWR VPWR wire4197/X sky130_fd_sc_hd__clkbuf_1
Xwire3463 _5255_/A1 VGND VGND VPWR VPWR _5309_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3474 _5480_/A0 VGND VGND VPWR VPWR _4305_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2740 _6335_/B1 VGND VGND VPWR VPWR _6290_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_77_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3485 wire3486/X VGND VGND VPWR VPWR wire3485/X sky130_fd_sc_hd__clkbuf_1
Xwire2751 wire2752/X VGND VGND VPWR VPWR _6340_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire2762 _6093_/A2 VGND VGND VPWR VPWR _6330_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire2773 _6127_/A2 VGND VGND VPWR VPWR _6150_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2784 _5992_/X VGND VGND VPWR VPWR _6184_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2795 _6200_/A2 VGND VGND VPWR VPWR _6103_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_92_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3730_ _6460_/Q _6445_/Q _6811_/Q VGND VGND VPWR VPWR _3730_/X sky130_fd_sc_hd__or3_2
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3661_ wire364/X _6784_/Q _3791_/A VGND VGND VPWR VPWR _3661_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5400_ hold535/X _5517_/A0 _5400_/S VGND VGND VPWR VPWR _6975_/D sky130_fd_sc_hd__mux2_1
X_6380_ _6379_/X _7202_/Q _6386_/S VGND VGND VPWR VPWR _7202_/D sky130_fd_sc_hd__mux2_1
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3592_ input6/X _3777_/A2 _3763_/A2 input29/X wire784/X VGND VGND VPWR VPWR _3593_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5331_ _5331_/A _5562_/B VGND VGND VPWR VPWR _5331_/Y sky130_fd_sc_hd__nand2_1
X_5262_ _5352_/A0 hold447/X _5264_/S VGND VGND VPWR VPWR _6852_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7001_ _7001_/CLK _7001_/D wire3996/A VGND VGND VPWR VPWR _7001_/Q sky130_fd_sc_hd__dfrtp_1
X_4213_ hold394/X _4237_/A0 _4215_/S VGND VGND VPWR VPWR _6667_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5193_ _5193_/A _5193_/B VGND VGND VPWR VPWR _5199_/S sky130_fd_sc_hd__nand2_2
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4144_ _4255_/A1 _6608_/Q _4146_/S VGND VGND VPWR VPWR _4144_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4075_ hold589/X _5208_/A1 _4079_/S VGND VGND VPWR VPWR _4075_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_4_0_csclk clkbuf_3_5_0_csclk/A VGND VGND VPWR VPWR _7059_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_51_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4977_ _5094_/B _4971_/Y _4976_/X VGND VGND VPWR VPWR _5145_/A sky130_fd_sc_hd__o21ai_1
XFILLER_149_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6716_ _7036_/CLK _6716_/D wire3974/X VGND VGND VPWR VPWR _6716_/Q sky130_fd_sc_hd__dfrtp_1
X_3928_ _3928_/A0 _3928_/A1 _3928_/S VGND VGND VPWR VPWR _3928_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6647_ _7206_/CLK _6647_/D VGND VGND VPWR VPWR _6647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3859_ _3859_/A1 _3856_/B _3853_/B _6453_/Q _3858_/X VGND VGND VPWR VPWR _6453_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_164_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6578_ _6939_/CLK hold17/X _6923_/SET_B VGND VGND VPWR VPWR _6578_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5529_ _5529_/A _5529_/B VGND VGND VPWR VPWR _5533_/S sky130_fd_sc_hd__and2_1
XFILLER_133_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2014 _5831_/A1 VGND VGND VPWR VPWR wire2014/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2025 _6197_/B2 VGND VGND VPWR VPWR wire2025/X sky130_fd_sc_hd__clkbuf_1
Xwire2036 hold96/A VGND VGND VPWR VPWR _6100_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1302 _3595_/A2 VGND VGND VPWR VPWR _3682_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_115_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2047 _6870_/Q VGND VGND VPWR VPWR wire2047/X sky130_fd_sc_hd__clkbuf_1
Xwire1313 wire1314/X VGND VGND VPWR VPWR wire1313/X sky130_fd_sc_hd__clkbuf_1
Xwire2058 _6866_/Q VGND VGND VPWR VPWR _6010_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2069 _6860_/Q VGND VGND VPWR VPWR _6077_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1324 _5878_/X VGND VGND VPWR VPWR _5879_/D sky130_fd_sc_hd__clkbuf_1
Xwire1335 wire1336/X VGND VGND VPWR VPWR wire1335/X sky130_fd_sc_hd__clkbuf_1
XFILLER_75_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1346 _5003_/A VGND VGND VPWR VPWR _4743_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_115_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1357 wire1358/X VGND VGND VPWR VPWR wire1357/X sky130_fd_sc_hd__clkbuf_1
Xwire1368 hold70/X VGND VGND VPWR VPWR _4070_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1379 wire1379/A VGND VGND VPWR VPWR _3417_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_86_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire610 _5498_/S VGND VGND VPWR VPWR _5495_/S sky130_fd_sc_hd__dlymetal6s2s_1
Xwire621 _5484_/Y VGND VGND VPWR VPWR wire621/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire632 _5474_/S VGND VGND VPWR VPWR _5471_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_11_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire643 wire644/X VGND VGND VPWR VPWR _5450_/S sky130_fd_sc_hd__clkbuf_1
XFILLER_128_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire654 wire654/A VGND VGND VPWR VPWR _5440_/S sky130_fd_sc_hd__clkbuf_2
Xmax_length3972 wire3970/A VGND VGND VPWR VPWR _6685_/RESET_B sky130_fd_sc_hd__clkbuf_2
XFILLER_183_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire676 _5402_/S VGND VGND VPWR VPWR _5400_/S sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_length3983 wire3984/X VGND VGND VPWR VPWR _7185_/RESET_B sky130_fd_sc_hd__clkbuf_2
Xmax_length3994 wire3996/A VGND VGND VPWR VPWR _7141_/RESET_B sky130_fd_sc_hd__clkbuf_2
Xwire698 _5339_/S VGND VGND VPWR VPWR _5338_/S sky130_fd_sc_hd__clkbuf_1
XFILLER_109_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3260 wire3260/A VGND VGND VPWR VPWR _4282_/B sky130_fd_sc_hd__clkbuf_1
Xwire3271 _5553_/B VGND VGND VPWR VPWR _5580_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3282 _4222_/B VGND VGND VPWR VPWR _5223_/B sky130_fd_sc_hd__clkbuf_2
Xwire3293 wire3294/X VGND VGND VPWR VPWR wire3293/X sky130_fd_sc_hd__clkbuf_1
XFILLER_172_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2570 _6075_/B1 VGND VGND VPWR VPWR _6197_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2581 _6023_/A VGND VGND VPWR VPWR _6183_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2592 _5028_/X VGND VGND VPWR VPWR _5029_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_93_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1880 _6067_/B2 VGND VGND VPWR VPWR _3672_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire1891 _6949_/Q VGND VGND VPWR VPWR _3221_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_65_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4900_ _5023_/B _5016_/A VGND VGND VPWR VPWR _4900_/X sky130_fd_sc_hd__and2_1
X_5880_ _6243_/A1 _5946_/A2 _5869_/X _5879_/X _5946_/C1 VGND VGND VPWR VPWR _5880_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4831_ _4940_/B _4831_/A2 _4524_/Y VGND VGND VPWR VPWR _5162_/A sky130_fd_sc_hd__o21ai_1
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4762_ _4763_/A1 _4460_/A _4984_/B _4761_/X VGND VGND VPWR VPWR _4762_/X sky130_fd_sc_hd__a211o_1
X_6501_ _7134_/CLK _6501_/D _6833_/RESET_B VGND VGND VPWR VPWR _6501_/Q sky130_fd_sc_hd__dfrtp_1
X_3713_ _6064_/A1 wire935/X wire919/X _6064_/B2 wire755/X VGND VGND VPWR VPWR _3721_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4693_ _4693_/A _4694_/A _4693_/C VGND VGND VPWR VPWR _4698_/B sky130_fd_sc_hd__or3_1
X_6432_ _6432_/A _6432_/B VGND VGND VPWR VPWR _6432_/X sky130_fd_sc_hd__and2_1
X_3644_ _6800_/Q _3417_/Y _4016_/A _6513_/Q _3643_/X VGND VGND VPWR VPWR _3644_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_106_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6363_ _4228_/B _6363_/A2 _6363_/B1 _4228_/Y VGND VGND VPWR VPWR _6363_/X sky130_fd_sc_hd__a22o_1
X_3575_ _3575_/A1 _3338_/Y wire808/X _3575_/B2 wire775/X VGND VGND VPWR VPWR _3575_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_136_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5314_ _5314_/A0 hold607/X _5314_/S VGND VGND VPWR VPWR _6898_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6294_ _7184_/Q _6343_/A2 _5650_/Y VGND VGND VPWR VPWR _6294_/X sky130_fd_sc_hd__o21ba_1
XFILLER_114_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5245_ _5389_/A0 hold228/X _5248_/S VGND VGND VPWR VPWR _6837_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold17 hold17/A VGND VGND VPWR VPWR hold17/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 hold28/A VGND VGND VPWR VPWR hold28/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 hold39/A VGND VGND VPWR VPWR hold39/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5176_ _4655_/B _5027_/B _5108_/B _4679_/B VGND VGND VPWR VPWR _5176_/X sky130_fd_sc_hd__o22a_1
XFILLER_152_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4127_ _4127_/A0 hold246/X _4127_/S VGND VGND VPWR VPWR _6594_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4058_ hold554/X _4114_/A0 _4060_/S VGND VGND VPWR VPWR _4058_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_5_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A VGND VGND VPWR VPWR _7193_/CLK sky130_fd_sc_hd__clkbuf_8
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length2512 _6006_/Y VGND VGND VPWR VPWR wire2506/A sky130_fd_sc_hd__clkbuf_1
XFILLER_138_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length3268 _4159_/B VGND VGND VPWR VPWR _4240_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_153_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1110 _3384_/B1 VGND VGND VPWR VPWR _3366_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire1121 _3340_/Y VGND VGND VPWR VPWR _3777_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1143 wire1144/X VGND VGND VPWR VPWR _3401_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire1154 wire1155/X VGND VGND VPWR VPWR _3635_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire1165 _3612_/A2 VGND VGND VPWR VPWR _3746_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1176 _3769_/B1 VGND VGND VPWR VPWR _5466_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1187 _3322_/Y VGND VGND VPWR VPWR _3581_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire1198 _3562_/B1 VGND VGND VPWR VPWR _5376_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire440 _3352_/X VGND VGND VPWR VPWR _3355_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_7_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire451 _6169_/X VGND VGND VPWR VPWR wire451/X sky130_fd_sc_hd__clkbuf_1
XFILLER_156_554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire462 _5902_/X VGND VGND VPWR VPWR wire462/X sky130_fd_sc_hd__clkbuf_1
XFILLER_171_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire484 _5550_/S VGND VGND VPWR VPWR _5547_/S sky130_fd_sc_hd__dlymetal6s2s_1
Xhold509 _6997_/Q VGND VGND VPWR VPWR hold509/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3360_ _7102_/Q _3421_/A2 _3357_/X _3359_/X VGND VGND VPWR VPWR _3360_/X sky130_fd_sc_hd__a211o_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3291_ _3303_/A _3293_/A VGND VGND VPWR VPWR _3339_/B sky130_fd_sc_hd__nand2_2
XFILLER_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5030_ _5030_/A _5073_/B _5079_/B _5029_/X VGND VGND VPWR VPWR _5030_/X sky130_fd_sc_hd__or4b_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3090 wire3091/X VGND VGND VPWR VPWR _5930_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_66_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6981_ _7140_/CLK _6981_/D wire4065/X VGND VGND VPWR VPWR _6981_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_80_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5932_ _6303_/A1 _5932_/A2 _5931_/X VGND VGND VPWR VPWR _5935_/C sky130_fd_sc_hd__a21o_1
XFILLER_18_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5863_ _6236_/A1 _5941_/A2 _5929_/B1 _6238_/A1 VGND VGND VPWR VPWR _5863_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4814_ _4814_/A _4814_/B _4814_/C VGND VGND VPWR VPWR _4814_/X sky130_fd_sc_hd__or3_1
X_5794_ _6121_/A1 _7165_/Q _5793_/X VGND VGND VPWR VPWR _5794_/X sky130_fd_sc_hd__a21o_1
XFILLER_193_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4745_ _4745_/A _4745_/B VGND VGND VPWR VPWR _4875_/B sky130_fd_sc_hd__nor2_1
XFILLER_21_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4676_ _4842_/A1 _4676_/A2 _4680_/B _4589_/B VGND VGND VPWR VPWR _4676_/X sky130_fd_sc_hd__o22a_1
XFILLER_174_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6415_ _6433_/A _6433_/B VGND VGND VPWR VPWR _6415_/X sky130_fd_sc_hd__and2_1
X_3627_ _3627_/A _3627_/B _3627_/C _3627_/D VGND VGND VPWR VPWR _3633_/C sky130_fd_sc_hd__or4_1
XFILLER_134_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6346_ _6346_/A _6697_/Q VGND VGND VPWR VPWR _6346_/Y sky130_fd_sc_hd__nand2_1
X_3558_ _6114_/A1 _3667_/A2 _3625_/B1 _3558_/B2 VGND VGND VPWR VPWR _3583_/A sky130_fd_sc_hd__a22o_1
XFILLER_1_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6277_ _6277_/A1 _6277_/A2 _6303_/B1 _6277_/B2 VGND VGND VPWR VPWR _6277_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3489_ _3538_/A _3489_/B VGND VGND VPWR VPWR _3489_/Y sky130_fd_sc_hd__nor2_1
Xinput107 wb_adr_i[17] VGND VGND VPWR VPWR _4337_/A sky130_fd_sc_hd__clkbuf_1
Xinput118 wb_adr_i[27] VGND VGND VPWR VPWR _3885_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_103_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5228_ hold511/X _5269_/A0 _5228_/S VGND VGND VPWR VPWR _6823_/D sky130_fd_sc_hd__mux2_1
Xinput129 wb_adr_i[8] VGND VGND VPWR VPWR _4339_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_56_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5159_ _5159_/A _5159_/B _5159_/C VGND VGND VPWR VPWR _5160_/C sky130_fd_sc_hd__nand3_1
XFILLER_29_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_1_0_csclk clkbuf_2_1_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_3_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length2320 _6614_/Q VGND VGND VPWR VPWR _5931_/A1 sky130_fd_sc_hd__clkbuf_1
XANTENNA_80 wire2240/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_91 _5990_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_579 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length1685 hold95/A VGND VGND VPWR VPWR wire1684/A sky130_fd_sc_hd__clkbuf_1
XFILLER_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4530_ _4530_/A _4530_/B _4530_/C _4530_/D VGND VGND VPWR VPWR _4530_/X sky130_fd_sc_hd__and4_1
XFILLER_117_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold306 _6611_/Q VGND VGND VPWR VPWR hold306/X sky130_fd_sc_hd__dlygate4sd3_1
X_4461_ _4461_/A _4461_/B VGND VGND VPWR VPWR _5126_/A sky130_fd_sc_hd__nor2_1
Xhold317 _4024_/X VGND VGND VPWR VPWR _6517_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold328 _7058_/Q VGND VGND VPWR VPWR hold328/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 _6672_/Q VGND VGND VPWR VPWR hold339/X sky130_fd_sc_hd__dlygate4sd3_1
X_6200_ _6905_/Q _6200_/A2 _6200_/B1 _6200_/B2 VGND VGND VPWR VPWR _6216_/B sky130_fd_sc_hd__a22o_1
X_3412_ _3411_/X _6789_/Q _3791_/B VGND VGND VPWR VPWR _6789_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_719 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7180_ _7180_/CLK _7180_/D _7185_/RESET_B VGND VGND VPWR VPWR _7180_/Q sky130_fd_sc_hd__dfrtp_1
X_4392_ _4390_/C _4390_/D _4467_/A _4389_/Y VGND VGND VPWR VPWR _4560_/A sky130_fd_sc_hd__a31o_1
XFILLER_171_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6131_ _6958_/Q _6131_/A2 _6131_/B1 _7062_/Q VGND VGND VPWR VPWR _6131_/X sky130_fd_sc_hd__a22o_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ _3466_/A _3546_/B VGND VGND VPWR VPWR _3343_/Y sky130_fd_sc_hd__nor2_1
XFILLER_97_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _6062_/A1 _6062_/A2 _6062_/B1 _6062_/B2 _6061_/X VGND VGND VPWR VPWR _6068_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ _3293_/A _3414_/B VGND VGND VPWR VPWR _3320_/A sky130_fd_sc_hd__nand2_2
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _5013_/A _5013_/B VGND VGND VPWR VPWR _5013_/X sky130_fd_sc_hd__or2_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6964_ _7046_/CLK _6964_/D wire4052/X VGND VGND VPWR VPWR hold91/A sky130_fd_sc_hd__dfrtp_1
XFILLER_81_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5915_ _5915_/A1 _5915_/A2 _5932_/A2 _6277_/A1 _5914_/X VGND VGND VPWR VPWR _5923_/A
+ sky130_fd_sc_hd__a221o_1
X_6895_ _7110_/CLK _6895_/D wire4004/X VGND VGND VPWR VPWR _6895_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5846_ _6213_/B2 _5846_/A2 _5846_/B1 _6212_/A1 _5845_/X VGND VGND VPWR VPWR _5846_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_167_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5777_ _5777_/A1 _5777_/A2 _5777_/B1 _6129_/A1 VGND VGND VPWR VPWR _5777_/X sky130_fd_sc_hd__a22o_1
Xmax_length807 wire808/X VGND VGND VPWR VPWR _3692_/A2 sky130_fd_sc_hd__clkbuf_1
X_4728_ _4735_/A _4728_/B VGND VGND VPWR VPWR _4728_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4659_ _4659_/A _4659_/B VGND VGND VPWR VPWR _5065_/B sky130_fd_sc_hd__nor2_1
XFILLER_174_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3804 _4664_/B VGND VGND VPWR VPWR _4685_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire3826 _4657_/B VGND VGND VPWR VPWR _4999_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6329_ _6329_/A1 _6329_/A2 _6329_/B1 _6329_/B2 VGND VGND VPWR VPWR _6329_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3848 _3872_/Y VGND VGND VPWR VPWR wire3848/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3859 wire3860/X VGND VGND VPWR VPWR wire3859/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length2150 _6774_/Q VGND VGND VPWR VPWR wire2148/A sky130_fd_sc_hd__clkbuf_1
XFILLER_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_32_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7129_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_180_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_47_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7064_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_75_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3961_ _6825_/Q _3961_/B VGND VGND VPWR VPWR _3961_/X sky130_fd_sc_hd__and2_1
XFILLER_63_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5700_ _7152_/Q _5706_/B _5700_/C VGND VGND VPWR VPWR _5700_/X sky130_fd_sc_hd__and3_1
XFILLER_188_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6680_ _7206_/CLK _6680_/D _6348_/B VGND VGND VPWR VPWR _6680_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3892_ _6698_/Q _3876_/X _6693_/Q VGND VGND VPWR VPWR _6698_/D sky130_fd_sc_hd__a21o_1
XFILLER_149_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5631_ _7155_/Q _5624_/B _5637_/B VGND VGND VPWR VPWR _5631_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_188_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5562_ _5562_/A _5562_/B VGND VGND VPWR VPWR _5569_/S sky130_fd_sc_hd__nand2_1
XFILLER_117_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4513_ _4516_/B _4521_/A VGND VGND VPWR VPWR _4515_/C sky130_fd_sc_hd__nand2_1
Xhold103 _7128_/Q VGND VGND VPWR VPWR hold103/X sky130_fd_sc_hd__dlygate4sd3_1
X_5493_ _5493_/A _5493_/B VGND VGND VPWR VPWR _5501_/S sky130_fd_sc_hd__nand2_1
Xhold114 _3807_/B VGND VGND VPWR VPWR hold114/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 _7118_/Q VGND VGND VPWR VPWR hold125/X sky130_fd_sc_hd__dlygate4sd3_1
X_4444_ _4434_/B _4444_/B VGND VGND VPWR VPWR _4444_/Y sky130_fd_sc_hd__nand2b_1
Xhold136 _6948_/Q VGND VGND VPWR VPWR hold136/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold147 _6677_/Q VGND VGND VPWR VPWR hold147/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 _3242_/X VGND VGND VPWR VPWR hold158/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold169 _5227_/X VGND VGND VPWR VPWR _6822_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7163_ _7185_/CLK _7163_/D _7176_/RESET_B VGND VGND VPWR VPWR _7163_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_125_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4375_ _4846_/A _4846_/B _4538_/A VGND VGND VPWR VPWR _4951_/B sky130_fd_sc_hd__nor3b_2
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6114_ _6114_/A1 _6114_/A2 _6211_/B1 _6114_/B2 _6113_/X VGND VGND VPWR VPWR _6119_/C
+ sky130_fd_sc_hd__a221o_1
X_3326_ _3714_/A _3534_/A VGND VGND VPWR VPWR _3326_/Y sky130_fd_sc_hd__nor2_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7094_ _7094_/CLK _7094_/D fanout3964/A VGND VGND VPWR VPWR _7094_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_100_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1709 _6113_/B2 VGND VGND VPWR VPWR wire1709/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _6045_/A _6045_/B _6045_/C VGND VGND VPWR VPWR _6045_/X sky130_fd_sc_hd__or3_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ hold24/X hold66/X _3820_/A VGND VGND VPWR VPWR _3257_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3188_ _6691_/Q VGND VGND VPWR VPWR _6346_/A sky130_fd_sc_hd__inv_2
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6947_ _7135_/CLK _6947_/D _7042_/SET_B VGND VGND VPWR VPWR _6947_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_156_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6878_ _7135_/CLK hold76/X wire4056/X VGND VGND VPWR VPWR hold75/A sky130_fd_sc_hd__dfrtp_1
XFILLER_139_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5829_ _6920_/Q _5829_/A2 _5829_/B1 _5829_/B2 VGND VGND VPWR VPWR _5829_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length604 _5506_/S VGND VGND VPWR VPWR _5505_/S sky130_fd_sc_hd__clkbuf_1
Xmax_length615 _5487_/S VGND VGND VPWR VPWR _5489_/S sky130_fd_sc_hd__clkbuf_1
Xmax_length626 _5483_/S VGND VGND VPWR VPWR wire625/A sky130_fd_sc_hd__clkbuf_1
XFILLER_108_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire4302 wire4302/A VGND VGND VPWR VPWR _4951_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_163_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout3517 wire3525/X VGND VGND VPWR VPWR wire3523/A sky130_fd_sc_hd__clkbuf_1
XFILLER_190_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3623 _6393_/A0 VGND VGND VPWR VPWR _4130_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold670 _7022_/Q VGND VGND VPWR VPWR hold670/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold681 _6846_/Q VGND VGND VPWR VPWR hold681/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 _6599_/Q VGND VGND VPWR VPWR hold692/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3645 _5476_/A0 VGND VGND VPWR VPWR _5554_/A0 sky130_fd_sc_hd__clkbuf_2
Xwire2900 _5696_/X VGND VGND VPWR VPWR _5698_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_78_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2911 _5840_/B1 VGND VGND VPWR VPWR _5811_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire3656 wire3656/A VGND VGND VPWR VPWR _5269_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_89_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3667 wire3668/X VGND VGND VPWR VPWR wire3667/X sky130_fd_sc_hd__clkbuf_1
Xwire2922 _5754_/A2 VGND VGND VPWR VPWR _5786_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire2933 _5690_/X VGND VGND VPWR VPWR wire2933/X sky130_fd_sc_hd__clkbuf_1
Xwire3689 _5705_/A VGND VGND VPWR VPWR wire3689/X sky130_fd_sc_hd__clkbuf_1
Xwire2966 wire2967/X VGND VGND VPWR VPWR _5934_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2977 wire2977/A VGND VGND VPWR VPWR _5931_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire2988 _5885_/B1 VGND VGND VPWR VPWR _5963_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2999 _5830_/A2 VGND VGND VPWR VPWR wire2999/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput208 _3229_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[5] sky130_fd_sc_hd__buf_12
XFILLER_154_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput219 _3936_/X VGND VGND VPWR VPWR mgmt_gpio_out[15] sky130_fd_sc_hd__clkbuf_1
XFILLER_126_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4160_ hold409/X _4211_/A1 _4162_/S VGND VGND VPWR VPWR _6621_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4091_ hold275/X _4090_/X _4101_/S VGND VGND VPWR VPWR _6567_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6801_ _6803_/CLK _6801_/D wire3950/A VGND VGND VPWR VPWR _6801_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_90_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4993_ _4993_/A _4993_/B VGND VGND VPWR VPWR _5036_/B sky130_fd_sc_hd__nor2_1
XFILLER_51_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6732_ _6803_/CLK _6732_/D fanout3952/X VGND VGND VPWR VPWR _6732_/Q sky130_fd_sc_hd__dfrtp_1
X_3944_ _6460_/Q _3946_/B VGND VGND VPWR VPWR _3944_/Y sky130_fd_sc_hd__nor2_1
XFILLER_177_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6663_ _6701_/CLK _6663_/D wire3945/A VGND VGND VPWR VPWR _6663_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3875_ _7160_/Q _6813_/Q _3940_/S VGND VGND VPWR VPWR _5592_/B sky130_fd_sc_hd__mux2_2
XFILLER_149_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5614_ _7149_/Q _7148_/Q VGND VGND VPWR VPWR _5706_/B sky130_fd_sc_hd__and2_2
XFILLER_149_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6594_ _6811_/CLK _6594_/D wire3948/A VGND VGND VPWR VPWR _6594_/Q sky130_fd_sc_hd__dfrtp_1
X_5545_ _5545_/A0 _7103_/Q _5547_/S VGND VGND VPWR VPWR _5545_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5476_ _5476_/A0 hold176/X _5480_/S VGND VGND VPWR VPWR _7042_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_3_0_0_csclk clkbuf_3_1_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_0_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_105_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7215_ _7215_/A VGND VGND VPWR VPWR _7215_/X sky130_fd_sc_hd__clkbuf_1
X_4427_ _4354_/A _4354_/B _4355_/Y _4350_/B VGND VGND VPWR VPWR _4427_/X sky130_fd_sc_hd__a211o_1
XFILLER_132_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2207 hold377/X VGND VGND VPWR VPWR _6228_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
X_7146_ _7180_/CLK _7146_/D _7161_/RESET_B VGND VGND VPWR VPWR _7146_/Q sky130_fd_sc_hd__dfrtp_1
X_4358_ _4407_/A _4359_/B VGND VGND VPWR VPWR _4360_/B sky130_fd_sc_hd__and2_1
Xwire2218 _6281_/A1 VGND VGND VPWR VPWR _3612_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_101_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2229 wire2230/X VGND VGND VPWR VPWR _5872_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_113_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1506 _3413_/X VGND VGND VPWR VPWR wire1506/X sky130_fd_sc_hd__clkbuf_1
X_3309_ hold62/X hold26/X _3301_/C VGND VGND VPWR VPWR hold63/A sky130_fd_sc_hd__or3b_1
Xwire1517 _3511_/A VGND VGND VPWR VPWR wire1517/X sky130_fd_sc_hd__clkbuf_1
XFILLER_98_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1528 _7211_/Q VGND VGND VPWR VPWR _3486_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_86_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7077_ _7124_/CLK _7077_/D wire4049/A VGND VGND VPWR VPWR _7077_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_86_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4289_ _5224_/A0 hold366/X _4293_/S VGND VGND VPWR VPWR _6736_/D sky130_fd_sc_hd__mux2_1
Xwire1539 _6123_/A1 VGND VGND VPWR VPWR wire1539/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6028_ _6040_/B _6029_/B _6029_/C _6029_/D VGND VGND VPWR VPWR _6028_/Y sky130_fd_sc_hd__nor4_1
XFILLER_100_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire803 _3528_/Y VGND VGND VPWR VPWR _4159_/A sky130_fd_sc_hd__clkbuf_1
Xwire814 _3504_/Y VGND VGND VPWR VPWR _4147_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xwire825 _3474_/Y VGND VGND VPWR VPWR wire825/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire836 _4174_/A VGND VGND VPWR VPWR wire836/X sky130_fd_sc_hd__dlymetal6s2s_1
Xwire847 wire848/X VGND VGND VPWR VPWR wire847/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire858 wire858/A VGND VGND VPWR VPWR wire858/X sky130_fd_sc_hd__clkbuf_1
XFILLER_108_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire869 wire871/X VGND VGND VPWR VPWR _5286_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_155_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4110 input68/X VGND VGND VPWR VPWR wire4110/X sky130_fd_sc_hd__clkbuf_1
Xwire4121 wire4122/X VGND VGND VPWR VPWR wire4121/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4132 wire4133/X VGND VGND VPWR VPWR wire4132/X sky130_fd_sc_hd__clkbuf_1
Xwire4143 wire4144/X VGND VGND VPWR VPWR wire4143/X sky130_fd_sc_hd__clkbuf_1
Xwire4154 wire4155/X VGND VGND VPWR VPWR wire4154/X sky130_fd_sc_hd__clkbuf_1
XFILLER_150_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3420 _5490_/A0 VGND VGND VPWR VPWR _5586_/A0 sky130_fd_sc_hd__clkbuf_2
Xwire4165 wire4166/X VGND VGND VPWR VPWR _3494_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire4176 input53/X VGND VGND VPWR VPWR wire4176/X sky130_fd_sc_hd__clkbuf_1
Xwire3431 _5541_/A1 VGND VGND VPWR VPWR _5427_/A0 sky130_fd_sc_hd__clkbuf_1
Xwire3442 wire3443/X VGND VGND VPWR VPWR wire3442/X sky130_fd_sc_hd__clkbuf_1
Xwire4187 wire4188/X VGND VGND VPWR VPWR wire4187/X sky130_fd_sc_hd__clkbuf_1
Xwire3453 _4033_/A1 VGND VGND VPWR VPWR _4323_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire4198 input46/X VGND VGND VPWR VPWR wire4198/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3464 _5540_/A1 VGND VGND VPWR VPWR _5255_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2730 _6009_/X VGND VGND VPWR VPWR wire2730/X sky130_fd_sc_hd__clkbuf_1
Xwire3475 _5567_/A0 VGND VGND VPWR VPWR _4281_/A0 sky130_fd_sc_hd__clkbuf_1
Xwire2741 _6225_/A2 VGND VGND VPWR VPWR _6335_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire3486 wire3486/A VGND VGND VPWR VPWR wire3486/X sky130_fd_sc_hd__clkbuf_1
Xwire2752 _6027_/B VGND VGND VPWR VPWR wire2752/X sky130_fd_sc_hd__clkbuf_1
Xwire3497 wire3498/X VGND VGND VPWR VPWR _3974_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_77_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2763 _6202_/A2 VGND VGND VPWR VPWR _6093_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2774 _6201_/A2 VGND VGND VPWR VPWR _6127_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_77_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2796 _6174_/A2 VGND VGND VPWR VPWR _6126_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3660_ _3660_/A _3660_/B _3660_/C VGND VGND VPWR VPWR _3660_/X sky130_fd_sc_hd__or3_1
XFILLER_9_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3591_ _6477_/Q _3966_/A _3992_/A _6493_/Q wire779/X VGND VGND VPWR VPWR _3593_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5330_ hold608/X _5339_/A0 _5330_/S VGND VGND VPWR VPWR _6913_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5261_ _5342_/A0 hold155/X _5263_/S VGND VGND VPWR VPWR _6851_/D sky130_fd_sc_hd__mux2_1
X_7000_ _7001_/CLK _7000_/D wire3992/X VGND VGND VPWR VPWR _7000_/Q sky130_fd_sc_hd__dfrtp_1
X_4212_ hold407/X _4248_/A0 _4215_/S VGND VGND VPWR VPWR _6666_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5192_ _5198_/A0 hold474/X _5192_/S VGND VGND VPWR VPWR _6797_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4143_ _6394_/A0 hold239/X _4146_/S VGND VGND VPWR VPWR _6607_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4074_ hold485/X _4073_/X _4084_/S VGND VGND VPWR VPWR _6555_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4976_ _4976_/A1 _4688_/B _4976_/B1 VGND VGND VPWR VPWR _4976_/X sky130_fd_sc_hd__a21o_1
X_6715_ _7208_/CLK _6715_/D _7112_/SET_B VGND VGND VPWR VPWR _6715_/Q sky130_fd_sc_hd__dfrtp_1
X_3927_ _3927_/A0 _3927_/A1 _3927_/S VGND VGND VPWR VPWR _3927_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3858_ _6541_/Q _3858_/B VGND VGND VPWR VPWR _3858_/X sky130_fd_sc_hd__and2b_1
X_6646_ _7193_/CLK _6646_/D VGND VGND VPWR VPWR _6646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length2705 _6203_/B1 VGND VGND VPWR VPWR _6111_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_192_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length2727 _6187_/B1 VGND VGND VPWR VPWR wire2726/A sky130_fd_sc_hd__clkbuf_1
X_3789_ _3789_/A _3789_/B _3789_/C _3789_/D VGND VGND VPWR VPWR _3789_/X sky130_fd_sc_hd__or4_1
X_6577_ _6701_/CLK _6577_/D wire3945/X VGND VGND VPWR VPWR _6577_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_117_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5528_ _5528_/A0 hold149/X _5528_/S VGND VGND VPWR VPWR _5528_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5459_ _5459_/A0 hold596/X _5462_/S VGND VGND VPWR VPWR _7027_/D sky130_fd_sc_hd__mux2_1
XFILLER_105_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2004 _6893_/Q VGND VGND VPWR VPWR _5758_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire2015 _6888_/Q VGND VGND VPWR VPWR _5831_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2026 _6881_/Q VGND VGND VPWR VPWR _6197_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2037 hold434/X VGND VGND VPWR VPWR _6075_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
X_7129_ _7129_/CLK _7129_/D wire4056/X VGND VGND VPWR VPWR _7129_/Q sky130_fd_sc_hd__dfrtp_1
Xwire1303 _3647_/A2 VGND VGND VPWR VPWR _3595_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire2048 wire2049/X VGND VGND VPWR VPWR _3189_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_59_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2059 _6865_/Q VGND VGND VPWR VPWR _5842_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1314 _6173_/X VGND VGND VPWR VPWR wire1314/X sky130_fd_sc_hd__clkbuf_1
XFILLER_47_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1325 _5846_/X VGND VGND VPWR VPWR _5847_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1336 wire1337/X VGND VGND VPWR VPWR wire1336/X sky130_fd_sc_hd__clkbuf_1
Xwire1347 _4486_/A VGND VGND VPWR VPWR _4753_/B sky130_fd_sc_hd__clkbuf_2
Xwire1358 wire1359/X VGND VGND VPWR VPWR wire1358/X sky130_fd_sc_hd__clkbuf_1
Xwire1369 _3489_/B VGND VGND VPWR VPWR _4120_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire600 _5514_/S VGND VGND VPWR VPWR wire600/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire611 wire613/A VGND VGND VPWR VPWR _5498_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire633 _5474_/S VGND VGND VPWR VPWR _5469_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire644 _5456_/S VGND VGND VPWR VPWR wire644/X sky130_fd_sc_hd__clkbuf_1
Xmax_length3951 wire3950/A VGND VGND VPWR VPWR _6495_/SET_B sky130_fd_sc_hd__buf_4
Xmax_length3962 _6437_/A VGND VGND VPWR VPWR _6438_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire677 _5391_/S VGND VGND VPWR VPWR _5388_/S sky130_fd_sc_hd__clkbuf_2
Xwire688 _5363_/S VGND VGND VPWR VPWR _5361_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_40_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire699 _5331_/Y VGND VGND VPWR VPWR _5339_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_170_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3250 _6392_/B VGND VGND VPWR VPWR _5229_/B sky130_fd_sc_hd__clkbuf_2
Xwire3261 _4318_/B VGND VGND VPWR VPWR wire3261/X sky130_fd_sc_hd__clkbuf_1
Xwire3272 _5520_/B VGND VGND VPWR VPWR _5571_/B sky130_fd_sc_hd__buf_2
Xwire3283 _4234_/B VGND VGND VPWR VPWR _4222_/B sky130_fd_sc_hd__clkbuf_2
Xwire3294 _3850_/X VGND VGND VPWR VPWR wire3294/X sky130_fd_sc_hd__clkbuf_1
XFILLER_93_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2560 _6328_/A2 VGND VGND VPWR VPWR _6264_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire2571 _6296_/B1 VGND VGND VPWR VPWR _6075_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2582 _5968_/A2 VGND VGND VPWR VPWR _5902_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_77_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2593 _4963_/B VGND VGND VPWR VPWR _4923_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_37_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1870 _6200_/B2 VGND VGND VPWR VPWR _5849_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1881 _6963_/Q VGND VGND VPWR VPWR _6067_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1892 _5766_/A1 VGND VGND VPWR VPWR _3568_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_92_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4830_ _4369_/X _4832_/B _4940_/A VGND VGND VPWR VPWR _4830_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4761_ _4761_/A _4761_/B _4761_/C _4760_/X VGND VGND VPWR VPWR _4761_/X sky130_fd_sc_hd__or4b_1
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3712_ _3712_/A1 _3547_/Y _3711_/Y _3712_/B2 VGND VGND VPWR VPWR _3712_/X sky130_fd_sc_hd__a22o_1
X_6500_ _7074_/CLK _6500_/D fanout3976/X VGND VGND VPWR VPWR _6500_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4692_ _4704_/A _4692_/B VGND VGND VPWR VPWR _4863_/B sky130_fd_sc_hd__or2_1
XFILLER_174_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6431_ _6441_/A _6431_/B VGND VGND VPWR VPWR _6431_/X sky130_fd_sc_hd__and2_1
X_3643_ _7209_/Q _6392_/A _5187_/A _6795_/Q VGND VGND VPWR VPWR _3643_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6362_ _6362_/A _6362_/B _6362_/C _6360_/X VGND VGND VPWR VPWR _6386_/S sky130_fd_sc_hd__or4b_4
X_3574_ _6684_/Q _3574_/A2 _3676_/A2 _3574_/B2 VGND VGND VPWR VPWR _3574_/X sky130_fd_sc_hd__a22o_1
X_5313_ _5313_/A _5553_/B VGND VGND VPWR VPWR _5320_/S sky130_fd_sc_hd__nand2_1
XFILLER_114_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6293_ _6293_/A1 wire977/X _6280_/X _6292_/X _6293_/C1 VGND VGND VPWR VPWR _6293_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_142_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5244_ _5244_/A0 hold611/X _5248_/S VGND VGND VPWR VPWR _6836_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold18 hold18/A VGND VGND VPWR VPWR hold18/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 hold29/A VGND VGND VPWR VPWR hold29/X sky130_fd_sc_hd__dlygate4sd3_1
X_5175_ _5137_/D _5174_/X _5148_/Y VGND VGND VPWR VPWR _5183_/B sky130_fd_sc_hd__o21a_1
XFILLER_69_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4126_ _5508_/A0 hold512/X _4128_/S VGND VGND VPWR VPWR _6593_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4057_ hold163/X _4056_/X _4061_/S VGND VGND VPWR VPWR _6547_/D sky130_fd_sc_hd__mux2_1
XFILLER_37_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4959_ _5123_/A _5163_/A _5163_/B VGND VGND VPWR VPWR _4959_/X sky130_fd_sc_hd__and3_1
XFILLER_184_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3203 _4496_/B VGND VGND VPWR VPWR _5094_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_177_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6629_ _7193_/CLK _6629_/D VGND VGND VPWR VPWR _6629_/Q sky130_fd_sc_hd__dfxtp_1
Xmax_length2546 _5999_/A2 VGND VGND VPWR VPWR _6277_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_193_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1100 _3501_/B1 VGND VGND VPWR VPWR _3403_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire1111 _3344_/Y VGND VGND VPWR VPWR _3384_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1122 _3340_/Y VGND VGND VPWR VPWR _3494_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1133 _3498_/A2 VGND VGND VPWR VPWR _3668_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire1144 _3329_/Y VGND VGND VPWR VPWR wire1144/X sky130_fd_sc_hd__clkbuf_1
Xwire1155 _3736_/B1 VGND VGND VPWR VPWR wire1155/X sky130_fd_sc_hd__clkbuf_1
XFILLER_75_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1166 _3436_/A2 VGND VGND VPWR VPWR _5358_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1177 _3323_/Y VGND VGND VPWR VPWR _3769_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1188 wire1189/X VGND VGND VPWR VPWR _3428_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire1199 _3615_/B1 VGND VGND VPWR VPWR _3562_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_142_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire430 _3572_/X VGND VGND VPWR VPWR wire430/X sky130_fd_sc_hd__clkbuf_1
XFILLER_156_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire441 wire442/X VGND VGND VPWR VPWR wire441/X sky130_fd_sc_hd__clkbuf_1
Xwire452 _6120_/X VGND VGND VPWR VPWR wire452/X sky130_fd_sc_hd__clkbuf_1
XFILLER_156_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire463 _5814_/X VGND VGND VPWR VPWR wire463/X sky130_fd_sc_hd__clkbuf_1
Xwire474 wire475/X VGND VGND VPWR VPWR _5560_/S sky130_fd_sc_hd__clkbuf_2
Xwire485 wire485/A VGND VGND VPWR VPWR _5550_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_7_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire496 wire497/X VGND VGND VPWR VPWR _5307_/S sky130_fd_sc_hd__buf_2
XFILLER_171_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3290_ _3472_/A _3536_/B VGND VGND VPWR VPWR _3290_/Y sky130_fd_sc_hd__nor2_1
XFILLER_97_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire3080 _5962_/A2 VGND VGND VPWR VPWR _5890_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire3091 _5821_/A2 VGND VGND VPWR VPWR wire3091/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2390 _6519_/Q VGND VGND VPWR VPWR _6314_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_93_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6980_ _7046_/CLK hold90/X wire4052/X VGND VGND VPWR VPWR hold89/A sky130_fd_sc_hd__dfrtp_1
XFILLER_81_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5931_ _5931_/A1 _5931_/A2 _5931_/B1 _5931_/B2 VGND VGND VPWR VPWR _5931_/X sky130_fd_sc_hd__a22o_1
XFILLER_81_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5862_ _7207_/Q _5943_/A2 _5963_/B1 _6223_/A1 _5861_/X VGND VGND VPWR VPWR _5869_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4813_ _4985_/C _4813_/B _4813_/C _4813_/D VGND VGND VPWR VPWR _4815_/C sky130_fd_sc_hd__or4_1
XFILLER_61_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5793_ _6846_/Q _5793_/A2 _5785_/X wire588/X _6095_/C1 VGND VGND VPWR VPWR _5793_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_178_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4744_ _4758_/A _4758_/B _4744_/C VGND VGND VPWR VPWR _4744_/X sky130_fd_sc_hd__and3_1
XFILLER_159_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4675_ _4675_/A _4675_/B VGND VGND VPWR VPWR _4675_/Y sky130_fd_sc_hd__nor2_1
XFILLER_147_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6414_ _6433_/A _6433_/B VGND VGND VPWR VPWR _6414_/X sky130_fd_sc_hd__and2_1
X_3626_ _3626_/A1 _4052_/B _4300_/A _3626_/B2 _3614_/X VGND VGND VPWR VPWR _3626_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6345_ _6346_/A _3888_/B _6692_/Q VGND VGND VPWR VPWR _6345_/X sky130_fd_sc_hd__o21a_1
X_3557_ _6108_/B2 _3557_/A2 _3557_/B1 _5755_/A1 VGND VGND VPWR VPWR _3557_/X sky130_fd_sc_hd__a22o_1
X_6276_ _6276_/A1 _6302_/A2 _6302_/B1 _6276_/B2 _6272_/X VGND VGND VPWR VPWR _6280_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_163_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3488_ hold75/A _5286_/A wire851/X _7214_/A VGND VGND VPWR VPWR _3488_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput108 wb_adr_i[18] VGND VGND VPWR VPWR _4337_/D sky130_fd_sc_hd__clkbuf_1
X_5227_ _5227_/A0 _5513_/A0 _5228_/S VGND VGND VPWR VPWR _5227_/X sky130_fd_sc_hd__mux2_1
Xinput119 wb_adr_i[28] VGND VGND VPWR VPWR _3885_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_102_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5158_ _5158_/A _5158_/B _5158_/C VGND VGND VPWR VPWR _5159_/C sky130_fd_sc_hd__nor3_1
XFILLER_186_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4109_ hold16/X _6578_/Q _4109_/S VGND VGND VPWR VPWR hold17/A sky130_fd_sc_hd__mux2_1
XFILLER_57_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5089_ _4753_/B _4871_/B _4659_/B _5089_/B2 VGND VGND VPWR VPWR _5089_/X sky130_fd_sc_hd__o22a_1
XFILLER_44_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_70 _6088_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_81 _3629_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmax_length3055 _5852_/A2 VGND VGND VPWR VPWR _5761_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_153_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_92 _5955_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length3099 _5664_/X VGND VGND VPWR VPWR _5821_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_153_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length2376 hold697/X VGND VGND VPWR VPWR _4039_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_180_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length4290 _4605_/A VGND VGND VPWR VPWR _4342_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_156_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4460_ _4460_/A _4514_/B VGND VGND VPWR VPWR _4860_/A sky130_fd_sc_hd__nand2_2
Xhold307 _6924_/Q VGND VGND VPWR VPWR hold307/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold318 _6874_/Q VGND VGND VPWR VPWR hold318/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold329 _6520_/Q VGND VGND VPWR VPWR hold329/X sky130_fd_sc_hd__dlygate4sd3_1
X_3411_ wire374/X _6788_/Q _3791_/A VGND VGND VPWR VPWR _3411_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_558 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4391_ _4390_/C _4390_/D _4467_/A _4389_/Y VGND VGND VPWR VPWR _4391_/Y sky130_fd_sc_hd__a31oi_1
X_6130_ _6130_/A1 _6130_/A2 _6339_/A2 _6130_/B2 _6129_/X VGND VGND VPWR VPWR _6130_/X
+ sky130_fd_sc_hd__a221o_1
X_3342_ _3546_/A _3342_/B VGND VGND VPWR VPWR _3342_/Y sky130_fd_sc_hd__nor2_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _6915_/Q _6061_/A2 _6082_/A2 _6061_/B2 VGND VGND VPWR VPWR _6061_/X sky130_fd_sc_hd__a22o_1
X_3273_ hold68/X _3282_/A VGND VGND VPWR VPWR _3414_/B sky130_fd_sc_hd__and2b_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5012_ _4657_/A _4657_/B _4387_/B _5130_/B VGND VGND VPWR VPWR _5012_/X sky130_fd_sc_hd__a31o_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6963_ _6963_/CLK _6963_/D _6401_/A VGND VGND VPWR VPWR _6963_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_81_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5914_ _6273_/B2 _5943_/A2 _5943_/B1 _5914_/B2 VGND VGND VPWR VPWR _5914_/X sky130_fd_sc_hd__a22o_1
X_6894_ _6989_/CLK _6894_/D wire3995/X VGND VGND VPWR VPWR _6894_/Q sky130_fd_sc_hd__dfrtp_1
X_5845_ _6199_/B2 _5845_/A2 _5845_/B1 _6215_/A1 VGND VGND VPWR VPWR _5845_/X sky130_fd_sc_hd__a22o_1
XFILLER_167_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5776_ _5776_/A1 _5776_/A2 _5776_/B1 _7078_/Q VGND VGND VPWR VPWR _5776_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4727_ _4739_/A _4724_/A _4726_/Y _4727_/B1 VGND VGND VPWR VPWR _4992_/C sky130_fd_sc_hd__o31a_1
XFILLER_107_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4658_ _5021_/A _4784_/B VGND VGND VPWR VPWR _4713_/A sky130_fd_sc_hd__or2_1
XFILLER_190_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput90 spimemio_flash_io2_oeb VGND VGND VPWR VPWR input90/X sky130_fd_sc_hd__clkbuf_1
XFILLER_123_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3609_ _3609_/A1 _3709_/A2 _3609_/B1 _6677_/Q VGND VGND VPWR VPWR _3609_/X sky130_fd_sc_hd__a22o_1
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4589_ _4613_/A _4589_/B VGND VGND VPWR VPWR _4673_/A sky130_fd_sc_hd__or2_2
Xwire3805 _4912_/A1 VGND VGND VPWR VPWR _4696_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_150_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6328_ _6328_/A1 _6328_/A2 _6328_/B1 _6328_/B2 _6327_/X VGND VGND VPWR VPWR _6331_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_1_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3849 _4610_/A VGND VGND VPWR VPWR _4575_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_67_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6259_ _6259_/A1 _6322_/B1 _6321_/B1 _6259_/B2 _6258_/X VGND VGND VPWR VPWR _6267_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_748 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3960_ _6824_/Q _3960_/B VGND VGND VPWR VPWR _3960_/X sky130_fd_sc_hd__and2_1
XFILLER_51_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3891_ _6541_/Q _3890_/A _3890_/Y _6543_/Q VGND VGND VPWR VPWR _6541_/D sky130_fd_sc_hd__a22o_1
XFILLER_149_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5630_ _5650_/B _6014_/A _6040_/A _5610_/X _7154_/Q VGND VGND VPWR VPWR _7154_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_149_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5561_ _5561_/A0 hold125/X _5561_/S VGND VGND VPWR VPWR _7118_/D sky130_fd_sc_hd__mux2_1
XFILLER_163_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4512_ _4516_/A _4512_/B VGND VGND VPWR VPWR _4515_/B sky130_fd_sc_hd__nand2_1
XFILLER_157_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5492_ _5588_/A0 hold656/X _5492_/S VGND VGND VPWR VPWR _7057_/D sky130_fd_sc_hd__mux2_1
XFILLER_156_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold104 _6832_/Q VGND VGND VPWR VPWR hold104/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold115 _3262_/X VGND VGND VPWR VPWR hold115/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 _6958_/Q VGND VGND VPWR VPWR hold126/X sky130_fd_sc_hd__dlygate4sd3_1
X_4443_ _4445_/A _4443_/B VGND VGND VPWR VPWR _5003_/A sky130_fd_sc_hd__or2_1
XFILLER_132_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold137 _7131_/Q VGND VGND VPWR VPWR hold137/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 _6923_/Q VGND VGND VPWR VPWR hold148/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold159 _3243_/Y VGND VGND VPWR VPWR hold159/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4374_ _4745_/A _4532_/B VGND VGND VPWR VPWR _5112_/A sky130_fd_sc_hd__nor2_1
X_7162_ _3937_/A1 _7162_/D wire4007/A VGND VGND VPWR VPWR _7162_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3325_ _3339_/B _3465_/B VGND VGND VPWR VPWR _3325_/Y sky130_fd_sc_hd__nor2_1
X_6113_ _6113_/A1 _6113_/A2 _6113_/B1 _6113_/B2 VGND VGND VPWR VPWR _6113_/X sky130_fd_sc_hd__a22o_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7093_ _7093_/CLK _7093_/D wire3959/A VGND VGND VPWR VPWR _7093_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3256_ _3314_/A VGND VGND VPWR VPWR _3256_/Y sky130_fd_sc_hd__inv_2
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ _6069_/A _6044_/B _6044_/C _6044_/D VGND VGND VPWR VPWR _6045_/C sky130_fd_sc_hd__or4_1
XFILLER_140_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3187_ _4654_/A VGND VGND VPWR VPWR _4546_/A sky130_fd_sc_hd__clkinv_2
XFILLER_27_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6946_ _7135_/CLK _6946_/D wire4052/X VGND VGND VPWR VPWR _6946_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_42_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6877_ _7134_/CLK _6877_/D _7134_/RESET_B VGND VGND VPWR VPWR hold96/A sky130_fd_sc_hd__dfrtp_1
XFILLER_50_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5828_ _6976_/Q _5850_/B VGND VGND VPWR VPWR _5828_/X sky130_fd_sc_hd__or2_1
XFILLER_10_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5759_ _5759_/A1 _5759_/A2 _5759_/B1 _6112_/B2 VGND VGND VPWR VPWR _5759_/X sky130_fd_sc_hd__a22o_1
Xmax_length627 _5472_/S VGND VGND VPWR VPWR _5468_/S sky130_fd_sc_hd__clkbuf_1
XFILLER_185_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold660 _6961_/Q VGND VGND VPWR VPWR hold660/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3613 _5537_/A1 VGND VGND VPWR VPWR _5459_/A0 sky130_fd_sc_hd__clkbuf_1
Xhold671 _7008_/Q VGND VGND VPWR VPWR hold671/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3624 _4295_/A0 VGND VGND VPWR VPWR _5211_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold682 _6558_/Q VGND VGND VPWR VPWR hold682/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3646 _5476_/A0 VGND VGND VPWR VPWR _5359_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2901 _5777_/A2 VGND VGND VPWR VPWR _5742_/B1 sky130_fd_sc_hd__clkbuf_1
Xhold693 _7091_/Q VGND VGND VPWR VPWR hold693/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2912 _5757_/B1 VGND VGND VPWR VPWR _5896_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3668 wire3669/X VGND VGND VPWR VPWR wire3668/X sky130_fd_sc_hd__clkbuf_1
Xwire2923 _5852_/B1 VGND VGND VPWR VPWR _5754_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire3679 _5872_/B VGND VGND VPWR VPWR _5960_/B sky130_fd_sc_hd__clkbuf_1
Xwire2934 _5961_/B2 VGND VGND VPWR VPWR _5895_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_89_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2945 _5950_/B1 VGND VGND VPWR VPWR _5910_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2956 _5949_/B1 VGND VGND VPWR VPWR _5921_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2967 wire2967/A VGND VGND VPWR VPWR wire2967/X sky130_fd_sc_hd__clkbuf_1
Xwire2978 _5714_/B1 VGND VGND VPWR VPWR _5684_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire2989 _5748_/B1 VGND VGND VPWR VPWR _5885_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput209 _3228_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[6] sky130_fd_sc_hd__buf_12
XFILLER_126_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4090_ hold217/X _5351_/A0 _4100_/S VGND VGND VPWR VPWR _4090_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6800_ _6803_/CLK _6800_/D wire3950/A VGND VGND VPWR VPWR _6800_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_91_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4992_ _4875_/X _4992_/B _4992_/C VGND VGND VPWR VPWR _5050_/C sky130_fd_sc_hd__and3b_1
XFILLER_63_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6731_ _6755_/CLK _6731_/D fanout3952/X VGND VGND VPWR VPWR _6731_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_189_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3943_ _3943_/A0 _3943_/A1 _3951_/S VGND VGND VPWR VPWR _3943_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6662_ _6701_/CLK _6662_/D wire3945/X VGND VGND VPWR VPWR _6662_/Q sky130_fd_sc_hd__dfstp_1
X_3874_ _6457_/Q hold5/A _6543_/Q _3834_/B VGND VGND VPWR VPWR _6442_/D sky130_fd_sc_hd__o211a_1
XFILLER_31_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5613_ _6564_/Q _5705_/B VGND VGND VPWR VPWR _5618_/B sky130_fd_sc_hd__nand2_1
X_6593_ _7109_/CLK _6593_/D wire3999/A VGND VGND VPWR VPWR _6593_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_191_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5544_ _5544_/A _5553_/B VGND VGND VPWR VPWR _5544_/Y sky130_fd_sc_hd__nand2_1
XFILLER_191_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5475_ _5475_/A _5475_/B VGND VGND VPWR VPWR _5483_/S sky130_fd_sc_hd__nand2_1
XFILLER_145_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7214_ _7214_/A VGND VGND VPWR VPWR _7214_/X sky130_fd_sc_hd__clkbuf_1
X_4426_ _4462_/B _4426_/B VGND VGND VPWR VPWR _4947_/A sky130_fd_sc_hd__nand2_1
XFILLER_160_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7145_ _7180_/CLK _7145_/D wire3996/X VGND VGND VPWR VPWR _7145_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_59_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2208 _6725_/Q VGND VGND VPWR VPWR _6328_/B2 sky130_fd_sc_hd__clkbuf_2
X_4357_ _4407_/A _4359_/B VGND VGND VPWR VPWR _4360_/A sky130_fd_sc_hd__nor2_1
Xwire2219 _6718_/Q VGND VGND VPWR VPWR _6281_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1507 wire1507/A VGND VGND VPWR VPWR _3403_/B2 sky130_fd_sc_hd__clkbuf_1
X_3308_ _5241_/A _4111_/B VGND VGND VPWR VPWR _3308_/Y sky130_fd_sc_hd__nor2_1
X_7076_ _7076_/CLK _7076_/D wire3981/X VGND VGND VPWR VPWR _7076_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1518 _3307_/Y VGND VGND VPWR VPWR _3511_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4288_ _4288_/A _4300_/B VGND VGND VPWR VPWR _4293_/S sky130_fd_sc_hd__nand2_2
Xwire1529 _7210_/Q VGND VGND VPWR VPWR _6305_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_100_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3239_ _4342_/B VGND VGND VPWR VPWR _4793_/A sky130_fd_sc_hd__inv_2
X_6027_ _6027_/A _6027_/B _6027_/C _6027_/D VGND VGND VPWR VPWR _6029_/D sky130_fd_sc_hd__or4_1
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6929_ _6973_/CLK hold80/X fanout4078/X VGND VGND VPWR VPWR hold79/A sky130_fd_sc_hd__dfrtp_1
XFILLER_168_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_31_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7084_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_168_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire804 _3528_/Y VGND VGND VPWR VPWR wire804/X sky130_fd_sc_hd__dlymetal6s2s_1
Xwire815 _3503_/Y VGND VGND VPWR VPWR _4198_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length402 _4101_/S VGND VGND VPWR VPWR _4097_/S sky130_fd_sc_hd__clkbuf_2
Xwire826 _3474_/Y VGND VGND VPWR VPWR _4264_/A sky130_fd_sc_hd__clkbuf_2
Xwire837 _3451_/Y VGND VGND VPWR VPWR _4174_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xwire848 _3420_/X VGND VGND VPWR VPWR wire848/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_46_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7031_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_136_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout4005 fanout4005/A VGND VGND VPWR VPWR fanout4005/X sky130_fd_sc_hd__buf_6
XFILLER_129_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length468 _5588_/S VGND VGND VPWR VPWR _5583_/S sky130_fd_sc_hd__clkbuf_1
XFILLER_89_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout4027 wire4029/X VGND VGND VPWR VPWR fanout4027/X sky130_fd_sc_hd__buf_6
Xwire4100 input71/X VGND VGND VPWR VPWR wire4100/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout4038 wire4086/A VGND VGND VPWR VPWR wire4042/A sky130_fd_sc_hd__buf_6
XFILLER_108_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4111 input68/X VGND VGND VPWR VPWR _3437_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire4122 wire4123/X VGND VGND VPWR VPWR wire4122/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4133 _3623_/A1 VGND VGND VPWR VPWR wire4133/X sky130_fd_sc_hd__clkbuf_1
Xwire4144 input61/X VGND VGND VPWR VPWR wire4144/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3410 _5551_/A0 VGND VGND VPWR VPWR _5410_/A0 sky130_fd_sc_hd__clkbuf_2
Xwire4155 input58/X VGND VGND VPWR VPWR wire4155/X sky130_fd_sc_hd__clkbuf_1
Xwire4166 wire4167/X VGND VGND VPWR VPWR wire4166/X sky130_fd_sc_hd__clkbuf_1
Xwire4177 input52/X VGND VGND VPWR VPWR _3732_/A1 sky130_fd_sc_hd__clkbuf_1
Xhold490 _6663_/Q VGND VGND VPWR VPWR hold490/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3432 _5541_/A1 VGND VGND VPWR VPWR _5508_/A0 sky130_fd_sc_hd__clkbuf_2
Xwire4188 input49/X VGND VGND VPWR VPWR wire4188/X sky130_fd_sc_hd__clkbuf_1
Xwire3443 hold107/X VGND VGND VPWR VPWR wire3443/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_1_0_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_89_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire4199 wire4200/X VGND VGND VPWR VPWR _3619_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2720 _6187_/B1 VGND VGND VPWR VPWR wire2720/X sky130_fd_sc_hd__clkbuf_1
Xwire3465 wire3466/X VGND VGND VPWR VPWR _5540_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2731 _6256_/A2 VGND VGND VPWR VPWR _6057_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3476 _5381_/A0 VGND VGND VPWR VPWR _5567_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2742 wire2743/X VGND VGND VPWR VPWR _6225_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire3498 _5533_/A1 VGND VGND VPWR VPWR wire3498/X sky130_fd_sc_hd__clkbuf_2
Xwire2753 _6003_/X VGND VGND VPWR VPWR _6027_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2764 _6151_/A2 VGND VGND VPWR VPWR _6049_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2775 _5994_/X VGND VGND VPWR VPWR _6201_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_65_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2786 _6092_/B1 VGND VGND VPWR VPWR _6258_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2797 _6200_/A2 VGND VGND VPWR VPWR _6174_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_92_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3590_ _3590_/A1 _3321_/Y _3496_/Y _6317_/B2 _3561_/X VGND VGND VPWR VPWR _3593_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_186_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length991 wire992/X VGND VGND VPWR VPWR wire990/A sky130_fd_sc_hd__clkbuf_1
X_5260_ _5359_/A0 hold321/X _5263_/S VGND VGND VPWR VPWR _6850_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4211_ hold405/X _4211_/A1 _4215_/S VGND VGND VPWR VPWR _6665_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5191_ _5197_/A0 hold471/X _5192_/S VGND VGND VPWR VPWR _6796_/D sky130_fd_sc_hd__mux2_1
X_4142_ _4259_/A1 _4142_/A1 _4146_/S VGND VGND VPWR VPWR _6606_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4073_ hold248/X _4122_/A0 _4083_/S VGND VGND VPWR VPWR _4073_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4975_ _4971_/A _4797_/A _4607_/D _4974_/Y _4574_/Y VGND VGND VPWR VPWR _5095_/C
+ sky130_fd_sc_hd__a311o_1
XFILLER_189_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6714_ _7208_/CLK _6714_/D _7112_/SET_B VGND VGND VPWR VPWR _6714_/Q sky130_fd_sc_hd__dfrtp_1
Xmax_length4119 input67/X VGND VGND VPWR VPWR wire4118/A sky130_fd_sc_hd__clkbuf_1
X_3926_ _3926_/A0 _3926_/A1 _3928_/S VGND VGND VPWR VPWR _3926_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6645_ _7193_/CLK _6645_/D VGND VGND VPWR VPWR _6645_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3857_ _3858_/B _3857_/B VGND VGND VPWR VPWR _6454_/D sky130_fd_sc_hd__xnor2_1
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length2728 _6027_/C VGND VGND VPWR VPWR _6187_/B1 sky130_fd_sc_hd__clkbuf_2
X_6576_ _7017_/CLK _6576_/D fanout4078/X VGND VGND VPWR VPWR _6576_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_166_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3788_ _3788_/A _3788_/B _3788_/C _3788_/D VGND VGND VPWR VPWR _3789_/D sky130_fd_sc_hd__or4_1
XFILLER_117_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5527_ _5527_/A0 hold221/X _5528_/S VGND VGND VPWR VPWR _7088_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5458_ _5485_/A0 hold601/X _5462_/S VGND VGND VPWR VPWR _7026_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4409_ _4412_/A1 _4538_/B _4408_/Y VGND VGND VPWR VPWR _4433_/C sky130_fd_sc_hd__a21o_1
XFILLER_182_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2005 _3606_/A1 VGND VGND VPWR VPWR _5739_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_132_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5389_ _5389_/A0 hold235/X _5393_/S VGND VGND VPWR VPWR _6965_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2016 _6886_/Q VGND VGND VPWR VPWR _5775_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2027 wire2028/X VGND VGND VPWR VPWR _6183_/B2 sky130_fd_sc_hd__clkbuf_2
X_7128_ _7129_/CLK _7128_/D wire4056/X VGND VGND VPWR VPWR _7128_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_86_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2038 hold93/A VGND VGND VPWR VPWR _6059_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1304 _3268_/Y VGND VGND VPWR VPWR _3647_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2049 wire2050/X VGND VGND VPWR VPWR wire2049/X sky130_fd_sc_hd__clkbuf_1
Xwire1315 _6127_/X VGND VGND VPWR VPWR _6144_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_101_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1326 _5834_/X VGND VGND VPWR VPWR _5835_/D sky130_fd_sc_hd__clkbuf_1
Xwire1337 _5687_/X VGND VGND VPWR VPWR wire1337/X sky130_fd_sc_hd__clkbuf_1
XFILLER_74_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7059_ _7059_/CLK _7059_/D fanout4027/X VGND VGND VPWR VPWR _7059_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_74_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1359 wire1360/X VGND VGND VPWR VPWR wire1359/X sky130_fd_sc_hd__clkbuf_1
XFILLER_74_448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire601 _5519_/S VGND VGND VPWR VPWR _5514_/S sky130_fd_sc_hd__clkbuf_2
Xwire612 _5499_/S VGND VGND VPWR VPWR _5497_/S sky130_fd_sc_hd__dlymetal6s2s_1
Xwire623 _5479_/S VGND VGND VPWR VPWR _5480_/S sky130_fd_sc_hd__dlymetal6s2s_1
Xwire634 wire635/X VGND VGND VPWR VPWR _5461_/S sky130_fd_sc_hd__clkbuf_1
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length3941 _6429_/A VGND VGND VPWR VPWR _6441_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire645 wire646/X VGND VGND VPWR VPWR _5456_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_7_747 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire667 _5411_/S VGND VGND VPWR VPWR _5408_/S sky130_fd_sc_hd__clkbuf_1
Xwire678 _5393_/S VGND VGND VPWR VPWR _5391_/S sky130_fd_sc_hd__clkbuf_2
Xwire689 _5363_/S VGND VGND VPWR VPWR _5366_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_171_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3240 _5071_/A VGND VGND VPWR VPWR _5033_/A sky130_fd_sc_hd__clkbuf_1
Xwire3262 wire3262/A VGND VGND VPWR VPWR _5448_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_123_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3284 _4276_/B VGND VGND VPWR VPWR _5562_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2550 _6203_/A2 VGND VGND VPWR VPWR _6175_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3295 hold141/X VGND VGND VPWR VPWR _3282_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2561 _6314_/A2 VGND VGND VPWR VPWR _6328_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2572 _6320_/B1 VGND VGND VPWR VPWR _6296_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire2583 _5968_/A2 VGND VGND VPWR VPWR _5946_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2594 _4900_/X VGND VGND VPWR VPWR _4901_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_65_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1860 hold89/A VGND VGND VPWR VPWR wire1860/X sky130_fd_sc_hd__clkbuf_1
Xwire1871 _6969_/Q VGND VGND VPWR VPWR _6200_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1882 _6962_/Q VGND VGND VPWR VPWR _3747_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire1893 _6101_/A1 VGND VGND VPWR VPWR _5766_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4760_ _4760_/A1 _5113_/A1 _4734_/B _5135_/A1 _4758_/Y VGND VGND VPWR VPWR _4760_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_159_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3711_ _3711_/A _3711_/B VGND VGND VPWR VPWR _3711_/Y sky130_fd_sc_hd__nor2_1
XFILLER_174_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4691_ _4707_/A _4704_/B VGND VGND VPWR VPWR _4708_/B sky130_fd_sc_hd__or2_1
XFILLER_119_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6430_ _6430_/A _6432_/B VGND VGND VPWR VPWR _6430_/X sky130_fd_sc_hd__and2_1
X_3642_ _3642_/A _3642_/B _3642_/C _3642_/D VGND VGND VPWR VPWR _3660_/B sky130_fd_sc_hd__or4_1
X_6361_ _6358_/A _6389_/A2 _4228_/A VGND VGND VPWR VPWR _6362_/B sky130_fd_sc_hd__a21boi_1
XFILLER_174_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3573_ _3573_/A _3573_/B _3573_/C _3573_/D VGND VGND VPWR VPWR _3583_/C sky130_fd_sc_hd__or4_1
XFILLER_127_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5312_ _5339_/A0 hold581/X _5312_/S VGND VGND VPWR VPWR _6897_/D sky130_fd_sc_hd__mux2_1
X_6292_ _6292_/A _6292_/B _6292_/C VGND VGND VPWR VPWR _6292_/X sky130_fd_sc_hd__or3_1
XFILLER_114_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5243_ _5351_/A0 hold217/X _5248_/S VGND VGND VPWR VPWR _6835_/D sky130_fd_sc_hd__mux2_1
XFILLER_69_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold19 hold19/A VGND VGND VPWR VPWR hold19/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5174_ _5174_/A _5174_/B _5174_/C _5173_/X VGND VGND VPWR VPWR _5174_/X sky130_fd_sc_hd__or4b_1
XFILLER_68_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4125_ _5309_/A0 hold609/X _4125_/S VGND VGND VPWR VPWR _6592_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4056_ hold102/X _4113_/A0 _4060_/S VGND VGND VPWR VPWR _4056_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4958_ _4958_/A1 _4526_/B _4958_/B1 _5108_/A _4957_/Y VGND VGND VPWR VPWR _5163_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_184_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3909_ _5650_/A _3908_/B _3906_/X _5590_/A2 _6562_/Q VGND VGND VPWR VPWR _6564_/D
+ sky130_fd_sc_hd__a32o_1
Xmax_length3215 _5035_/B VGND VGND VPWR VPWR _4717_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_177_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4889_ _4486_/A _5003_/A _4872_/B VGND VGND VPWR VPWR _4890_/D sky130_fd_sc_hd__a21oi_1
XFILLER_137_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length3248 _5210_/B VGND VGND VPWR VPWR _5193_/B sky130_fd_sc_hd__clkbuf_2
X_6628_ _7193_/CLK _6628_/D VGND VGND VPWR VPWR _6628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6559_ _7109_/CLK _6559_/D wire3999/X VGND VGND VPWR VPWR _6559_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1101 _5221_/B VGND VGND VPWR VPWR _3501_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1112 _3341_/Y VGND VGND VPWR VPWR _3384_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_101_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1134 _3550_/B1 VGND VGND VPWR VPWR _5475_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_47_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1156 _3736_/B1 VGND VGND VPWR VPWR _5448_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1167 _3548_/B1 VGND VGND VPWR VPWR _3436_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_74_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1178 _3700_/A2 VGND VGND VPWR VPWR _3443_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire1189 _3684_/A2 VGND VGND VPWR VPWR wire1189/X sky130_fd_sc_hd__clkbuf_1
XFILLER_62_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire420 _3751_/X VGND VGND VPWR VPWR wire420/X sky130_fd_sc_hd__clkbuf_1
XFILLER_168_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire431 _3570_/X VGND VGND VPWR VPWR _3573_/C sky130_fd_sc_hd__clkbuf_1
Xwire442 _6342_/X VGND VGND VPWR VPWR wire442/X sky130_fd_sc_hd__clkbuf_1
Xwire453 _6095_/X VGND VGND VPWR VPWR wire453/X sky130_fd_sc_hd__clkbuf_1
Xwire464 _5751_/X VGND VGND VPWR VPWR wire464/X sky130_fd_sc_hd__clkbuf_1
XFILLER_156_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire475 wire476/X VGND VGND VPWR VPWR wire475/X sky130_fd_sc_hd__clkbuf_1
XFILLER_156_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire497 wire498/X VGND VGND VPWR VPWR wire497/X sky130_fd_sc_hd__clkbuf_1
XFILLER_171_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3070 _5959_/A2 VGND VGND VPWR VPWR _5927_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire3081 _5915_/A2 VGND VGND VPWR VPWR _5962_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3092 wire3092/A VGND VGND VPWR VPWR _5799_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2380 _6527_/Q VGND VGND VPWR VPWR _3686_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_66_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2391 _6518_/Q VGND VGND VPWR VPWR _6288_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1690 _6063_/B2 VGND VGND VPWR VPWR _3668_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_19_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5930_ _6302_/B2 _5930_/A2 _5930_/B1 _6306_/B2 _5929_/X VGND VGND VPWR VPWR _5935_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_53_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5861_ _6230_/A1 _5953_/B1 _5965_/A2 _6224_/B2 VGND VGND VPWR VPWR _5861_/X sky130_fd_sc_hd__a22o_1
X_4812_ _4984_/C _5090_/A _4805_/X _4811_/X VGND VGND VPWR VPWR _4813_/D sky130_fd_sc_hd__or4bb_1
XFILLER_34_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5792_ _5792_/A _5792_/B _5792_/C VGND VGND VPWR VPWR _5792_/X sky130_fd_sc_hd__or3_1
XFILLER_33_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4743_ _4753_/A _4743_/B VGND VGND VPWR VPWR _4764_/A sky130_fd_sc_hd__nor2_1
XFILLER_147_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4674_ _4674_/A _4684_/A VGND VGND VPWR VPWR _4692_/B sky130_fd_sc_hd__nand2_1
XFILLER_147_578 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6413_ _6432_/A _6428_/B VGND VGND VPWR VPWR _6413_/X sky130_fd_sc_hd__and2_1
X_3625_ _6086_/A1 _3625_/A2 _3625_/B1 _3625_/B2 wire774/X VGND VGND VPWR VPWR _3627_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_135_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6344_ _7187_/Q _6319_/S wire441/X _6343_/X VGND VGND VPWR VPWR _7187_/D sky130_fd_sc_hd__o22a_1
XFILLER_115_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3556_ _3556_/A1 _3770_/A2 _4312_/A _6759_/Q VGND VGND VPWR VPWR _3556_/X sky130_fd_sc_hd__a22o_1
XFILLER_1_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6275_ _6523_/Q _6324_/A2 _6324_/B1 _6763_/Q _6274_/X VGND VGND VPWR VPWR _6275_/X
+ sky130_fd_sc_hd__a221o_1
X_3487_ _3487_/A1 _3654_/B1 wire886/X _3487_/B2 _3486_/X VGND VGND VPWR VPWR _3499_/A
+ sky130_fd_sc_hd__a221o_2
Xinput109 wb_adr_i[19] VGND VGND VPWR VPWR _4337_/C sky130_fd_sc_hd__clkbuf_1
X_5226_ hold546/X _5523_/A0 _5228_/S VGND VGND VPWR VPWR _6821_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5157_ _5110_/C _5153_/X _5178_/C _5156_/Y VGND VGND VPWR VPWR _5157_/X sky130_fd_sc_hd__o31a_1
XFILLER_29_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4108_ _4139_/A1 hold622/X _4108_/S VGND VGND VPWR VPWR _6577_/D sky130_fd_sc_hd__mux2_1
X_5088_ _5088_/A1 _5071_/A _5070_/Y _5087_/X VGND VGND VPWR VPWR _5104_/C sky130_fd_sc_hd__a22o_1
XFILLER_84_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4039_ _4039_/A0 _4134_/A1 _4039_/S VGND VGND VPWR VPWR _6530_/D sky130_fd_sc_hd__mux2_1
XFILLER_44_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_60 _3590_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_71 _5692_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_82 _4199_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_93 _5715_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmax_length2333 hold237/X VGND VGND VPWR VPWR _4142_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_138_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3089 _5666_/X VGND VGND VPWR VPWR wire3088/A sky130_fd_sc_hd__clkbuf_1
XFILLER_21_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length2399 _6514_/Q VGND VGND VPWR VPWR _3587_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_134_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold308 _6673_/Q VGND VGND VPWR VPWR hold308/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold319 _6946_/Q VGND VGND VPWR VPWR hold319/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3410_ _3410_/A _3410_/B VGND VGND VPWR VPWR _3410_/X sky130_fd_sc_hd__or2_1
X_4390_ _4390_/A _4654_/A _4390_/C _4390_/D VGND VGND VPWR VPWR _4390_/X sky130_fd_sc_hd__or4_1
XFILLER_98_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3341_ _3507_/B _3342_/B VGND VGND VPWR VPWR _3341_/Y sky130_fd_sc_hd__nor2_1
XFILLER_98_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6060_ _7112_/Q _6060_/A2 _6060_/B1 _6060_/B2 _6059_/X VGND VGND VPWR VPWR _6069_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ hold83/X _3288_/A VGND VGND VPWR VPWR _3293_/A sky130_fd_sc_hd__and2b_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _4873_/Y _5130_/B _5010_/X _5050_/C VGND VGND VPWR VPWR _5033_/B sky130_fd_sc_hd__o31a_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6962_ _7083_/CLK _6962_/D wire4037/X VGND VGND VPWR VPWR _6962_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_19_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5913_ _5913_/A _5913_/B _5913_/C _5913_/D VGND VGND VPWR VPWR _5913_/X sky130_fd_sc_hd__or4_1
XFILLER_179_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6893_ _7110_/CLK _6893_/D wire4004/X VGND VGND VPWR VPWR _6893_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5844_ _5844_/A1 _5844_/A2 _5843_/X VGND VGND VPWR VPWR _5847_/C sky130_fd_sc_hd__a21o_1
XFILLER_61_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5775_ _5775_/A1 _5775_/A2 _5775_/B1 _5775_/B2 VGND VGND VPWR VPWR _5775_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4726_ _5001_/C VGND VGND VPWR VPWR _4726_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4657_ _4657_/A _4657_/B _4657_/C VGND VGND VPWR VPWR _5130_/A sky130_fd_sc_hd__and3_1
XFILLER_175_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput80 spi_sck VGND VGND VPWR VPWR input80/X sky130_fd_sc_hd__clkbuf_1
X_3608_ _6083_/B2 wire965/X wire889/X _7121_/Q VGND VGND VPWR VPWR _3608_/X sky130_fd_sc_hd__a22o_1
XFILLER_135_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput91 spimemio_flash_io3_do VGND VGND VPWR VPWR input91/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4588_ _4588_/A _4588_/B _4621_/B _4935_/A VGND VGND VPWR VPWR _4589_/B sky130_fd_sc_hd__or4bb_2
XFILLER_89_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3806 _4666_/B VGND VGND VPWR VPWR _4912_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
X_6327_ _6327_/A1 _6327_/A2 _6327_/B1 _6327_/B2 VGND VGND VPWR VPWR _6327_/X sky130_fd_sc_hd__a22o_1
X_3539_ _5786_/B2 wire878/A _3539_/B1 _3539_/B2 VGND VGND VPWR VPWR _3539_/X sky130_fd_sc_hd__a22o_1
Xwire3817 _4814_/A VGND VGND VPWR VPWR _4693_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3828 _4781_/A VGND VGND VPWR VPWR _4359_/B sky130_fd_sc_hd__buf_2
XFILLER_89_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3839 wire3840/X VGND VGND VPWR VPWR _3934_/S sky130_fd_sc_hd__clkbuf_1
XFILLER_88_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6258_ _6258_/A1 _6258_/A2 _6258_/B1 _6258_/B2 _6246_/X VGND VGND VPWR VPWR _6258_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5209_ hold683/X _5216_/A0 _5209_/S VGND VGND VPWR VPWR _6810_/D sky130_fd_sc_hd__mux2_1
XFILLER_57_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6189_ _6189_/A1 _5977_/X _6189_/B1 _7117_/Q _6188_/X VGND VGND VPWR VPWR _6192_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_29_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3890_ _3890_/A _3890_/B VGND VGND VPWR VPWR _3890_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5560_ _5587_/A0 hold690/X _5560_/S VGND VGND VPWR VPWR _7117_/D sky130_fd_sc_hd__mux2_1
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4511_ _4871_/A _4743_/B _4508_/X _4510_/X VGND VGND VPWR VPWR _4515_/A sky130_fd_sc_hd__o211a_1
XFILLER_129_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5491_ _5491_/A0 hold595/X _5491_/S VGND VGND VPWR VPWR _7056_/D sky130_fd_sc_hd__mux2_1
XFILLER_8_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold105 _6840_/Q VGND VGND VPWR VPWR hold105/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold116 _3284_/A VGND VGND VPWR VPWR _3288_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4442_ _4445_/A _4443_/B VGND VGND VPWR VPWR _4512_/B sky130_fd_sc_hd__nor2_1
Xhold127 _6739_/Q VGND VGND VPWR VPWR hold127/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 _6908_/Q VGND VGND VPWR VPWR hold138/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 _7089_/Q VGND VGND VPWR VPWR hold149/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7161_ _7180_/CLK _7161_/D _7161_/RESET_B VGND VGND VPWR VPWR _7161_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_144_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4373_ _4570_/C _4781_/B VGND VGND VPWR VPWR _4532_/B sky130_fd_sc_hd__or2_1
XFILLER_98_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6112_ _6112_/A1 _6198_/A2 _6112_/B1 _6112_/B2 _6111_/X VGND VGND VPWR VPWR _6119_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3324_ _3324_/A _3465_/B VGND VGND VPWR VPWR _3324_/Y sky130_fd_sc_hd__nor2_1
X_7092_ _7092_/CLK _7092_/D fanout3944/X VGND VGND VPWR VPWR _7092_/Q sky130_fd_sc_hd__dfstp_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ _6954_/Q _6056_/A2 _6037_/X _6042_/X VGND VGND VPWR VPWR _6044_/D sky130_fd_sc_hd__a211o_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ _3301_/C hold62/X hold26/X VGND VGND VPWR VPWR _3255_/X sky130_fd_sc_hd__or3b_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3186_ _6445_/Q VGND VGND VPWR VPWR _3868_/A sky130_fd_sc_hd__inv_2
XFILLER_54_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6945_ _6945_/CLK _6945_/D fanout4078/X VGND VGND VPWR VPWR _6945_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_81_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
X_6876_ _7129_/CLK _6876_/D wire4056/A VGND VGND VPWR VPWR _6876_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5827_ _6191_/B2 _5827_/A2 _5827_/B1 _6181_/B2 _5826_/X VGND VGND VPWR VPWR _5835_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_139_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5758_ _5758_/A1 _5758_/A2 _5756_/X _5757_/X VGND VGND VPWR VPWR _5771_/A sky130_fd_sc_hd__a211o_1
X_4709_ _4709_/A1 _4677_/B _5054_/B _4708_/X VGND VGND VPWR VPWR _4709_/X sky130_fd_sc_hd__o211a_1
X_5689_ _5705_/B _5703_/B VGND VGND VPWR VPWR _5691_/B sky130_fd_sc_hd__and2_1
XFILLER_135_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire4304 _4846_/A VGND VGND VPWR VPWR _4396_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_135_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold650 _7142_/Q VGND VGND VPWR VPWR hold650/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3614 _4266_/A1 VGND VGND VPWR VPWR _5537_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold661 _6919_/Q VGND VGND VPWR VPWR hold661/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold672 _6905_/Q VGND VGND VPWR VPWR hold672/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3625 _6393_/A0 VGND VGND VPWR VPWR _4295_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold683 _6810_/Q VGND VGND VPWR VPWR hold683/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 _6557_/Q VGND VGND VPWR VPWR hold694/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3636 _5485_/A0 VGND VGND VPWR VPWR _5206_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire3647 _5476_/A0 VGND VGND VPWR VPWR _5581_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2902 _5827_/B1 VGND VGND VPWR VPWR _5777_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_131_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3658 _5350_/A0 VGND VGND VPWR VPWR _5242_/A0 sky130_fd_sc_hd__clkbuf_2
Xwire2913 _5776_/B1 VGND VGND VPWR VPWR _5715_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_131_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2924 _5852_/B1 VGND VGND VPWR VPWR _5817_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3669 _3953_/X VGND VGND VPWR VPWR wire3669/X sky130_fd_sc_hd__clkbuf_1
Xwire2935 _5917_/B1 VGND VGND VPWR VPWR _5961_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2957 _5821_/B1 VGND VGND VPWR VPWR _5949_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2968 wire2968/A VGND VGND VPWR VPWR _5736_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire2979 _5737_/A2 VGND VGND VPWR VPWR _5714_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_182_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length1270 _3605_/A2 VGND VGND VPWR VPWR _3421_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_141_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4991_ _5103_/A _4991_/B VGND VGND VPWR VPWR _4991_/Y sky130_fd_sc_hd__nor2_1
XFILLER_91_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6730_ _7059_/CLK _6730_/D wire4042/A VGND VGND VPWR VPWR _6730_/Q sky130_fd_sc_hd__dfstp_1
X_3942_ _3963_/B _3942_/A2 _6440_/B _3941_/Y VGND VGND VPWR VPWR _3942_/X sky130_fd_sc_hd__a22o_2
XFILLER_149_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6661_ _6701_/CLK _6661_/D wire3945/X VGND VGND VPWR VPWR _6661_/Q sky130_fd_sc_hd__dfrtp_1
X_3873_ _6429_/A _6431_/B VGND VGND VPWR VPWR _3873_/X sky130_fd_sc_hd__and2_1
XFILLER_32_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5612_ _7149_/Q _7148_/Q VGND VGND VPWR VPWR _5705_/B sky130_fd_sc_hd__nor2_4
X_6592_ _7072_/CLK _6592_/D wire4001/X VGND VGND VPWR VPWR _6592_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_191_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5543_ hold591/X _5543_/A1 _5543_/S VGND VGND VPWR VPWR _7102_/D sky130_fd_sc_hd__mux2_1
X_5474_ hold668/X _5519_/A0 _5474_/S VGND VGND VPWR VPWR _7041_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7213_ _7213_/A VGND VGND VPWR VPWR _7213_/X sky130_fd_sc_hd__clkbuf_2
X_4425_ _4524_/A _4425_/B VGND VGND VPWR VPWR _4425_/Y sky130_fd_sc_hd__nand2_1
XFILLER_132_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7144_ _7187_/CLK _7144_/D _7161_/RESET_B VGND VGND VPWR VPWR _7144_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_99_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4356_ _4354_/A _4354_/B _4355_/Y _4350_/B VGND VGND VPWR VPWR _4944_/A sky130_fd_sc_hd__o2bb2ai_2
XFILLER_98_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2209 wire2210/X VGND VGND VPWR VPWR _6306_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3307_ _3414_/B _3378_/B VGND VGND VPWR VPWR _3307_/Y sky130_fd_sc_hd__nand2_1
XFILLER_140_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7075_ _7075_/CLK _7075_/D _7075_/SET_B VGND VGND VPWR VPWR _7075_/Q sky130_fd_sc_hd__dfstp_1
X_4287_ _4311_/A0 hold376/X _4287_/S VGND VGND VPWR VPWR _6735_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6026_ _6026_/A _6026_/B _6026_/C _6026_/D VGND VGND VPWR VPWR _6029_/C sky130_fd_sc_hd__or4_1
X_3238_ _4376_/A VGND VGND VPWR VPWR _4533_/A sky130_fd_sc_hd__inv_2
XFILLER_27_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6928_ _7017_/CLK _6928_/D wire4081/X VGND VGND VPWR VPWR hold99/A sky130_fd_sc_hd__dfrtp_1
XFILLER_167_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6859_ _7127_/CLK _6859_/D _6407_/A VGND VGND VPWR VPWR _6859_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_168_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire805 wire806/X VGND VGND VPWR VPWR wire805/X sky130_fd_sc_hd__clkbuf_1
Xwire816 _3502_/Y VGND VGND VPWR VPWR _4153_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire849 wire849/A VGND VGND VPWR VPWR wire849/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout4017 input75/X VGND VGND VPWR VPWR wire4018/A sky130_fd_sc_hd__buf_6
Xfanout4028 wire4092/A VGND VGND VPWR VPWR fanout4028/X sky130_fd_sc_hd__buf_6
XFILLER_108_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4101 wire4102/X VGND VGND VPWR VPWR _3960_/B sky130_fd_sc_hd__clkbuf_1
Xwire4112 input67/X VGND VGND VPWR VPWR _3928_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_108_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire4123 wire4123/A VGND VGND VPWR VPWR wire4123/X sky130_fd_sc_hd__clkbuf_1
Xwire4134 wire4135/X VGND VGND VPWR VPWR _3623_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4145 input60/X VGND VGND VPWR VPWR _3352_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3400 _5392_/A0 VGND VGND VPWR VPWR _5464_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3411 wire3412/X VGND VGND VPWR VPWR _5551_/A0 sky130_fd_sc_hd__clkbuf_2
Xwire4156 wire4157/X VGND VGND VPWR VPWR _3967_/A0 sky130_fd_sc_hd__clkbuf_1
Xwire3422 _5490_/A0 VGND VGND VPWR VPWR _5481_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire4167 wire4168/X VGND VGND VPWR VPWR wire4167/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold480 _6795_/Q VGND VGND VPWR VPWR hold480/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3433 _5568_/A0 VGND VGND VPWR VPWR _5541_/A1 sky130_fd_sc_hd__clkbuf_2
Xhold491 _7039_/Q VGND VGND VPWR VPWR hold491/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire4178 wire4179/X VGND VGND VPWR VPWR _3358_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire4189 wire4190/X VGND VGND VPWR VPWR _3461_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2710 _6087_/B1 VGND VGND VPWR VPWR _6255_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire3466 wire3466/A VGND VGND VPWR VPWR wire3466/X sky130_fd_sc_hd__clkbuf_1
Xwire2721 _6210_/A2 VGND VGND VPWR VPWR _6115_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2732 _6086_/A2 VGND VGND VPWR VPWR _6256_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire3477 _5381_/A0 VGND VGND VPWR VPWR _5246_/A0 sky130_fd_sc_hd__clkbuf_1
Xwire2743 _6023_/C VGND VGND VPWR VPWR wire2743/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3499 _5533_/A1 VGND VGND VPWR VPWR _4322_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_77_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2754 _6114_/A2 VGND VGND VPWR VPWR _6074_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire2765 wire2765/A VGND VGND VPWR VPWR _6151_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire2776 _6327_/A2 VGND VGND VPWR VPWR _6247_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire2787 _6208_/B1 VGND VGND VPWR VPWR _6157_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire2798 wire2799/X VGND VGND VPWR VPWR _6200_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_18_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_3_0_mgmt_gpio_in[4] clkbuf_2_3_0_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR _3927_/A1
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_146_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4210_ _4210_/A _4240_/B VGND VGND VPWR VPWR _4215_/S sky130_fd_sc_hd__and2_2
X_5190_ _5196_/A0 hold480/X _5192_/S VGND VGND VPWR VPWR _6795_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4141_ _4141_/A _5223_/B VGND VGND VPWR VPWR _4146_/S sky130_fd_sc_hd__nand2_2
XFILLER_110_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4072_ hold483/X _4071_/X _4084_/S VGND VGND VPWR VPWR _6554_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4974_ _4981_/B _5021_/B _4560_/Y _4981_/A VGND VGND VPWR VPWR _4974_/Y sky130_fd_sc_hd__a211oi_1
X_3925_ _6577_/Q _3925_/A1 _3958_/B VGND VGND VPWR VPWR _3925_/X sky130_fd_sc_hd__mux2_1
X_6713_ _7112_/CLK hold71/X _7112_/SET_B VGND VGND VPWR VPWR _6713_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_149_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6644_ _7193_/CLK _6644_/D VGND VGND VPWR VPWR _6644_/Q sky130_fd_sc_hd__dfxtp_1
Xmax_length3419 _5586_/A0 VGND VGND VPWR VPWR _5526_/A0 sky130_fd_sc_hd__clkbuf_1
X_3856_ _6454_/Q _3856_/B VGND VGND VPWR VPWR _3857_/B sky130_fd_sc_hd__nor2_1
XFILLER_165_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6575_ _6701_/CLK _6575_/D wire3945/X VGND VGND VPWR VPWR _6575_/Q sky130_fd_sc_hd__dfrtp_1
X_3787_ _3787_/A1 _3315_/Y _3727_/Y _6812_/Q _3734_/X VGND VGND VPWR VPWR _3788_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5526_ _5526_/A0 hold624/X _5528_/S VGND VGND VPWR VPWR _7087_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5457_ _5457_/A _5511_/B VGND VGND VPWR VPWR _5465_/S sky130_fd_sc_hd__nand2_1
XFILLER_160_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4408_ _4407_/A _4538_/B _4591_/A VGND VGND VPWR VPWR _4408_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_182_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5388_ _5406_/A0 hold91/X _5388_/S VGND VGND VPWR VPWR _6964_/D sky130_fd_sc_hd__mux2_1
Xwire2006 _6077_/B2 VGND VGND VPWR VPWR _3606_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2017 _5756_/A1 VGND VGND VPWR VPWR _3229_/A sky130_fd_sc_hd__clkbuf_1
X_7127_ _7127_/CLK _7127_/D wire4056/X VGND VGND VPWR VPWR _7127_/Q sky130_fd_sc_hd__dfstp_1
Xwire2028 _3381_/B2 VGND VGND VPWR VPWR wire2028/X sky130_fd_sc_hd__clkbuf_1
X_4339_ _4339_/A _4339_/B _4339_/C _4339_/D VGND VGND VPWR VPWR _4348_/C sky130_fd_sc_hd__and4_1
XFILLER_101_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2039 _6874_/Q VGND VGND VPWR VPWR _5986_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1305 _6339_/X VGND VGND VPWR VPWR _6340_/C1 sky130_fd_sc_hd__clkbuf_1
Xwire1316 wire1317/X VGND VGND VPWR VPWR _6012_/B sky130_fd_sc_hd__clkbuf_1
Xwire1327 wire1328/X VGND VGND VPWR VPWR _5835_/C sky130_fd_sc_hd__clkbuf_1
Xwire1338 _5592_/Y VGND VGND VPWR VPWR _6343_/A2 sky130_fd_sc_hd__clkbuf_2
X_7058_ _7083_/CLK _7058_/D wire4037/X VGND VGND VPWR VPWR _7058_/Q sky130_fd_sc_hd__dfstp_1
Xwire1349 _4425_/Y VGND VGND VPWR VPWR _4504_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6009_ _6040_/B _6039_/C _6030_/C VGND VGND VPWR VPWR _6009_/X sky130_fd_sc_hd__and3_1
XFILLER_55_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire602 _5507_/S VGND VGND VPWR VPWR _5503_/S sky130_fd_sc_hd__clkbuf_1
XFILLER_183_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire613 wire613/A VGND VGND VPWR VPWR _5499_/S sky130_fd_sc_hd__clkbuf_1
Xwire624 _5482_/S VGND VGND VPWR VPWR _5479_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_10_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire635 _5463_/S VGND VGND VPWR VPWR wire635/X sky130_fd_sc_hd__clkbuf_1
Xwire646 _5448_/Y VGND VGND VPWR VPWR wire646/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire657 _5438_/S VGND VGND VPWR VPWR _5434_/S sky130_fd_sc_hd__clkbuf_2
Xmax_length3975 fanout3973/X VGND VGND VPWR VPWR wire3974/A sky130_fd_sc_hd__buf_4
Xwire668 _5411_/S VGND VGND VPWR VPWR _5410_/S sky130_fd_sc_hd__clkbuf_1
XFILLER_108_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire679 wire679/A VGND VGND VPWR VPWR _5379_/S sky130_fd_sc_hd__clkbuf_1
Xmax_length3997 fanout3993/X VGND VGND VPWR VPWR wire3996/A sky130_fd_sc_hd__clkbuf_2
XFILLER_124_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3230 _4759_/A VGND VGND VPWR VPWR _4488_/A sky130_fd_sc_hd__clkbuf_2
Xwire3241 _5182_/A2 VGND VGND VPWR VPWR _5071_/A sky130_fd_sc_hd__clkbuf_2
Xwire3252 _4135_/B VGND VGND VPWR VPWR _5529_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_49_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3274 _5225_/B VGND VGND VPWR VPWR _5553_/B sky130_fd_sc_hd__buf_2
Xwire3285 hold57/X VGND VGND VPWR VPWR _4276_/B sky130_fd_sc_hd__clkbuf_2
Xwire2540 _6201_/B1 VGND VGND VPWR VPWR _6127_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire3296 wire3297/X VGND VGND VPWR VPWR _3934_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2551 wire2552/X VGND VGND VPWR VPWR _6203_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire2562 wire2563/X VGND VGND VPWR VPWR _6314_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire2573 wire2574/X VGND VGND VPWR VPWR _6320_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire2584 _5709_/A2 VGND VGND VPWR VPWR _5968_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire2595 _4731_/X VGND VGND VPWR VPWR _4741_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1850 wire1851/X VGND VGND VPWR VPWR wire1850/X sky130_fd_sc_hd__clkbuf_1
Xwire1861 _6977_/Q VGND VGND VPWR VPWR _6206_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1872 wire1873/X VGND VGND VPWR VPWR _5823_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire1883 _6961_/Q VGND VGND VPWR VPWR _6205_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1894 _6949_/Q VGND VGND VPWR VPWR _6101_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_45_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3710_ _3710_/A _3710_/B _3710_/C _3710_/D VGND VGND VPWR VPWR _3722_/C sky130_fd_sc_hd__or4_1
XFILLER_41_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4690_ _4707_/A _4692_/B VGND VGND VPWR VPWR _4708_/A sky130_fd_sc_hd__or2_1
X_3641_ _3641_/A1 _3641_/A2 _4040_/A _6533_/Q _3640_/X VGND VGND VPWR VPWR _3642_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6360_ _6358_/A _6360_/A2 wire3754/X VGND VGND VPWR VPWR _6360_/X sky130_fd_sc_hd__a21bo_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3572_ _3572_/A1 _3312_/Y wire813/X _3572_/B2 _3571_/X VGND VGND VPWR VPWR _3572_/X
+ sky130_fd_sc_hd__a221o_1
X_5311_ _5509_/A0 hold488/X _5311_/S VGND VGND VPWR VPWR _6896_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6291_ _6291_/A _6291_/B _6291_/C _6291_/D VGND VGND VPWR VPWR _6291_/X sky130_fd_sc_hd__or4_1
XFILLER_142_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5242_ _5242_/A0 hold330/X _5248_/S VGND VGND VPWR VPWR _6834_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_30_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7139_/CLK sky130_fd_sc_hd__clkbuf_16
Xfanout3691 _3195_/Y VGND VGND VPWR VPWR _3907_/A sky130_fd_sc_hd__buf_6
X_5173_ _4753_/A _5003_/A _5003_/B _4996_/A _4510_/C VGND VGND VPWR VPWR _5173_/X
+ sky130_fd_sc_hd__o221a_1
X_4124_ _5416_/A0 hold590/X _4125_/S VGND VGND VPWR VPWR _6591_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput1 debug_mode VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__clkbuf_1
X_4055_ hold417/X _4054_/X _4061_/S VGND VGND VPWR VPWR _6546_/D sky130_fd_sc_hd__mux2_1
XFILLER_49_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_45_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7079_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_36_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4957_ _4957_/A _4957_/B VGND VGND VPWR VPWR _4957_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3908_ _5593_/B _3908_/B VGND VGND VPWR VPWR _3908_/Y sky130_fd_sc_hd__nand2_1
XFILLER_165_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4888_ _4460_/A _4871_/Y _4984_/B _5065_/A VGND VGND VPWR VPWR _4890_/C sky130_fd_sc_hd__a211o_1
XFILLER_138_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length3238 _4232_/X VGND VGND VPWR VPWR _6391_/A3 sky130_fd_sc_hd__clkbuf_1
Xmax_length2504 _6025_/B VGND VGND VPWR VPWR _6181_/A2 sky130_fd_sc_hd__clkbuf_2
X_3839_ _6471_/Q _3839_/B VGND VGND VPWR VPWR _3840_/S sky130_fd_sc_hd__nor2_1
X_6627_ _7196_/CLK _6627_/D VGND VGND VPWR VPWR _6627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6558_ _7072_/CLK _6558_/D wire4001/X VGND VGND VPWR VPWR _6558_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_152_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5509_ _5509_/A0 hold542/X _5509_/S VGND VGND VPWR VPWR _7072_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6489_ _7027_/CLK _6489_/D fanout3976/X VGND VGND VPWR VPWR _6489_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1102 _5221_/B VGND VGND VPWR VPWR _5214_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_87_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1113 _3699_/A2 VGND VGND VPWR VPWR _5403_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_75_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1124 _3564_/A2 VGND VGND VPWR VPWR _5331_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_75_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1135 _3498_/A2 VGND VGND VPWR VPWR _3550_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_101_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1146 wire1146/A VGND VGND VPWR VPWR _3684_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire1157 _3327_/Y VGND VGND VPWR VPWR _3736_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1168 wire1168/A VGND VGND VPWR VPWR _3548_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_75_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1179 _3537_/A2 VGND VGND VPWR VPWR _3700_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_142_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire410 _4086_/S VGND VGND VPWR VPWR _4082_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire421 _3696_/X VGND VGND VPWR VPWR _3701_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_156_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire432 wire433/X VGND VGND VPWR VPWR wire432/X sky130_fd_sc_hd__clkbuf_1
XFILLER_156_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire443 _6317_/X VGND VGND VPWR VPWR wire443/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire454 wire455/X VGND VGND VPWR VPWR wire454/X sky130_fd_sc_hd__clkbuf_1
Xwire465 _5581_/S VGND VGND VPWR VPWR _5582_/S sky130_fd_sc_hd__clkbuf_1
XFILLER_171_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length3772 _5859_/A1 VGND VGND VPWR VPWR _6194_/C1 sky130_fd_sc_hd__clkbuf_1
Xwire476 _5553_/Y VGND VGND VPWR VPWR wire476/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire498 wire499/X VGND VGND VPWR VPWR wire498/X sky130_fd_sc_hd__clkbuf_1
XFILLER_124_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3060 _5670_/X VGND VGND VPWR VPWR wire3060/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire3071 _5878_/A2 VGND VGND VPWR VPWR _5959_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire3082 wire3083/X VGND VGND VPWR VPWR _5915_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_66_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3093 _5759_/A2 VGND VGND VPWR VPWR _5956_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2370 _6532_/Q VGND VGND VPWR VPWR wire2370/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2381 wire2382/X VGND VGND VPWR VPWR _6262_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire2392 _6517_/Q VGND VGND VPWR VPWR _3687_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_19_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1680 _7046_/Q VGND VGND VPWR VPWR wire1680/X sky130_fd_sc_hd__clkbuf_1
Xwire1691 hold94/A VGND VGND VPWR VPWR _6063_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5860_ _5860_/A0 wire399/X _5860_/S VGND VGND VPWR VPWR _7169_/D sky130_fd_sc_hd__mux2_1
X_4811_ _4712_/B _4673_/A _4759_/Y _4786_/Y _4810_/X VGND VGND VPWR VPWR _4811_/X
+ sky130_fd_sc_hd__o2111a_1
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5791_ _6140_/B2 _5791_/A2 _5791_/B1 _6127_/B2 _5790_/X VGND VGND VPWR VPWR _5792_/C
+ sky130_fd_sc_hd__a221o_1
X_4742_ _4742_/A _4742_/B _4742_/C VGND VGND VPWR VPWR _5134_/A sky130_fd_sc_hd__and3_1
XFILLER_147_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4673_ _4673_/A _5016_/B VGND VGND VPWR VPWR _5107_/C sky130_fd_sc_hd__nor2_1
X_6412_ _6432_/A _6428_/B VGND VGND VPWR VPWR _6412_/X sky130_fd_sc_hd__and2_1
X_3624_ _6090_/A1 wire860/X wire813/X _3624_/B2 _3611_/X VGND VGND VPWR VPWR _3627_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6343_ _7186_/Q _6343_/A2 _5650_/Y VGND VGND VPWR VPWR _6343_/X sky130_fd_sc_hd__o21ba_1
XFILLER_127_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3555_ _3555_/A1 _3302_/Y _3555_/B1 _5933_/B2 VGND VGND VPWR VPWR _3555_/X sky130_fd_sc_hd__a22o_1
XFILLER_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6274_ _6274_/A1 _6274_/A2 _6323_/B1 _6274_/B2 VGND VGND VPWR VPWR _6274_/X sky130_fd_sc_hd__a22o_1
X_3486_ _6982_/Q _3486_/A2 _3486_/B1 _3486_/B2 VGND VGND VPWR VPWR _3486_/X sky130_fd_sc_hd__a22o_1
XFILLER_102_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5225_ _5225_/A _5225_/B VGND VGND VPWR VPWR _5228_/S sky130_fd_sc_hd__and2_1
XFILLER_142_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5156_ _5156_/A _5156_/B _5156_/C VGND VGND VPWR VPWR _5156_/Y sky130_fd_sc_hd__nor3_1
XFILLER_111_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4107_ _4114_/A0 hold553/X _4107_/S VGND VGND VPWR VPWR _6576_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5087_ _5155_/B _5087_/B VGND VGND VPWR VPWR _5087_/X sky130_fd_sc_hd__or2_1
X_4038_ hold635/X _4298_/A0 _4039_/S VGND VGND VPWR VPWR _6529_/D sky130_fd_sc_hd__mux2_1
XFILLER_25_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5989_ _6000_/A _6033_/A _6020_/C VGND VGND VPWR VPWR _6022_/B sky130_fd_sc_hd__and3_1
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_50 _6132_/C1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_61 _5734_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_72 wire1904/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_83 _6330_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_94 _5959_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput190 _3211_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[23] sky130_fd_sc_hd__buf_12
XFILLER_153_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold309 _6674_/Q VGND VGND VPWR VPWR hold309/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3340_ _3344_/A hold85/A VGND VGND VPWR VPWR _3340_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_3_4_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A VGND VGND VPWR VPWR _7206_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _3297_/A hold27/X VGND VGND VPWR VPWR hold28/A sky130_fd_sc_hd__or2_1
XFILLER_140_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _5042_/C _5148_/B _5134_/B _5010_/D VGND VGND VPWR VPWR _5010_/X sky130_fd_sc_hd__or4_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6961_ _7109_/CLK _6961_/D wire3999/A VGND VGND VPWR VPWR _6961_/Q sky130_fd_sc_hd__dfrtp_1
X_5912_ _6285_/B2 _5936_/B1 _5912_/B1 _6603_/Q _5911_/X VGND VGND VPWR VPWR _5913_/D
+ sky130_fd_sc_hd__a221o_1
X_6892_ _7127_/CLK _6892_/D wire4061/A VGND VGND VPWR VPWR _6892_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5843_ _7025_/Q _5843_/A2 _5843_/B1 _6198_/A1 VGND VGND VPWR VPWR _5843_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5774_ _7165_/Q _5773_/X _6171_/S VGND VGND VPWR VPWR _7165_/D sky130_fd_sc_hd__mux2_1
X_4725_ _4731_/C _4731_/B _4444_/Y _4378_/B VGND VGND VPWR VPWR _5001_/C sky130_fd_sc_hd__a211oi_4
XFILLER_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4656_ _4668_/A _4942_/A VGND VGND VPWR VPWR _4656_/Y sky130_fd_sc_hd__nor2_1
XFILLER_147_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3607_ _3711_/A _3607_/B VGND VGND VPWR VPWR _3607_/Y sky130_fd_sc_hd__nor2_1
Xinput70 mgmt_gpio_in[7] VGND VGND VPWR VPWR input70/X sky130_fd_sc_hd__clkbuf_1
Xinput81 spi_sdo VGND VGND VPWR VPWR input81/X sky130_fd_sc_hd__clkbuf_1
X_4587_ _4632_/A _4587_/B VGND VGND VPWR VPWR _4965_/A sky130_fd_sc_hd__nor2_1
Xinput92 spimemio_flash_io3_oeb VGND VGND VPWR VPWR input92/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6326_ _6326_/A1 _6326_/A2 _6326_/B1 _7211_/Q _6325_/X VGND VGND VPWR VPWR _6331_/B
+ sky130_fd_sc_hd__a221o_1
X_3538_ _3538_/A _3538_/B VGND VGND VPWR VPWR _4222_/A sky130_fd_sc_hd__nor2_1
Xwire3807 _4749_/B VGND VGND VPWR VPWR _4876_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_107_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3818 _4629_/A VGND VGND VPWR VPWR _4814_/A sky130_fd_sc_hd__clkbuf_2
Xwire3829 _4819_/C VGND VGND VPWR VPWR _4544_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_88_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6257_ _6257_/A _6257_/B _6257_/C _6257_/D VGND VGND VPWR VPWR _6257_/X sky130_fd_sc_hd__or4_1
X_3469_ _6846_/Q _3605_/B1 _3469_/B1 _3469_/B2 VGND VGND VPWR VPWR _3469_/X sky130_fd_sc_hd__a22o_1
XFILLER_67_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5208_ hold699/X _5208_/A1 _5209_/S VGND VGND VPWR VPWR _6809_/D sky130_fd_sc_hd__mux2_1
XFILLER_190_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6188_ _6188_/A1 _6188_/A2 _6188_/B1 _6188_/B2 VGND VGND VPWR VPWR _6188_/X sky130_fd_sc_hd__a22o_1
XFILLER_69_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5139_ _5139_/A _5139_/B _5139_/C _5139_/D VGND VGND VPWR VPWR _5139_/X sky130_fd_sc_hd__or4_1
XFILLER_184_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length2197 _6738_/Q VGND VGND VPWR VPWR _3618_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4510_ _4510_/A _4510_/B _4510_/C VGND VGND VPWR VPWR _4510_/X sky130_fd_sc_hd__and3_1
XFILLER_117_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5490_ _5490_/A0 hold487/X _5490_/S VGND VGND VPWR VPWR _7055_/D sky130_fd_sc_hd__mux2_1
XFILLER_184_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold106 _6450_/Q VGND VGND VPWR VPWR hold106/X sky130_fd_sc_hd__dlygate4sd3_1
X_4441_ _4441_/A _4443_/B VGND VGND VPWR VPWR _4994_/A sky130_fd_sc_hd__or2_2
Xhold117 _3267_/Y VGND VGND VPWR VPWR hold117/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 _4292_/X VGND VGND VPWR VPWR _6739_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 _6749_/Q VGND VGND VPWR VPWR hold139/X sky130_fd_sc_hd__dlygate4sd3_1
X_7160_ _7180_/CLK _7160_/D fanout3986/X VGND VGND VPWR VPWR _7160_/Q sky130_fd_sc_hd__dfrtp_1
X_4372_ _4570_/C _4781_/B VGND VGND VPWR VPWR _4372_/Y sky130_fd_sc_hd__nor2_1
XFILLER_171_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6111_ _6111_/A1 _6111_/A2 _6111_/B1 _6111_/B2 VGND VGND VPWR VPWR _6111_/X sky130_fd_sc_hd__a22o_1
XFILLER_113_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3323_ _3546_/B _3476_/A VGND VGND VPWR VPWR _3323_/Y sky130_fd_sc_hd__nor2_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7091_ _7091_/CLK _7091_/D fanout4028/X VGND VGND VPWR VPWR _7091_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_112_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6042_ _6978_/Q _6042_/A2 _6042_/B1 _6042_/B2 _6041_/X VGND VGND VPWR VPWR _6042_/X
+ sky130_fd_sc_hd__a221o_1
X_3254_ hold166/X _3254_/A1 _3941_/A VGND VGND VPWR VPWR _3270_/B sky130_fd_sc_hd__mux2_1
XFILLER_98_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3185_ hold81/A VGND VGND VPWR VPWR _3830_/A sky130_fd_sc_hd__inv_2
XFILLER_39_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6944_ _7017_/CLK _6944_/D fanout4078/X VGND VGND VPWR VPWR _6944_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6875_ _7135_/CLK _6875_/D wire4056/A VGND VGND VPWR VPWR hold93/A sky130_fd_sc_hd__dfstp_1
X_5826_ _6936_/Q _5826_/A2 _5826_/B1 _6179_/A1 VGND VGND VPWR VPWR _5826_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5757_ _6115_/B2 _5757_/A2 _5757_/B1 _5757_/B2 _5754_/X VGND VGND VPWR VPWR _5757_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4708_ _4708_/A _4708_/B _4708_/C _4850_/B VGND VGND VPWR VPWR _4708_/X sky130_fd_sc_hd__and4_1
X_5688_ _5688_/A _5703_/B _5699_/B VGND VGND VPWR VPWR _5688_/X sky130_fd_sc_hd__and3_1
XFILLER_175_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4639_ _4639_/A _4639_/B VGND VGND VPWR VPWR _4985_/A sky130_fd_sc_hd__nor2_1
Xwire4305 _4570_/A VGND VGND VPWR VPWR _4846_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_162_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold640 _7009_/Q VGND VGND VPWR VPWR hold640/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_118_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold651 _6937_/Q VGND VGND VPWR VPWR hold651/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 _6597_/Q VGND VGND VPWR VPWR hold662/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3604 _5513_/A0 VGND VGND VPWR VPWR _5450_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3615 wire3616/X VGND VGND VPWR VPWR _4266_/A1 sky130_fd_sc_hd__clkbuf_1
Xhold673 _6498_/Q VGND VGND VPWR VPWR hold673/X sky130_fd_sc_hd__dlygate4sd3_1
X_6309_ _6309_/A1 _6309_/A2 _6309_/B1 _6744_/Q _6309_/C1 VGND VGND VPWR VPWR _6316_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold684 _6936_/Q VGND VGND VPWR VPWR hold684/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 _6600_/Q VGND VGND VPWR VPWR hold695/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2903 _5763_/A2 VGND VGND VPWR VPWR _5721_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire2914 _5757_/B1 VGND VGND VPWR VPWR _5776_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2925 wire2926/X VGND VGND VPWR VPWR _5852_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire2936 wire2937/X VGND VGND VPWR VPWR _5917_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire2947 wire2948/X VGND VGND VPWR VPWR _5929_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_131_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2958 _5686_/X VGND VGND VPWR VPWR _5821_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_134_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length1282 _3290_/Y VGND VGND VPWR VPWR wire1277/A sky130_fd_sc_hd__clkbuf_1
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4990_ _4979_/X _4990_/B VGND VGND VPWR VPWR _4991_/B sky130_fd_sc_hd__and2b_1
XFILLER_23_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3941_ _3941_/A _3941_/B VGND VGND VPWR VPWR _3941_/Y sky130_fd_sc_hd__nor2_2
XFILLER_90_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6660_ _7092_/CLK _6660_/D wire3945/A VGND VGND VPWR VPWR _6660_/Q sky130_fd_sc_hd__dfrtp_1
X_3872_ _6820_/Q _3872_/B _3872_/C VGND VGND VPWR VPWR _3872_/Y sky130_fd_sc_hd__nor3_1
XFILLER_149_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5611_ _6564_/Q _5609_/Y _7148_/Q VGND VGND VPWR VPWR _7148_/D sky130_fd_sc_hd__mux2_1
XFILLER_149_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6591_ _6989_/CLK _6591_/D wire3995/X VGND VGND VPWR VPWR _6591_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5542_ hold567/X _5587_/A0 _5542_/S VGND VGND VPWR VPWR _7101_/D sky130_fd_sc_hd__mux2_1
XFILLER_157_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5473_ hold617/X _5491_/A0 _5474_/S VGND VGND VPWR VPWR _7040_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4424_ _4758_/A _4758_/B _4758_/C VGND VGND VPWR VPWR _4424_/Y sky130_fd_sc_hd__nand3_1
X_4355_ _4544_/B _4359_/B _4402_/A VGND VGND VPWR VPWR _4355_/Y sky130_fd_sc_hd__a21oi_1
X_7143_ _7187_/CLK _7143_/D _6562_/SET_B VGND VGND VPWR VPWR _7143_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3306_ _3518_/B _3318_/B VGND VGND VPWR VPWR _3306_/Y sky130_fd_sc_hd__nor2_1
X_7074_ _7074_/CLK _7074_/D fanout3976/X VGND VGND VPWR VPWR _7074_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_101_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4286_ _4286_/A0 hold378/X _4287_/S VGND VGND VPWR VPWR _6734_/D sky130_fd_sc_hd__mux2_1
XFILLER_100_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1509 _3460_/B VGND VGND VPWR VPWR _3538_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_140_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6025_ _6025_/A _6025_/B _6025_/C _6025_/D VGND VGND VPWR VPWR _6026_/D sky130_fd_sc_hd__or4_1
X_3237_ _4450_/A VGND VGND VPWR VPWR _4667_/C sky130_fd_sc_hd__inv_2
XFILLER_39_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6927_ _6973_/CLK _6927_/D fanout4078/X VGND VGND VPWR VPWR _6927_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6858_ _7121_/CLK _6858_/D wire4041/X VGND VGND VPWR VPWR _6858_/Q sky130_fd_sc_hd__dfstp_1
Xwire806 _3527_/X VGND VGND VPWR VPWR wire806/X sky130_fd_sc_hd__clkbuf_1
X_5809_ _6887_/Q _5831_/A2 _5831_/B1 _5809_/B2 VGND VGND VPWR VPWR _5809_/X sky130_fd_sc_hd__a22o_1
XFILLER_183_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire817 wire818/X VGND VGND VPWR VPWR wire817/X sky130_fd_sc_hd__clkbuf_1
X_6789_ _3487_/B2 _6789_/D _6440_/X VGND VGND VPWR VPWR _6789_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_167_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire839 wire840/X VGND VGND VPWR VPWR wire839/X sky130_fd_sc_hd__clkbuf_1
XFILLER_129_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire4102 wire4103/X VGND VGND VPWR VPWR wire4102/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4113 wire4114/X VGND VGND VPWR VPWR _3943_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire4124 input66/X VGND VGND VPWR VPWR _3427_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_151_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire4135 wire4136/X VGND VGND VPWR VPWR wire4135/X sky130_fd_sc_hd__clkbuf_1
XFILLER_150_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4146 wire4147/X VGND VGND VPWR VPWR _3407_/B2 sky130_fd_sc_hd__clkbuf_1
Xhold470 _7104_/Q VGND VGND VPWR VPWR hold470/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3412 wire3413/X VGND VGND VPWR VPWR wire3412/X sky130_fd_sc_hd__clkbuf_1
Xwire4157 wire4158/X VGND VGND VPWR VPWR wire4157/X sky130_fd_sc_hd__clkbuf_1
Xwire4168 input56/X VGND VGND VPWR VPWR wire4168/X sky130_fd_sc_hd__clkbuf_1
Xhold481 _7112_/Q VGND VGND VPWR VPWR hold481/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3434 _5568_/A0 VGND VGND VPWR VPWR _5517_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire4179 wire4180/X VGND VGND VPWR VPWR wire4179/X sky130_fd_sc_hd__clkbuf_1
XFILLER_150_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2700 _6024_/C VGND VGND VPWR VPWR _6303_/B1 sky130_fd_sc_hd__clkbuf_2
Xhold492 _6662_/Q VGND VGND VPWR VPWR hold492/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire2711 _6205_/A2 VGND VGND VPWR VPWR _6087_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_131_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2722 _6136_/A2 VGND VGND VPWR VPWR _6061_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3478 _5291_/A0 VGND VGND VPWR VPWR _5381_/A0 sky130_fd_sc_hd__clkbuf_2
Xwire2744 _6008_/X VGND VGND VPWR VPWR _6023_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3489 _4208_/A1 VGND VGND VPWR VPWR _4139_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2755 _6211_/A2 VGND VGND VPWR VPWR _6114_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2777 _6298_/B1 VGND VGND VPWR VPWR _6327_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire2788 _6092_/B1 VGND VGND VPWR VPWR _6208_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_38_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2799 wire2799/A VGND VGND VPWR VPWR wire2799/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4140_ hold592/X _4251_/A0 _4140_/S VGND VGND VPWR VPWR _6605_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4071_ hold241/X _4130_/A1 _4083_/S VGND VGND VPWR VPWR _4071_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4973_ _5140_/A _4973_/B VGND VGND VPWR VPWR _4979_/C sky130_fd_sc_hd__or2_1
XFILLER_51_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6712_ _7112_/CLK _6712_/D wire4026/X VGND VGND VPWR VPWR _6712_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_177_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3924_ _6575_/Q _3924_/A1 _3958_/B VGND VGND VPWR VPWR _3924_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6643_ _7206_/CLK _6643_/D VGND VGND VPWR VPWR _6643_/Q sky130_fd_sc_hd__dfxtp_1
X_3855_ _6455_/Q _3856_/B _3854_/Y _6454_/Q VGND VGND VPWR VPWR _6455_/D sky130_fd_sc_hd__o22a_1
XFILLER_164_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3786_ _5999_/A1 _3298_/Y _3786_/B1 _6761_/Q _3785_/X VGND VGND VPWR VPWR _3788_/C
+ sky130_fd_sc_hd__a221o_1
X_6574_ _6705_/CLK _6574_/D _6437_/A VGND VGND VPWR VPWR _6574_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_117_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5525_ _5585_/A0 hold292/X _5525_/S VGND VGND VPWR VPWR _7086_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5456_ _5456_/A0 hold689/X _5456_/S VGND VGND VPWR VPWR _7025_/D sky130_fd_sc_hd__mux2_1
XFILLER_105_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4407_ _4407_/A _4538_/B VGND VGND VPWR VPWR _4436_/B sky130_fd_sc_hd__xnor2_2
XFILLER_99_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5387_ _5387_/A0 hold269/X _5388_/S VGND VGND VPWR VPWR _6963_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2007 _6892_/Q VGND VGND VPWR VPWR _6077_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_160_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2018 _3577_/A1 VGND VGND VPWR VPWR _5756_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
X_7126_ _7126_/CLK _7126_/D wire4046/A VGND VGND VPWR VPWR _7126_/Q sky130_fd_sc_hd__dfrtp_1
X_4338_ _4338_/A _4338_/B _4338_/C _4338_/D VGND VGND VPWR VPWR _4348_/B sky130_fd_sc_hd__and4_1
Xwire2029 _6880_/Q VGND VGND VPWR VPWR _3381_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1306 _6308_/X VGND VGND VPWR VPWR _6309_/C1 sky130_fd_sc_hd__clkbuf_1
XFILLER_113_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1317 _5999_/X VGND VGND VPWR VPWR wire1317/X sky130_fd_sc_hd__clkbuf_1
XFILLER_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4269_ hold579/X _4329_/A1 _4269_/S VGND VGND VPWR VPWR _6720_/D sky130_fd_sc_hd__mux2_1
X_7057_ _7125_/CLK _7057_/D wire4046/A VGND VGND VPWR VPWR _7057_/Q sky130_fd_sc_hd__dfrtp_2
Xwire1328 _5832_/X VGND VGND VPWR VPWR wire1328/X sky130_fd_sc_hd__clkbuf_1
Xwire1339 _4830_/Y VGND VGND VPWR VPWR _5126_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_46_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6008_ _6033_/A _6020_/C _6030_/C VGND VGND VPWR VPWR _6008_/X sky130_fd_sc_hd__and3_1
XFILLER_67_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire603 _5506_/S VGND VGND VPWR VPWR _5504_/S sky130_fd_sc_hd__clkbuf_1
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire625 wire625/A VGND VGND VPWR VPWR _5482_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_168_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire636 _5464_/S VGND VGND VPWR VPWR _5463_/S sky130_fd_sc_hd__dlymetal6s2s_1
Xwire658 _5429_/S VGND VGND VPWR VPWR _5424_/S sky130_fd_sc_hd__clkbuf_2
Xwire669 wire670/X VGND VGND VPWR VPWR _5411_/S sky130_fd_sc_hd__clkbuf_2
Xmax_length3987 fanout3986/X VGND VGND VPWR VPWR _6562_/SET_B sky130_fd_sc_hd__buf_2
XFILLER_6_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3220 _4453_/C VGND VGND VPWR VPWR _4443_/B sky130_fd_sc_hd__buf_2
XFILLER_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3231 _4759_/A VGND VGND VPWR VPWR _4735_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3242 _4231_/Y VGND VGND VPWR VPWR _5182_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2530 _6185_/B1 VGND VGND VPWR VPWR _6213_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire2541 _6187_/A2 VGND VGND VPWR VPWR _6201_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire3286 hold56/X VGND VGND VPWR VPWR hold57/A sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3297 _6443_/Q VGND VGND VPWR VPWR wire3297/X sky130_fd_sc_hd__clkbuf_1
Xwire2552 _5997_/Y VGND VGND VPWR VPWR wire2552/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2563 _6027_/A VGND VGND VPWR VPWR wire2563/X sky130_fd_sc_hd__clkbuf_1
XFILLER_172_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2574 _6183_/B1 VGND VGND VPWR VPWR wire2574/X sky130_fd_sc_hd__clkbuf_1
Xwire1840 _6994_/Q VGND VGND VPWR VPWR wire1840/X sky130_fd_sc_hd__clkbuf_1
Xwire2585 _5836_/A2 VGND VGND VPWR VPWR _5709_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_93_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1851 _5416_/A1 VGND VGND VPWR VPWR wire1851/X sky130_fd_sc_hd__clkbuf_1
Xwire2596 _4770_/A VGND VGND VPWR VPWR _4822_/A sky130_fd_sc_hd__clkbuf_1
Xwire1862 wire1862/A VGND VGND VPWR VPWR _6132_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire1873 wire1874/X VGND VGND VPWR VPWR wire1873/X sky130_fd_sc_hd__clkbuf_1
XFILLER_46_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1884 _6960_/Q VGND VGND VPWR VPWR _6188_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1895 hold136/X VGND VGND VPWR VPWR _5735_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3640_ _3640_/A1 _3315_/Y _4282_/A _6733_/Q VGND VGND VPWR VPWR _3640_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3571_ _3571_/A1 _3571_/A2 _3528_/Y _6624_/Q VGND VGND VPWR VPWR _3571_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5310_ _5508_/A0 hold530/X _5310_/S VGND VGND VPWR VPWR _6895_/D sky130_fd_sc_hd__mux2_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6290_ _6613_/Q _6290_/A2 _6327_/B1 _6290_/B2 _6289_/X VGND VGND VPWR VPWR _6291_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_114_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5241_ _5241_/A _5241_/B _5241_/C _5241_/D VGND VGND VPWR VPWR hold8/A sky130_fd_sc_hd__or4_1
XFILLER_170_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5172_ _5172_/A _5172_/B _5172_/C _5172_/D VGND VGND VPWR VPWR _5183_/A sky130_fd_sc_hd__nor4_1
XFILLER_68_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4123_ _5208_/A1 hold589/X _4125_/S VGND VGND VPWR VPWR _6590_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4054_ hold341/X _5242_/A0 _4060_/S VGND VGND VPWR VPWR _4054_/X sky130_fd_sc_hd__mux2_1
Xinput2 debug_oeb VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_opt_1_0_csclk _7117_/CLK VGND VGND VPWR VPWR clkbuf_opt_1_0_csclk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_37_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4956_ _4997_/A _4526_/B _4935_/C _4944_/X _4916_/B VGND VGND VPWR VPWR _5163_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_189_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3907_ _3907_/A _5592_/B VGND VGND VPWR VPWR _5651_/A sky130_fd_sc_hd__nor2_1
XFILLER_32_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4887_ _4885_/X _4887_/B _4887_/C _4887_/D VGND VGND VPWR VPWR _4890_/B sky130_fd_sc_hd__nand4b_1
XFILLER_138_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6626_ _7193_/CLK _6626_/D VGND VGND VPWR VPWR _6626_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3838_ _6541_/Q _3838_/B VGND VGND VPWR VPWR _3839_/B sky130_fd_sc_hd__nand2_1
XFILLER_192_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length2527 _6139_/A2 VGND VGND VPWR VPWR _6064_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_118_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6557_ _6989_/CLK _6557_/D wire3995/X VGND VGND VPWR VPWR _6557_/Q sky130_fd_sc_hd__dfrtp_1
X_3769_ _3769_/A1 _3314_/Y _3769_/B1 _3769_/B2 wire744/X VGND VGND VPWR VPWR _3769_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_106_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5508_ _5508_/A0 hold536/X _5510_/S VGND VGND VPWR VPWR _7071_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6488_ _7027_/CLK _6488_/D fanout3976/X VGND VGND VPWR VPWR _6488_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5439_ _5439_/A _5553_/B VGND VGND VPWR VPWR _5439_/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7109_ _7109_/CLK _7109_/D wire3999/A VGND VGND VPWR VPWR _7109_/Q sky130_fd_sc_hd__dfrtp_1
Xwire1103 wire1103/A VGND VGND VPWR VPWR _3692_/C1 sky130_fd_sc_hd__clkbuf_1
XFILLER_75_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1114 _3652_/A2 VGND VGND VPWR VPWR _3699_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1125 _3564_/A2 VGND VGND VPWR VPWR _3442_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1136 _3331_/Y VGND VGND VPWR VPWR _3498_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_142_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1147 _3654_/B1 VGND VGND VPWR VPWR _3426_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_101_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1158 _3452_/A2 VGND VGND VPWR VPWR _3685_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_28_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire400 _5050_/X VGND VGND VPWR VPWR wire400/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire411 wire412/X VGND VGND VPWR VPWR _4086_/S sky130_fd_sc_hd__clkbuf_2
Xwire422 _3651_/X VGND VGND VPWR VPWR _3659_/A sky130_fd_sc_hd__clkbuf_1
Xwire433 _3563_/X VGND VGND VPWR VPWR wire433/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire444 _6293_/X VGND VGND VPWR VPWR wire444/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire455 _6070_/X VGND VGND VPWR VPWR wire455/X sky130_fd_sc_hd__clkbuf_1
XFILLER_144_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire466 _5586_/S VGND VGND VPWR VPWR _5581_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire477 wire478/X VGND VGND VPWR VPWR _5555_/S sky130_fd_sc_hd__clkbuf_2
Xwire488 _5327_/S VGND VGND VPWR VPWR _5325_/S sky130_fd_sc_hd__clkbuf_2
Xwire499 wire500/X VGND VGND VPWR VPWR wire499/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_606 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3050 wire3051/X VGND VGND VPWR VPWR _5943_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire3061 _5956_/B1 VGND VGND VPWR VPWR _5944_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3072 wire3073/X VGND VGND VPWR VPWR _5878_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire3083 _5666_/X VGND VGND VPWR VPWR wire3083/X sky130_fd_sc_hd__clkbuf_1
Xwire3094 _5788_/A2 VGND VGND VPWR VPWR _5716_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2371 _6531_/Q VGND VGND VPWR VPWR _6222_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2382 wire2383/X VGND VGND VPWR VPWR wire2382/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2393 wire2394/X VGND VGND VPWR VPWR _6264_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire1670 hold602/X VGND VGND VPWR VPWR _5990_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1681 _6138_/B2 VGND VGND VPWR VPWR _5775_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1692 wire1693/X VGND VGND VPWR VPWR _3784_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_81_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4810_ _4806_/X _4810_/B _4810_/C _4810_/D VGND VGND VPWR VPWR _4810_/X sky130_fd_sc_hd__and4b_1
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5790_ _6135_/B2 _5790_/A2 _5790_/B1 _7062_/Q VGND VGND VPWR VPWR _5790_/X sky130_fd_sc_hd__a22o_1
XFILLER_187_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4741_ _4931_/B _4742_/C _4741_/C VGND VGND VPWR VPWR _4741_/X sky130_fd_sc_hd__and3_1
XFILLER_147_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4672_ _4672_/A _4686_/B VGND VGND VPWR VPWR _4672_/X sky130_fd_sc_hd__or2_1
X_6411_ _6432_/A _6428_/B VGND VGND VPWR VPWR _6411_/X sky130_fd_sc_hd__and2_1
XFILLER_135_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3623_ _3623_/A1 _3415_/Y _3466_/Y _3623_/B2 _3612_/X VGND VGND VPWR VPWR _3627_/A
+ sky130_fd_sc_hd__a221o_1
X_6342_ _6342_/A1 _6342_/A2 _6332_/X _6341_/X _6342_/C1 VGND VGND VPWR VPWR _6342_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_162_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3554_ _6744_/Q _4294_/A _4034_/A _3554_/B2 VGND VGND VPWR VPWR _3554_/X sky130_fd_sc_hd__a22o_1
XFILLER_155_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3485_ _3525_/A _3485_/B VGND VGND VPWR VPWR _6392_/A sky130_fd_sc_hd__nor2_1
X_6273_ _6273_/A1 _6336_/A2 _6273_/B1 _6273_/B2 VGND VGND VPWR VPWR _6273_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5224_ _5224_/A0 hold375/X _5224_/S VGND VGND VPWR VPWR _6820_/D sky130_fd_sc_hd__mux2_1
X_5155_ _5155_/A _5155_/B _5155_/C _4681_/X VGND VGND VPWR VPWR _5178_/C sky130_fd_sc_hd__or4b_1
XFILLER_57_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4106_ _4206_/A1 hold625/X _4108_/S VGND VGND VPWR VPWR _6575_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5086_ _5156_/B _5178_/A _5106_/C _5086_/D VGND VGND VPWR VPWR _5087_/B sky130_fd_sc_hd__or4_1
XFILLER_84_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4037_ hold688/X _6395_/A0 _4039_/S VGND VGND VPWR VPWR _6528_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5988_ _6014_/A _6040_/B _6040_/C VGND VGND VPWR VPWR _5988_/X sky130_fd_sc_hd__and3_1
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4939_ _5065_/D _5124_/C _4939_/C VGND VGND VPWR VPWR _4961_/A sky130_fd_sc_hd__or3_1
XFILLER_178_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_40 _6144_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_51 wire1428/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_62 _3487_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 _3667_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmax_length3058 _5671_/X VGND VGND VPWR VPWR _5824_/B1 sky130_fd_sc_hd__clkbuf_1
XANTENNA_84 _6204_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6609_ _7208_/CLK _6609_/D wire4026/A VGND VGND VPWR VPWR _6609_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_95 _5789_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput180 _3220_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[14] sky130_fd_sc_hd__buf_12
Xoutput191 _3210_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[24] sky130_fd_sc_hd__buf_12
XFILLER_153_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length4282 _4553_/A VGND VGND VPWR VPWR _4564_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_117_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length4293 _4342_/C VGND VGND VPWR VPWR _4565_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_184_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3581 _4122_/A0 VGND VGND VPWR VPWR _4131_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_116_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_44_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7089_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_137_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3270_ hold26/X _3270_/B VGND VGND VPWR VPWR hold27/A sky130_fd_sc_hd__nand2_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_59_csclk _7117_/CLK VGND VGND VPWR VPWR _7072_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_85_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2190 wire2191/X VGND VGND VPWR VPWR _6323_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_66_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6960_ _7109_/CLK _6960_/D wire3999/X VGND VGND VPWR VPWR _6960_/Q sky130_fd_sc_hd__dfrtp_1
X_5911_ _5911_/A1 _5953_/A2 _5963_/A2 _5911_/B2 VGND VGND VPWR VPWR _5911_/X sky130_fd_sc_hd__a22o_1
X_6891_ _7127_/CLK _6891_/D _6923_/SET_B VGND VGND VPWR VPWR _6891_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_62_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5842_ _5842_/A1 _5842_/A2 _5842_/B1 _6215_/B2 _5841_/X VGND VGND VPWR VPWR _5847_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_179_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5773_ _6121_/A1 _7164_/Q _5772_/X VGND VGND VPWR VPWR _5773_/X sky130_fd_sc_hd__a21o_1
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4724_ _4724_/A _4724_/B VGND VGND VPWR VPWR _4742_/C sky130_fd_sc_hd__nor2_1
XFILLER_174_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4655_ _4694_/A _4655_/B VGND VGND VPWR VPWR _5177_/B sky130_fd_sc_hd__nor2_1
Xinput60 mgmt_gpio_in[31] VGND VGND VPWR VPWR input60/X sky130_fd_sc_hd__clkbuf_1
X_3606_ _3606_/A1 wire956/X wire935/X _6077_/A1 VGND VGND VPWR VPWR _3606_/X sky130_fd_sc_hd__a22o_1
XFILLER_190_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput71 mgmt_gpio_in[8] VGND VGND VPWR VPWR input71/X sky130_fd_sc_hd__clkbuf_1
Xinput82 spi_sdoenb VGND VGND VPWR VPWR input82/X sky130_fd_sc_hd__clkbuf_1
X_4586_ _4629_/A _5018_/C VGND VGND VPWR VPWR _4587_/B sky130_fd_sc_hd__or2_1
Xinput93 trap VGND VGND VPWR VPWR input93/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6325_ _6659_/Q _6325_/A2 _6325_/B1 _6325_/B2 VGND VGND VPWR VPWR _6325_/X sky130_fd_sc_hd__a22o_1
X_3537_ _5777_/A1 _3537_/A2 _3536_/Y _6339_/A1 _3535_/X VGND VGND VPWR VPWR _3541_/C
+ sky130_fd_sc_hd__a221o_1
Xwire3808 _4971_/B VGND VGND VPWR VPWR _4749_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3819 _4638_/A VGND VGND VPWR VPWR _4629_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6256_ _6712_/Q _6256_/A2 _6256_/B1 _6256_/B2 _6255_/X VGND VGND VPWR VPWR _6257_/D
+ sky130_fd_sc_hd__a221o_1
X_3468_ _3468_/A _3468_/B _3468_/C _3468_/D VGND VGND VPWR VPWR _3543_/A sky130_fd_sc_hd__or4_1
XFILLER_103_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5207_ hold702/X _5220_/A0 _5209_/S VGND VGND VPWR VPWR _6808_/D sky130_fd_sc_hd__mux2_1
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6187_ _7016_/Q _6187_/A2 _6187_/B1 _6187_/B2 _6186_/X VGND VGND VPWR VPWR _6192_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3399_ _7101_/Q _3399_/A2 wire951/X _7141_/Q _3398_/X VGND VGND VPWR VPWR _3399_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5138_ _5148_/C _5138_/B VGND VGND VPWR VPWR _5139_/D sky130_fd_sc_hd__and2b_1
XFILLER_29_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5069_ _5069_/A _5160_/A VGND VGND VPWR VPWR _5104_/B sky130_fd_sc_hd__nor2_1
XFILLER_84_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length2154 _6254_/A1 VGND VGND VPWR VPWR wire2152/A sky130_fd_sc_hd__clkbuf_1
XFILLER_165_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length1497 _3416_/Y VGND VGND VPWR VPWR wire1496/A sky130_fd_sc_hd__clkbuf_1
XFILLER_106_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4440_ _4441_/A _4443_/B VGND VGND VPWR VPWR _4516_/B sky130_fd_sc_hd__nor2_4
Xhold107 _3977_/X VGND VGND VPWR VPWR hold107/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold118 _4279_/X VGND VGND VPWR VPWR _6728_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 _7046_/Q VGND VGND VPWR VPWR hold129/X sky130_fd_sc_hd__dlygate4sd3_1
X_4371_ _4570_/A _4570_/B VGND VGND VPWR VPWR _4781_/B sky130_fd_sc_hd__nand2_1
XFILLER_171_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6110_ _6110_/A _6110_/B VGND VGND VPWR VPWR _6110_/X sky130_fd_sc_hd__or2_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3322_ _3322_/A _3511_/B VGND VGND VPWR VPWR _3322_/Y sky130_fd_sc_hd__nor2_1
X_7090_ _7090_/CLK _7090_/D fanout3944/X VGND VGND VPWR VPWR _7090_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6041_ _6962_/Q _6078_/A2 _6063_/B1 _7042_/Q VGND VGND VPWR VPWR _6041_/X sky130_fd_sc_hd__a22o_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ hold165/X _3820_/A _3818_/A VGND VGND VPWR VPWR _3253_/X sky130_fd_sc_hd__a21bo_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3184_ _6472_/Q VGND VGND VPWR VPWR _3184_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6943_ _7017_/CLK _6943_/D fanout4078/X VGND VGND VPWR VPWR _6943_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_81_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6874_ _7135_/CLK _6874_/D wire4056/X VGND VGND VPWR VPWR _6874_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_62_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5825_ _5825_/A _5825_/B _5825_/C _5825_/D VGND VGND VPWR VPWR _5825_/X sky130_fd_sc_hd__or4_1
X_5756_ _5756_/A1 _5756_/A2 _5756_/B1 _5756_/B2 VGND VGND VPWR VPWR _5756_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length608 _5507_/S VGND VGND VPWR VPWR wire605/A sky130_fd_sc_hd__clkbuf_1
X_4707_ _4707_/A _4707_/B VGND VGND VPWR VPWR _4850_/B sky130_fd_sc_hd__or2_1
XFILLER_108_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5687_ _6031_/A1 _5721_/A2 _5723_/A2 _7010_/Q _5684_/X VGND VGND VPWR VPWR _5687_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4638_ _4638_/A _4638_/B VGND VGND VPWR VPWR _4638_/X sky130_fd_sc_hd__or2_1
XFILLER_162_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4306 wire4307/X VGND VGND VPWR VPWR _3780_/A1 sky130_fd_sc_hd__clkbuf_1
Xhold630 _6481_/Q VGND VGND VPWR VPWR hold630/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold641 _6719_/Q VGND VGND VPWR VPWR hold641/X sky130_fd_sc_hd__dlygate4sd3_1
X_4569_ _4569_/A _4569_/B VGND VGND VPWR VPWR _4569_/Y sky130_fd_sc_hd__nor2_1
Xwire3605 _5468_/A1 VGND VGND VPWR VPWR _5513_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold652 _6849_/Q VGND VGND VPWR VPWR hold652/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 _6920_/Q VGND VGND VPWR VPWR hold663/X sky130_fd_sc_hd__dlygate4sd3_1
X_6308_ _6308_/A1 _6308_/A2 _6308_/B1 _6769_/Q _6308_/C1 VGND VGND VPWR VPWR _6308_/X
+ sky130_fd_sc_hd__a221o_1
Xwire3616 wire3617/X VGND VGND VPWR VPWR wire3616/X sky130_fd_sc_hd__clkbuf_1
Xhold674 _6707_/Q VGND VGND VPWR VPWR hold674/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 _6943_/Q VGND VGND VPWR VPWR hold685/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3649 _4259_/A1 VGND VGND VPWR VPWR _4223_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2904 _5800_/A2 VGND VGND VPWR VPWR _5763_/A2 sky130_fd_sc_hd__clkbuf_1
Xhold696 _6887_/Q VGND VGND VPWR VPWR hold696/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2915 _5840_/B1 VGND VGND VPWR VPWR _5757_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_103_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6239_ _7090_/Q _6298_/A2 _6298_/B1 _6239_/B2 VGND VGND VPWR VPWR _6239_/X sky130_fd_sc_hd__a22o_1
Xwire2926 _5693_/X VGND VGND VPWR VPWR wire2926/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2937 wire2937/A VGND VGND VPWR VPWR wire2937/X sky130_fd_sc_hd__clkbuf_1
Xwire2948 _5820_/A2 VGND VGND VPWR VPWR wire2948/X sky130_fd_sc_hd__clkbuf_1
Xwire2959 wire2959/A VGND VGND VPWR VPWR _5762_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length1272 _3294_/Y VGND VGND VPWR VPWR wire1271/A sky130_fd_sc_hd__clkbuf_1
XFILLER_4_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3940_ _7161_/Q _6814_/Q _3940_/S VGND VGND VPWR VPWR _3940_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3871_ _3951_/A1 _3840_/S _3870_/X _6444_/Q VGND VGND VPWR VPWR _6444_/D sky130_fd_sc_hd__a22o_1
X_5610_ _6562_/Q _6564_/Q VGND VGND VPWR VPWR _5610_/X sky130_fd_sc_hd__or2_1
X_6590_ _6989_/CLK _6590_/D _7161_/RESET_B VGND VGND VPWR VPWR _6590_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5541_ hold498/X _5541_/A1 _5543_/S VGND VGND VPWR VPWR _7100_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5472_ hold491/X _5490_/A0 _5472_/S VGND VGND VPWR VPWR _7039_/D sky130_fd_sc_hd__mux2_1
X_7211_ _7211_/CLK _7211_/D wire4021/X VGND VGND VPWR VPWR _7211_/Q sky130_fd_sc_hd__dfrtp_1
X_4423_ _4758_/A _4758_/B _4758_/C VGND VGND VPWR VPWR _4485_/A sky130_fd_sc_hd__and3_1
XFILLER_160_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7142_ _7142_/CLK _7142_/D wire4046/A VGND VGND VPWR VPWR _7142_/Q sky130_fd_sc_hd__dfrtp_1
X_4354_ _4354_/A _4354_/B VGND VGND VPWR VPWR _4935_/B sky130_fd_sc_hd__nand2_1
XFILLER_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3305_ _3414_/B hold84/X VGND VGND VPWR VPWR _3305_/Y sky130_fd_sc_hd__nand2_1
X_7073_ _7110_/CLK _7073_/D _7110_/RESET_B VGND VGND VPWR VPWR _7073_/Q sky130_fd_sc_hd__dfrtp_2
X_4285_ _4285_/A0 hold381/X _4287_/S VGND VGND VPWR VPWR _6733_/D sky130_fd_sc_hd__mux2_1
XFILLER_98_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6024_ _6024_/A _6024_/B _6024_/C _6024_/D VGND VGND VPWR VPWR _6026_/C sky130_fd_sc_hd__or4_1
XFILLER_140_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3236_ _4396_/A VGND VGND VPWR VPWR _4420_/A sky130_fd_sc_hd__inv_2
XFILLER_73_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6926_ _7130_/CLK _6926_/D wire4061/X VGND VGND VPWR VPWR _6926_/Q sky130_fd_sc_hd__dfrtp_1
X_6857_ _7132_/CLK _6857_/D fanout4077/X VGND VGND VPWR VPWR _6857_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5808_ _6165_/A1 _5817_/B1 _5808_/B1 _6155_/B2 _5807_/X VGND VGND VPWR VPWR _5813_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6788_ _3487_/B2 _6788_/D _6439_/X VGND VGND VPWR VPWR _6788_/Q sky130_fd_sc_hd__dfrtn_1
Xwire818 _3497_/X VGND VGND VPWR VPWR wire818/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire829 wire830/X VGND VGND VPWR VPWR _4288_/A sky130_fd_sc_hd__clkbuf_2
X_5739_ _5739_/A1 _5739_/A2 _5739_/B1 _5739_/B2 _5738_/X VGND VGND VPWR VPWR _5740_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_136_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire4103 _3359_/B2 VGND VGND VPWR VPWR wire4103/X sky130_fd_sc_hd__clkbuf_1
XFILLER_151_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire4114 _3598_/A1 VGND VGND VPWR VPWR wire4114/X sky130_fd_sc_hd__clkbuf_1
Xwire4136 wire4137/X VGND VGND VPWR VPWR wire4136/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4147 wire4148/X VGND VGND VPWR VPWR wire4147/X sky130_fd_sc_hd__clkbuf_1
Xhold460 _6904_/Q VGND VGND VPWR VPWR hold460/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire4158 _3616_/A1 VGND VGND VPWR VPWR wire4158/X sky130_fd_sc_hd__clkbuf_1
Xwire3413 _5527_/A0 VGND VGND VPWR VPWR wire3413/X sky130_fd_sc_hd__clkbuf_1
Xwire3424 _5550_/A0 VGND VGND VPWR VPWR _5577_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold471 _6796_/Q VGND VGND VPWR VPWR hold471/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold482 _6998_/Q VGND VGND VPWR VPWR hold482/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4169 wire4170/X VGND VGND VPWR VPWR _3579_/A1 sky130_fd_sc_hd__clkbuf_1
Xhold493 _6560_/Q VGND VGND VPWR VPWR hold493/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3435 wire3436/X VGND VGND VPWR VPWR _5568_/A0 sky130_fd_sc_hd__clkbuf_2
Xwire2701 _6015_/X VGND VGND VPWR VPWR _6024_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3446 _5198_/A0 VGND VGND VPWR VPWR _4311_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_150_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2712 _6131_/A2 VGND VGND VPWR VPWR _6056_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3468 _5585_/A0 VGND VGND VPWR VPWR _5489_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2723 _6159_/A2 VGND VGND VPWR VPWR _6136_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire2734 _6206_/A2 VGND VGND VPWR VPWR _6086_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_131_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2745 _6166_/A2 VGND VGND VPWR VPWR _6067_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2756 _6160_/A2 VGND VGND VPWR VPWR _6062_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire2767 _6186_/A2 VGND VGND VPWR VPWR _6202_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2778 _5993_/B1 VGND VGND VPWR VPWR _6298_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_161_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2789 _6338_/B1 VGND VGND VPWR VPWR _6092_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_92_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3980 wire3981/X VGND VGND VPWR VPWR wire3980/X sky130_fd_sc_hd__buf_2
XFILLER_96_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3991 wire3992/X VGND VGND VPWR VPWR wire3991/X sky130_fd_sc_hd__buf_2
X_4070_ _4070_/A1 _4070_/A2 wire536/X wire886/X _4276_/B VGND VGND VPWR VPWR _4070_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_96_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4972_ _4783_/A _4794_/C _4971_/Y _4781_/Y _5013_/A VGND VGND VPWR VPWR _4973_/B
+ sky130_fd_sc_hd__o32ai_2
XFILLER_91_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6711_ _7208_/CLK _6711_/D _7112_/SET_B VGND VGND VPWR VPWR _6711_/Q sky130_fd_sc_hd__dfrtp_1
X_3923_ _6574_/Q _3923_/A1 _3958_/B VGND VGND VPWR VPWR _3923_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6642_ _7193_/CLK _6642_/D VGND VGND VPWR VPWR _6642_/Q sky130_fd_sc_hd__dfxtp_1
X_3854_ _3856_/B _3858_/B VGND VGND VPWR VPWR _3854_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6573_ _7084_/CLK hold11/X fanout4057/X VGND VGND VPWR VPWR hold10/A sky130_fd_sc_hd__dfrtp_1
X_3785_ _3785_/A1 _3256_/Y _3286_/Y _4282_/A _6731_/Q VGND VGND VPWR VPWR _3785_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_164_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5524_ _5584_/A0 hold191/X _5525_/S VGND VGND VPWR VPWR _7085_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR clkbuf_2_3_0_mgmt_gpio_in[4]/A
+ sky130_fd_sc_hd__clkbuf_8
X_5455_ _5518_/A0 hold678/X _5455_/S VGND VGND VPWR VPWR _7024_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4406_ _4560_/A _4731_/C _4731_/B VGND VGND VPWR VPWR _4453_/A sky130_fd_sc_hd__nand3_2
XFILLER_160_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5386_ _5554_/A0 hold327/X _5388_/S VGND VGND VPWR VPWR _6962_/D sky130_fd_sc_hd__mux2_1
XFILLER_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7125_ _7125_/CLK _7125_/D wire4049/A VGND VGND VPWR VPWR _7125_/Q sky130_fd_sc_hd__dfrtp_1
Xwire2008 _6062_/B2 VGND VGND VPWR VPWR _3664_/A1 sky130_fd_sc_hd__clkbuf_1
X_4337_ _4337_/A _4337_/B _4337_/C _4337_/D VGND VGND VPWR VPWR _4348_/A sky130_fd_sc_hd__and4_1
Xwire2019 wire2020/X VGND VGND VPWR VPWR _3577_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_87_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1307 _6288_/X VGND VGND VPWR VPWR _6291_/C sky130_fd_sc_hd__clkbuf_1
X_7056_ _7056_/CLK _7056_/D fanout3976/X VGND VGND VPWR VPWR _7056_/Q sky130_fd_sc_hd__dfrtp_1
Xwire1318 wire1319/X VGND VGND VPWR VPWR _6012_/A sky130_fd_sc_hd__clkbuf_1
X_4268_ hold641/X _5452_/A0 _4268_/S VGND VGND VPWR VPWR _6719_/D sky130_fd_sc_hd__mux2_1
Xwire1329 wire1330/X VGND VGND VPWR VPWR _5785_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6007_ _6019_/A _6038_/B VGND VGND VPWR VPWR _6025_/B sky130_fd_sc_hd__nor2_1
X_3219_ _6965_/Q VGND VGND VPWR VPWR _3219_/Y sky130_fd_sc_hd__inv_2
X_4199_ _4199_/A0 _4235_/A0 _4203_/S VGND VGND VPWR VPWR _6655_/D sky130_fd_sc_hd__mux2_1
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6909_ _7079_/CLK _6909_/D wire4044/X VGND VGND VPWR VPWR _6909_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire637 wire638/X VGND VGND VPWR VPWR _5464_/S sky130_fd_sc_hd__clkbuf_2
Xwire648 _5447_/S VGND VGND VPWR VPWR _5444_/S sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_length3955 wire3956/X VGND VGND VPWR VPWR _6483_/SET_B sky130_fd_sc_hd__buf_2
XFILLER_108_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire659 _5418_/S VGND VGND VPWR VPWR _5420_/S sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_length3966 wire3965/A VGND VGND VPWR VPWR _6672_/SET_B sky130_fd_sc_hd__buf_2
Xmax_length3988 _7159_/RESET_B VGND VGND VPWR VPWR _7161_/RESET_B sky130_fd_sc_hd__clkbuf_2
XFILLER_40_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3210 _4477_/X VGND VGND VPWR VPWR _5105_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3221 _4491_/B VGND VGND VPWR VPWR _4871_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_123_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3232 wire3233/X VGND VGND VPWR VPWR _4709_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold290 _6624_/Q VGND VGND VPWR VPWR hold290/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3243 wire3244/X VGND VGND VPWR VPWR _5241_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3254 _4324_/B VGND VGND VPWR VPWR _5203_/B sky130_fd_sc_hd__clkbuf_2
Xwire2520 _6002_/Y VGND VGND VPWR VPWR _6176_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3265 _4318_/B VGND VGND VPWR VPWR _5502_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3276 _4300_/B VGND VGND VPWR VPWR _5403_/B sky130_fd_sc_hd__clkbuf_2
Xwire2542 _5998_/Y VGND VGND VPWR VPWR _6187_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire3287 wire3288/X VGND VGND VPWR VPWR _3888_/B sky130_fd_sc_hd__clkbuf_2
Xwire2553 _6023_/B VGND VGND VPWR VPWR _6308_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire3298 _6353_/S VGND VGND VPWR VPWR _6356_/S sky130_fd_sc_hd__clkbuf_2
Xwire2564 _5980_/Y VGND VGND VPWR VPWR _6027_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2575 _6022_/A VGND VGND VPWR VPWR _6183_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1830 _5761_/A1 VGND VGND VPWR VPWR _6116_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2586 _5858_/A2 VGND VGND VPWR VPWR _5814_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire1841 _6991_/Q VGND VGND VPWR VPWR _6153_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire2597 _4686_/X VGND VGND VPWR VPWR _4882_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1852 hold642/X VGND VGND VPWR VPWR _5416_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire1874 _6968_/Q VGND VGND VPWR VPWR wire1874/X sky130_fd_sc_hd__clkbuf_1
XFILLER_105_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1885 wire1886/X VGND VGND VPWR VPWR _3437_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire1896 _6947_/Q VGND VGND VPWR VPWR _6063_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_130 hold112/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3570_ _6116_/A1 _3570_/A2 wire870/X _3570_/B2 _3569_/X VGND VGND VPWR VPWR _3570_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_155_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5240_ _5240_/A0 hold40/X _5240_/S VGND VGND VPWR VPWR hold41/A sky130_fd_sc_hd__mux2_1
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5171_ _5171_/A _5171_/B VGND VGND VPWR VPWR _5172_/D sky130_fd_sc_hd__nor2_1
XFILLER_123_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4122_ _4122_/A0 hold248/X _4127_/S VGND VGND VPWR VPWR _6589_/D sky130_fd_sc_hd__mux2_1
X_4053_ _4111_/B _5241_/C _4052_/X _3308_/Y _5286_/B VGND VGND VPWR VPWR _4053_/X
+ sky130_fd_sc_hd__o221a_1
Xinput3 debug_out VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4955_ _4955_/A1 _4933_/Y _4828_/X VGND VGND VPWR VPWR _5123_/A sky130_fd_sc_hd__a21oi_1
X_3906_ _6019_/A _6018_/A VGND VGND VPWR VPWR _3906_/X sky130_fd_sc_hd__or2_1
XFILLER_177_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4886_ _5135_/A1 _4872_/B _4758_/Y _4504_/B VGND VGND VPWR VPWR _4887_/B sky130_fd_sc_hd__o211a_1
X_6625_ _7093_/CLK _6625_/D wire3959/X VGND VGND VPWR VPWR _6625_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_137_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3229 _4387_/Y VGND VGND VPWR VPWR _4760_/A1 sky130_fd_sc_hd__clkbuf_2
X_3837_ _3850_/B _6542_/Q _3836_/Y _6461_/Q VGND VGND VPWR VPWR _6461_/D sky130_fd_sc_hd__a31o_1
XFILLER_192_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6556_ _6989_/CLK _6556_/D wire3995/X VGND VGND VPWR VPWR _6556_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3768_ _6227_/A1 _4010_/A _4022_/A _6516_/Q VGND VGND VPWR VPWR _3768_/X sky130_fd_sc_hd__a22o_1
Xmax_length1805 _7005_/Q VGND VGND VPWR VPWR wire1804/A sky130_fd_sc_hd__clkbuf_1
XFILLER_192_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5507_ _5558_/A0 hold383/X _5507_/S VGND VGND VPWR VPWR _7070_/D sky130_fd_sc_hd__mux2_1
X_6487_ _7074_/CLK _6487_/D fanout3976/X VGND VGND VPWR VPWR _6487_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_145_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3699_ _6979_/Q _3699_/A2 _3699_/B1 _7208_/Q VGND VGND VPWR VPWR _3699_/X sky130_fd_sc_hd__a22o_1
XFILLER_10_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5438_ _5519_/A0 hold640/X _5438_/S VGND VGND VPWR VPWR _7009_/D sky130_fd_sc_hd__mux2_1
Xoutput340 _6649_/Q VGND VGND VPWR VPWR wb_dat_o[2] sky130_fd_sc_hd__buf_12
XFILLER_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5369_ _5396_/A1 hold210/X _5369_/S VGND VGND VPWR VPWR _6947_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7108_ _7132_/CLK _7108_/D fanout4077/X VGND VGND VPWR VPWR _7108_/Q sky130_fd_sc_hd__dfrtp_1
Xwire1104 _3473_/C1 VGND VGND VPWR VPWR _3409_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_101_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1115 _3358_/B1 VGND VGND VPWR VPWR _3557_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1126 _3334_/Y VGND VGND VPWR VPWR _3564_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1137 wire1138/X VGND VGND VPWR VPWR _3716_/A2 sky130_fd_sc_hd__clkbuf_1
X_7039_ _7133_/CLK _7039_/D fanout4073/X VGND VGND VPWR VPWR _7039_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_101_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1159 _3423_/B1 VGND VGND VPWR VPWR _3557_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire401 _4925_/X VGND VGND VPWR VPWR wire401/X sky130_fd_sc_hd__clkbuf_1
XFILLER_129_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire412 _4070_/X VGND VGND VPWR VPWR wire412/X sky130_fd_sc_hd__clkbuf_1
XFILLER_168_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire423 _3631_/X VGND VGND VPWR VPWR _3632_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire434 _3524_/X VGND VGND VPWR VPWR _3542_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_128_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire445 wire446/X VGND VGND VPWR VPWR wire445/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire456 wire457/X VGND VGND VPWR VPWR wire456/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire467 _5588_/S VGND VGND VPWR VPWR _5587_/S sky130_fd_sc_hd__clkbuf_1
Xwire478 _5553_/Y VGND VGND VPWR VPWR wire478/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire489 _5322_/X VGND VGND VPWR VPWR _5327_/S sky130_fd_sc_hd__clkbuf_1
XFILLER_124_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_618 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire3051 _5671_/X VGND VGND VPWR VPWR wire3051/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3062 _5897_/B1 VGND VGND VPWR VPWR _5956_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire3073 _5667_/X VGND VGND VPWR VPWR wire3073/X sky130_fd_sc_hd__clkbuf_1
Xwire3084 _5805_/B1 VGND VGND VPWR VPWR _5735_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3095 _5759_/A2 VGND VGND VPWR VPWR _5788_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire2350 _6567_/Q VGND VGND VPWR VPWR wire2350/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2361 wire2362/X VGND VGND VPWR VPWR _3671_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire2372 _6530_/Q VGND VGND VPWR VPWR _3508_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_93_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2383 _6527_/Q VGND VGND VPWR VPWR wire2383/X sky130_fd_sc_hd__clkbuf_1
XFILLER_93_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2394 _4024_/A0 VGND VGND VPWR VPWR wire2394/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1660 _6124_/A1 VGND VGND VPWR VPWR wire1660/X sky130_fd_sc_hd__clkbuf_1
Xwire1671 _5483_/A1 VGND VGND VPWR VPWR _5848_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire1682 _7046_/Q VGND VGND VPWR VPWR _6138_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire1693 wire1694/X VGND VGND VPWR VPWR wire1693/X sky130_fd_sc_hd__clkbuf_1
XFILLER_46_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4740_ _4931_/B _4742_/C VGND VGND VPWR VPWR _4740_/Y sky130_fd_sc_hd__nand2_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4671_ _4672_/A _4686_/B VGND VGND VPWR VPWR _4671_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6410_ _6432_/A _6437_/B VGND VGND VPWR VPWR _6410_/X sky130_fd_sc_hd__and2_1
X_3622_ _6728_/Q _4276_/A _3616_/X wire426/X _3621_/X VGND VGND VPWR VPWR _3633_/B
+ sky130_fd_sc_hd__a2111o_1
X_6341_ _6341_/A _6341_/B _6341_/C _6341_/D VGND VGND VPWR VPWR _6341_/X sky130_fd_sc_hd__or4_1
X_3553_ _3553_/A1 _3553_/A2 _4282_/A _6303_/A1 VGND VGND VPWR VPWR _3553_/X sky130_fd_sc_hd__a22o_1
Xwire990 wire990/A VGND VGND VPWR VPWR _6217_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_143_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6272_ _6533_/Q _6272_/B VGND VGND VPWR VPWR _6272_/X sky130_fd_sc_hd__and2_1
XFILLER_170_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3484_ _3484_/A _3484_/B _3484_/C _3484_/D VGND VGND VPWR VPWR _3543_/B sky130_fd_sc_hd__or4_1
XFILLER_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5223_ _5223_/A _5223_/B VGND VGND VPWR VPWR _5224_/S sky130_fd_sc_hd__nand2_1
XFILLER_170_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5154_ _5076_/B _4630_/A _5017_/A VGND VGND VPWR VPWR _5155_/C sky130_fd_sc_hd__a21oi_1
X_4105_ _4247_/A0 hold614/X _4108_/S VGND VGND VPWR VPWR _6574_/D sky130_fd_sc_hd__mux2_1
XFILLER_111_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5085_ _4420_/A _5106_/A _5109_/C _5107_/B _5153_/B VGND VGND VPWR VPWR _5086_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_56_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4036_ hold664/X _4122_/A0 _4039_/S VGND VGND VPWR VPWR _6527_/D sky130_fd_sc_hd__mux2_1
XFILLER_71_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5987_ _7155_/Q _7156_/Q VGND VGND VPWR VPWR _6040_/C sky130_fd_sc_hd__and2b_1
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4938_ _4938_/A1 _4428_/B _4957_/B _5177_/B _4506_/Y VGND VGND VPWR VPWR _4939_/C
+ sky130_fd_sc_hd__a311o_1
XFILLER_178_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_30 _3464_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmax_length3015 _5757_/A2 VGND VGND VPWR VPWR _5776_/A2 sky130_fd_sc_hd__clkbuf_1
X_4869_ _4930_/C _4868_/X _4930_/A VGND VGND VPWR VPWR _4928_/B sky130_fd_sc_hd__o21ba_1
XANTENNA_41 wire1319/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_52 wire1456/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_63 _3387_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6608_ _7091_/CLK _6608_/D wire4026/A VGND VGND VPWR VPWR _6608_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA_74 _3691_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_85 _6204_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_96 _5776_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6539_ _7090_/CLK _6539_/D wire3943/A VGND VGND VPWR VPWR _6539_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput181 _3219_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[15] sky130_fd_sc_hd__buf_12
Xoutput192 _3209_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[25] sky130_fd_sc_hd__buf_12
XFILLER_121_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length4294 _4566_/A VGND VGND VPWR VPWR _4569_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_183_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_551 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2180 _6746_/Q VGND VGND VPWR VPWR _3758_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2191 _6740_/Q VGND VGND VPWR VPWR wire2191/X sky130_fd_sc_hd__clkbuf_1
XFILLER_93_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1490 wire1491/X VGND VGND VPWR VPWR wire1490/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5910_ _6286_/A1 _5910_/A2 _5909_/X VGND VGND VPWR VPWR _5910_/X sky130_fd_sc_hd__a21o_1
X_6890_ _7127_/CLK _6890_/D fanout4054/A VGND VGND VPWR VPWR _6890_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5841_ _6205_/A1 _5841_/A2 _5841_/B1 _6210_/B2 VGND VGND VPWR VPWR _5841_/X sky130_fd_sc_hd__a22o_1
X_5772_ _6120_/A1 _5772_/A2 wire994/X _5771_/X _6120_/C1 VGND VGND VPWR VPWR _5772_/X
+ sky130_fd_sc_hd__o221a_1
X_4723_ _4650_/Y _4722_/X _6362_/A _4648_/Y VGND VGND VPWR VPWR _4723_/X sky130_fd_sc_hd__a211o_1
XFILLER_175_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4654_ _4654_/A _4654_/B _4390_/A VGND VGND VPWR VPWR _4654_/X sky130_fd_sc_hd__or3b_1
Xinput50 mgmt_gpio_in[22] VGND VGND VPWR VPWR input50/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3605_ _6092_/B2 _3605_/A2 _3605_/B1 _6844_/Q VGND VGND VPWR VPWR _3605_/X sky130_fd_sc_hd__a22o_1
Xinput61 mgmt_gpio_in[32] VGND VGND VPWR VPWR input61/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4585_ _4588_/A _4935_/A _4412_/A1 VGND VGND VPWR VPWR _4585_/X sky130_fd_sc_hd__or3b_1
Xinput72 mgmt_gpio_in[9] VGND VGND VPWR VPWR input72/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput83 spimemio_flash_clk VGND VGND VPWR VPWR input83/X sky130_fd_sc_hd__clkbuf_1
Xinput94 uart_enabled VGND VGND VPWR VPWR _3957_/B sky130_fd_sc_hd__clkbuf_1
X_6324_ _6324_/A1 _6324_/A2 _6324_/B1 _6765_/Q _6323_/X VGND VGND VPWR VPWR _6331_/A
+ sky130_fd_sc_hd__a221o_1
X_3536_ _3536_/A _3536_/B VGND VGND VPWR VPWR _3536_/Y sky130_fd_sc_hd__nor2_1
XFILLER_131_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6255_ _6255_/A1 _6255_/A2 _6255_/B1 _7208_/Q VGND VGND VPWR VPWR _6255_/X sky130_fd_sc_hd__a22o_1
X_3467_ _6325_/B2 _3574_/A2 _4210_/A _6333_/B2 _3464_/X VGND VGND VPWR VPWR _3468_/D
+ sky130_fd_sc_hd__a221o_1
X_5206_ hold701/X _5206_/A1 _5209_/S VGND VGND VPWR VPWR _6807_/D sky130_fd_sc_hd__mux2_1
X_6186_ _6186_/A1 _6186_/A2 _6186_/B1 _7072_/Q VGND VGND VPWR VPWR _6186_/X sky130_fd_sc_hd__a22o_1
X_3398_ _7000_/Q _5421_/A _3425_/B1 _3398_/B2 VGND VGND VPWR VPWR _3398_/X sky130_fd_sc_hd__a22o_1
XFILLER_111_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5137_ _5148_/A _5151_/B _5148_/D _5137_/D VGND VGND VPWR VPWR _5138_/B sky130_fd_sc_hd__or4_1
XFILLER_57_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5068_ _5068_/A _5068_/B VGND VGND VPWR VPWR _5068_/X sky130_fd_sc_hd__or2_1
XFILLER_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4019_ _6395_/A0 hold262/X _4021_/S VGND VGND VPWR VPWR _6513_/D sky130_fd_sc_hd__mux2_1
XFILLER_37_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold108 hold108/A VGND VGND VPWR VPWR hold108/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_156_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold119 _7201_/Q VGND VGND VPWR VPWR hold119/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_125_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4370_ _4745_/A _4497_/A _4228_/C VGND VGND VPWR VPWR _4930_/A sky130_fd_sc_hd__o21ai_1
XFILLER_98_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3321_ _3510_/A _3674_/B VGND VGND VPWR VPWR _3321_/Y sky130_fd_sc_hd__nor2_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _6040_/A _6040_/B _6040_/C VGND VGND VPWR VPWR _6040_/X sky130_fd_sc_hd__and3_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _6468_/Q _3252_/B VGND VGND VPWR VPWR _3818_/A sky130_fd_sc_hd__nand2_1
XFILLER_39_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6942_ _7131_/CLK _6942_/D wire4058/A VGND VGND VPWR VPWR _6942_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6873_ _7133_/CLK hold86/X fanout4073/X VGND VGND VPWR VPWR _6873_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_62_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5824_ _5824_/A1 _5824_/A2 _5824_/B1 _6188_/B2 _5823_/X VGND VGND VPWR VPWR _5825_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5755_ _5755_/A1 _5808_/B1 _5755_/B1 _5755_/B2 VGND VGND VPWR VPWR _5755_/X sky130_fd_sc_hd__a22o_1
XFILLER_175_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4706_ _4707_/A _4683_/B _4863_/B _4705_/X VGND VGND VPWR VPWR _4708_/C sky130_fd_sc_hd__o211a_1
X_5686_ _7152_/Q _5700_/C _5703_/C VGND VGND VPWR VPWR _5686_/X sky130_fd_sc_hd__and3_1
XFILLER_108_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4637_ _4637_/A1 _4752_/B _4799_/B1 _5027_/A _4636_/X VGND VGND VPWR VPWR _4642_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_190_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire4307 input11/X VGND VGND VPWR VPWR wire4307/X sky130_fd_sc_hd__clkbuf_1
XFILLER_163_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold620 _6758_/Q VGND VGND VPWR VPWR hold620/X sky130_fd_sc_hd__dlygate4sd3_1
X_4568_ _4666_/B _4688_/B VGND VGND VPWR VPWR _4568_/X sky130_fd_sc_hd__or2_1
Xhold631 _6480_/Q VGND VGND VPWR VPWR hold631/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold642 _6989_/Q VGND VGND VPWR VPWR hold642/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold653 _6865_/Q VGND VGND VPWR VPWR hold653/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3606 hold38/A VGND VGND VPWR VPWR _5468_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
X_6307_ _6534_/Q _6307_/A2 _6302_/X _6304_/X _6306_/X VGND VGND VPWR VPWR _6307_/X
+ sky130_fd_sc_hd__a2111o_1
Xhold664 _6527_/Q VGND VGND VPWR VPWR hold664/X sky130_fd_sc_hd__dlygate4sd3_1
X_3519_ _3531_/A _3519_/B VGND VGND VPWR VPWR _3519_/Y sky130_fd_sc_hd__nor2_1
Xwire3617 wire3618/X VGND VGND VPWR VPWR wire3617/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold675 _7023_/Q VGND VGND VPWR VPWR hold675/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3628 wire3628/A VGND VGND VPWR VPWR _5212_/C sky130_fd_sc_hd__clkbuf_2
Xhold686 _7016_/Q VGND VGND VPWR VPWR hold686/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4499_ _4420_/A _4450_/A _4498_/X _4489_/X _4484_/X VGND VGND VPWR VPWR _4503_/D
+ sky130_fd_sc_hd__o311a_1
Xhold697 _6530_/Q VGND VGND VPWR VPWR hold697/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3639 _5251_/A1 VGND VGND VPWR VPWR _5536_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_104_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2905 _5842_/B1 VGND VGND VPWR VPWR _5800_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
X_6238_ _6238_/A1 _6238_/A2 _6313_/B1 _6238_/B2 _6237_/X VGND VGND VPWR VPWR _6241_/C
+ sky130_fd_sc_hd__a221o_1
Xwire2916 _5820_/B1 VGND VGND VPWR VPWR _5840_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_76_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2938 _5783_/A2 VGND VGND VPWR VPWR _5744_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_103_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2949 wire2949/A VGND VGND VPWR VPWR _5812_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_134_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ _6169_/A1 wire980/X _6156_/X _6168_/X _6169_/C1 VGND VGND VPWR VPWR _6169_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_43_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7088_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_58_csclk _7117_/CLK VGND VGND VPWR VPWR _7109_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_193_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3870_ _6471_/Q _6445_/Q _3839_/B VGND VGND VPWR VPWR _3870_/X sky130_fd_sc_hd__a21o_1
XFILLER_71_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5540_ hold557/X _5540_/A1 _5543_/S VGND VGND VPWR VPWR _7099_/D sky130_fd_sc_hd__mux2_1
XFILLER_192_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5471_ hold615/X _5558_/A0 _5471_/S VGND VGND VPWR VPWR _7038_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_646 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7210_ _7210_/CLK _7210_/D fanout3952/X VGND VGND VPWR VPWR _7210_/Q sky130_fd_sc_hd__dfrtp_1
X_4422_ _4758_/A _4758_/C VGND VGND VPWR VPWR _4441_/A sky130_fd_sc_hd__nand2_1
XFILLER_145_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7141_ _7141_/CLK _7141_/D _7141_/RESET_B VGND VGND VPWR VPWR _7141_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4353_ _4412_/A1 _4359_/B _4379_/A VGND VGND VPWR VPWR _4354_/B sky130_fd_sc_hd__a21o_1
X_3304_ _3344_/A _3528_/B VGND VGND VPWR VPWR _3304_/Y sky130_fd_sc_hd__nor2_1
X_7072_ _7072_/CLK _7072_/D wire4001/X VGND VGND VPWR VPWR _7072_/Q sky130_fd_sc_hd__dfrtp_1
X_4284_ _4284_/A0 hold380/X _4287_/S VGND VGND VPWR VPWR _6732_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6023_ _6023_/A _6023_/B _6023_/C _6023_/D VGND VGND VPWR VPWR _6026_/B sky130_fd_sc_hd__or4_1
X_3235_ _7152_/Q VGND VGND VPWR VPWR _3235_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6925_ _6973_/CLK _6925_/D fanout4078/X VGND VGND VPWR VPWR _6925_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6856_ _7017_/CLK _6856_/D fanout4077/X VGND VGND VPWR VPWR hold98/A sky130_fd_sc_hd__dfrtp_1
XFILLER_120_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5807_ _6147_/B2 _5807_/A2 _5807_/B1 _6967_/Q VGND VGND VPWR VPWR _5807_/X sky130_fd_sc_hd__a22o_1
X_3999_ hold571/X _3999_/A1 _4000_/S VGND VGND VPWR VPWR _6496_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6787_ _3487_/B2 _6787_/D _6438_/X VGND VGND VPWR VPWR _6787_/Q sky130_fd_sc_hd__dfrtn_1
Xwire808 _3519_/Y VGND VGND VPWR VPWR wire808/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_167_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire819 wire820/X VGND VGND VPWR VPWR _4300_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5738_ _6087_/A1 _5738_/A2 _5738_/B1 _5738_/B2 VGND VGND VPWR VPWR _5738_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5669_ _7150_/Q _7151_/Q VGND VGND VPWR VPWR _5699_/C sky130_fd_sc_hd__and2b_1
XFILLER_135_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout3308 _5021_/B VGND VGND VPWR VPWR _5074_/A2 sky130_fd_sc_hd__buf_6
Xwire4104 input70/X VGND VGND VPWR VPWR _3359_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire4115 wire4116/X VGND VGND VPWR VPWR _3872_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire4126 wire4127/X VGND VGND VPWR VPWR _7214_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_123_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire4137 wire4138/X VGND VGND VPWR VPWR wire4137/X sky130_fd_sc_hd__clkbuf_1
Xhold450 _6803_/Q VGND VGND VPWR VPWR hold450/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 _6932_/Q VGND VGND VPWR VPWR hold461/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire4148 wire4149/X VGND VGND VPWR VPWR wire4148/X sky130_fd_sc_hd__clkbuf_1
Xwire3414 _5248_/A0 VGND VGND VPWR VPWR _5527_/A0 sky130_fd_sc_hd__clkbuf_1
Xhold472 _6793_/Q VGND VGND VPWR VPWR hold472/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire4159 wire4160/X VGND VGND VPWR VPWR _3616_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire3425 _5247_/A0 VGND VGND VPWR VPWR _5550_/A0 sky130_fd_sc_hd__clkbuf_1
Xhold483 _6554_/Q VGND VGND VPWR VPWR hold483/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3436 wire3437/X VGND VGND VPWR VPWR wire3436/X sky130_fd_sc_hd__clkbuf_1
Xwire3447 _4134_/A1 VGND VGND VPWR VPWR _5198_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold494 _6894_/Q VGND VGND VPWR VPWR hold494/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2702 _6203_/B1 VGND VGND VPWR VPWR _6153_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2713 _6154_/A2 VGND VGND VPWR VPWR _6131_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3469 _5576_/A0 VGND VGND VPWR VPWR _5585_/A0 sky130_fd_sc_hd__clkbuf_2
Xwire2724 wire2725/X VGND VGND VPWR VPWR _6159_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire2735 _6206_/A2 VGND VGND VPWR VPWR _6190_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire2746 _6174_/B1 VGND VGND VPWR VPWR _6166_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2757 _6211_/A2 VGND VGND VPWR VPWR _6160_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire2768 _6000_/X VGND VGND VPWR VPWR _6186_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_161_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2779 _6024_/B VGND VGND VPWR VPWR _5993_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_180_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_79_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3970 wire3970/A VGND VGND VPWR VPWR wire3970/X sky130_fd_sc_hd__clkbuf_2
Xwire3981 wire3981/A VGND VGND VPWR VPWR wire3981/X sky130_fd_sc_hd__buf_2
Xwire3992 wire3992/A VGND VGND VPWR VPWR wire3992/X sky130_fd_sc_hd__buf_2
XFILLER_110_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4971_ _4971_/A _4971_/B VGND VGND VPWR VPWR _4971_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6710_ _7208_/CLK _6710_/D wire4026/X VGND VGND VPWR VPWR _6710_/Q sky130_fd_sc_hd__dfrtp_1
X_3922_ _3199_/Y _3922_/A1 _3958_/B VGND VGND VPWR VPWR _3922_/X sky130_fd_sc_hd__mux2_1
X_3853_ _6453_/Q _3853_/B VGND VGND VPWR VPWR _3858_/B sky130_fd_sc_hd__nor2_1
X_6641_ _7206_/CLK _6641_/D VGND VGND VPWR VPWR _6641_/Q sky130_fd_sc_hd__dfxtp_1
X_6572_ _6973_/CLK _6572_/D _7087_/RESET_B VGND VGND VPWR VPWR _6572_/Q sky130_fd_sc_hd__dfrtp_1
X_3784_ _3784_/A1 _3331_/Y _3784_/B1 _3784_/B2 wire738/X VGND VGND VPWR VPWR _3788_/B
+ sky130_fd_sc_hd__a221o_1
X_5523_ _5523_/A0 hold544/X _5523_/S VGND VGND VPWR VPWR _7084_/D sky130_fd_sc_hd__mux2_1
XFILLER_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5454_ _5454_/A0 hold675/X _5455_/S VGND VGND VPWR VPWR _7023_/D sky130_fd_sc_hd__mux2_1
X_4405_ _4560_/A _4731_/C _4731_/B VGND VGND VPWR VPWR _4742_/B sky130_fd_sc_hd__and3_1
XFILLER_132_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5385_ _5385_/A _5520_/B VGND VGND VPWR VPWR _5393_/S sky130_fd_sc_hd__nand2_1
X_4336_ _4390_/A _4390_/C _4390_/D VGND VGND VPWR VPWR _4547_/A sky130_fd_sc_hd__or3_1
X_7124_ _7124_/CLK _7124_/D wire4049/A VGND VGND VPWR VPWR _7124_/Q sky130_fd_sc_hd__dfrtp_1
Xwire2009 _6891_/Q VGND VGND VPWR VPWR _6062_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7055_ _7133_/CLK _7055_/D _7134_/RESET_B VGND VGND VPWR VPWR _7055_/Q sky130_fd_sc_hd__dfrtp_1
X_4267_ hold638/X _5469_/A1 _4268_/S VGND VGND VPWR VPWR _6718_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1308 _6275_/X VGND VGND VPWR VPWR _6280_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_86_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1319 wire1320/X VGND VGND VPWR VPWR wire1319/X sky130_fd_sc_hd__clkbuf_1
X_6006_ _6038_/A _6006_/B VGND VGND VPWR VPWR _6006_/Y sky130_fd_sc_hd__nor2_1
X_3218_ _6973_/Q VGND VGND VPWR VPWR _3218_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4198_ _4198_/A _4234_/B VGND VGND VPWR VPWR _4203_/S sky130_fd_sc_hd__and2_2
XFILLER_39_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6908_ _7135_/CLK _6908_/D _6404_/A VGND VGND VPWR VPWR _6908_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_24_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6839_ _7084_/CLK _6839_/D wire4056/A VGND VGND VPWR VPWR _6839_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire605 wire605/A VGND VGND VPWR VPWR _5506_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_183_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire616 _5490_/S VGND VGND VPWR VPWR _5487_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire638 wire639/X VGND VGND VPWR VPWR wire638/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire649 _5439_/Y VGND VGND VPWR VPWR _5447_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_109_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length3989 fanout3986/X VGND VGND VPWR VPWR _7159_/RESET_B sky130_fd_sc_hd__clkbuf_2
XFILLER_136_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3200 _4971_/A VGND VGND VPWR VPWR _4798_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3211 _4670_/B VGND VGND VPWR VPWR _4672_/A sky130_fd_sc_hd__clkbuf_2
Xhold280 _7014_/Q VGND VGND VPWR VPWR hold280/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3233 _4367_/Y VGND VGND VPWR VPWR wire3233/X sky130_fd_sc_hd__clkbuf_1
Xhold291 _6538_/Q VGND VGND VPWR VPWR hold291/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3244 wire3245/X VGND VGND VPWR VPWR wire3244/X sky130_fd_sc_hd__clkbuf_1
Xwire3255 _5535_/B VGND VGND VPWR VPWR _5511_/B sky130_fd_sc_hd__clkbuf_2
Xwire2510 _6202_/B1 VGND VGND VPWR VPWR _6151_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire2521 _6326_/A2 VGND VGND VPWR VPWR _6286_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2532 _6001_/Y VGND VGND VPWR VPWR _6185_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire3277 _4270_/B VGND VGND VPWR VPWR _4300_/B sky130_fd_sc_hd__clkbuf_2
Xwire2543 _6277_/A2 VGND VGND VPWR VPWR _6334_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3288 wire3289/X VGND VGND VPWR VPWR wire3288/X sky130_fd_sc_hd__clkbuf_1
Xwire3299 _4654_/X VGND VGND VPWR VPWR _5021_/C sky130_fd_sc_hd__clkbuf_2
Xwire2554 _6258_/A2 VGND VGND VPWR VPWR _5985_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire1820 _7001_/Q VGND VGND VPWR VPWR wire1820/X sky130_fd_sc_hd__clkbuf_1
XFILLER_93_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2565 _6141_/A2 VGND VGND VPWR VPWR _6065_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire1831 wire1832/X VGND VGND VPWR VPWR _5761_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2576 _6075_/A2 VGND VGND VPWR VPWR _6197_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2587 _5793_/A2 VGND VGND VPWR VPWR _5729_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire2598 _4672_/X VGND VGND VPWR VPWR _5128_/B sky130_fd_sc_hd__clkbuf_1
Xwire1853 wire1853/A VGND VGND VPWR VPWR _6087_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_92_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1864 _6973_/Q VGND VGND VPWR VPWR _6116_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire1875 wire1876/X VGND VGND VPWR VPWR _3441_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_45_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1886 _6959_/Q VGND VGND VPWR VPWR wire1886/X sky130_fd_sc_hd__clkbuf_1
XFILLER_73_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1897 _5985_/A1 VGND VGND VPWR VPWR _3754_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_18_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_120 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_131 input63/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5170_ _5170_/A _5170_/B _5170_/C _5169_/X VGND VGND VPWR VPWR _5171_/B sky130_fd_sc_hd__or4b_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4121_ _4130_/A1 hold241/X _4127_/S VGND VGND VPWR VPWR _4121_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4052_ _5241_/C _4052_/B VGND VGND VPWR VPWR _4052_/X sky130_fd_sc_hd__and2b_1
XFILLER_83_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput4 mask_rev_in[0] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4954_ _5158_/B _4954_/B _4954_/C _5158_/C VGND VGND VPWR VPWR _4960_/B sky130_fd_sc_hd__or4_1
XFILLER_189_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3905_ _6014_/A _6000_/A VGND VGND VPWR VPWR _6018_/A sky130_fd_sc_hd__nand2_1
XFILLER_32_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4885_ _5039_/A _4885_/B _4885_/C _4885_/D VGND VGND VPWR VPWR _4885_/X sky130_fd_sc_hd__or4_1
XFILLER_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6624_ _7093_/CLK _6624_/D wire3959/X VGND VGND VPWR VPWR _6624_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3836_ _3850_/A _6541_/Q _6545_/Q VGND VGND VPWR VPWR _3836_/Y sky130_fd_sc_hd__nor3_1
XFILLER_165_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3767_ _6766_/Q _3767_/A2 _3767_/B1 _5877_/B2 VGND VGND VPWR VPWR _3767_/X sky130_fd_sc_hd__a22o_1
X_6555_ _6811_/CLK _6555_/D _6430_/A VGND VGND VPWR VPWR _6555_/Q sky130_fd_sc_hd__dfrtp_1
X_5506_ _5506_/A0 hold506/X _5506_/S VGND VGND VPWR VPWR _7069_/D sky130_fd_sc_hd__mux2_1
X_6486_ _6824_/CLK _6486_/D wire3956/X VGND VGND VPWR VPWR _6486_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_10_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3698_ _5711_/B2 _3698_/A2 _3698_/B1 _6055_/A1 _3697_/X VGND VGND VPWR VPWR _3701_/C
+ sky130_fd_sc_hd__a221o_1
X_5437_ _5437_/A0 hold671/X _5438_/S VGND VGND VPWR VPWR _7008_/D sky130_fd_sc_hd__mux2_1
Xoutput330 wire3768/X VGND VGND VPWR VPWR wb_dat_o[20] sky130_fd_sc_hd__buf_12
XFILLER_161_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput341 _7195_/Q VGND VGND VPWR VPWR wb_dat_o[30] sky130_fd_sc_hd__buf_12
XFILLER_160_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5368_ _5581_/A0 hold319/X _5369_/S VGND VGND VPWR VPWR _6946_/D sky130_fd_sc_hd__mux2_1
XFILLER_126_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7107_ _7130_/CLK _7107_/D wire4061/X VGND VGND VPWR VPWR _7107_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4319_ hold345/X _5503_/A0 _4323_/S VGND VGND VPWR VPWR _6761_/D sky130_fd_sc_hd__mux2_1
X_5299_ _5584_/A0 hold193/X _5303_/S VGND VGND VPWR VPWR _6885_/D sky130_fd_sc_hd__mux2_1
Xwire1116 _3486_/A2 VGND VGND VPWR VPWR _3358_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
X_7038_ _7115_/CLK _7038_/D wire3980/X VGND VGND VPWR VPWR _7038_/Q sky130_fd_sc_hd__dfrtp_1
Xwire1138 _3634_/A2 VGND VGND VPWR VPWR wire1138/X sky130_fd_sc_hd__clkbuf_1
Xwire1149 _3561_/A2 VGND VGND VPWR VPWR _3654_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_74_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire413 _4069_/S VGND VGND VPWR VPWR _4061_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_11_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire424 wire425/X VGND VGND VPWR VPWR _3627_/D sky130_fd_sc_hd__clkbuf_1
Xwire435 _3506_/X VGND VGND VPWR VPWR _3515_/B sky130_fd_sc_hd__clkbuf_1
Xwire446 wire447/X VGND VGND VPWR VPWR wire446/X sky130_fd_sc_hd__clkbuf_1
Xwire457 wire458/X VGND VGND VPWR VPWR wire457/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire479 _5561_/S VGND VGND VPWR VPWR _5557_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3030 _5680_/A2 VGND VGND VPWR VPWR _5784_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire3041 _5778_/A2 VGND VGND VPWR VPWR _5955_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_78_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3052 _5852_/A2 VGND VGND VPWR VPWR _5797_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire3063 _5736_/A2 VGND VGND VPWR VPWR _5897_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire2340 _6599_/Q VGND VGND VPWR VPWR _6317_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3085 _5832_/A2 VGND VGND VPWR VPWR _5805_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2351 wire2352/X VGND VGND VPWR VPWR _3928_/A0 sky130_fd_sc_hd__clkbuf_1
Xwire3096 _5848_/A2 VGND VGND VPWR VPWR _5759_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2362 _6537_/Q VGND VGND VPWR VPWR wire2362/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2373 _5952_/A1 VGND VGND VPWR VPWR _6339_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire2384 _6237_/B2 VGND VGND VPWR VPWR _3784_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_19_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1650 _5673_/A1 VGND VGND VPWR VPWR wire1650/X sky130_fd_sc_hd__clkbuf_1
Xwire1661 _7054_/Q VGND VGND VPWR VPWR _6124_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1683 _6103_/B2 VGND VGND VPWR VPWR _5756_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire1694 _5680_/B2 VGND VGND VPWR VPWR wire1694/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4670_ _4739_/A _4670_/B VGND VGND VPWR VPWR _4670_/Y sky130_fd_sc_hd__nor2_1
XFILLER_159_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3621_ _3621_/A1 _3672_/B1 hold64/A _3621_/B2 wire773/X VGND VGND VPWR VPWR _3621_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3552_ _7098_/Q _5535_/A _5214_/A _5216_/A1 VGND VGND VPWR VPWR _3552_/X sky130_fd_sc_hd__a22o_1
X_6340_ _6340_/A1 _6340_/A2 _6337_/X _6340_/C1 VGND VGND VPWR VPWR _6341_/D sky130_fd_sc_hd__a211o_1
Xwire980 wire981/X VGND VGND VPWR VPWR wire980/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_700 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6271_ _6728_/Q _6320_/A2 _6320_/B1 _6271_/B2 VGND VGND VPWR VPWR _6271_/X sky130_fd_sc_hd__a22o_1
XFILLER_142_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3483_ _3483_/A1 _3292_/Y _3656_/B1 _3483_/B2 wire822/X VGND VGND VPWR VPWR _3484_/D
+ sky130_fd_sc_hd__a221o_1
X_5222_ _3711_/A _3379_/B _5422_/A0 _5221_/X _5203_/B VGND VGND VPWR VPWR _6819_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_88_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5153_ _5153_/A _5153_/B _5152_/X VGND VGND VPWR VPWR _5153_/X sky130_fd_sc_hd__or3b_1
XFILLER_111_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4104_ _4104_/A _5580_/B VGND VGND VPWR VPWR _4104_/Y sky130_fd_sc_hd__nand2_1
XFILLER_84_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5084_ _5108_/A _5027_/B _5108_/B _5152_/A1 _4909_/Y VGND VGND VPWR VPWR _5153_/B
+ sky130_fd_sc_hd__o221ai_2
X_4035_ hold634/X _4130_/A1 _4039_/S VGND VGND VPWR VPWR _6526_/D sky130_fd_sc_hd__mux2_1
XFILLER_2_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5986_ _5986_/A1 _6075_/A2 _6075_/B1 _5986_/B2 _5985_/X VGND VGND VPWR VPWR _6045_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4937_ _4955_/A1 _4957_/B _4864_/D VGND VGND VPWR VPWR _5124_/C sky130_fd_sc_hd__a21o_1
XFILLER_33_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_20 _3701_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_31 _3692_/C1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4868_ _4868_/A _5068_/A _4868_/C _4868_/D VGND VGND VPWR VPWR _4868_/X sky130_fd_sc_hd__or4_1
Xmax_length3016 _5856_/A2 VGND VGND VPWR VPWR _5757_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_42 wire1320/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_53 wire1476/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_64 wire1687/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6607_ _7208_/CLK _6607_/D wire4026/A VGND VGND VPWR VPWR _6607_/Q sky130_fd_sc_hd__dfrtp_2
X_3819_ _3818_/Y _6468_/Q _3828_/S VGND VGND VPWR VPWR _6468_/D sky130_fd_sc_hd__mux2_1
XANTENNA_75 _3388_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_86 _6213_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4799_ _4753_/B _4805_/B2 _4799_/B1 _4655_/B VGND VGND VPWR VPWR _4799_/X sky130_fd_sc_hd__o22a_1
XANTENNA_97 _5776_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6538_ _7090_/CLK _6538_/D wire3948/X VGND VGND VPWR VPWR _6538_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_146_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6469_ _3487_/B2 _6469_/D _6424_/X VGND VGND VPWR VPWR hold60/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput171 _3959_/X VGND VGND VPWR VPWR debug_in sky130_fd_sc_hd__buf_12
XFILLER_121_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput182 _3218_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[16] sky130_fd_sc_hd__buf_12
Xoutput193 _3208_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[26] sky130_fd_sc_hd__buf_12
XFILLER_121_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_663 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2170 wire2171/X VGND VGND VPWR VPWR _3549_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_78_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2181 _6745_/Q VGND VGND VPWR VPWR _6321_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_66_558 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1480 wire1481/X VGND VGND VPWR VPWR wire1480/X sky130_fd_sc_hd__clkbuf_2
Xwire1491 wire1492/X VGND VGND VPWR VPWR wire1491/X sky130_fd_sc_hd__clkbuf_1
XFILLER_47_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5840_ _6211_/A1 _5840_/A2 _5840_/B1 _6201_/A1 _5839_/X VGND VGND VPWR VPWR _5847_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5771_ _5771_/A _5771_/B _5771_/C VGND VGND VPWR VPWR _5771_/X sky130_fd_sc_hd__or3_1
X_4722_ _5130_/A _4722_/B _4722_/C VGND VGND VPWR VPWR _4722_/X sky130_fd_sc_hd__or3_1
XFILLER_159_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4653_ _4693_/A _4694_/A _4653_/C VGND VGND VPWR VPWR _4653_/X sky130_fd_sc_hd__or3_1
XFILLER_147_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput40 mgmt_gpio_in[13] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__clkbuf_1
X_3604_ _7137_/Q wire953/X wire795/A _3604_/B2 VGND VGND VPWR VPWR _3604_/X sky130_fd_sc_hd__a22o_1
Xinput51 mgmt_gpio_in[23] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__clkbuf_1
Xinput62 mgmt_gpio_in[33] VGND VGND VPWR VPWR input62/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4584_ _5105_/A1 _5105_/A2 _4842_/A1 _4623_/A VGND VGND VPWR VPWR _4584_/X sky130_fd_sc_hd__o22a_1
Xinput73 pad_flash_io0_di VGND VGND VPWR VPWR _3952_/B sky130_fd_sc_hd__clkbuf_1
Xinput84 spimemio_flash_csb VGND VGND VPWR VPWR input84/X sky130_fd_sc_hd__clkbuf_1
Xinput95 usr1_vcc_pwrgood VGND VGND VPWR VPWR input95/X sky130_fd_sc_hd__clkbuf_1
X_6323_ _6323_/A1 _6323_/A2 _6323_/B1 _6323_/B2 VGND VGND VPWR VPWR _6323_/X sky130_fd_sc_hd__a22o_1
X_3535_ _3535_/A1 _3325_/Y _3665_/B1 _3535_/B2 VGND VGND VPWR VPWR _3535_/X sky130_fd_sc_hd__a22o_1
XFILLER_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6254_ _6254_/A1 _6304_/A2 _6304_/B1 _6757_/Q _6253_/X VGND VGND VPWR VPWR _6254_/X
+ sky130_fd_sc_hd__a221o_1
X_3466_ _3466_/A _3536_/B VGND VGND VPWR VPWR _3466_/Y sky130_fd_sc_hd__nor2_1
XFILLER_131_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5205_ _5205_/A _5511_/B VGND VGND VPWR VPWR _5209_/S sky130_fd_sc_hd__and2_1
XFILLER_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3397_ _7117_/Q wire961/X _5268_/A _6185_/B2 VGND VGND VPWR VPWR _3397_/X sky130_fd_sc_hd__a22o_1
X_6185_ _6185_/A1 _6185_/A2 _6185_/B1 _6185_/B2 _6184_/X VGND VGND VPWR VPWR _6192_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_97_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5136_ _5136_/A _5136_/B _4759_/Y VGND VGND VPWR VPWR _5137_/D sky130_fd_sc_hd__or3b_1
XFILLER_84_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5067_ _5067_/A _5067_/B _5067_/C VGND VGND VPWR VPWR _5069_/A sky130_fd_sc_hd__nor3_1
X_4018_ _4308_/A0 hold256/X _4021_/S VGND VGND VPWR VPWR _6512_/D sky130_fd_sc_hd__mux2_1
XFILLER_37_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5969_ _5969_/A1 _7173_/Q wire459/X VGND VGND VPWR VPWR _5969_/X sky130_fd_sc_hd__a21o_1
XFILLER_166_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length2112 _6818_/Q VGND VGND VPWR VPWR _3940_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_148_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xnet4299_2 _3487_/B2 VGND VGND VPWR VPWR _3941_/B sky130_fd_sc_hd__inv_2
XFILLER_156_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold109 _4117_/X VGND VGND VPWR VPWR _6585_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3320_ _3320_/A _3465_/B VGND VGND VPWR VPWR _3320_/Y sky130_fd_sc_hd__nor2_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _3941_/A hold25/X _3250_/Y VGND VGND VPWR VPWR hold26/A sky130_fd_sc_hd__o21ai_2
XFILLER_113_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6941_ _6973_/CLK _6941_/D fanout4078/X VGND VGND VPWR VPWR hold97/A sky130_fd_sc_hd__dfrtp_1
X_6872_ _7017_/CLK _6872_/D fanout4078/X VGND VGND VPWR VPWR _6872_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_179_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5823_ _5823_/A1 _5849_/A2 _5702_/X _6984_/Q VGND VGND VPWR VPWR _5823_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5754_ _6103_/A1 _5754_/A2 _5754_/B1 _5754_/B2 VGND VGND VPWR VPWR _5754_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4705_ _4704_/A _4707_/B _4703_/X _4704_/X VGND VGND VPWR VPWR _4705_/X sky130_fd_sc_hd__o211a_1
XFILLER_147_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5685_ _5693_/A _5705_/B _5699_/C VGND VGND VPWR VPWR _5685_/X sky130_fd_sc_hd__and3_1
XFILLER_190_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4636_ _5027_/A _4635_/B _4679_/B _4799_/B1 VGND VGND VPWR VPWR _4636_/X sky130_fd_sc_hd__o22a_1
XFILLER_148_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold610 _6912_/Q VGND VGND VPWR VPWR hold610/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 _7096_/Q VGND VGND VPWR VPWR hold621/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire4308 input10/X VGND VGND VPWR VPWR _3350_/A1 sky130_fd_sc_hd__clkbuf_1
X_4567_ _4607_/B _4567_/B VGND VGND VPWR VPWR _4567_/X sky130_fd_sc_hd__or2_1
Xhold632 _7007_/Q VGND VGND VPWR VPWR hold632/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold643 _6848_/Q VGND VGND VPWR VPWR hold643/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold654 _7047_/Q VGND VGND VPWR VPWR hold654/X sky130_fd_sc_hd__dlygate4sd3_1
X_6306_ _5938_/A _6333_/A2 _6306_/B1 _6306_/B2 _6305_/X VGND VGND VPWR VPWR _6306_/X
+ sky130_fd_sc_hd__a221o_1
Xwire3607 _4113_/A0 VGND VGND VPWR VPWR _5351_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold665 _7110_/Q VGND VGND VPWR VPWR hold665/X sky130_fd_sc_hd__dlygate4sd3_1
X_3518_ _3518_/A _3518_/B VGND VGND VPWR VPWR _4276_/A sky130_fd_sc_hd__nor2_2
Xhold676 _7093_/Q VGND VGND VPWR VPWR hold676/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3618 wire3619/X VGND VGND VPWR VPWR wire3618/X sky130_fd_sc_hd__clkbuf_1
X_4498_ _4947_/A _4944_/B _4933_/A _4566_/A _4932_/A VGND VGND VPWR VPWR _4498_/X
+ sky130_fd_sc_hd__a2111o_1
Xhold687 _7077_/Q VGND VGND VPWR VPWR hold687/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2906 _5827_/B1 VGND VGND VPWR VPWR _5842_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold698 _6993_/Q VGND VGND VPWR VPWR hold698/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6237_ _6686_/Q _6237_/A2 _6312_/B1 _6237_/B2 VGND VGND VPWR VPWR _6237_/X sky130_fd_sc_hd__a22o_1
XFILLER_104_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2917 _5694_/X VGND VGND VPWR VPWR _5820_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
X_3449_ _3448_/X _6788_/Q _3791_/B VGND VGND VPWR VPWR _6788_/D sky130_fd_sc_hd__mux2_1
Xwire2928 _5783_/C1 VGND VGND VPWR VPWR _5722_/C1 sky130_fd_sc_hd__clkbuf_1
Xwire2939 _5768_/A2 VGND VGND VPWR VPWR _5783_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ _6168_/A _6168_/B _6168_/C VGND VGND VPWR VPWR _6168_/X sky130_fd_sc_hd__or3_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5119_ _5119_/A _5119_/B _5119_/C VGND VGND VPWR VPWR _5119_/Y sky130_fd_sc_hd__nor3_1
XFILLER_84_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6099_ _6099_/A1 _6152_/B1 _6099_/B1 _6099_/B2 _6098_/X VGND VGND VPWR VPWR _6099_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_85_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A VGND VGND VPWR VPWR _3937_/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length1241 _3302_/Y VGND VGND VPWR VPWR _3783_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_4_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5470_ _3210_/A _5584_/A0 _5472_/S VGND VGND VPWR VPWR _7037_/D sky130_fd_sc_hd__mux2_1
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4421_ _4591_/A _4436_/B VGND VGND VPWR VPWR _4758_/C sky130_fd_sc_hd__nor2_2
XFILLER_172_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7140_ _7140_/CLK _7140_/D wire4071/A VGND VGND VPWR VPWR _7140_/Q sky130_fd_sc_hd__dfrtp_1
X_4352_ _4378_/B _4352_/B VGND VGND VPWR VPWR _4474_/A sky130_fd_sc_hd__or2_1
XFILLER_113_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3303_ _3303_/A _3378_/B VGND VGND VPWR VPWR _3303_/Y sky130_fd_sc_hd__nand2_1
X_4283_ _4295_/A0 _6228_/A1 _4287_/S VGND VGND VPWR VPWR _6731_/D sky130_fd_sc_hd__mux2_1
X_7071_ _7110_/CLK _7071_/D _7110_/RESET_B VGND VGND VPWR VPWR _7071_/Q sky130_fd_sc_hd__dfrtp_1
X_6022_ _6022_/A _6022_/B _6022_/C _6022_/D VGND VGND VPWR VPWR _6026_/A sky130_fd_sc_hd__or4_1
XFILLER_86_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6924_ _7127_/CLK _6924_/D _7051_/SET_B VGND VGND VPWR VPWR _6924_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_81_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6855_ _7133_/CLK _6855_/D fanout4077/X VGND VGND VPWR VPWR _6855_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5806_ _6166_/A1 _5806_/A2 _5806_/B1 _6163_/A1 _5805_/X VGND VGND VPWR VPWR _5813_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_167_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6786_ _3945_/A1 _6786_/D _6437_/X VGND VGND VPWR VPWR _6786_/Q sky130_fd_sc_hd__dfrtn_1
X_3998_ hold564/X _5199_/A0 _4000_/S VGND VGND VPWR VPWR _6495_/D sky130_fd_sc_hd__mux2_1
Xwire809 _3513_/X VGND VGND VPWR VPWR wire809/X sky130_fd_sc_hd__clkbuf_1
XFILLER_176_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5737_ _6089_/B2 _5737_/A2 _5736_/X VGND VGND VPWR VPWR _5740_/C sky130_fd_sc_hd__a21o_1
XFILLER_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5668_ _5985_/A1 _5735_/B1 _5724_/B1 _5986_/B2 _5665_/X VGND VGND VPWR VPWR _5681_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_163_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4619_ _4632_/A _4655_/B VGND VGND VPWR VPWR _4986_/A sky130_fd_sc_hd__nor2_1
XFILLER_191_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5599_ _5606_/A _5599_/B _5599_/C VGND VGND VPWR VPWR _7144_/D sky130_fd_sc_hd__and3_1
Xwire4105 input7/X VGND VGND VPWR VPWR _3500_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_151_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4116 wire4117/X VGND VGND VPWR VPWR wire4116/X sky130_fd_sc_hd__clkbuf_1
Xwire4127 input65/X VGND VGND VPWR VPWR wire4127/X sky130_fd_sc_hd__clkbuf_1
Xhold440 _7059_/Q VGND VGND VPWR VPWR hold440/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4138 input63/X VGND VGND VPWR VPWR wire4138/X sky130_fd_sc_hd__clkbuf_1
Xwire3404 _4118_/A0 VGND VGND VPWR VPWR _5365_/A0 sky130_fd_sc_hd__clkbuf_2
Xwire4149 input59/X VGND VGND VPWR VPWR wire4149/X sky130_fd_sc_hd__clkbuf_1
Xhold451 _6801_/Q VGND VGND VPWR VPWR hold451/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3415 _5578_/A0 VGND VGND VPWR VPWR _5248_/A0 sky130_fd_sc_hd__clkbuf_1
Xhold462 _6616_/Q VGND VGND VPWR VPWR hold462/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold473 _6737_/Q VGND VGND VPWR VPWR hold473/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3426 _4110_/A0 VGND VGND VPWR VPWR _5247_/A0 sky130_fd_sc_hd__clkbuf_2
Xhold484 _6664_/Q VGND VGND VPWR VPWR hold484/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3437 wire3438/X VGND VGND VPWR VPWR wire3437/X sky130_fd_sc_hd__clkbuf_1
Xhold495 _6794_/Q VGND VGND VPWR VPWR hold495/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3448 _4134_/A1 VGND VGND VPWR VPWR _4045_/A0 sky130_fd_sc_hd__clkbuf_1
Xwire2703 _6090_/A2 VGND VGND VPWR VPWR _6054_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire3459 _5462_/A0 VGND VGND VPWR VPWR _5453_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2714 _6205_/A2 VGND VGND VPWR VPWR _6154_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_77_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2725 _6210_/A2 VGND VGND VPWR VPWR wire2725/X sky130_fd_sc_hd__clkbuf_1
Xwire2736 wire2737/X VGND VGND VPWR VPWR _6206_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2747 _6199_/B1 VGND VGND VPWR VPWR _6174_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire2758 wire2759/X VGND VGND VPWR VPWR _6211_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2769 _6301_/A2 VGND VGND VPWR VPWR _6324_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_92_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length952 wire953/X VGND VGND VPWR VPWR _3354_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_181_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout3832 _6435_/B VGND VGND VPWR VPWR _6441_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_48_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length1093 _3450_/Y VGND VGND VPWR VPWR _3594_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_68_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4970_ _4488_/A _4846_/D _5127_/A _5158_/A VGND VGND VPWR VPWR _5140_/A sky130_fd_sc_hd__a211o_1
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3921_ _3198_/Y _3921_/A1 _3921_/S VGND VGND VPWR VPWR _3921_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6640_ _7206_/CLK _6640_/D VGND VGND VPWR VPWR _6640_/Q sky130_fd_sc_hd__dfxtp_1
X_3852_ _3850_/X _3851_/Y _3856_/B VGND VGND VPWR VPWR _3853_/B sky130_fd_sc_hd__o21ba_1
XFILLER_32_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6571_ _7084_/CLK _6571_/D _7035_/SET_B VGND VGND VPWR VPWR _6571_/Q sky130_fd_sc_hd__dfrtp_1
X_3783_ _6842_/Q _3783_/A2 _3783_/B1 _3783_/B2 VGND VGND VPWR VPWR _3783_/X sky130_fd_sc_hd__a22o_1
XFILLER_192_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5522_ _5522_/A0 hold180/X _5523_/S VGND VGND VPWR VPWR _7083_/D sky130_fd_sc_hd__mux2_1
XFILLER_157_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5453_ _5453_/A0 hold670/X _5453_/S VGND VGND VPWR VPWR _7022_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4404_ _4546_/A _4404_/B _4415_/A VGND VGND VPWR VPWR _4731_/B sky130_fd_sc_hd__nand3_2
Xclkbuf_leaf_42_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _6973_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_133_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5384_ _5456_/A0 hold660/X _5384_/S VGND VGND VPWR VPWR _6961_/D sky130_fd_sc_hd__mux2_1
XFILLER_132_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7123_ _7126_/CLK _7123_/D wire4042/X VGND VGND VPWR VPWR _7123_/Q sky130_fd_sc_hd__dfrtp_1
X_4335_ _4335_/A0 hold382/X _4335_/S VGND VGND VPWR VPWR _6775_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7054_ _7084_/CLK _7054_/D _7035_/SET_B VGND VGND VPWR VPWR _7054_/Q sky130_fd_sc_hd__dfrtp_1
X_4266_ hold525/X _4266_/A1 _4269_/S VGND VGND VPWR VPWR _6717_/D sky130_fd_sc_hd__mux2_1
Xwire1309 _6254_/X VGND VGND VPWR VPWR _6257_/C sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_57_csclk clkbuf_opt_1_0_csclk/X VGND VGND VPWR VPWR _7110_/CLK sky130_fd_sc_hd__clkbuf_16
X_6005_ _6005_/A1 _6049_/B _6005_/B1 _6858_/Q _6004_/X VGND VGND VPWR VPWR _6012_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_101_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3217_ _3217_/A VGND VGND VPWR VPWR _3217_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4197_ _6654_/Q wire379/X _4197_/S VGND VGND VPWR VPWR _6654_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6907_ _6939_/CLK _6907_/D _6404_/A VGND VGND VPWR VPWR _6907_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6838_ _7088_/CLK _6838_/D wire4069/A VGND VGND VPWR VPWR _6838_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire606 _5509_/S VGND VGND VPWR VPWR _5510_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_6769_ _7115_/CLK _6769_/D wire3981/X VGND VGND VPWR VPWR _6769_/Q sky130_fd_sc_hd__dfrtp_1
Xwire617 wire618/X VGND VGND VPWR VPWR _5490_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_7_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire628 wire629/X VGND VGND VPWR VPWR _5472_/S sky130_fd_sc_hd__clkbuf_2
Xwire639 wire640/X VGND VGND VPWR VPWR wire639/X sky130_fd_sc_hd__clkbuf_1
Xmax_length3946 fanout3944/X VGND VGND VPWR VPWR wire3945/A sky130_fd_sc_hd__buf_2
XFILLER_6_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3979 wire3981/X VGND VGND VPWR VPWR _7030_/RESET_B sky130_fd_sc_hd__clkbuf_2
XFILLER_109_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3201 _5113_/A2 VGND VGND VPWR VPWR _4871_/B sky130_fd_sc_hd__clkbuf_2
Xwire3212 _4477_/X VGND VGND VPWR VPWR _4670_/B sky130_fd_sc_hd__clkbuf_1
Xhold270 _6741_/Q VGND VGND VPWR VPWR hold270/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3223 _4427_/X VGND VGND VPWR VPWR _4933_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold281 _6918_/Q VGND VGND VPWR VPWR hold281/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 _7086_/Q VGND VGND VPWR VPWR hold292/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3245 wire3246/X VGND VGND VPWR VPWR wire3245/X sky130_fd_sc_hd__clkbuf_1
Xwire2511 _6006_/Y VGND VGND VPWR VPWR _6202_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2522 _6238_/A2 VGND VGND VPWR VPWR _6326_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3267 _4159_/B VGND VGND VPWR VPWR _4318_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_77_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3289 _3887_/Y VGND VGND VPWR VPWR wire3289/X sky130_fd_sc_hd__clkbuf_1
Xwire2544 _6129_/A2 VGND VGND VPWR VPWR _6087_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire1810 wire1811/X VGND VGND VPWR VPWR _6053_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire2555 _6092_/A2 VGND VGND VPWR VPWR _6258_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire1821 _7000_/Q VGND VGND VPWR VPWR _6191_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2566 _6164_/A2 VGND VGND VPWR VPWR _6141_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1832 _6997_/Q VGND VGND VPWR VPWR wire1832/X sky130_fd_sc_hd__clkbuf_1
Xwire2577 _6296_/A2 VGND VGND VPWR VPWR _6075_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1843 _6990_/Q VGND VGND VPWR VPWR _6129_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire2588 _5772_/A2 VGND VGND VPWR VPWR _5793_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2599 _4671_/Y VGND VGND VPWR VPWR _5158_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1865 _5743_/A VGND VGND VPWR VPWR _6086_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_45_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1876 wire1877/X VGND VGND VPWR VPWR wire1876/X sky130_fd_sc_hd__clkbuf_1
XFILLER_46_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1887 _6957_/Q VGND VGND VPWR VPWR _6098_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire1898 _6946_/Q VGND VGND VPWR VPWR _5985_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_110 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_121 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_132 input62/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4120_ hold29/A _4120_/B _4120_/C hold7/X VGND VGND VPWR VPWR _4120_/X sky130_fd_sc_hd__or4_1
XFILLER_110_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3790 wire3791/X VGND VGND VPWR VPWR wire3790/X sky130_fd_sc_hd__clkbuf_1
X_4051_ _4134_/A1 hold277/X _4051_/S VGND VGND VPWR VPWR _6540_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput5 mask_rev_in[10] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4953_ _4387_/B _4475_/A _4487_/B VGND VGND VPWR VPWR _5158_/C sky130_fd_sc_hd__o21a_1
XFILLER_101_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3904_ _7156_/Q _7155_/Q VGND VGND VPWR VPWR _6000_/A sky130_fd_sc_hd__and2b_1
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4884_ _4931_/B _4870_/B _4876_/B _4744_/X VGND VGND VPWR VPWR _4885_/D sky130_fd_sc_hd__o31a_1
X_6623_ _7094_/CLK _6623_/D _6672_/SET_B VGND VGND VPWR VPWR _6623_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_138_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3835_ _6444_/Q _6462_/Q _3835_/S VGND VGND VPWR VPWR _6462_/D sky130_fd_sc_hd__mux2_1
Xmax_length3209 _4482_/B VGND VGND VPWR VPWR _5105_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_177_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6554_ _6811_/CLK _6554_/D _6430_/A VGND VGND VPWR VPWR _6554_/Q sky130_fd_sc_hd__dfrtp_1
X_3766_ _7095_/Q _5535_/A _3766_/B1 _3766_/B2 _3736_/X VGND VGND VPWR VPWR _3789_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length2519 _6176_/B1 VGND VGND VPWR VPWR _6130_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_118_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5505_ _5505_/A0 hold298/X _5505_/S VGND VGND VPWR VPWR _7068_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6485_ _6825_/CLK _6485_/D wire3956/X VGND VGND VPWR VPWR _6485_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_106_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3697_ _3697_/A1 _3697_/A2 _5225_/A _5227_/A0 VGND VGND VPWR VPWR _3697_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5436_ _5436_/A0 hold632/X _5438_/S VGND VGND VPWR VPWR _7007_/D sky130_fd_sc_hd__mux2_1
Xoutput320 _6642_/Q VGND VGND VPWR VPWR wb_dat_o[11] sky130_fd_sc_hd__buf_12
XFILLER_133_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput331 _6631_/Q VGND VGND VPWR VPWR wb_dat_o[21] sky130_fd_sc_hd__buf_12
Xoutput342 wire3714/X VGND VGND VPWR VPWR wb_dat_o[31] sky130_fd_sc_hd__buf_12
X_5367_ _5367_/A _5403_/B VGND VGND VPWR VPWR _5369_/S sky130_fd_sc_hd__nand2_1
XFILLER_160_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7106_ _7130_/CLK _7106_/D fanout4077/X VGND VGND VPWR VPWR _7106_/Q sky130_fd_sc_hd__dfrtp_1
X_4318_ _4318_/A _4318_/B VGND VGND VPWR VPWR _4323_/S sky130_fd_sc_hd__and2_1
XFILLER_59_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5298_ _5487_/A0 hold448/X _5298_/S VGND VGND VPWR VPWR _6884_/D sky130_fd_sc_hd__mux2_1
Xwire1106 _3658_/A VGND VGND VPWR VPWR _3473_/C1 sky130_fd_sc_hd__dlymetal6s2s_1
X_7037_ _7134_/CLK _7037_/D fanout4057/X VGND VGND VPWR VPWR _7037_/Q sky130_fd_sc_hd__dfrtp_1
Xwire1128 _3763_/B1 VGND VGND VPWR VPWR _5430_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4249_ _4249_/A0 hold225/X _4251_/S VGND VGND VPWR VPWR _6703_/D sky130_fd_sc_hd__mux2_1
Xwire1139 _3771_/A2 VGND VGND VPWR VPWR _3634_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_75_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire403 _4103_/S VGND VGND VPWR VPWR _4101_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3710 _3191_/Y VGND VGND VPWR VPWR wire3709/A sky130_fd_sc_hd__clkbuf_1
Xwire414 _4053_/X VGND VGND VPWR VPWR _4069_/S sky130_fd_sc_hd__buf_2
XFILLER_156_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire425 _3626_/X VGND VGND VPWR VPWR wire425/X sky130_fd_sc_hd__clkbuf_1
Xwire436 _3494_/X VGND VGND VPWR VPWR _3499_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_149_580 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire447 _6268_/X VGND VGND VPWR VPWR wire447/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire458 _6045_/X VGND VGND VPWR VPWR wire458/X sky130_fd_sc_hd__clkbuf_1
Xwire469 wire470/X VGND VGND VPWR VPWR _5588_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_109_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length3798 hold5/X VGND VGND VPWR VPWR hold6/A sky130_fd_sc_hd__clkbuf_1
XFILLER_164_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3020 _5936_/B1 VGND VGND VPWR VPWR _5952_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire3031 _5741_/A2 VGND VGND VPWR VPWR _5807_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3042 _5826_/B1 VGND VGND VPWR VPWR _5778_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire3053 _5790_/B1 VGND VGND VPWR VPWR _5715_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3064 _5853_/B1 VGND VGND VPWR VPWR _5736_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2330 _6608_/Q VGND VGND VPWR VPWR _6286_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3075 _5807_/A2 VGND VGND VPWR VPWR _5784_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2341 _5924_/A1 VGND VGND VPWR VPWR _6293_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3086 _5846_/B1 VGND VGND VPWR VPWR _5832_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire2352 _6566_/Q VGND VGND VPWR VPWR wire2352/X sky130_fd_sc_hd__clkbuf_1
Xwire2363 wire2364/X VGND VGND VPWR VPWR _6249_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2374 wire2375/X VGND VGND VPWR VPWR _5952_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2385 _6526_/Q VGND VGND VPWR VPWR _6237_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire1640 _7064_/Q VGND VGND VPWR VPWR _6188_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire2396 _6334_/A1 VGND VGND VPWR VPWR _3493_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1651 _7058_/Q VGND VGND VPWR VPWR _5673_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire1662 wire1663/X VGND VGND VPWR VPWR _3561_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire1673 _6173_/B2 VGND VGND VPWR VPWR _3387_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire1684 wire1684/A VGND VGND VPWR VPWR _6103_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_74_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1695 _7042_/Q VGND VGND VPWR VPWR _5680_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3620_ _5906_/A1 _3676_/A2 _4198_/A _6657_/Q wire556/X VGND VGND VPWR VPWR _3620_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_159_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3551_ _3551_/A1 _3769_/B1 _3687_/B1 _5934_/B2 VGND VGND VPWR VPWR _3551_/X sky130_fd_sc_hd__a22o_1
Xwire970 _3275_/Y VGND VGND VPWR VPWR wire970/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire981 _6046_/B VGND VGND VPWR VPWR wire981/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire992 _6028_/Y VGND VGND VPWR VPWR wire992/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6270_ _7184_/Q _6319_/S wire445/X _6269_/X VGND VGND VPWR VPWR _7184_/D sky130_fd_sc_hd__o22a_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3482_ _3482_/A _3482_/B VGND VGND VPWR VPWR _4022_/A sky130_fd_sc_hd__nor2_1
XFILLER_115_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5221_ _5221_/A _5221_/B VGND VGND VPWR VPWR _5221_/X sky130_fd_sc_hd__or2_1
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5152_ _5152_/A1 _5027_/B _5108_/B _5152_/B2 VGND VGND VPWR VPWR _5152_/X sky130_fd_sc_hd__o22a_1
XFILLER_57_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4103_ hold10/X _4102_/X _4103_/S VGND VGND VPWR VPWR hold11/A sky130_fd_sc_hd__mux2_1
XFILLER_29_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5083_ _5083_/A _5083_/B _5083_/C _5083_/D VGND VGND VPWR VPWR _5107_/B sky130_fd_sc_hd__or4_1
XFILLER_84_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4034_ _4034_/A _5210_/B VGND VGND VPWR VPWR _4039_/S sky130_fd_sc_hd__and2_2
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5985_ _5985_/A1 _5985_/A2 _5985_/B1 _7135_/Q _5981_/X VGND VGND VPWR VPWR _5985_/X
+ sky130_fd_sc_hd__a221o_1
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4936_ _4947_/B VGND VGND VPWR VPWR _4957_/B sky130_fd_sc_hd__inv_2
XFILLER_178_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_10 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4867_ _4465_/X _4488_/B _4830_/Y _4847_/Y _4866_/X VGND VGND VPWR VPWR _4868_/D
+ sky130_fd_sc_hd__a2111o_1
XANTENNA_21 _5588_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_32 _3684_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_43 _5913_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_54 _3509_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6606_ _7208_/CLK _6606_/D wire4026/A VGND VGND VPWR VPWR _6606_/Q sky130_fd_sc_hd__dfrtp_1
X_3818_ _3818_/A _3818_/B VGND VGND VPWR VPWR _3818_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_193_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_65 _5747_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 wire2121/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4798_ _4569_/A _4561_/Y _4800_/A2 _4759_/B _4798_/B2 VGND VGND VPWR VPWR _4984_/C
+ sky130_fd_sc_hd__a32o_1
XANTENNA_87 _6211_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_98 wire3153/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6537_ _7090_/CLK _6537_/D _6430_/A VGND VGND VPWR VPWR _6537_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3749_ _3749_/A _3749_/B _3749_/C _3749_/D VGND VGND VPWR VPWR _3790_/A sky130_fd_sc_hd__or4_1
XFILLER_134_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6468_ _3487_/B2 _6468_/D _6423_/X VGND VGND VPWR VPWR _6468_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_97_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5419_ _5464_/A0 hold628/X _5420_/S VGND VGND VPWR VPWR _6992_/D sky130_fd_sc_hd__mux2_1
X_6399_ _6433_/A _6433_/B VGND VGND VPWR VPWR _6399_/X sky130_fd_sc_hd__and2_1
Xoutput172 wire2117/X VGND VGND VPWR VPWR irq[0] sky130_fd_sc_hd__buf_12
Xoutput183 _3217_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[17] sky130_fd_sc_hd__buf_12
Xoutput194 _3207_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[27] sky130_fd_sc_hd__buf_12
XFILLER_99_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length3540 _5532_/A1 VGND VGND VPWR VPWR wire3539/A sky130_fd_sc_hd__clkbuf_1
XFILLER_109_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2160 _6755_/Q VGND VGND VPWR VPWR wire2160/X sky130_fd_sc_hd__clkbuf_1
XFILLER_120_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2171 _6749_/Q VGND VGND VPWR VPWR wire2171/X sky130_fd_sc_hd__clkbuf_1
Xwire2182 _6743_/Q VGND VGND VPWR VPWR _3636_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_93_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2193 wire2194/X VGND VGND VPWR VPWR _6299_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire1470 wire1471/X VGND VGND VPWR VPWR wire1470/X sky130_fd_sc_hd__clkbuf_1
Xwire1481 wire1482/X VGND VGND VPWR VPWR wire1481/X sky130_fd_sc_hd__clkbuf_1
Xwire1492 _3918_/X VGND VGND VPWR VPWR wire1492/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5770_ _5770_/A _5770_/B _5770_/C _5770_/D VGND VGND VPWR VPWR _5770_/X sky130_fd_sc_hd__or4_1
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4721_ _4721_/A _4981_/A _4721_/C VGND VGND VPWR VPWR _4992_/B sky130_fd_sc_hd__or3_1
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4652_ _4652_/A _4652_/B VGND VGND VPWR VPWR _4652_/X sky130_fd_sc_hd__or2_1
XFILLER_30_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput30 mask_rev_in[4] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__clkbuf_1
X_3603_ _3602_/X _6786_/Q _3917_/A VGND VGND VPWR VPWR _6786_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput41 mgmt_gpio_in[14] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__clkbuf_1
Xinput52 mgmt_gpio_in[24] VGND VGND VPWR VPWR input52/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4583_ _4814_/A _4814_/B VGND VGND VPWR VPWR _4623_/A sky130_fd_sc_hd__or2_1
Xinput63 mgmt_gpio_in[34] VGND VGND VPWR VPWR input63/X sky130_fd_sc_hd__clkbuf_1
Xinput74 pad_flash_io1_di VGND VGND VPWR VPWR input74/X sky130_fd_sc_hd__clkbuf_1
X_6322_ _6322_/A1 _6322_/A2 _6322_/B1 _6322_/B2 _6321_/X VGND VGND VPWR VPWR _6332_/B
+ sky130_fd_sc_hd__a221o_1
Xinput85 spimemio_flash_io0_do VGND VGND VPWR VPWR input85/X sky130_fd_sc_hd__clkbuf_1
X_3534_ _3534_/A _3729_/B VGND VGND VPWR VPWR _4330_/A sky130_fd_sc_hd__nor2_1
XFILLER_116_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput96 usr1_vdd_pwrgood VGND VGND VPWR VPWR input96/X sky130_fd_sc_hd__clkbuf_1
XFILLER_115_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6253_ _6253_/A1 _6334_/B1 _6329_/A2 _6661_/Q VGND VGND VPWR VPWR _6253_/X sky130_fd_sc_hd__a22o_1
X_3465_ _3518_/A _3465_/B VGND VGND VPWR VPWR _3465_/Y sky130_fd_sc_hd__nor2_1
XFILLER_107_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5204_ _5422_/A0 hold418/X _5204_/S VGND VGND VPWR VPWR _6806_/D sky130_fd_sc_hd__mux2_1
XFILLER_103_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6184_ _6936_/Q _6184_/A2 _6184_/B1 _6184_/B2 VGND VGND VPWR VPWR _6184_/X sky130_fd_sc_hd__a22o_1
X_3396_ _6936_/Q _3396_/A2 wire911/X _3396_/B2 _3395_/X VGND VGND VPWR VPWR _3409_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_97_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5135_ _5135_/A1 _5003_/B _4758_/Y _4860_/A _4504_/B VGND VGND VPWR VPWR _5136_/B
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_84_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5066_ _5066_/A _5125_/A _5066_/C VGND VGND VPWR VPWR _5067_/C sky130_fd_sc_hd__or3_1
XFILLER_38_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4017_ _6393_/A0 hold304/X _4021_/S VGND VGND VPWR VPWR _6511_/D sky130_fd_sc_hd__mux2_1
XFILLER_44_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5968_ _6342_/A1 _5968_/A2 _5957_/X _5967_/X _6342_/C1 VGND VGND VPWR VPWR _5968_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4919_ _5021_/A _4633_/B _4665_/Y VGND VGND VPWR VPWR _4919_/X sky130_fd_sc_hd__o21ba_1
XFILLER_166_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5899_ _5899_/A1 _5964_/A2 _5955_/B1 _5899_/B2 VGND VGND VPWR VPWR _5899_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length2102 _6823_/Q VGND VGND VPWR VPWR wire2101/A sky130_fd_sc_hd__clkbuf_1
XFILLER_138_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length1401 _3472_/A VGND VGND VPWR VPWR _3344_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_165_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length1434 _4797_/A VGND VGND VPWR VPWR _4749_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_180_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_662 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length4093 wire4092/A VGND VGND VPWR VPWR wire4088/A sky130_fd_sc_hd__clkbuf_1
XFILLER_184_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_length1990 hold220/X VGND VGND VPWR VPWR _6066_/B2 sky130_fd_sc_hd__clkbuf_2
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ wire3728/X _3941_/A VGND VGND VPWR VPWR _3250_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_98_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6940_ _7129_/CLK _6940_/D wire4056/X VGND VGND VPWR VPWR _6940_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6871_ _7133_/CLK _6871_/D _7047_/RESET_B VGND VGND VPWR VPWR _6871_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5822_ _6182_/A1 _5822_/A2 _5821_/X VGND VGND VPWR VPWR _5825_/C sky130_fd_sc_hd__a21o_1
XFILLER_179_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5753_ _7164_/Q _5752_/X _6122_/S VGND VGND VPWR VPWR _7164_/D sky130_fd_sc_hd__mux2_1
X_4704_ _4704_/A _4704_/B VGND VGND VPWR VPWR _4704_/X sky130_fd_sc_hd__or2_1
XFILLER_148_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5684_ _7082_/Q _5684_/A2 _5684_/B1 _6866_/Q VGND VGND VPWR VPWR _5684_/X sky130_fd_sc_hd__a22o_1
XFILLER_175_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4635_ _5027_/A _4635_/B VGND VGND VPWR VPWR _4635_/Y sky130_fd_sc_hd__nor2_1
XFILLER_175_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold600 _7116_/Q VGND VGND VPWR VPWR hold600/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold611 _6836_/Q VGND VGND VPWR VPWR hold611/X sky130_fd_sc_hd__dlygate4sd3_1
X_4566_ _4566_/A _4596_/B VGND VGND VPWR VPWR _4567_/B sky130_fd_sc_hd__or2_1
Xhold622 _6577_/Q VGND VGND VPWR VPWR hold622/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold633 _6503_/Q VGND VGND VPWR VPWR hold633/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold644 _7004_/Q VGND VGND VPWR VPWR hold644/X sky130_fd_sc_hd__dlygate4sd3_1
X_6305_ _6305_/A1 _6336_/A2 _6326_/B1 _6305_/B2 VGND VGND VPWR VPWR _6305_/X sky130_fd_sc_hd__a22o_1
XFILLER_150_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3517_ _7139_/Q wire948/X _3548_/A2 _6140_/B2 _3516_/X VGND VGND VPWR VPWR _3524_/A
+ sky130_fd_sc_hd__a221o_1
Xwire3608 _5234_/A0 VGND VGND VPWR VPWR _4113_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_171_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold655 _6770_/Q VGND VGND VPWR VPWR hold655/X sky130_fd_sc_hd__dlygate4sd3_1
X_4497_ _4497_/A _4687_/B VGND VGND VPWR VPWR _4882_/A sky130_fd_sc_hd__or2_1
Xhold666 _7036_/Q VGND VGND VPWR VPWR hold666/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold677 _7005_/Q VGND VGND VPWR VPWR hold677/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3619 wire3620/X VGND VGND VPWR VPWR wire3619/X sky130_fd_sc_hd__clkbuf_1
Xhold688 _6528_/Q VGND VGND VPWR VPWR hold688/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6236_ _6236_/A1 _6340_/A2 _6337_/B1 _6236_/B2 _6235_/X VGND VGND VPWR VPWR _6242_/C
+ sky130_fd_sc_hd__a221o_1
Xhold699 _6809_/Q VGND VGND VPWR VPWR hold699/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire2907 _5696_/X VGND VGND VPWR VPWR _5827_/B1 sky130_fd_sc_hd__clkbuf_2
X_3448_ wire369/X _6787_/Q _3791_/A VGND VGND VPWR VPWR _3448_/X sky130_fd_sc_hd__mux2_1
Xwire2918 _5965_/A2 VGND VGND VPWR VPWR _5909_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_134_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6167_ _6167_/A _6167_/B _6167_/C _6167_/D VGND VGND VPWR VPWR _6168_/C sky130_fd_sc_hd__or4_1
X_3379_ _3711_/A _3379_/B VGND VGND VPWR VPWR _5221_/B sky130_fd_sc_hd__nor2_2
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5118_ _4538_/B _4478_/Y _4644_/B _4829_/Y _5117_/X VGND VGND VPWR VPWR _5119_/C
+ sky130_fd_sc_hd__a2111o_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6098_ _6098_/A1 _6131_/A2 _6149_/B1 _7122_/Q VGND VGND VPWR VPWR _6098_/X sky130_fd_sc_hd__a22o_1
XFILLER_84_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5049_ _5049_/A _5049_/B _5049_/C _5049_/D VGND VGND VPWR VPWR _5151_/A sky130_fd_sc_hd__or4_1
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4420_ _4420_/A _4450_/A _4566_/A VGND VGND VPWR VPWR _4738_/A sky130_fd_sc_hd__or3_2
XFILLER_132_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4351_ _4351_/A _4351_/B VGND VGND VPWR VPWR _4352_/B sky130_fd_sc_hd__nand2_1
XFILLER_99_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3302_ _3546_/B _3512_/B VGND VGND VPWR VPWR _3302_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7070_ _7115_/CLK _7070_/D wire3980/X VGND VGND VPWR VPWR _7070_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4282_ _4282_/A _4282_/B VGND VGND VPWR VPWR _4287_/S sky130_fd_sc_hd__nand2_2
XFILLER_98_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6021_ _6021_/A _6021_/B VGND VGND VPWR VPWR _6027_/D sky130_fd_sc_hd__nor2_1
XFILLER_86_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3233_ _3233_/A VGND VGND VPWR VPWR _3233_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_101_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_1_1_csclk clkbuf_1_1_1_csclk/A VGND VGND VPWR VPWR clkbuf_2_3_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_39_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6923_ _6939_/CLK _6923_/D _6923_/SET_B VGND VGND VPWR VPWR _6923_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_82_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6854_ _7131_/CLK _6854_/D wire4058/A VGND VGND VPWR VPWR _6854_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5805_ _6152_/A1 _5805_/A2 _5805_/B1 _6951_/Q VGND VGND VPWR VPWR _5805_/X sky130_fd_sc_hd__a22o_1
X_6785_ _3945_/A1 _6785_/D _6436_/X VGND VGND VPWR VPWR _6785_/Q sky130_fd_sc_hd__dfrtn_1
X_3997_ hold565/X _4311_/A0 _4000_/S VGND VGND VPWR VPWR _6494_/D sky130_fd_sc_hd__mux2_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5736_ _5736_/A1 _5736_/A2 _5736_/B1 _5736_/B2 VGND VGND VPWR VPWR _5736_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5667_ _5688_/A _5705_/B _5700_/C VGND VGND VPWR VPWR _5667_/X sky130_fd_sc_hd__and3_1
XFILLER_136_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4618_ _5107_/A _4916_/A _4618_/C _4618_/D VGND VGND VPWR VPWR _4642_/A sky130_fd_sc_hd__and4b_1
XFILLER_190_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5598_ _7144_/Q _5604_/D VGND VGND VPWR VPWR _5599_/C sky130_fd_sc_hd__or2_1
XFILLER_190_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4106 wire4107/X VGND VGND VPWR VPWR _3957_/A sky130_fd_sc_hd__clkbuf_1
Xwire4117 _3598_/A1 VGND VGND VPWR VPWR wire4117/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold430 _6534_/Q VGND VGND VPWR VPWR hold430/X sky130_fd_sc_hd__dlygate4sd3_1
X_4549_ _4963_/A VGND VGND VPWR VPWR _4549_/Y sky130_fd_sc_hd__inv_2
Xwire4128 wire4129/X VGND VGND VPWR VPWR _3581_/B2 sky130_fd_sc_hd__clkbuf_1
Xhold441 _6909_/Q VGND VGND VPWR VPWR hold441/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 _7054_/Q VGND VGND VPWR VPWR hold452/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4139 wire4140/X VGND VGND VPWR VPWR _3718_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_150_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold463 _6617_/Q VGND VGND VPWR VPWR hold463/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3416 hold45/X VGND VGND VPWR VPWR _5578_/A0 sky130_fd_sc_hd__clkbuf_1
Xhold474 _6797_/Q VGND VGND VPWR VPWR hold474/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3438 wire3438/A VGND VGND VPWR VPWR wire3438/X sky130_fd_sc_hd__clkbuf_1
Xhold485 _6555_/Q VGND VGND VPWR VPWR hold485/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 _6561_/Q VGND VGND VPWR VPWR hold496/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3449 _4209_/A1 VGND VGND VPWR VPWR _4134_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire2704 _6111_/B1 VGND VGND VPWR VPWR _6090_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2715 _6188_/A2 VGND VGND VPWR VPWR _6205_/A2 sky130_fd_sc_hd__clkbuf_2
X_6219_ _7181_/Q wire449/X _6219_/S VGND VGND VPWR VPWR _6219_/X sky130_fd_sc_hd__mux2_1
Xwire2726 wire2726/A VGND VGND VPWR VPWR _6210_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_89_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2737 _6009_/X VGND VGND VPWR VPWR wire2737/X sky130_fd_sc_hd__clkbuf_1
X_7199_ _7204_/CLK _7199_/D wire4260/X VGND VGND VPWR VPWR hold77/A sky130_fd_sc_hd__dfrtp_1
Xwire2748 wire2749/X VGND VGND VPWR VPWR _6199_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_58_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2759 _6003_/X VGND VGND VPWR VPWR wire2759/X sky130_fd_sc_hd__clkbuf_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length931 _3317_/Y VGND VGND VPWR VPWR wire929/A sky130_fd_sc_hd__clkbuf_2
XFILLER_127_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3950 wire3950/A VGND VGND VPWR VPWR wire3950/X sky130_fd_sc_hd__clkbuf_4
XFILLER_68_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3961 wire3963/A VGND VGND VPWR VPWR wire3961/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3920_ _3197_/Y _3920_/A1 _3921_/S VGND VGND VPWR VPWR _3920_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3851_ _6455_/Q _6454_/Q _3834_/B VGND VGND VPWR VPWR _3851_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_177_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6570_ _7088_/CLK _6570_/D wire4069/A VGND VGND VPWR VPWR _6570_/Q sky130_fd_sc_hd__dfrtp_1
X_3782_ _6474_/Q _3782_/A2 _3674_/Y _3782_/B2 _3735_/X VGND VGND VPWR VPWR _3788_/A
+ sky130_fd_sc_hd__a221o_1
X_5521_ _5554_/A0 hold326/X _5523_/S VGND VGND VPWR VPWR _7082_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5452_ _5452_/A0 hold648/X _5453_/S VGND VGND VPWR VPWR _7021_/D sky130_fd_sc_hd__mux2_1
XFILLER_8_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4403_ _4404_/B _4415_/A _4546_/A VGND VGND VPWR VPWR _4731_/C sky130_fd_sc_hd__a21o_1
XFILLER_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5383_ _5551_/A0 hold573/X _5384_/S VGND VGND VPWR VPWR _6960_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7122_ _7126_/CLK _7122_/D wire4039/X VGND VGND VPWR VPWR _7122_/Q sky130_fd_sc_hd__dfrtp_1
X_4334_ _4334_/A0 hold379/X _4335_/S VGND VGND VPWR VPWR _6774_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7053_ _7134_/CLK _7053_/D _7134_/RESET_B VGND VGND VPWR VPWR _7053_/Q sky130_fd_sc_hd__dfrtp_1
X_4265_ hold637/X _5422_/A0 _4268_/S VGND VGND VPWR VPWR _6716_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6004_ _6004_/A1 _6074_/A2 _6074_/B1 _6004_/B2 VGND VGND VPWR VPWR _6004_/X sky130_fd_sc_hd__a22o_1
XFILLER_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3216_ _3216_/A VGND VGND VPWR VPWR _3216_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4196_ _6653_/Q wire374/X _4196_/S VGND VGND VPWR VPWR _6653_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6906_ _6963_/CLK _6906_/D _7042_/SET_B VGND VGND VPWR VPWR _6906_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_23_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6837_ _6973_/CLK _6837_/D wire4069/X VGND VGND VPWR VPWR _6837_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire607 _5507_/S VGND VGND VPWR VPWR _5509_/S sky130_fd_sc_hd__clkbuf_1
X_6768_ _6775_/CLK _6768_/D wire3978/X VGND VGND VPWR VPWR _6768_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_149_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire618 _5492_/S VGND VGND VPWR VPWR wire618/X sky130_fd_sc_hd__clkbuf_1
Xwire629 wire630/X VGND VGND VPWR VPWR wire629/X sky130_fd_sc_hd__clkbuf_1
Xmax_length3936 wire3935/A VGND VGND VPWR VPWR _6743_/SET_B sky130_fd_sc_hd__clkbuf_2
XFILLER_109_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5719_ _5719_/A _5719_/B _5719_/C _5719_/D VGND VGND VPWR VPWR _5719_/X sky130_fd_sc_hd__or4_1
X_6699_ _7206_/CLK _6699_/D _6348_/B VGND VGND VPWR VPWR _6699_/Q sky130_fd_sc_hd__dfrtp_1
Xmax_length3969 wire3970/X VGND VGND VPWR VPWR wire3968/A sky130_fd_sc_hd__clkbuf_2
XFILLER_148_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3202 _5094_/A VGND VGND VPWR VPWR _5113_/A2 sky130_fd_sc_hd__clkbuf_2
Xhold260 _6638_/Q VGND VGND VPWR VPWR hold260/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 _4295_/X VGND VGND VPWR VPWR _6741_/D sky130_fd_sc_hd__dlygate4sd3_1
Xwire3213 _4526_/B VGND VGND VPWR VPWR _4506_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_104_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3224 _4524_/A VGND VGND VPWR VPWR _4516_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold282 _7139_/Q VGND VGND VPWR VPWR hold282/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3235 wire3236/X VGND VGND VPWR VPWR _5034_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_172_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3246 hold7/X VGND VGND VPWR VPWR wire3246/X sky130_fd_sc_hd__clkbuf_1
Xwire2501 _6152_/B1 VGND VGND VPWR VPWR _6055_/B1 sky130_fd_sc_hd__clkbuf_2
Xhold293 _6747_/Q VGND VGND VPWR VPWR hold293/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3257 _4324_/B VGND VGND VPWR VPWR _5535_/B sky130_fd_sc_hd__buf_2
Xwire2523 wire2524/X VGND VGND VPWR VPWR _6238_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire2534 _6301_/B1 VGND VGND VPWR VPWR _6324_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3279 wire3280/X VGND VGND VPWR VPWR _5475_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2545 _5999_/A2 VGND VGND VPWR VPWR _6129_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1800 wire1801/X VGND VGND VPWR VPWR wire1800/X sky130_fd_sc_hd__clkbuf_1
Xwire1811 wire1812/X VGND VGND VPWR VPWR wire1811/X sky130_fd_sc_hd__clkbuf_1
Xwire2556 _6208_/A2 VGND VGND VPWR VPWR _6157_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_131_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1822 wire1823/X VGND VGND VPWR VPWR _6158_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire2567 _6215_/A2 VGND VGND VPWR VPWR _6164_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire1833 _6996_/Q VGND VGND VPWR VPWR _6086_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire2578 _6320_/A2 VGND VGND VPWR VPWR _6296_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire1844 wire1845/X VGND VGND VPWR VPWR _3560_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2589 _5858_/A2 VGND VGND VPWR VPWR _5772_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire1855 _6986_/Q VGND VGND VPWR VPWR _5999_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_18_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1866 _6972_/Q VGND VGND VPWR VPWR _5743_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_65_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1877 _6967_/Q VGND VGND VPWR VPWR wire1877/X sky130_fd_sc_hd__clkbuf_1
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1888 hold230/X VGND VGND VPWR VPWR _5377_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_65_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1899 wire1900/X VGND VGND VPWR VPWR _6210_/B2 sky130_fd_sc_hd__clkbuf_2
XANTENNA_100 _4114_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_111 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_122 wb_clk_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_133 input61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length794 wire795/X VGND VGND VPWR VPWR _3757_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_142_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3780 _6544_/Q VGND VGND VPWR VPWR _3850_/A sky130_fd_sc_hd__buf_2
XFILLER_122_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4050_ _4139_/A1 hold276/X _4051_/S VGND VGND VPWR VPWR _6539_/D sky130_fd_sc_hd__mux2_1
Xwire3791 wire3792/X VGND VGND VPWR VPWR wire3791/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput6 mask_rev_in[11] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4952_ _4952_/A _5031_/B _5059_/B VGND VGND VPWR VPWR _4954_/C sky130_fd_sc_hd__or3_1
XFILLER_45_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3903_ _7153_/Q _7154_/Q VGND VGND VPWR VPWR _6014_/A sky130_fd_sc_hd__and2b_1
X_4883_ _4931_/B _4450_/Y _4870_/B _4417_/X VGND VGND VPWR VPWR _4885_/C sky130_fd_sc_hd__o31a_1
X_3834_ _6541_/Q _3834_/B VGND VGND VPWR VPWR _3835_/S sky130_fd_sc_hd__nand2_1
X_6622_ _7094_/CLK _6622_/D _6672_/SET_B VGND VGND VPWR VPWR _6622_/Q sky130_fd_sc_hd__dfrtp_1
X_6553_ _7131_/CLK hold13/X wire4058/X VGND VGND VPWR VPWR hold12/A sky130_fd_sc_hd__dfrtp_1
X_3765_ _3765_/A1 wire813/X wire395/X wire415/X _3472_/Y VGND VGND VPWR VPWR _3765_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_192_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5504_ _5504_/A0 hold503/X _5504_/S VGND VGND VPWR VPWR _7067_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6484_ _7036_/CLK _6484_/D wire3974/A VGND VGND VPWR VPWR _6484_/Q sky130_fd_sc_hd__dfstp_2
X_3696_ _3696_/A1 wire942/X wire905/X input72/X _3695_/X VGND VGND VPWR VPWR _3696_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5435_ _5453_/A0 hold659/X _5438_/S VGND VGND VPWR VPWR _7006_/D sky130_fd_sc_hd__mux2_1
Xoutput310 _3940_/X VGND VGND VPWR VPWR serial_load sky130_fd_sc_hd__buf_12
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput321 _6643_/Q VGND VGND VPWR VPWR wb_dat_o[12] sky130_fd_sc_hd__buf_12
Xoutput332 _6632_/Q VGND VGND VPWR VPWR wb_dat_o[22] sky130_fd_sc_hd__buf_12
XFILLER_160_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput343 _6650_/Q VGND VGND VPWR VPWR wb_dat_o[3] sky130_fd_sc_hd__buf_12
XFILLER_161_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5366_ _5375_/A0 hold348/X _5366_/S VGND VGND VPWR VPWR _6945_/D sky130_fd_sc_hd__mux2_1
X_7105_ _7135_/CLK _7105_/D wire4056/X VGND VGND VPWR VPWR _7105_/Q sky130_fd_sc_hd__dfrtp_1
X_4317_ hold537/X _5558_/A0 _4317_/S VGND VGND VPWR VPWR _6760_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5297_ _5396_/A1 hold207/X _5298_/S VGND VGND VPWR VPWR _6883_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1107 _3735_/A2 VGND VGND VPWR VPWR _3983_/A sky130_fd_sc_hd__clkbuf_1
X_7036_ _7036_/CLK _7036_/D wire3985/X VGND VGND VPWR VPWR _7036_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1118 _3341_/Y VGND VGND VPWR VPWR _3652_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
X_4248_ _4248_/A0 hold218/X _4251_/S VGND VGND VPWR VPWR _6702_/D sky130_fd_sc_hd__mux2_1
Xwire1129 _3553_/A2 VGND VGND VPWR VPWR _3763_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_142_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4179_ _4179_/A0 hold260/X _4179_/S VGND VGND VPWR VPWR _6638_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire404 _4087_/X VGND VGND VPWR VPWR _4103_/S sky130_fd_sc_hd__clkbuf_2
Xwire415 wire416/X VGND VGND VPWR VPWR wire415/X sky130_fd_sc_hd__clkbuf_1
Xwire426 _3620_/X VGND VGND VPWR VPWR wire426/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire437 wire438/X VGND VGND VPWR VPWR _3499_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_183_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire448 _6243_/X VGND VGND VPWR VPWR wire448/X sky130_fd_sc_hd__clkbuf_1
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire459 _5968_/X VGND VGND VPWR VPWR wire459/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3010 wire3011/X VGND VGND VPWR VPWR wire3010/X sky130_fd_sc_hd__clkbuf_1
XFILLER_105_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3021 wire3022/X VGND VGND VPWR VPWR _5936_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_151_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3032 _5680_/A2 VGND VGND VPWR VPWR _5741_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_183_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3043 _5764_/A2 VGND VGND VPWR VPWR _5745_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_104_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3054 _5761_/B1 VGND VGND VPWR VPWR _5790_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire3065 _5791_/A2 VGND VGND VPWR VPWR _5797_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_132_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2331 wire2332/X VGND VGND VPWR VPWR _6238_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_116_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3076 wire3077/X VGND VGND VPWR VPWR _5807_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire2342 _6598_/Q VGND VGND VPWR VPWR _5924_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_78_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3087 wire3088/X VGND VGND VPWR VPWR _5846_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire2353 _6560_/Q VGND VGND VPWR VPWR _3929_/A0 sky130_fd_sc_hd__clkbuf_1
Xwire3098 _5664_/X VGND VGND VPWR VPWR _5848_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2364 wire2365/X VGND VGND VPWR VPWR wire2364/X sky130_fd_sc_hd__clkbuf_1
Xwire2375 _4039_/A0 VGND VGND VPWR VPWR wire2375/X sky130_fd_sc_hd__clkbuf_1
Xwire1630 _7070_/Q VGND VGND VPWR VPWR _3483_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire1641 _7063_/Q VGND VGND VPWR VPWR _6154_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire2386 hold518/X VGND VGND VPWR VPWR _6324_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1652 wire1653/X VGND VGND VPWR VPWR _6172_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2397 _6515_/Q VGND VGND VPWR VPWR _6334_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1663 wire1664/X VGND VGND VPWR VPWR wire1663/X sky130_fd_sc_hd__clkbuf_1
Xwire1674 _7048_/Q VGND VGND VPWR VPWR _6173_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1696 wire1697/X VGND VGND VPWR VPWR _6215_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _6945_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_56_csclk _7117_/CLK VGND VGND VPWR VPWR _7016_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_186_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire960 _3280_/Y VGND VGND VPWR VPWR wire960/X sky130_fd_sc_hd__clkbuf_2
X_3550_ _7069_/Q _3550_/A2 _3550_/B1 _5756_/B2 VGND VGND VPWR VPWR _3550_/X sky130_fd_sc_hd__a22o_1
XFILLER_128_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire971 _3275_/Y VGND VGND VPWR VPWR wire971/X sky130_fd_sc_hd__dlymetal6s2s_1
Xwire982 _6029_/X VGND VGND VPWR VPWR _6046_/B sky130_fd_sc_hd__clkbuf_2
Xwire993 _5813_/X VGND VGND VPWR VPWR wire993/X sky130_fd_sc_hd__clkbuf_1
X_3481_ _6478_/Q _3782_/A2 _3992_/A _6494_/Q VGND VGND VPWR VPWR _3481_/X sky130_fd_sc_hd__a22o_1
XFILLER_6_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5220_ _5220_/A0 hold522/X _5220_/S VGND VGND VPWR VPWR _6818_/D sky130_fd_sc_hd__mux2_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout3471 hold15/X VGND VGND VPWR VPWR hold16/A sky130_fd_sc_hd__buf_6
X_5151_ _5151_/A _5151_/B _5151_/C _5174_/C VGND VGND VPWR VPWR _5151_/X sky130_fd_sc_hd__or4_1
XFILLER_69_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4102_ _6841_/Q hold3/X _4102_/S VGND VGND VPWR VPWR _4102_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5082_ _4673_/A _5108_/B _5015_/B VGND VGND VPWR VPWR _5083_/D sky130_fd_sc_hd__o21bai_1
XFILLER_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4033_ _6324_/A1 _4033_/A1 _4033_/S VGND VGND VPWR VPWR _6525_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5984_ _6019_/A _6021_/B VGND VGND VPWR VPWR _6023_/B sky130_fd_sc_hd__nor2_1
XFILLER_40_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4935_ _4935_/A _4935_/B _4935_/C VGND VGND VPWR VPWR _4947_/B sky130_fd_sc_hd__or3_1
Xclkbuf_3_7_0_csclk clkbuf_3_7_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_7_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_33_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_11 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 wire630/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4866_ _5126_/A _5162_/A _4866_/C _4866_/D VGND VGND VPWR VPWR _4866_/X sky130_fd_sc_hd__or4_1
XFILLER_177_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_33 _3625_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmax_length3029 _5676_/X VGND VGND VPWR VPWR wire3022/A sky130_fd_sc_hd__clkbuf_1
X_6605_ _6702_/CLK _6605_/D wire3958/X VGND VGND VPWR VPWR _6605_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA_44 wire1328/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3817_ _3820_/A _3821_/S _6467_/Q VGND VGND VPWR VPWR _3818_/B sky130_fd_sc_hd__o21a_1
XANTENNA_55 wire1539/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4797_ _4797_/A _4797_/B VGND VGND VPWR VPWR _4810_/D sky130_fd_sc_hd__nand2_1
XFILLER_165_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_66 _6089_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_77 _6282_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_88 _6211_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6536_ _7090_/CLK _6536_/D wire3943/A VGND VGND VPWR VPWR _6536_/Q sky130_fd_sc_hd__dfrtp_1
X_3748_ _3748_/A1 wire963/X wire836/X _3748_/B2 _3747_/X VGND VGND VPWR VPWR _3749_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA_99 _5566_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6467_ _3487_/B2 _6467_/D _6422_/X VGND VGND VPWR VPWR _6467_/Q sky130_fd_sc_hd__dfrtp_1
X_3679_ _3679_/A _3679_/B _3679_/C _3679_/D VGND VGND VPWR VPWR _3689_/A sky130_fd_sc_hd__or4_1
XFILLER_134_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5418_ _5508_/A0 hold531/X _5418_/S VGND VGND VPWR VPWR _6991_/D sky130_fd_sc_hd__mux2_1
X_6398_ _6429_/A _6431_/B VGND VGND VPWR VPWR _6398_/X sky130_fd_sc_hd__and2_1
Xoutput173 wire1450/X VGND VGND VPWR VPWR irq[1] sky130_fd_sc_hd__buf_12
XFILLER_161_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput184 _3216_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[18] sky130_fd_sc_hd__buf_12
X_5349_ _5349_/A _5553_/B VGND VGND VPWR VPWR _5353_/S sky130_fd_sc_hd__nand2_1
Xoutput195 _3206_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[28] sky130_fd_sc_hd__buf_12
XFILLER_102_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7019_ _7121_/CLK _7019_/D wire4042/X VGND VGND VPWR VPWR _7019_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length3541 _5532_/A1 VGND VGND VPWR VPWR _4049_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length2840 _5707_/A2 VGND VGND VPWR VPWR wire2836/A sky130_fd_sc_hd__clkbuf_1
XFILLER_137_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2161 _6754_/Q VGND VGND VPWR VPWR _6302_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2172 wire2173/X VGND VGND VPWR VPWR _6282_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2183 _5911_/B2 VGND VGND VPWR VPWR _6282_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_93_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2194 _6739_/Q VGND VGND VPWR VPWR wire2194/X sky130_fd_sc_hd__clkbuf_1
Xwire1460 wire1461/X VGND VGND VPWR VPWR wire1460/X sky130_fd_sc_hd__clkbuf_1
Xwire1471 _3925_/X VGND VGND VPWR VPWR wire1471/X sky130_fd_sc_hd__clkbuf_1
Xwire1482 wire1483/X VGND VGND VPWR VPWR wire1482/X sky130_fd_sc_hd__clkbuf_1
Xwire1493 _3730_/X VGND VGND VPWR VPWR _3735_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4720_ _5031_/B _4899_/B _4720_/C VGND VGND VPWR VPWR _4722_/C sky130_fd_sc_hd__or3_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4651_ _4693_/A _4660_/B VGND VGND VPWR VPWR _4651_/X sky130_fd_sc_hd__or2_1
XFILLER_187_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput20 mask_rev_in[24] VGND VGND VPWR VPWR input20/X sky130_fd_sc_hd__clkbuf_1
X_3602_ wire367/X _6785_/Q _3791_/A VGND VGND VPWR VPWR _3602_/X sky130_fd_sc_hd__mux2_1
Xinput31 mask_rev_in[5] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__clkbuf_1
X_4582_ _4632_/A _4582_/B VGND VGND VPWR VPWR _4984_/A sky130_fd_sc_hd__nor2_1
Xinput42 mgmt_gpio_in[15] VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__clkbuf_1
Xinput53 mgmt_gpio_in[25] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__clkbuf_1
Xinput64 mgmt_gpio_in[35] VGND VGND VPWR VPWR input64/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire790 wire791/X VGND VGND VPWR VPWR _5205_/A sky130_fd_sc_hd__clkbuf_1
Xinput75 porb VGND VGND VPWR VPWR input75/X sky130_fd_sc_hd__clkbuf_1
X_3533_ _3533_/A1 _3533_/A2 _3342_/Y _6130_/B2 wire562/X VGND VGND VPWR VPWR _3541_/B
+ sky130_fd_sc_hd__a221o_1
X_6321_ _6321_/A1 _6321_/A2 _6321_/B1 _6321_/B2 VGND VGND VPWR VPWR _6321_/X sky130_fd_sc_hd__a22o_1
XFILLER_128_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput86 spimemio_flash_io0_oeb VGND VGND VPWR VPWR input86/X sky130_fd_sc_hd__clkbuf_1
Xinput97 usr2_vcc_pwrgood VGND VGND VPWR VPWR input97/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6252_ _6252_/A1 _6330_/A2 _6322_/A2 _6252_/B2 _6248_/X VGND VGND VPWR VPWR _6257_/B
+ sky130_fd_sc_hd__a221o_1
X_3464_ _6322_/A1 _3707_/B1 _3464_/B1 _6321_/B2 VGND VGND VPWR VPWR _3464_/X sky130_fd_sc_hd__a22o_1
XFILLER_107_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5203_ _5203_/A _5203_/B VGND VGND VPWR VPWR _5204_/S sky130_fd_sc_hd__nand2_1
X_6183_ _6183_/A1 _6183_/A2 _6183_/B1 _6183_/B2 _6182_/X VGND VGND VPWR VPWR _6193_/B
+ sky130_fd_sc_hd__a221o_1
X_3395_ _5823_/A1 _3441_/A2 _3393_/X wire573/X VGND VGND VPWR VPWR _3395_/X sky130_fd_sc_hd__a211o_1
XFILLER_130_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5134_ _5134_/A _5134_/B _5134_/C _5134_/D VGND VGND VPWR VPWR _5148_/D sky130_fd_sc_hd__or4_1
XFILLER_69_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5065_ _5065_/A _5065_/B _5065_/C _5065_/D VGND VGND VPWR VPWR _5066_/C sky130_fd_sc_hd__or4_1
XFILLER_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4016_ _4016_/A _5529_/B VGND VGND VPWR VPWR _4021_/S sky130_fd_sc_hd__nand2_2
XFILLER_72_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5967_ _5967_/A _5967_/B _5967_/C _5967_/D VGND VGND VPWR VPWR _5967_/X sky130_fd_sc_hd__or4_1
X_4918_ _4492_/A _4721_/C _4719_/A VGND VGND VPWR VPWR _4963_/B sky130_fd_sc_hd__a21oi_1
XFILLER_21_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5898_ _6635_/Q _5898_/A2 _5910_/A2 _6607_/Q _5897_/X VGND VGND VPWR VPWR _5901_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_193_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4849_ _4520_/B _4506_/B _4708_/A VGND VGND VPWR VPWR _4865_/C sky130_fd_sc_hd__o21ai_1
XFILLER_165_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6519_ _7090_/CLK _6519_/D wire3945/A VGND VGND VPWR VPWR _6519_/Q sky130_fd_sc_hd__dfrtp_1
Xmax_length1446 _4417_/X VGND VGND VPWR VPWR _4418_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_106_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length4072 wire4071/A VGND VGND VPWR VPWR _7138_/RESET_B sky130_fd_sc_hd__clkbuf_2
XFILLER_8_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length3393 _5491_/A0 VGND VGND VPWR VPWR _5437_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_125_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1290 _3531_/A VGND VGND VPWR VPWR _3504_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6870_ _7129_/CLK _6870_/D fanout4057/X VGND VGND VPWR VPWR _6870_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5821_ _6177_/A1 _5821_/A2 _5821_/B1 _7016_/Q VGND VGND VPWR VPWR _5821_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5752_ _6121_/A1 _7163_/Q wire464/X VGND VGND VPWR VPWR _5752_/X sky130_fd_sc_hd__a21o_1
XFILLER_148_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4703_ _4624_/B _4704_/B _4701_/X _4702_/X VGND VGND VPWR VPWR _4703_/X sky130_fd_sc_hd__o211a_1
XFILLER_187_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5683_ _5683_/A _5706_/B _5703_/B VGND VGND VPWR VPWR _5683_/X sky130_fd_sc_hd__and3_1
XFILLER_30_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4634_ _4634_/A _4915_/A _4987_/A _4634_/D VGND VGND VPWR VPWR _4642_/B sky130_fd_sc_hd__nor4_1
XFILLER_147_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4565_ _4565_/A _4666_/B VGND VGND VPWR VPWR _4565_/X sky130_fd_sc_hd__or2_2
Xhold601 _7026_/Q VGND VGND VPWR VPWR hold601/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold612 _6759_/Q VGND VGND VPWR VPWR hold612/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold623 _6863_/Q VGND VGND VPWR VPWR hold623/X sky130_fd_sc_hd__dlygate4sd3_1
X_6304_ _6304_/A1 _6304_/A2 _6304_/B1 _6759_/Q _6303_/X VGND VGND VPWR VPWR _6304_/X
+ sky130_fd_sc_hd__a221o_1
Xhold634 _6526_/Q VGND VGND VPWR VPWR hold634/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 _7015_/Q VGND VGND VPWR VPWR hold645/X sky130_fd_sc_hd__dlygate4sd3_1
X_3516_ _6958_/Q _5376_/A _3516_/B1 _6966_/Q VGND VGND VPWR VPWR _3516_/X sky130_fd_sc_hd__a22o_1
X_4496_ _4745_/A _4496_/B VGND VGND VPWR VPWR _5050_/A sky130_fd_sc_hd__or2_1
Xhold656 _7057_/Q VGND VGND VPWR VPWR hold656/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3609 hold38/X VGND VGND VPWR VPWR _5234_/A0 sky130_fd_sc_hd__clkbuf_2
Xhold667 _7115_/Q VGND VGND VPWR VPWR hold667/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold678 _7024_/Q VGND VGND VPWR VPWR hold678/X sky130_fd_sc_hd__dlygate4sd3_1
X_6235_ _6235_/A1 _6310_/A2 _6310_/B1 _6235_/B2 VGND VGND VPWR VPWR _6235_/X sky130_fd_sc_hd__a22o_1
Xhold689 _7025_/Q VGND VGND VPWR VPWR hold689/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3447_ _3447_/A _3447_/B _3447_/C _3447_/D VGND VGND VPWR VPWR _3447_/X sky130_fd_sc_hd__or4_1
Xwire2908 _5940_/A2 VGND VGND VPWR VPWR _5964_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2919 _5695_/A2 VGND VGND VPWR VPWR _5965_/A2 sky130_fd_sc_hd__clkbuf_2
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3378_ _3416_/B _3378_/B VGND VGND VPWR VPWR _3378_/Y sky130_fd_sc_hd__nand2_1
X_6166_ _6166_/A1 _6166_/A2 _6166_/B1 _6967_/Q _6165_/X VGND VGND VPWR VPWR _6167_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5117_ _4971_/A _4783_/Y _4973_/B VGND VGND VPWR VPWR _5117_/X sky130_fd_sc_hd__a21o_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6097_ _7177_/Q _6096_/X _6122_/S VGND VGND VPWR VPWR _7177_/D sky130_fd_sc_hd__mux2_1
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5048_ _5134_/C _5132_/A _5048_/C VGND VGND VPWR VPWR _5048_/X sky130_fd_sc_hd__or3_1
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6999_ _7001_/CLK _6999_/D _7141_/RESET_B VGND VGND VPWR VPWR _6999_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length1221 _3346_/A2 VGND VGND VPWR VPWR _3695_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_107_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4350_ _4654_/A _4350_/B _4542_/A VGND VGND VPWR VPWR _4351_/B sky130_fd_sc_hd__nand3_1
XFILLER_125_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3301_ hold62/X hold26/X _3301_/C VGND VGND VPWR VPWR _3301_/X sky130_fd_sc_hd__or3_1
X_4281_ _4281_/A0 hold486/X _4281_/S VGND VGND VPWR VPWR _6730_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6020_ _6033_/A _6039_/A _6020_/C VGND VGND VPWR VPWR _6020_/X sky130_fd_sc_hd__and3_1
X_3232_ _3232_/A VGND VGND VPWR VPWR _3232_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_113_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6922_ _7127_/CLK _6922_/D _6923_/SET_B VGND VGND VPWR VPWR _6922_/Q sky130_fd_sc_hd__dfstp_1
X_6853_ _6939_/CLK _6853_/D _6407_/A VGND VGND VPWR VPWR hold51/A sky130_fd_sc_hd__dfrtp_1
XFILLER_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5804_ _6158_/B2 _5804_/A2 _5799_/X _5803_/X VGND VGND VPWR VPWR _5804_/X sky130_fd_sc_hd__a211o_1
X_6784_ _6545_/CLK _6784_/D _6435_/X VGND VGND VPWR VPWR _6784_/Q sky130_fd_sc_hd__dfrtn_1
X_3996_ hold562/X _4286_/A0 _4000_/S VGND VGND VPWR VPWR _6493_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5735_ _6884_/Q _5735_/A2 _5735_/B1 _5735_/B2 _5734_/X VGND VGND VPWR VPWR _5735_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5666_ _5683_/A _5706_/C _5703_/C VGND VGND VPWR VPWR _5666_/X sky130_fd_sc_hd__and3_1
XFILLER_136_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4617_ _4420_/A _4667_/C _4569_/A _4800_/A2 _5019_/A VGND VGND VPWR VPWR _5107_/A
+ sky130_fd_sc_hd__a41o_1
X_5597_ _7144_/Q _5604_/D VGND VGND VPWR VPWR _5599_/B sky130_fd_sc_hd__nand2_1
Xhold420 _6601_/Q VGND VGND VPWR VPWR hold420/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire4107 wire4108/X VGND VGND VPWR VPWR wire4107/X sky130_fd_sc_hd__clkbuf_1
Xhold431 _6792_/Q VGND VGND VPWR VPWR hold431/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire4118 wire4118/A VGND VGND VPWR VPWR _3598_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_190_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4548_ _4780_/A _4802_/B _4548_/B1 VGND VGND VPWR VPWR _4963_/A sky130_fd_sc_hd__o21ai_2
Xwire4129 wire4130/X VGND VGND VPWR VPWR wire4129/X sky130_fd_sc_hd__clkbuf_1
Xhold442 _6532_/Q VGND VGND VPWR VPWR hold442/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 _6950_/Q VGND VGND VPWR VPWR hold453/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3406 _3999_/A1 VGND VGND VPWR VPWR _4127_/A0 sky130_fd_sc_hd__clkbuf_1
Xhold464 _6985_/Q VGND VGND VPWR VPWR hold464/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3417 hold43/X VGND VGND VPWR VPWR hold44/A sky130_fd_sc_hd__clkbuf_1
Xhold475 _6722_/Q VGND VGND VPWR VPWR hold475/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3428 _5436_/A0 VGND VGND VPWR VPWR _5199_/A0 sky130_fd_sc_hd__clkbuf_1
Xhold486 _6730_/Q VGND VGND VPWR VPWR hold486/X sky130_fd_sc_hd__dlygate4sd3_1
X_4479_ _4497_/A _4672_/A VGND VGND VPWR VPWR _4823_/A sky130_fd_sc_hd__nor2_1
Xwire3439 _5463_/A0 VGND VGND VPWR VPWR _5256_/A1 sky130_fd_sc_hd__clkbuf_1
Xhold497 _6711_/Q VGND VGND VPWR VPWR hold497/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire2716 _6014_/X VGND VGND VPWR VPWR _6188_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_131_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6218_ _6201_/X _6207_/X _6217_/X wire980/X _6218_/B2 VGND VGND VPWR VPWR _6218_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_58_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7198_ _7204_/CLK _7198_/D wire4260/X VGND VGND VPWR VPWR _7198_/Q sky130_fd_sc_hd__dfrtp_1
Xwire2738 wire2739/X VGND VGND VPWR VPWR _6089_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_38_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2749 _6008_/X VGND VGND VPWR VPWR wire2749/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6149_ _6149_/A1 _6149_/A2 _6149_/B1 _7124_/Q VGND VGND VPWR VPWR _6149_/X sky130_fd_sc_hd__a22o_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length976 wire977/X VGND VGND VPWR VPWR _6342_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_154_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length1073 _3476_/Y VGND VGND VPWR VPWR _3656_/A2 sky130_fd_sc_hd__clkbuf_1
Xfanout3845 wire3848/X VGND VGND VPWR VPWR wire3847/A sky130_fd_sc_hd__clkbuf_2
Xmax_length1084 _3463_/Y VGND VGND VPWR VPWR _4294_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_150_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_728 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3984 wire3985/X VGND VGND VPWR VPWR wire3984/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3995 wire3996/X VGND VGND VPWR VPWR wire3995/X sky130_fd_sc_hd__buf_2
XFILLER_49_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3850_ _3850_/A _3850_/B _6541_/Q VGND VGND VPWR VPWR _3850_/X sky130_fd_sc_hd__or3_1
X_3781_ _3781_/A _3781_/B _3781_/C _3781_/D VGND VGND VPWR VPWR _3789_/C sky130_fd_sc_hd__or4_1
X_5520_ _5520_/A _5520_/B VGND VGND VPWR VPWR _5528_/S sky130_fd_sc_hd__nand2_1
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5451_ _5451_/A0 hold627/X _5453_/S VGND VGND VPWR VPWR _7020_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4402_ _4402_/A _4544_/B _4538_/B VGND VGND VPWR VPWR _4415_/A sky130_fd_sc_hd__and3_1
X_5382_ _5517_/A0 hold520/X _5382_/S VGND VGND VPWR VPWR _6959_/D sky130_fd_sc_hd__mux2_1
X_7121_ _7121_/CLK hold78/X wire4086/X VGND VGND VPWR VPWR _7121_/Q sky130_fd_sc_hd__dfrtp_1
X_4333_ _4333_/A0 hold365/X _4335_/S VGND VGND VPWR VPWR _6773_/D sky130_fd_sc_hd__mux2_1
XFILLER_5_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7052_ _7129_/CLK _7052_/D wire4055/X VGND VGND VPWR VPWR _7052_/Q sky130_fd_sc_hd__dfrtp_1
X_4264_ _4264_/A _4324_/B VGND VGND VPWR VPWR _4269_/S sky130_fd_sc_hd__and2_1
XFILLER_101_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3215_ _3215_/A VGND VGND VPWR VPWR _3215_/Y sky130_fd_sc_hd__inv_2
X_6003_ _6014_/A _6020_/C _6040_/C VGND VGND VPWR VPWR _6003_/X sky130_fd_sc_hd__and3_1
X_4195_ _6652_/Q wire369/X _4196_/S VGND VGND VPWR VPWR _6652_/D sky130_fd_sc_hd__mux2_1
XFILLER_27_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6905_ _7064_/CLK _6905_/D wire4045/X VGND VGND VPWR VPWR _6905_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6836_ _7088_/CLK _6836_/D wire4069/A VGND VGND VPWR VPWR _6836_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6767_ _7066_/CLK _6767_/D _6767_/RESET_B VGND VGND VPWR VPWR _6767_/Q sky130_fd_sc_hd__dfrtp_1
X_3979_ hold42/X _7203_/Q _3979_/S VGND VGND VPWR VPWR hold43/A sky130_fd_sc_hd__mux2_1
Xwire619 wire620/X VGND VGND VPWR VPWR _5492_/S sky130_fd_sc_hd__clkbuf_2
X_5718_ _6067_/B2 _5784_/B1 _5718_/B1 _5718_/B2 _5717_/X VGND VGND VPWR VPWR _5719_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6698_ _7193_/CLK _6698_/D _6780_/RESET_B VGND VGND VPWR VPWR _6698_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_136_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5649_ _7145_/Q _5648_/X _5647_/S _7161_/Q VGND VGND VPWR VPWR _7161_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_164_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold250 _7123_/Q VGND VGND VPWR VPWR hold250/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 _7129_/Q VGND VGND VPWR VPWR hold261/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3214 _5035_/B VGND VGND VPWR VPWR _4526_/B sky130_fd_sc_hd__clkbuf_2
Xhold272 _6742_/Q VGND VGND VPWR VPWR hold272/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3225 _4742_/A VGND VGND VPWR VPWR _4524_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold283 _6537_/Q VGND VGND VPWR VPWR hold283/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold294 _6612_/Q VGND VGND VPWR VPWR hold294/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3236 wire3237/X VGND VGND VPWR VPWR wire3236/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2502 _6204_/B1 VGND VGND VPWR VPWR _6152_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire2513 _6304_/A2 VGND VGND VPWR VPWR _6321_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_78_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2524 _6025_/A VGND VGND VPWR VPWR wire2524/X sky130_fd_sc_hd__clkbuf_1
Xwire2535 _5999_/B1 VGND VGND VPWR VPWR _6301_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1801 _6111_/A1 VGND VGND VPWR VPWR wire1801/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1812 wire1813/X VGND VGND VPWR VPWR wire1812/X sky130_fd_sc_hd__clkbuf_1
Xwire2557 _6092_/A2 VGND VGND VPWR VPWR _6208_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire2568 _6185_/A2 VGND VGND VPWR VPWR _6215_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire1823 _3440_/A1 VGND VGND VPWR VPWR wire1823/X sky130_fd_sc_hd__clkbuf_1
Xwire2579 wire2580/X VGND VGND VPWR VPWR _6320_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire1834 wire1835/X VGND VGND VPWR VPWR _6060_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire1845 _5416_/A1 VGND VGND VPWR VPWR wire1845/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1856 _6983_/Q VGND VGND VPWR VPWR _6155_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1867 _6971_/Q VGND VGND VPWR VPWR _6057_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1878 _5769_/B2 VGND VGND VPWR VPWR _6118_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1889 _6953_/Q VGND VGND VPWR VPWR _6212_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_45_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_101 wire3875/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_112 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_123 input59/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_134 _3936_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_1_1_1_csclk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_167_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3770 _5593_/B VGND VGND VPWR VPWR _5650_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_122_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3781 hold113/X VGND VGND VPWR VPWR _3807_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_68_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire3792 wire3793/X VGND VGND VPWR VPWR wire3792/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput7 mask_rev_in[12] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4951_ _4951_/A _4951_/B _5060_/A VGND VGND VPWR VPWR _5059_/B sky130_fd_sc_hd__and3_1
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3902_ _7157_/Q _7158_/Q VGND VGND VPWR VPWR _6019_/A sky130_fd_sc_hd__nand2b_2
X_4882_ _4882_/A _4882_/B VGND VGND VPWR VPWR _4896_/B sky130_fd_sc_hd__nand2_1
XFILLER_177_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6621_ _7211_/CLK _6621_/D wire3959/X VGND VGND VPWR VPWR _6621_/Q sky130_fd_sc_hd__dfrtp_1
X_3833_ _3832_/X hold81/A _3833_/S VGND VGND VPWR VPWR _6463_/D sky130_fd_sc_hd__mux2_1
XFILLER_192_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6552_ _7131_/CLK hold88/X wire4058/X VGND VGND VPWR VPWR hold87/A sky130_fd_sc_hd__dfrtp_1
X_3764_ _6804_/Q _5200_/A _3761_/X _3763_/X VGND VGND VPWR VPWR _3764_/X sky130_fd_sc_hd__a211o_1
X_5503_ _5503_/A0 hold543/X _5503_/S VGND VGND VPWR VPWR _7066_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6483_ _6824_/CLK _6483_/D _6483_/SET_B VGND VGND VPWR VPWR _6483_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_173_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3695_ _3695_/A1 _3695_/A2 wire793/X _3695_/B2 VGND VGND VPWR VPWR _3695_/X sky130_fd_sc_hd__a22o_1
XFILLER_106_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput300 _6483_/Q VGND VGND VPWR VPWR pll_trim[9] sky130_fd_sc_hd__buf_12
X_5434_ _5452_/A0 hold677/X _5434_/S VGND VGND VPWR VPWR _7005_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput311 _3939_/X VGND VGND VPWR VPWR serial_resetn sky130_fd_sc_hd__buf_12
XFILLER_145_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput322 _6644_/Q VGND VGND VPWR VPWR wb_dat_o[13] sky130_fd_sc_hd__buf_12
Xoutput333 _6633_/Q VGND VGND VPWR VPWR wb_dat_o[23] sky130_fd_sc_hd__buf_12
XFILLER_133_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput344 _6651_/Q VGND VGND VPWR VPWR wb_dat_o[4] sky130_fd_sc_hd__buf_12
XFILLER_114_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5365_ _5365_/A0 hold101/X _5366_/S VGND VGND VPWR VPWR _6944_/D sky130_fd_sc_hd__mux2_1
XFILLER_126_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_3_0_csclk clkbuf_3_3_0_csclk/A VGND VGND VPWR VPWR _7117_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_99_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7104_ _7104_/CLK _7104_/D wire4042/X VGND VGND VPWR VPWR _7104_/Q sky130_fd_sc_hd__dfstp_1
X_4316_ hold612/X _4316_/A1 _4316_/S VGND VGND VPWR VPWR _6759_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5296_ _5554_/A0 hold305/X _5298_/S VGND VGND VPWR VPWR _6882_/D sky130_fd_sc_hd__mux2_1
X_7035_ _7084_/CLK hold73/X _7035_/SET_B VGND VGND VPWR VPWR hold72/A sky130_fd_sc_hd__dfstp_1
Xwire1108 _3650_/B1 VGND VGND VPWR VPWR _3735_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1119 _3777_/B1 VGND VGND VPWR VPWR _3682_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
X_4247_ _4247_/A0 hold172/X _4251_/S VGND VGND VPWR VPWR _6701_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4178_ _4178_/A0 hold257/X _4179_/S VGND VGND VPWR VPWR _6637_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_51_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6819_ _7036_/CLK _6819_/D wire3974/X VGND VGND VPWR VPWR _6819_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire405 wire406/X VGND VGND VPWR VPWR _4084_/S sky130_fd_sc_hd__clkbuf_2
Xwire416 _3764_/X VGND VGND VPWR VPWR wire416/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire427 _3619_/X VGND VGND VPWR VPWR _3633_/A sky130_fd_sc_hd__clkbuf_1
Xwire438 _3491_/X VGND VGND VPWR VPWR wire438/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire449 _6218_/X VGND VGND VPWR VPWR wire449/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3000 _5839_/A2 VGND VGND VPWR VPWR _5798_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_151_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3011 _5677_/X VGND VGND VPWR VPWR wire3011/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3022 wire3022/A VGND VGND VPWR VPWR wire3022/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3033 _5927_/B1 VGND VGND VPWR VPWR _5680_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3044 _5801_/A2 VGND VGND VPWR VPWR _5764_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire2310 _6620_/Q VGND VGND VPWR VPWR _6320_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2321 _6613_/Q VGND VGND VPWR VPWR _3624_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire3066 _5791_/A2 VGND VGND VPWR VPWR _5717_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2332 _4142_/A1 VGND VGND VPWR VPWR wire2332/X sky130_fd_sc_hd__clkbuf_1
Xwire3077 wire3078/X VGND VGND VPWR VPWR wire3077/X sky130_fd_sc_hd__clkbuf_1
Xwire2343 _3670_/A1 VGND VGND VPWR VPWR _6268_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire3088 wire3088/A VGND VGND VPWR VPWR wire3088/X sky130_fd_sc_hd__clkbuf_1
XFILLER_78_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2354 _6540_/Q VGND VGND VPWR VPWR _6335_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2365 _6537_/Q VGND VGND VPWR VPWR wire2365/X sky130_fd_sc_hd__clkbuf_1
Xwire1620 _7077_/Q VGND VGND VPWR VPWR wire1620/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1631 _6133_/A1 VGND VGND VPWR VPWR _5789_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2387 _6329_/B2 VGND VGND VPWR VPWR _3483_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire1642 wire1643/X VGND VGND VPWR VPWR _3594_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2398 _6514_/Q VGND VGND VPWR VPWR _6299_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_46_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1653 wire1654/X VGND VGND VPWR VPWR wire1653/X sky130_fd_sc_hd__clkbuf_1
Xwire1664 wire1665/X VGND VGND VPWR VPWR wire1664/X sky130_fd_sc_hd__clkbuf_1
Xwire1675 wire1676/X VGND VGND VPWR VPWR _3421_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire1686 wire1687/X VGND VGND VPWR VPWR _3639_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_73_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1697 wire1698/X VGND VGND VPWR VPWR wire1697/X sky130_fd_sc_hd__clkbuf_1
XFILLER_74_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire950 _3306_/Y VGND VGND VPWR VPWR wire950/X sky130_fd_sc_hd__dlymetal6s2s_1
Xwire961 wire962/X VGND VGND VPWR VPWR wire961/X sky130_fd_sc_hd__clkbuf_2
Xwire972 _6315_/X VGND VGND VPWR VPWR _6316_/C sky130_fd_sc_hd__clkbuf_1
Xwire983 _6292_/A VGND VGND VPWR VPWR _6316_/A sky130_fd_sc_hd__clkbuf_1
Xwire994 wire995/X VGND VGND VPWR VPWR wire994/X sky130_fd_sc_hd__clkbuf_1
XFILLER_115_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3480_ _6129_/A1 _3480_/A2 _3480_/B1 _6330_/A1 wire823/X VGND VGND VPWR VPWR _3484_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_170_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5150_ _4418_/B _5035_/Y _5036_/Y _4744_/X _5039_/X VGND VGND VPWR VPWR _5174_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4101_ hold386/X _4100_/X _4101_/S VGND VGND VPWR VPWR _6572_/D sky130_fd_sc_hd__mux2_1
XFILLER_69_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5081_ _4679_/B _5027_/B _5080_/X VGND VGND VPWR VPWR _5109_/C sky130_fd_sc_hd__o21ai_1
XFILLER_69_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4032_ hold411/X _4322_/A1 _4032_/S VGND VGND VPWR VPWR _6524_/D sky130_fd_sc_hd__mux2_1
XFILLER_37_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5983_ _6000_/A _6040_/A VGND VGND VPWR VPWR _6021_/B sky130_fd_sc_hd__nand2_1
XFILLER_80_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4934_ _4957_/A _4933_/Y _4842_/Y VGND VGND VPWR VPWR _5065_/D sky130_fd_sc_hd__a21o_1
XFILLER_178_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4865_ _5162_/B _4865_/B _4865_/C _4865_/D VGND VGND VPWR VPWR _4866_/D sky130_fd_sc_hd__or4_1
XANTENNA_12 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_23 wire631/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6604_ _6701_/CLK _6604_/D _6429_/A VGND VGND VPWR VPWR _6604_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA_34 _3625_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3816_ _3820_/A _3821_/S VGND VGND VPWR VPWR _3816_/Y sky130_fd_sc_hd__nor2_1
XFILLER_177_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_45 wire1330/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4796_ _4976_/A1 _4565_/X _4795_/Y _4971_/A VGND VGND VPWR VPWR _4797_/B sky130_fd_sc_hd__a2bb2o_1
XANTENNA_56 wire1544/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_67 _6089_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmax_length2307 _6634_/Q VGND VGND VPWR VPWR _3748_/B2 sky130_fd_sc_hd__clkbuf_1
XANTENNA_78 _6258_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6535_ _6755_/CLK _6535_/D wire3950/X VGND VGND VPWR VPWR _6535_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_89 _6211_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3747_ _3747_/A1 _3747_/A2 _3747_/B1 _3747_/B2 VGND VGND VPWR VPWR _3747_/X sky130_fd_sc_hd__a22o_1
Xmax_length2329 _6609_/Q VGND VGND VPWR VPWR _3575_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_119_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6466_ _3487_/B2 _6466_/D _6421_/X VGND VGND VPWR VPWR hold24/A sky130_fd_sc_hd__dfrtp_1
XFILLER_118_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3678_ _3678_/A1 _3678_/A2 _3678_/B1 _6666_/Q _3677_/X VGND VGND VPWR VPWR _3679_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5417_ _5462_/A0 hold477/X _5417_/S VGND VGND VPWR VPWR _6990_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6397_ _6397_/A0 hold552/X _6397_/S VGND VGND VPWR VPWR _7211_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput174 wire1448/X VGND VGND VPWR VPWR irq[2] sky130_fd_sc_hd__buf_12
X_5348_ _5348_/A0 hold79/X _5348_/S VGND VGND VPWR VPWR hold80/A sky130_fd_sc_hd__mux2_1
Xoutput185 _3215_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[19] sky130_fd_sc_hd__buf_12
Xoutput196 _3205_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[29] sky130_fd_sc_hd__buf_12
XFILLER_101_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5279_ _5522_/A0 hold144/X _5281_/S VGND VGND VPWR VPWR _6867_/D sky130_fd_sc_hd__mux2_1
X_7018_ _7036_/CLK _7018_/D wire3974/A VGND VGND VPWR VPWR _7018_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_28_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length4287 _4591_/A VGND VGND VPWR VPWR _4938_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_109_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2140 wire2141/X VGND VGND VPWR VPWR _3585_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_120_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2151 _6773_/Q VGND VGND VPWR VPWR _6278_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_78_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2162 _6753_/Q VGND VGND VPWR VPWR _6276_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2173 wire2174/X VGND VGND VPWR VPWR wire2173/X sky130_fd_sc_hd__clkbuf_1
Xwire2184 _6743_/Q VGND VGND VPWR VPWR _5911_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1450 wire1451/X VGND VGND VPWR VPWR wire1450/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2195 wire2196/X VGND VGND VPWR VPWR _6274_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire1461 wire1462/X VGND VGND VPWR VPWR wire1461/X sky130_fd_sc_hd__clkbuf_1
Xwire1472 wire1473/X VGND VGND VPWR VPWR wire1472/X sky130_fd_sc_hd__buf_6
Xwire1483 wire1484/X VGND VGND VPWR VPWR wire1483/X sky130_fd_sc_hd__clkbuf_1
XFILLER_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1494 _3416_/Y VGND VGND VPWR VPWR _3519_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_62_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4650_ _5031_/A VGND VGND VPWR VPWR _4650_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput10 mask_rev_in[15] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__clkbuf_1
X_3601_ _3601_/A _3601_/B _3601_/C _3601_/D VGND VGND VPWR VPWR _3601_/X sky130_fd_sc_hd__or4_1
Xinput21 mask_rev_in[25] VGND VGND VPWR VPWR input21/X sky130_fd_sc_hd__clkbuf_1
Xinput32 mask_rev_in[6] VGND VGND VPWR VPWR input32/X sky130_fd_sc_hd__clkbuf_1
X_4581_ _4693_/A _4581_/B VGND VGND VPWR VPWR _4581_/X sky130_fd_sc_hd__or2_2
Xinput43 mgmt_gpio_in[16] VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__clkbuf_1
Xinput54 mgmt_gpio_in[26] VGND VGND VPWR VPWR input54/X sky130_fd_sc_hd__clkbuf_1
X_6320_ _6730_/Q _6320_/A2 _6320_/B1 _6320_/B2 VGND VGND VPWR VPWR _6320_/X sky130_fd_sc_hd__a22o_1
Xinput65 mgmt_gpio_in[36] VGND VGND VPWR VPWR input65/X sky130_fd_sc_hd__clkbuf_1
X_3532_ _6328_/B2 _3532_/A2 wire801/X _6329_/A1 VGND VGND VPWR VPWR _3532_/X sky130_fd_sc_hd__a22o_1
Xwire780 wire781/X VGND VGND VPWR VPWR wire780/X sky130_fd_sc_hd__clkbuf_1
Xwire791 wire792/X VGND VGND VPWR VPWR wire791/X sky130_fd_sc_hd__clkbuf_1
Xinput76 qspi_enabled VGND VGND VPWR VPWR input76/X sky130_fd_sc_hd__clkbuf_1
Xinput87 spimemio_flash_io1_do VGND VGND VPWR VPWR input87/X sky130_fd_sc_hd__clkbuf_1
Xinput98 usr2_vdd_pwrgood VGND VGND VPWR VPWR input98/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6251_ _6522_/Q _6324_/A2 _6324_/B1 _6762_/Q _6250_/X VGND VGND VPWR VPWR _6257_/A
+ sky130_fd_sc_hd__a221o_1
X_3463_ _3482_/A _3485_/B VGND VGND VPWR VPWR _3463_/Y sky130_fd_sc_hd__nor2_1
XFILLER_143_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5202_ _5432_/A0 hold427/X _5202_/S VGND VGND VPWR VPWR _6805_/D sky130_fd_sc_hd__mux2_1
X_6182_ _6182_/A1 _6182_/A2 _6182_/B1 _6182_/B2 _6181_/X VGND VGND VPWR VPWR _6182_/X
+ sky130_fd_sc_hd__a221o_1
X_3394_ _3394_/A1 _3394_/A2 _5466_/A _3394_/B2 _3382_/X VGND VGND VPWR VPWR _3394_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5133_ _5133_/A1 _5133_/A2 _4670_/Y _4897_/C VGND VGND VPWR VPWR _5134_/D sky130_fd_sc_hd__a211o_1
XFILLER_111_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5064_ _5064_/A _5064_/B _5064_/C _5064_/D VGND VGND VPWR VPWR _5125_/A sky130_fd_sc_hd__or4_1
X_4015_ hold669/X _6397_/A0 _4015_/S VGND VGND VPWR VPWR _6510_/D sky130_fd_sc_hd__mux2_1
XFILLER_37_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5966_ _6625_/Q _5966_/A2 _5966_/B1 _6329_/B2 _5965_/X VGND VGND VPWR VPWR _5967_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4917_ _4694_/A _5027_/A _5115_/B VGND VGND VPWR VPWR _5109_/A sky130_fd_sc_hd__o21bai_1
XFILLER_178_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5897_ _6259_/B2 _5897_/A2 _5897_/B1 _6676_/Q VGND VGND VPWR VPWR _5897_/X sky130_fd_sc_hd__a22o_1
XFILLER_178_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4848_ _4848_/A1 _4677_/B _5049_/A VGND VGND VPWR VPWR _4865_/B sky130_fd_sc_hd__o21bai_1
XFILLER_165_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4779_ _4484_/A _5072_/A3 _4794_/A VGND VGND VPWR VPWR _5095_/B sky130_fd_sc_hd__a21oi_1
XFILLER_193_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6518_ _6701_/CLK _6518_/D wire3945/X VGND VGND VPWR VPWR _6518_/Q sky130_fd_sc_hd__dfstp_1
Xmax_length1403 _3255_/X VGND VGND VPWR VPWR _3657_/A1_N sky130_fd_sc_hd__clkbuf_1
Xmax_length1436 _5002_/A VGND VGND VPWR VPWR _4520_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_134_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length1447 _4417_/X VGND VGND VPWR VPWR _4876_/A sky130_fd_sc_hd__clkbuf_1
X_6449_ _3927_/A1 _6449_/D _6404_/X VGND VGND VPWR VPWR hold14/A sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_40_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7017_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_0_0_csclk clkbuf_2_1_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_1_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_75_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_55_csclk _7117_/CLK VGND VGND VPWR VPWR _7102_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4051 wire4052/X VGND VGND VPWR VPWR _7035_/SET_B sky130_fd_sc_hd__buf_2
Xmax_length4062 fanout4054/A VGND VGND VPWR VPWR wire4061/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length4084 _7075_/SET_B VGND VGND VPWR VPWR fanout4047/A sky130_fd_sc_hd__clkbuf_1
XFILLER_157_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length3350 _4451_/B VGND VGND VPWR VPWR _5043_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_184_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1280 _3646_/A2 VGND VGND VPWR VPWR _3420_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1291 _3531_/A VGND VGND VPWR VPWR _3502_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5820_ _6864_/Q _5820_/A2 _5820_/B1 _6191_/A1 _5819_/X VGND VGND VPWR VPWR _5825_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5751_ _6844_/Q _5793_/A2 _5740_/X _5750_/X _6095_/C1 VGND VGND VPWR VPWR _5751_/X
+ sky130_fd_sc_hd__o221a_1
X_4702_ _4704_/A _4683_/B _4920_/B1 _4624_/B VGND VGND VPWR VPWR _4702_/X sky130_fd_sc_hd__o22a_1
XFILLER_148_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5682_ _7152_/Q _5699_/B _5706_/C VGND VGND VPWR VPWR _5682_/X sky130_fd_sc_hd__and3_1
XFILLER_147_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4633_ _4638_/B _4633_/B VGND VGND VPWR VPWR _4982_/A sky130_fd_sc_hd__nor2_1
XFILLER_163_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4564_ _4476_/A _4564_/B _4588_/B VGND VGND VPWR VPWR _4666_/B sky130_fd_sc_hd__nand3b_2
Xhold602 _7050_/Q VGND VGND VPWR VPWR hold602/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold613 _6756_/Q VGND VGND VPWR VPWR hold613/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold624 _7087_/Q VGND VGND VPWR VPWR hold624/X sky130_fd_sc_hd__dlygate4sd3_1
X_6303_ _6303_/A1 _6334_/B1 _6303_/B1 _6303_/B2 VGND VGND VPWR VPWR _6303_/X sky130_fd_sc_hd__a22o_1
Xhold635 _6529_/Q VGND VGND VPWR VPWR hold635/X sky130_fd_sc_hd__dlygate4sd3_1
X_3515_ _3515_/A _3515_/B _3515_/C _3515_/D VGND VGND VPWR VPWR _3542_/B sky130_fd_sc_hd__or4_1
XFILLER_155_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold646 _6548_/Q VGND VGND VPWR VPWR hold646/X sky130_fd_sc_hd__dlygate4sd3_1
X_4495_ _4495_/A _4495_/B VGND VGND VPWR VPWR _4496_/B sky130_fd_sc_hd__nand2_1
XFILLER_89_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold657 _6598_/Q VGND VGND VPWR VPWR hold657/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold668 _7041_/Q VGND VGND VPWR VPWR hold668/X sky130_fd_sc_hd__dlygate4sd3_1
X_6234_ _6234_/A1 _6309_/A2 _6309_/B1 _6234_/B2 _6233_/X VGND VGND VPWR VPWR _6242_/B
+ sky130_fd_sc_hd__a221o_1
Xhold679 _6559_/Q VGND VGND VPWR VPWR hold679/X sky130_fd_sc_hd__dlygate4sd3_1
X_3446_ _3446_/A _3446_/B _3446_/C _3446_/D VGND VGND VPWR VPWR _3446_/X sky130_fd_sc_hd__or4_1
Xwire2909 _5695_/B1 VGND VGND VPWR VPWR _5940_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_131_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ _6165_/A1 _6172_/A2 _6174_/A2 _6903_/Q VGND VGND VPWR VPWR _6165_/X sky130_fd_sc_hd__a22o_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3377_ _3472_/A _3526_/A VGND VGND VPWR VPWR _3658_/A sky130_fd_sc_hd__nor2_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5116_ _4454_/Y _4729_/Y _4988_/D _5091_/X _5115_/X VGND VGND VPWR VPWR _5172_/A
+ sky130_fd_sc_hd__a2111o_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6096_ _6121_/A1 _7176_/Q wire453/X VGND VGND VPWR VPWR _6096_/X sky130_fd_sc_hd__a21o_1
XFILLER_57_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5047_ _5049_/A _5049_/B _5049_/C _5049_/D VGND VGND VPWR VPWR _5048_/C sky130_fd_sc_hd__or4_1
XFILLER_38_550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6998_ _7115_/CLK _6998_/D _7030_/RESET_B VGND VGND VPWR VPWR _6998_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_13_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5949_ _6336_/B2 _5949_/A2 _5949_/B1 _6765_/Q VGND VGND VPWR VPWR _5949_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length1266 _3295_/Y VGND VGND VPWR VPWR wire1265/A sky130_fd_sc_hd__clkbuf_1
XFILLER_134_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3300_ _3476_/A hold85/X VGND VGND VPWR VPWR _3300_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4280_ _5566_/A0 hold371/X _4281_/S VGND VGND VPWR VPWR _6729_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3231_ _3231_/A VGND VGND VPWR VPWR _3231_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6921_ _6921_/CLK _6921_/D wire4046/X VGND VGND VPWR VPWR _6921_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6852_ _7129_/CLK _6852_/D wire4055/X VGND VGND VPWR VPWR _6852_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5803_ _6153_/A1 _5803_/A2 _5800_/X _5802_/X VGND VGND VPWR VPWR _5803_/X sky130_fd_sc_hd__a211o_1
XFILLER_22_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6783_ _3487_/B2 _6783_/D _6434_/X VGND VGND VPWR VPWR _6783_/Q sky130_fd_sc_hd__dfrtn_1
X_3995_ hold572/X _5196_/A0 _4000_/S VGND VGND VPWR VPWR _6492_/D sky130_fd_sc_hd__mux2_1
X_5734_ _5734_/A1 _5790_/B1 _5734_/B1 _6077_/A1 VGND VGND VPWR VPWR _5734_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5665_ _6004_/A1 _5727_/A2 _5716_/A2 _6011_/A1 VGND VGND VPWR VPWR _5665_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4616_ _5023_/C _4673_/A VGND VGND VPWR VPWR _5019_/A sky130_fd_sc_hd__nor2_1
X_5596_ _6565_/Q _5596_/B _5651_/B VGND VGND VPWR VPWR _5606_/A sky130_fd_sc_hd__or3_1
Xhold410 _7097_/Q VGND VGND VPWR VPWR hold410/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire4108 wire4109/X VGND VGND VPWR VPWR wire4108/X sky130_fd_sc_hd__clkbuf_1
X_4547_ _4547_/A _4573_/B VGND VGND VPWR VPWR _4802_/B sky130_fd_sc_hd__or2_1
Xhold421 _6957_/Q VGND VGND VPWR VPWR hold421/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 _6688_/Q VGND VGND VPWR VPWR hold432/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 _6531_/Q VGND VGND VPWR VPWR hold443/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold454 _6886_/Q VGND VGND VPWR VPWR hold454/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3407 wire3408/X VGND VGND VPWR VPWR _3999_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_104_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold465 _6658_/Q VGND VGND VPWR VPWR hold465/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4478_ _4672_/A VGND VGND VPWR VPWR _4478_/Y sky130_fd_sc_hd__inv_2
Xwire3429 _5454_/A0 VGND VGND VPWR VPWR _5436_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold476 _6955_/Q VGND VGND VPWR VPWR hold476/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 _7055_/Q VGND VGND VPWR VPWR hold487/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold498 _7100_/Q VGND VGND VPWR VPWR hold498/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire2706 _6184_/B1 VGND VGND VPWR VPWR _6203_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6217_ _6217_/A _6217_/B _6217_/C _6217_/D VGND VGND VPWR VPWR _6217_/X sky130_fd_sc_hd__or4_1
Xwire2717 _6310_/A2 VGND VGND VPWR VPWR _6283_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
X_3429_ _6158_/A1 _5553_/A _5544_/A _6152_/B2 _3424_/X VGND VGND VPWR VPWR _3431_/C
+ sky130_fd_sc_hd__a221o_1
X_7197_ _7204_/CLK _7197_/D wire4260/X VGND VGND VPWR VPWR _7197_/Q sky130_fd_sc_hd__dfrtp_1
Xwire2739 _6023_/C VGND VGND VPWR VPWR wire2739/X sky130_fd_sc_hd__clkbuf_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6148_ _6148_/A _6148_/B VGND VGND VPWR VPWR _6148_/X sky130_fd_sc_hd__and2_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6079_ _6900_/Q _6126_/A2 _6079_/B1 _6079_/B2 _6078_/X VGND VGND VPWR VPWR _6084_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_523 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length1030 _4222_/A VGND VGND VPWR VPWR _3609_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_5_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3930 wire3931/X VGND VGND VPWR VPWR wire3930/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3963 wire3963/A VGND VGND VPWR VPWR _6437_/A sky130_fd_sc_hd__clkbuf_2
Xwire3974 wire3974/A VGND VGND VPWR VPWR wire3974/X sky130_fd_sc_hd__buf_2
XFILLER_1_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3985 wire3985/A VGND VGND VPWR VPWR wire3985/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3996 wire3996/A VGND VGND VPWR VPWR wire3996/X sky130_fd_sc_hd__buf_2
XFILLER_95_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3780_ _3780_/A1 _3268_/Y _3780_/B1 _6234_/B2 wire739/X VGND VGND VPWR VPWR _3781_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_9_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5450_ _5450_/A0 hold402/X _5450_/S VGND VGND VPWR VPWR _7019_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4401_ _4451_/A _4538_/B VGND VGND VPWR VPWR _4739_/A sky130_fd_sc_hd__nand2_2
XFILLER_145_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5381_ _5381_/A0 hold126/X _5381_/S VGND VGND VPWR VPWR _6958_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A VGND VGND VPWR VPWR _7180_/CLK sky130_fd_sc_hd__clkbuf_8
X_7120_ _7136_/CLK _7120_/D wire4086/X VGND VGND VPWR VPWR _7120_/Q sky130_fd_sc_hd__dfstp_1
X_4332_ _5231_/A0 hold364/X _4335_/S VGND VGND VPWR VPWR _6772_/D sky130_fd_sc_hd__mux2_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7051_ _7135_/CLK _7051_/D _7051_/SET_B VGND VGND VPWR VPWR _7051_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4263_ _4263_/A0 _4263_/A1 _4263_/S VGND VGND VPWR VPWR _6715_/D sky130_fd_sc_hd__mux2_1
XFILLER_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6002_ _6018_/A _6038_/A VGND VGND VPWR VPWR _6002_/Y sky130_fd_sc_hd__nor2_1
X_3214_ _3214_/A VGND VGND VPWR VPWR _3214_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4194_ _6651_/Q _4194_/A1 _4196_/S VGND VGND VPWR VPWR _6651_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6904_ _7088_/CLK _6904_/D wire4069/A VGND VGND VPWR VPWR _6904_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_82_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6835_ _6945_/CLK _6835_/D fanout4078/X VGND VGND VPWR VPWR _6835_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6766_ _6775_/CLK _6766_/D wire3981/A VGND VGND VPWR VPWR _6766_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3978_ hold626/X _5436_/A0 _3982_/S VGND VGND VPWR VPWR _6479_/D sky130_fd_sc_hd__mux2_1
Xwire609 _5495_/S VGND VGND VPWR VPWR _5494_/S sky130_fd_sc_hd__clkbuf_1
X_5717_ _6048_/B2 _5717_/A2 _5717_/B1 _6061_/B2 VGND VGND VPWR VPWR _5717_/X sky130_fd_sc_hd__a22o_1
XFILLER_164_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6697_ _7206_/CLK _6697_/D _4189_/B VGND VGND VPWR VPWR _6697_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5648_ _7146_/Q _7147_/Q _5648_/C _7144_/Q VGND VGND VPWR VPWR _5648_/X sky130_fd_sc_hd__or4b_1
XFILLER_108_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5579_ _5579_/A0 hold212/X _5579_/S VGND VGND VPWR VPWR _7134_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold240 _6819_/Q VGND VGND VPWR VPWR _5221_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold251 _7078_/Q VGND VGND VPWR VPWR hold251/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 _6513_/Q VGND VGND VPWR VPWR hold262/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3204 _4728_/B VGND VGND VPWR VPWR _4870_/B sky130_fd_sc_hd__clkbuf_2
Xhold273 _4296_/X VGND VGND VPWR VPWR _6742_/D sky130_fd_sc_hd__dlygate4sd3_1
Xwire3226 _4387_/Y VGND VGND VPWR VPWR _4981_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_132_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3237 _4232_/X VGND VGND VPWR VPWR wire3237/X sky130_fd_sc_hd__clkbuf_1
Xhold284 _6568_/Q VGND VGND VPWR VPWR hold284/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire2503 _6181_/A2 VGND VGND VPWR VPWR _6204_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold295 _6615_/Q VGND VGND VPWR VPWR hold295/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire2514 _6278_/A2 VGND VGND VPWR VPWR _6304_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3259 _4240_/B VGND VGND VPWR VPWR _4246_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2525 _6112_/B1 VGND VGND VPWR VPWR _6005_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire2536 _5998_/Y VGND VGND VPWR VPWR _5999_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2547 _5997_/Y VGND VGND VPWR VPWR _5999_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1802 _5759_/A1 VGND VGND VPWR VPWR _6111_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1813 _5432_/A1 VGND VGND VPWR VPWR wire1813/X sky130_fd_sc_hd__clkbuf_1
Xwire2558 _6338_/A2 VGND VGND VPWR VPWR _6092_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1824 _6999_/Q VGND VGND VPWR VPWR _3440_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2569 _5980_/Y VGND VGND VPWR VPWR _6185_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1835 wire1836/X VGND VGND VPWR VPWR wire1835/X sky130_fd_sc_hd__clkbuf_1
Xwire1846 wire1847/X VGND VGND VPWR VPWR _3216_/A sky130_fd_sc_hd__clkbuf_1
Xwire1857 _6981_/Q VGND VGND VPWR VPWR _3217_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_85_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1868 _6970_/Q VGND VGND VPWR VPWR _5692_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire1879 _6965_/Q VGND VGND VPWR VPWR _5769_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_102 _3937_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_113 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_124 _3658_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length796 _3546_/Y VGND VGND VPWR VPWR wire795/A sky130_fd_sc_hd__clkbuf_1
XFILLER_108_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout3610 hold36/X VGND VGND VPWR VPWR hold37/A sky130_fd_sc_hd__clkbuf_1
XFILLER_170_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout3621 wire3628/A VGND VGND VPWR VPWR _6393_/A0 sky130_fd_sc_hd__buf_6
XFILLER_5_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout3643 wire3652/A VGND VGND VPWR VPWR _5476_/A0 sky130_fd_sc_hd__buf_6
Xfanout3654 hold153/X VGND VGND VPWR VPWR wire3661/A sky130_fd_sc_hd__buf_6
XFILLER_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3760 _3963_/B VGND VGND VPWR VPWR _3941_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_150_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3771 _6194_/C1 VGND VGND VPWR VPWR _6121_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_96_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3782 wire3783/X VGND VGND VPWR VPWR _3928_/S sky130_fd_sc_hd__clkbuf_2
Xwire3793 _6461_/Q VGND VGND VPWR VPWR wire3793/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput8 mask_rev_in[13] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4950_ _4947_/Y _4950_/B _4950_/C VGND VGND VPWR VPWR _4954_/B sky130_fd_sc_hd__nand3b_1
X_3901_ _6564_/Q _5596_/B VGND VGND VPWR VPWR _6563_/D sky130_fd_sc_hd__or2_1
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4881_ _4396_/X _4740_/Y _4453_/A VGND VGND VPWR VPWR _4885_/B sky130_fd_sc_hd__a21oi_1
X_6620_ _7208_/CLK _6620_/D wire4026/X VGND VGND VPWR VPWR _6620_/Q sky130_fd_sc_hd__dfrtp_1
X_3832_ _3830_/A _3832_/A1 _3850_/A VGND VGND VPWR VPWR _3832_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6551_ _7131_/CLK _6551_/D wire4055/X VGND VGND VPWR VPWR _6551_/Q sky130_fd_sc_hd__dfrtp_1
X_3763_ input4/X _3763_/A2 _3763_/B1 _7002_/Q _3762_/X VGND VGND VPWR VPWR _3763_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5502_ _5502_/A _5502_/B VGND VGND VPWR VPWR _5507_/S sky130_fd_sc_hd__nand2_1
X_6482_ _6825_/CLK _6482_/D wire3956/X VGND VGND VPWR VPWR _6482_/Q sky130_fd_sc_hd__dfstp_1
X_3694_ _3694_/A1 wire970/X wire896/X _6059_/A1 wire762/X VGND VGND VPWR VPWR _3701_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_145_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5433_ _5469_/A1 hold644/X _5434_/S VGND VGND VPWR VPWR _7004_/D sky130_fd_sc_hd__mux2_1
Xoutput301 _6807_/Q VGND VGND VPWR VPWR pwr_ctrl_out[0] sky130_fd_sc_hd__buf_12
XFILLER_105_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput312 _3958_/X VGND VGND VPWR VPWR spi_sdi sky130_fd_sc_hd__buf_12
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput323 _6645_/Q VGND VGND VPWR VPWR wb_dat_o[14] sky130_fd_sc_hd__buf_12
XFILLER_160_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5364_ _5364_/A0 hold685/X _5366_/S VGND VGND VPWR VPWR _6943_/D sky130_fd_sc_hd__mux2_1
Xoutput334 _7189_/Q VGND VGND VPWR VPWR wb_dat_o[24] sky130_fd_sc_hd__buf_12
Xoutput345 _6652_/Q VGND VGND VPWR VPWR wb_dat_o[5] sky130_fd_sc_hd__buf_12
XFILLER_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7103_ _7127_/CLK _7103_/D wire4061/A VGND VGND VPWR VPWR _7103_/Q sky130_fd_sc_hd__dfstp_1
X_4315_ hold620/X _4327_/A1 _4316_/S VGND VGND VPWR VPWR _6758_/D sky130_fd_sc_hd__mux2_1
X_5295_ _5295_/A _5403_/B VGND VGND VPWR VPWR _5298_/S sky130_fd_sc_hd__nand2_2
XFILLER_99_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7034_ _7074_/CLK _7034_/D wire3974/X VGND VGND VPWR VPWR _7034_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_113_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4246_ _4246_/A _4246_/B VGND VGND VPWR VPWR _4251_/S sky130_fd_sc_hd__nand2_2
Xwire1109 _3344_/Y VGND VGND VPWR VPWR _3650_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_28_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4177_ _4255_/A1 _6636_/Q _4179_/S VGND VGND VPWR VPWR _4177_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6818_ _7080_/CLK _6818_/D wire3992/A VGND VGND VPWR VPWR _6818_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire406 wire407/X VGND VGND VPWR VPWR wire406/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire417 _3757_/X VGND VGND VPWR VPWR _3760_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_149_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6749_ _6963_/CLK _6749_/D _6401_/A VGND VGND VPWR VPWR _6749_/Q sky130_fd_sc_hd__dfrtp_1
Xwire428 _3593_/X VGND VGND VPWR VPWR _3601_/C sky130_fd_sc_hd__clkbuf_1
Xwire439 _3444_/X VGND VGND VPWR VPWR _3445_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3001 _5760_/A2 VGND VGND VPWR VPWR _5885_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire3012 _5856_/A2 VGND VGND VPWR VPWR _5811_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_183_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3023 _5756_/B1 VGND VGND VPWR VPWR _5775_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3034 _5962_/B1 VGND VGND VPWR VPWR _5927_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire2300 _6284_/B2 VGND VGND VPWR VPWR _5911_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire3045 _5840_/A2 VGND VGND VPWR VPWR _5801_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire3056 wire3057/X VGND VGND VPWR VPWR _5852_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire2311 _6619_/Q VGND VGND VPWR VPWR _6296_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire2322 _6612_/Q VGND VGND VPWR VPWR _6265_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3067 _5853_/B1 VGND VGND VPWR VPWR _5791_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3078 _5844_/A2 VGND VGND VPWR VPWR wire3078/X sky130_fd_sc_hd__clkbuf_1
XFILLER_120_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2344 _6597_/Q VGND VGND VPWR VPWR _3670_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire2355 _6300_/A1 VGND VGND VPWR VPWR _5933_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1610 _7084_/Q VGND VGND VPWR VPWR _6076_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2366 _6224_/A1 VGND VGND VPWR VPWR _5877_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire1621 wire1622/X VGND VGND VPWR VPWR _3590_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2377 _3554_/B2 VGND VGND VPWR VPWR _6312_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1632 _7070_/Q VGND VGND VPWR VPWR _6133_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1643 _5761_/B2 VGND VGND VPWR VPWR wire1643/X sky130_fd_sc_hd__clkbuf_1
Xwire2388 _6520_/Q VGND VGND VPWR VPWR _6329_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_74_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1654 wire1655/X VGND VGND VPWR VPWR wire1654/X sky130_fd_sc_hd__clkbuf_1
Xwire1665 _6105_/B2 VGND VGND VPWR VPWR wire1665/X sky130_fd_sc_hd__clkbuf_1
XFILLER_46_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1676 _5809_/B2 VGND VGND VPWR VPWR wire1676/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1687 _5747_/A1 VGND VGND VPWR VPWR wire1687/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1698 _7041_/Q VGND VGND VPWR VPWR wire1698/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire940 wire941/X VGND VGND VPWR VPWR wire940/X sky130_fd_sc_hd__clkbuf_1
Xwire951 wire953/X VGND VGND VPWR VPWR wire951/X sky130_fd_sc_hd__clkbuf_1
Xwire962 _3278_/Y VGND VGND VPWR VPWR wire962/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire973 wire974/X VGND VGND VPWR VPWR _6292_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_182_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire984 _6341_/A VGND VGND VPWR VPWR _6267_/A sky130_fd_sc_hd__clkbuf_1
Xwire995 _5770_/X VGND VGND VPWR VPWR wire995/X sky130_fd_sc_hd__clkbuf_1
XFILLER_170_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire4280 _4564_/B VGND VGND VPWR VPWR _4935_/A sky130_fd_sc_hd__clkbuf_2
Xwire4291 _4565_/A VGND VGND VPWR VPWR _4621_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4100_ hold105/X _5374_/A0 _4100_/S VGND VGND VPWR VPWR _4100_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5080_ _5027_/A _5108_/B _4922_/B VGND VGND VPWR VPWR _5080_/X sky130_fd_sc_hd__o21ba_1
Xwire3590 _4200_/A1 VGND VGND VPWR VPWR _5504_/A0 sky130_fd_sc_hd__clkbuf_2
X_4031_ hold396/X _4321_/A1 _4033_/S VGND VGND VPWR VPWR _6523_/D sky130_fd_sc_hd__mux2_1
XFILLER_111_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5982_ _6040_/A _6039_/A _6020_/C VGND VGND VPWR VPWR _5982_/X sky130_fd_sc_hd__and3_1
XFILLER_24_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4933_ _4933_/A _4935_/C VGND VGND VPWR VPWR _4933_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4864_ _5064_/A _5124_/B _4864_/C _4864_/D VGND VGND VPWR VPWR _4865_/D sky130_fd_sc_hd__or4_1
XFILLER_178_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_13 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_24 wire738/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6603_ _6701_/CLK _6603_/D wire3945/X VGND VGND VPWR VPWR _6603_/Q sky130_fd_sc_hd__dfrtp_1
X_3815_ _3814_/X hold60/A _3828_/S VGND VGND VPWR VPWR _6469_/D sky130_fd_sc_hd__mux2_1
XANTENNA_35 _3625_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4795_ _4802_/D _4795_/B VGND VGND VPWR VPWR _4795_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_46 _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_57 _6158_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6534_ _6755_/CLK _6534_/D wire3950/X VGND VGND VPWR VPWR _6534_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_68 wire1816/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_79 wire2225/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3746_ _3746_/A1 _3746_/A2 _4153_/A _6221_/B2 wire745/X VGND VGND VPWR VPWR _3749_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6465_ _3487_/B2 _6465_/D _6420_/X VGND VGND VPWR VPWR hold66/A sky130_fd_sc_hd__dfrtp_1
X_3677_ _6265_/A1 _4147_/A _3677_/B1 _6264_/A1 VGND VGND VPWR VPWR _3677_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5416_ _5416_/A0 _5416_/A1 _5416_/S VGND VGND VPWR VPWR _6989_/D sky130_fd_sc_hd__mux2_1
XFILLER_106_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6396_ _6396_/A0 _7210_/Q _6396_/S VGND VGND VPWR VPWR _6396_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5347_ _5365_/A0 hold99/X _5348_/S VGND VGND VPWR VPWR _6928_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput175 wire1350/X VGND VGND VPWR VPWR mgmt_gpio_oeb[0] sky130_fd_sc_hd__buf_12
XFILLER_99_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput186 wire1354/X VGND VGND VPWR VPWR mgmt_gpio_oeb[1] sky130_fd_sc_hd__buf_12
Xoutput197 _3231_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[2] sky130_fd_sc_hd__buf_12
XFILLER_114_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5278_ _5359_/A0 hold324/X _5281_/S VGND VGND VPWR VPWR _6866_/D sky130_fd_sc_hd__mux2_1
X_7017_ _7017_/CLK _7017_/D wire4081/X VGND VGND VPWR VPWR _7017_/Q sky130_fd_sc_hd__dfrtp_1
X_4229_ _6699_/Q _6698_/Q _6700_/Q VGND VGND VPWR VPWR _4232_/B sky130_fd_sc_hd__or3_1
XFILLER_28_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length3521 _5389_/A0 VGND VGND VPWR VPWR _5380_/A0 sky130_fd_sc_hd__clkbuf_1
Xmax_length3554 _5505_/A0 VGND VGND VPWR VPWR _5583_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_109_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length3576 hold21/X VGND VGND VPWR VPWR wire3575/A sky130_fd_sc_hd__clkbuf_1
XFILLER_164_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2130 wire2131/X VGND VGND VPWR VPWR _3757_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire2141 _6801_/Q VGND VGND VPWR VPWR wire2141/X sky130_fd_sc_hd__clkbuf_1
Xwire2152 wire2152/A VGND VGND VPWR VPWR _5887_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_38_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2163 wire2164/X VGND VGND VPWR VPWR _6252_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_78_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2174 _3626_/B2 VGND VGND VPWR VPWR wire2174/X sky130_fd_sc_hd__clkbuf_1
Xwire1440 _4434_/X VGND VGND VPWR VPWR _5113_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2185 _6259_/B2 VGND VGND VPWR VPWR _3664_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_120_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1451 _3960_/X VGND VGND VPWR VPWR wire1451/X sky130_fd_sc_hd__clkbuf_1
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2196 _6738_/Q VGND VGND VPWR VPWR wire2196/X sky130_fd_sc_hd__clkbuf_1
Xwire1462 _3929_/X VGND VGND VPWR VPWR wire1462/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1473 wire1474/X VGND VGND VPWR VPWR wire1473/X sky130_fd_sc_hd__clkbuf_1
Xwire1484 wire1485/X VGND VGND VPWR VPWR wire1484/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1495 _3456_/B VGND VGND VPWR VPWR _3525_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3600_ _3600_/A _3600_/B _3600_/C _3600_/D VGND VGND VPWR VPWR _3601_/D sky130_fd_sc_hd__or4_1
XFILLER_159_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput11 mask_rev_in[16] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__clkbuf_1
Xinput22 mask_rev_in[26] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__clkbuf_1
X_4580_ _4661_/B _4581_/B VGND VGND VPWR VPWR _4684_/B sky130_fd_sc_hd__nor2_1
Xinput33 mask_rev_in[7] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__clkbuf_1
Xinput44 mgmt_gpio_in[17] VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput55 mgmt_gpio_in[27] VGND VGND VPWR VPWR input55/X sky130_fd_sc_hd__clkbuf_1
X_3531_ _3531_/A _4120_/B VGND VGND VPWR VPWR _3531_/Y sky130_fd_sc_hd__nor2_1
Xwire770 wire771/X VGND VGND VPWR VPWR wire770/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire781 wire782/X VGND VGND VPWR VPWR wire781/X sky130_fd_sc_hd__clkbuf_1
Xinput66 mgmt_gpio_in[37] VGND VGND VPWR VPWR input66/X sky130_fd_sc_hd__clkbuf_1
Xinput77 ser_tx VGND VGND VPWR VPWR input77/X sky130_fd_sc_hd__clkbuf_1
Xwire792 _3546_/Y VGND VGND VPWR VPWR wire792/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput88 spimemio_flash_io1_oeb VGND VGND VPWR VPWR input88/X sky130_fd_sc_hd__clkbuf_1
Xinput99 wb_adr_i[0] VGND VGND VPWR VPWR input99/X sky130_fd_sc_hd__clkbuf_1
XFILLER_182_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6250_ _6250_/A1 _6274_/A2 _6323_/B1 _6250_/B2 VGND VGND VPWR VPWR _6250_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3462_ _3462_/A _3534_/A VGND VGND VPWR VPWR _4306_/A sky130_fd_sc_hd__nor2_2
X_5201_ _5467_/A1 hold414/X _5202_/S VGND VGND VPWR VPWR _6804_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6181_ _7109_/Q _6181_/A2 _6181_/B1 _6181_/B2 VGND VGND VPWR VPWR _6181_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3393_ _7072_/Q _3393_/A2 _3393_/B1 _6189_/A1 _3383_/X VGND VGND VPWR VPWR _3393_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5132_ _5132_/A _5132_/B VGND VGND VPWR VPWR _5151_/B sky130_fd_sc_hd__or2_1
XFILLER_97_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5063_ _4659_/A _5027_/A _4515_/C VGND VGND VPWR VPWR _5064_/D sky130_fd_sc_hd__o21ai_1
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4014_ hold555/X _4139_/A1 _4014_/S VGND VGND VPWR VPWR _6509_/D sky130_fd_sc_hd__mux2_1
XFILLER_37_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5965_ _6659_/Q _5965_/A2 _5965_/B1 _6510_/Q VGND VGND VPWR VPWR _5965_/X sky130_fd_sc_hd__a22o_1
XFILLER_52_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4916_ _4916_/A _4916_/B VGND VGND VPWR VPWR _5153_/A sky130_fd_sc_hd__nand2_1
X_5896_ _6762_/Q _5921_/A2 _5896_/B1 _6522_/Q _5895_/X VGND VGND VPWR VPWR _5901_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_138_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4847_ _4847_/A _4882_/B VGND VGND VPWR VPWR _4847_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4778_ _4778_/A _4778_/B VGND VGND VPWR VPWR _4778_/Y sky130_fd_sc_hd__nand2_1
XFILLER_165_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6517_ _7090_/CLK _6517_/D wire3945/A VGND VGND VPWR VPWR _6517_/Q sky130_fd_sc_hd__dfrtp_1
X_3729_ _5212_/A _3729_/B VGND VGND VPWR VPWR _5203_/A sky130_fd_sc_hd__nor2_1
XFILLER_134_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length1437 _5002_/A VGND VGND VPWR VPWR _4958_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_106_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6448_ _3927_/A1 _6448_/D _6403_/X VGND VGND VPWR VPWR hold47/A sky130_fd_sc_hd__dfrtp_1
XFILLER_164_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6379_ _4228_/C _6379_/A2 _6379_/B1 _4228_/A _6378_/X VGND VGND VPWR VPWR _6379_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length4030 fanout4028/X VGND VGND VPWR VPWR wire4029/A sky130_fd_sc_hd__buf_4
XFILLER_156_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length4063 fanout4060/X VGND VGND VPWR VPWR fanout4054/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length4074 fanout4073/X VGND VGND VPWR VPWR _7047_/RESET_B sky130_fd_sc_hd__clkbuf_2
Xmax_length4085 wire4086/X VGND VGND VPWR VPWR _7075_/SET_B sky130_fd_sc_hd__clkbuf_2
XFILLER_144_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_length1993 _6896_/Q VGND VGND VPWR VPWR _5824_/A1 sky130_fd_sc_hd__clkbuf_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1281 _3290_/Y VGND VGND VPWR VPWR _3646_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_35_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1292 _3451_/A VGND VGND VPWR VPWR _3531_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5750_ _5750_/A _5750_/B _5750_/C _5750_/D VGND VGND VPWR VPWR _5750_/X sky130_fd_sc_hd__or4_1
XFILLER_15_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4701_ _4709_/A1 _4661_/B _4624_/B _4699_/X _4700_/X VGND VGND VPWR VPWR _4701_/X
+ sky130_fd_sc_hd__o311a_1
X_5681_ _5681_/A _5681_/B _5681_/C _5681_/D VGND VGND VPWR VPWR _5681_/X sky130_fd_sc_hd__or4_1
X_4632_ _4632_/A _5027_/A VGND VGND VPWR VPWR _4987_/A sky130_fd_sc_hd__nor2_1
XFILLER_8_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4563_ _4846_/B _4563_/B VGND VGND VPWR VPWR _4718_/B sky130_fd_sc_hd__nand2_1
XFILLER_116_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold603 _6951_/Q VGND VGND VPWR VPWR hold603/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6302_ _6302_/A1 _6302_/A2 _6302_/B1 _6302_/B2 VGND VGND VPWR VPWR _6302_/X sky130_fd_sc_hd__a22o_1
XFILLER_7_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold614 _6574_/Q VGND VGND VPWR VPWR hold614/X sky130_fd_sc_hd__dlygate4sd3_1
X_3514_ _6132_/A1 _3316_/Y _3665_/A2 _6770_/Q wire809/X VGND VGND VPWR VPWR _3515_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold625 _6575_/Q VGND VGND VPWR VPWR hold625/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4494_ _4607_/B _4532_/B VGND VGND VPWR VPWR _4494_/Y sky130_fd_sc_hd__nor2_1
Xhold636 _6871_/Q VGND VGND VPWR VPWR hold636/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 _7049_/Q VGND VGND VPWR VPWR hold647/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 _7064_/Q VGND VGND VPWR VPWR hold658/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6233_ _6716_/Q _6308_/A2 _6308_/B1 _6766_/Q _6233_/C1 VGND VGND VPWR VPWR _6233_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_104_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold669 _6510_/Q VGND VGND VPWR VPWR hold669/X sky130_fd_sc_hd__dlygate4sd3_1
X_3445_ _3445_/A _3445_/B _3445_/C _3445_/D VGND VGND VPWR VPWR _3446_/D sky130_fd_sc_hd__or4_1
XFILLER_116_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6164_ _6164_/A1 _6164_/A2 _6164_/B1 _7039_/Q _6163_/X VGND VGND VPWR VPWR _6167_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ wire356/X _6790_/Q _3917_/A VGND VGND VPWR VPWR _6790_/D sky130_fd_sc_hd__mux2_1
XFILLER_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5115_ _5115_/A _5115_/B VGND VGND VPWR VPWR _5115_/X sky130_fd_sc_hd__or2_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6095_ _6844_/Q wire981/X wire587/X _6094_/X _6095_/C1 VGND VGND VPWR VPWR _6095_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5046_ _4516_/B _4514_/B _4746_/Y _4880_/X _5008_/C VGND VGND VPWR VPWR _5132_/A
+ sky130_fd_sc_hd__a2111o_1
XFILLER_38_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6997_ _7101_/CLK _6997_/D _7030_/RESET_B VGND VGND VPWR VPWR _6997_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_41_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5948_ _7173_/Q _5947_/X _5948_/S VGND VGND VPWR VPWR _7173_/D sky130_fd_sc_hd__mux2_1
XFILLER_159_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5879_ _5879_/A _5879_/B _5879_/C _5879_/D VGND VGND VPWR VPWR _5879_/X sky130_fd_sc_hd__or4_1
XFILLER_21_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length1245 _3300_/Y VGND VGND VPWR VPWR _3653_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_134_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length1278 _3782_/A2 VGND VGND VPWR VPWR _3966_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_108_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3181 _5108_/A VGND VGND VPWR VPWR _4913_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_138_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3230_ _3230_/A VGND VGND VPWR VPWR _3230_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6920_ _7109_/CLK _6920_/D wire3999/A VGND VGND VPWR VPWR _6920_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6851_ _6939_/CLK _6851_/D _6407_/A VGND VGND VPWR VPWR _6851_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_62_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5802_ _6959_/Q _5802_/A2 _5802_/B1 _6911_/Q _5801_/X VGND VGND VPWR VPWR _5802_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_90_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3994_ hold570/X _5195_/A0 _4000_/S VGND VGND VPWR VPWR _6491_/D sky130_fd_sc_hd__mux2_1
X_6782_ _7196_/CLK _6782_/D wire4264/X VGND VGND VPWR VPWR _6782_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5733_ _7068_/Q _5760_/A2 _5733_/B1 _6093_/A1 _5732_/X VGND VGND VPWR VPWR _5740_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_31_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5664_ _7152_/Q _5705_/B _5700_/C VGND VGND VPWR VPWR _5664_/X sky130_fd_sc_hd__and3_1
XFILLER_108_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_54_csclk _7117_/CLK VGND VGND VPWR VPWR _7137_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_135_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4615_ _4784_/B _4592_/A _5089_/B2 _4587_/B VGND VGND VPWR VPWR _4618_/D sky130_fd_sc_hd__o22a_1
X_5595_ _5604_/D VGND VGND VPWR VPWR _5595_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold400 _6678_/Q VGND VGND VPWR VPWR hold400/X sky130_fd_sc_hd__dlygate4sd3_1
X_4546_ _4546_/A _4546_/B VGND VGND VPWR VPWR _4573_/B sky130_fd_sc_hd__xnor2_1
Xhold411 _6524_/Q VGND VGND VPWR VPWR hold411/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 _6798_/Q VGND VGND VPWR VPWR hold422/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire4109 wire4110/X VGND VGND VPWR VPWR wire4109/X sky130_fd_sc_hd__clkbuf_1
Xhold433 _7052_/Q VGND VGND VPWR VPWR hold433/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold444 _7044_/Q VGND VGND VPWR VPWR hold444/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 _6802_/Q VGND VGND VPWR VPWR hold455/X sky130_fd_sc_hd__dlygate4sd3_1
X_4477_ _5018_/A _4664_/A VGND VGND VPWR VPWR _4477_/X sky130_fd_sc_hd__or2_2
Xwire3408 wire3409/X VGND VGND VPWR VPWR wire3408/X sky130_fd_sc_hd__clkbuf_1
Xhold466 _6659_/Q VGND VGND VPWR VPWR hold466/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 _6990_/Q VGND VGND VPWR VPWR hold477/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold488 _6896_/Q VGND VGND VPWR VPWR hold488/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold499 _6879_/Q VGND VGND VPWR VPWR hold499/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_69_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7036_/CLK sky130_fd_sc_hd__clkbuf_16
Xwire2707 _6015_/X VGND VGND VPWR VPWR _6184_/B1 sky130_fd_sc_hd__clkbuf_1
X_6216_ _6216_/A _6216_/B _6216_/C _6216_/D VGND VGND VPWR VPWR _6217_/D sky130_fd_sc_hd__or4_1
X_3428_ _6150_/B2 _5439_/A _3428_/B1 _7079_/Q _3419_/X VGND VGND VPWR VPWR _3431_/B
+ sky130_fd_sc_hd__a221o_1
X_7196_ _7196_/CLK _7196_/D VGND VGND VPWR VPWR _7196_/Q sky130_fd_sc_hd__dfxtp_1
Xwire2718 _6333_/B1 VGND VGND VPWR VPWR _6310_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2729 wire2730/X VGND VGND VPWR VPWR _6333_/A2 sky130_fd_sc_hd__clkbuf_2
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6147_ _6147_/A1 _6197_/A2 _6197_/B1 _6147_/B2 VGND VGND VPWR VPWR _6147_/X sky130_fd_sc_hd__a22o_1
X_3359_ _6202_/B2 _3533_/A2 wire885/X _3359_/B2 _3358_/X VGND VGND VPWR VPWR _3359_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6078_ hold91/A _6078_/A2 _6138_/B1 _6078_/B2 VGND VGND VPWR VPWR _6078_/X sky130_fd_sc_hd__a22o_1
X_5029_ _5109_/B _5029_/B _5029_/C _5029_/D VGND VGND VPWR VPWR _5029_/X sky130_fd_sc_hd__and4b_1
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length923 wire924/X VGND VGND VPWR VPWR wire920/A sky130_fd_sc_hd__clkbuf_1
XFILLER_127_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length945 _3308_/Y VGND VGND VPWR VPWR wire939/A sky130_fd_sc_hd__clkbuf_1
XFILLER_181_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length967 _3278_/Y VGND VGND VPWR VPWR wire966/A sky130_fd_sc_hd__clkbuf_1
XFILLER_119_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout3836 _6435_/B VGND VGND VPWR VPWR _6437_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_150_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length1097 _3417_/Y VGND VGND VPWR VPWR _5193_/A sky130_fd_sc_hd__clkbuf_2
Xwire3920 wire3921/X VGND VGND VPWR VPWR wire3920/X sky130_fd_sc_hd__clkbuf_1
Xwire3931 wire3932/X VGND VGND VPWR VPWR wire3931/X sky130_fd_sc_hd__clkbuf_1
Xwire3942 _6432_/A VGND VGND VPWR VPWR _6429_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_96_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4400_ _4450_/A _4400_/B VGND VGND VPWR VPWR _4742_/A sky130_fd_sc_hd__nor2_1
X_5380_ _5380_/A0 hold421/X _5382_/S VGND VGND VPWR VPWR _6957_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4331_ _5212_/C hold363/X _4335_/S VGND VGND VPWR VPWR _6771_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7050_ _7074_/CLK _7050_/D fanout3976/X VGND VGND VPWR VPWR _7050_/Q sky130_fd_sc_hd__dfstp_1
X_4262_ hold252/X _4274_/A1 _4263_/S VGND VGND VPWR VPWR _6714_/D sky130_fd_sc_hd__mux2_1
X_6001_ _6021_/A _6019_/B VGND VGND VPWR VPWR _6001_/Y sky130_fd_sc_hd__nor2_1
X_3213_ _7013_/Q VGND VGND VPWR VPWR _3213_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4193_ _6650_/Q wire367/X _4196_/S VGND VGND VPWR VPWR _6650_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6903_ _7116_/CLK _6903_/D wire4071/A VGND VGND VPWR VPWR _6903_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_70_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6834_ _6973_/CLK _6834_/D wire4069/X VGND VGND VPWR VPWR _6834_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6765_ _7066_/CLK _6765_/D wire3968/A VGND VGND VPWR VPWR _6765_/Q sky130_fd_sc_hd__dfrtp_1
X_3977_ hold106/X hold197/X _3979_/S VGND VGND VPWR VPWR _3977_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5716_ _6053_/A1 _5716_/A2 _5715_/X VGND VGND VPWR VPWR _5719_/C sky130_fd_sc_hd__a21o_1
XFILLER_31_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6696_ _7206_/CLK _6696_/D _6348_/B VGND VGND VPWR VPWR _6696_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_148_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5647_ _5651_/A _7160_/Q _5647_/S VGND VGND VPWR VPWR _7160_/D sky130_fd_sc_hd__mux2_1
XFILLER_40_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5578_ _5578_/A0 hold52/X _5579_/S VGND VGND VPWR VPWR hold53/A sky130_fd_sc_hd__mux2_1
XFILLER_151_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold230 _6954_/Q VGND VGND VPWR VPWR hold230/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 _6588_/Q VGND VGND VPWR VPWR hold241/X sky130_fd_sc_hd__dlygate4sd3_1
X_4529_ _4487_/B _4475_/A _5148_/A VGND VGND VPWR VPWR _4530_/D sky130_fd_sc_hd__a21oi_1
Xhold252 _6714_/Q VGND VGND VPWR VPWR hold252/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3205 _4494_/Y VGND VGND VPWR VPWR _4728_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold263 _6942_/Q VGND VGND VPWR VPWR hold263/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3216 _5001_/B VGND VGND VPWR VPWR _4514_/B sky130_fd_sc_hd__buf_2
Xhold274 _6536_/Q VGND VGND VPWR VPWR hold274/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3227 _4748_/A VGND VGND VPWR VPWR _4753_/A sky130_fd_sc_hd__clkbuf_2
Xhold285 _4093_/X VGND VGND VPWR VPWR _6568_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 _6583_/Q VGND VGND VPWR VPWR hold296/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3249 _4135_/B VGND VGND VPWR VPWR _5210_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_172_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2515 _6002_/Y VGND VGND VPWR VPWR _6278_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire2526 wire2526/A VGND VGND VPWR VPWR _6112_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_104_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2537 _6201_/B1 VGND VGND VPWR VPWR _6089_/A2 sky130_fd_sc_hd__clkbuf_1
X_7179_ _3937_/A1 _7179_/D wire4007/A VGND VGND VPWR VPWR _7179_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1803 wire1804/X VGND VGND VPWR VPWR _5759_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2548 _6104_/B1 VGND VGND VPWR VPWR _6054_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire1814 hold721/X VGND VGND VPWR VPWR _5432_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2559 _6023_/B VGND VGND VPWR VPWR _6338_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire1825 wire1826/X VGND VGND VPWR VPWR _6135_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire1836 _6995_/Q VGND VGND VPWR VPWR wire1836/X sky130_fd_sc_hd__clkbuf_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1847 _5763_/B2 VGND VGND VPWR VPWR wire1847/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1858 _6981_/Q VGND VGND VPWR VPWR _5755_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1869 _6970_/Q VGND VGND VPWR VPWR _6010_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_103 _3937_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_114 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_125 _6069_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3750 _4727_/B1 VGND VGND VPWR VPWR _4228_/B sky130_fd_sc_hd__clkbuf_4
Xwire3761 wire3762/X VGND VGND VPWR VPWR _3979_/S sky130_fd_sc_hd__clkbuf_2
Xwire3783 wire3784/X VGND VGND VPWR VPWR wire3783/X sky130_fd_sc_hd__clkbuf_1
XFILLER_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3794 _6460_/Q VGND VGND VPWR VPWR _3951_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput9 mask_rev_in[14] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3900_ _3907_/A _3908_/B VGND VGND VPWR VPWR _5596_/B sky130_fd_sc_hd__nor2_1
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4880_ _4516_/B _4521_/A _4985_/B VGND VGND VPWR VPWR _4880_/X sky130_fd_sc_hd__a21o_1
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3831_ _3831_/A _3831_/B VGND VGND VPWR VPWR _6464_/D sky130_fd_sc_hd__xnor2_1
XFILLER_177_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6550_ _7129_/CLK _6550_/D wire4055/X VGND VGND VPWR VPWR _6550_/Q sky130_fd_sc_hd__dfrtp_1
X_3762_ _6994_/Q _3762_/A2 _4330_/A _6771_/Q VGND VGND VPWR VPWR _3762_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5501_ _5501_/A0 hold538/X _5501_/S VGND VGND VPWR VPWR _7065_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6481_ _7027_/CLK _6481_/D fanout3976/X VGND VGND VPWR VPWR _6481_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_9_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3693_ _7067_/Q _3693_/A2 _3465_/Y _5899_/B2 VGND VGND VPWR VPWR _3693_/X sky130_fd_sc_hd__a22o_1
XFILLER_145_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5432_ _5432_/A0 _5432_/A1 _5434_/S VGND VGND VPWR VPWR _7003_/D sky130_fd_sc_hd__mux2_1
XFILLER_10_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput302 _6808_/Q VGND VGND VPWR VPWR pwr_ctrl_out[1] sky130_fd_sc_hd__buf_12
Xoutput313 wire3670/X VGND VGND VPWR VPWR spimemio_flash_io0_di sky130_fd_sc_hd__buf_12
X_5363_ _5585_/A0 hold263/X _5363_/S VGND VGND VPWR VPWR _6942_/D sky130_fd_sc_hd__mux2_1
Xoutput324 _6646_/Q VGND VGND VPWR VPWR wb_dat_o[15] sky130_fd_sc_hd__buf_12
Xoutput335 _7190_/Q VGND VGND VPWR VPWR wb_dat_o[25] sky130_fd_sc_hd__buf_12
Xoutput346 _6653_/Q VGND VGND VPWR VPWR wb_dat_o[6] sky130_fd_sc_hd__buf_12
X_7102_ _7102_/CLK _7102_/D wire4004/A VGND VGND VPWR VPWR _7102_/Q sky130_fd_sc_hd__dfrtp_1
X_4314_ hold618/X _4314_/A1 _4316_/S VGND VGND VPWR VPWR _6757_/D sky130_fd_sc_hd__mux2_1
X_5294_ _5579_/A0 hold211/X _5294_/S VGND VGND VPWR VPWR _6881_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7033_ _7080_/CLK _7033_/D _6562_/SET_B VGND VGND VPWR VPWR _7033_/Q sky130_fd_sc_hd__dfrtp_1
X_4245_ hold437/X _4251_/A0 _4245_/S VGND VGND VPWR VPWR _6690_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4176_ _5531_/A1 hold264/X _4179_/S VGND VGND VPWR VPWR _6635_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6817_ _7080_/CLK _6817_/D wire3991/X VGND VGND VPWR VPWR _6817_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire407 wire408/X VGND VGND VPWR VPWR wire407/X sky130_fd_sc_hd__clkbuf_1
X_6748_ _6963_/CLK hold32/X _6401_/A VGND VGND VPWR VPWR _6748_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_7_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire418 wire419/X VGND VGND VPWR VPWR _3755_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_183_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire429 wire430/X VGND VGND VPWR VPWR _3573_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6679_ _7208_/CLK _6679_/D wire4026/A VGND VGND VPWR VPWR _6679_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_3_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3002 _5789_/A2 VGND VGND VPWR VPWR _5727_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire3013 _5747_/B1 VGND VGND VPWR VPWR _5718_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3024 _5848_/B1 VGND VGND VPWR VPWR _5756_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3035 _5918_/A2 VGND VGND VPWR VPWR _5962_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_105_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2301 _6636_/Q VGND VGND VPWR VPWR _6284_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3046 _5826_/B1 VGND VGND VPWR VPWR _5840_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire3057 _5824_/B1 VGND VGND VPWR VPWR wire3057/X sky130_fd_sc_hd__clkbuf_1
Xwire2312 _5906_/B2 VGND VGND VPWR VPWR _6271_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_105_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2323 _6611_/Q VGND VGND VPWR VPWR _3765_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire3068 _5826_/A2 VGND VGND VPWR VPWR _5853_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3079 _5667_/X VGND VGND VPWR VPWR _5844_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2334 _6605_/Q VGND VGND VPWR VPWR _6328_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2345 _6596_/Q VGND VGND VPWR VPWR _6243_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1600 wire1601/X VGND VGND VPWR VPWR wire1600/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2356 _6539_/Q VGND VGND VPWR VPWR _6300_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_120_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1611 _6051_/A1 VGND VGND VPWR VPWR _5714_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2367 _6536_/Q VGND VGND VPWR VPWR _6224_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire1622 wire1623/X VGND VGND VPWR VPWR wire1622/X sky130_fd_sc_hd__clkbuf_1
XFILLER_120_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1633 _6099_/B2 VGND VGND VPWR VPWR _3206_/A sky130_fd_sc_hd__clkbuf_1
Xwire2378 _6529_/Q VGND VGND VPWR VPWR _3554_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2389 _6519_/Q VGND VGND VPWR VPWR _5934_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1644 _6101_/B2 VGND VGND VPWR VPWR _5761_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire1655 wire1656/X VGND VGND VPWR VPWR wire1655/X sky130_fd_sc_hd__clkbuf_1
Xwire1666 _7053_/Q VGND VGND VPWR VPWR _6105_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_18_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1677 _7047_/Q VGND VGND VPWR VPWR _5809_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_46_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1688 _6078_/B2 VGND VGND VPWR VPWR _5747_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire1699 _3394_/B2 VGND VGND VPWR VPWR _6181_/B2 sky130_fd_sc_hd__clkbuf_2
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire930 _3317_/Y VGND VGND VPWR VPWR wire930/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire941 wire944/X VGND VGND VPWR VPWR wire941/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire963 wire966/A VGND VGND VPWR VPWR wire963/X sky130_fd_sc_hd__dlymetal6s2s_1
Xwire974 _6291_/X VGND VGND VPWR VPWR wire974/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire985 _6292_/A VGND VGND VPWR VPWR _6341_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_115_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire996 _5728_/X VGND VGND VPWR VPWR wire996/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length583 _6396_/S VGND VGND VPWR VPWR _6395_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_127_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4270 wire4271/X VGND VGND VPWR VPWR _3475_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_69_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire4281 _4553_/A VGND VGND VPWR VPWR _4402_/A sky130_fd_sc_hd__clkbuf_2
Xwire4292 _4342_/C VGND VGND VPWR VPWR _4407_/A sky130_fd_sc_hd__buf_2
Xfanout3496 wire3511/A VGND VGND VPWR VPWR _4178_/A0 sky130_fd_sc_hd__clkbuf_1
Xwire3580 _4131_/A1 VGND VGND VPWR VPWR _4308_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
X_4030_ hold504/X _5504_/A0 _4033_/S VGND VGND VPWR VPWR _6522_/D sky130_fd_sc_hd__mux2_1
XFILLER_2_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2890 _5777_/B1 VGND VGND VPWR VPWR _5738_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5981_ _7082_/Q _6076_/A2 _6065_/A2 _5981_/B2 VGND VGND VPWR VPWR _5981_/X sky130_fd_sc_hd__a22o_1
XFILLER_52_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4932_ _4932_/A _4932_/B VGND VGND VPWR VPWR _4935_/C sky130_fd_sc_hd__or2_1
XFILLER_17_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4863_ _4863_/A _4863_/B VGND VGND VPWR VPWR _4864_/D sky130_fd_sc_hd__nand2_1
X_6602_ _6702_/CLK _6602_/D _6440_/A VGND VGND VPWR VPWR _6602_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_14 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3814_ _3252_/B _3811_/S _3813_/X _3244_/X VGND VGND VPWR VPWR _3814_/X sky130_fd_sc_hd__a31o_1
XANTENNA_25 wire813/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4794_ _4794_/A _4795_/B _4794_/C VGND VGND VPWR VPWR _5094_/B sky130_fd_sc_hd__or3_1
XFILLER_20_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_36 wire1255/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_47 _5740_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 _6134_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6533_ _6755_/CLK _6533_/D wire3954/X VGND VGND VPWR VPWR _6533_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA_69 _3560_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3745_ _6686_/Q _4240_/A _4246_/A _6701_/Q VGND VGND VPWR VPWR _3745_/X sky130_fd_sc_hd__a22o_1
XFILLER_192_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6464_ _3945_/A1 _6464_/D _6419_/X VGND VGND VPWR VPWR _6464_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_137_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3676_ _5900_/A1 _3676_/A2 hold30/A _6259_/A1 wire767/X VGND VGND VPWR VPWR _3679_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_106_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5415_ _5538_/A1 hold413/X _5415_/S VGND VGND VPWR VPWR _6988_/D sky130_fd_sc_hd__mux2_1
X_6395_ _6395_/A0 hold384/X _6395_/S VGND VGND VPWR VPWR _7209_/D sky130_fd_sc_hd__mux2_1
X_5346_ _5364_/A0 hold680/X _5348_/S VGND VGND VPWR VPWR _6927_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput176 _3224_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[10] sky130_fd_sc_hd__buf_12
Xoutput187 _3214_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[20] sky130_fd_sc_hd__buf_12
Xoutput198 _3204_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[30] sky130_fd_sc_hd__buf_12
XFILLER_153_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5277_ _5277_/A _5571_/B VGND VGND VPWR VPWR _5285_/S sky130_fd_sc_hd__nand2_1
XFILLER_141_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7016_ _7016_/CLK _7016_/D wire4001/A VGND VGND VPWR VPWR _7016_/Q sky130_fd_sc_hd__dfrtp_1
X_4228_ _4228_/A _4228_/B _4228_/C VGND VGND VPWR VPWR _4228_/Y sky130_fd_sc_hd__nor3_4
XFILLER_101_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4159_ _4159_/A _4159_/B VGND VGND VPWR VPWR _4164_/S sky130_fd_sc_hd__and2_1
XFILLER_95_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3533 hold48/X VGND VGND VPWR VPWR wire3532/A sky130_fd_sc_hd__clkbuf_1
XFILLER_109_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length4289 _4342_/B VGND VGND VPWR VPWR _4379_/C sky130_fd_sc_hd__clkbuf_2
Xmax_length3544 _4249_/A0 VGND VGND VPWR VPWR wire3543/A sky130_fd_sc_hd__clkbuf_1
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length3566 _5406_/A0 VGND VGND VPWR VPWR _5547_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_125_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length2887 _5932_/A2 VGND VGND VPWR VPWR _5954_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_127_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2120 wire2121/X VGND VGND VPWR VPWR wire2120/X sky130_fd_sc_hd__clkbuf_1
Xwire2131 wire2132/X VGND VGND VPWR VPWR wire2131/X sky130_fd_sc_hd__clkbuf_1
Xwire2142 _6796_/Q VGND VGND VPWR VPWR _3587_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_66_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2153 _6254_/A1 VGND VGND VPWR VPWR _3665_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire2164 _6752_/Q VGND VGND VPWR VPWR wire2164/X sky130_fd_sc_hd__clkbuf_1
XFILLER_93_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1430 _4919_/X VGND VGND VPWR VPWR _4920_/C1 sky130_fd_sc_hd__clkbuf_1
Xwire2175 _6748_/Q VGND VGND VPWR VPWR _3626_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1441 _4759_/B VGND VGND VPWR VPWR _4460_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_2_1_0_mgmt_gpio_in[4] clkbuf_2_1_0_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR _6545_/CLK
+ sky130_fd_sc_hd__clkbuf_8
Xwire2186 wire2187/X VGND VGND VPWR VPWR _6259_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire1452 _3938_/X VGND VGND VPWR VPWR wire1452/X sky130_fd_sc_hd__clkbuf_2
Xwire1463 wire1464/X VGND VGND VPWR VPWR wire1463/X sky130_fd_sc_hd__buf_6
XFILLER_74_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1474 wire1475/X VGND VGND VPWR VPWR wire1474/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1485 wire1486/X VGND VGND VPWR VPWR wire1485/X sky130_fd_sc_hd__clkbuf_1
XFILLER_46_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1496 wire1496/A VGND VGND VPWR VPWR _3456_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_74_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput12 mask_rev_in[17] VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__clkbuf_1
Xinput23 mask_rev_in[27] VGND VGND VPWR VPWR input23/X sky130_fd_sc_hd__clkbuf_1
XFILLER_168_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput34 mask_rev_in[8] VGND VGND VPWR VPWR input34/X sky130_fd_sc_hd__clkbuf_1
Xinput45 mgmt_gpio_in[18] VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire760 wire761/X VGND VGND VPWR VPWR wire760/X sky130_fd_sc_hd__clkbuf_1
X_3530_ _3726_/B _3538_/A VGND VGND VPWR VPWR hold64/A sky130_fd_sc_hd__nor2_1
XFILLER_128_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput56 mgmt_gpio_in[28] VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__clkbuf_1
Xwire771 _3665_/X VGND VGND VPWR VPWR wire771/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput67 mgmt_gpio_in[3] VGND VGND VPWR VPWR input67/X sky130_fd_sc_hd__buf_6
Xwire782 _3557_/X VGND VGND VPWR VPWR wire782/X sky130_fd_sc_hd__clkbuf_1
Xinput78 spi_csb VGND VGND VPWR VPWR input78/X sky130_fd_sc_hd__clkbuf_1
Xwire793 wire795/X VGND VGND VPWR VPWR wire793/X sky130_fd_sc_hd__clkbuf_1
Xinput89 spimemio_flash_io2_do VGND VGND VPWR VPWR input89/X sky130_fd_sc_hd__clkbuf_1
XFILLER_182_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3461_ _3461_/A1 _3308_/Y _4288_/A _3461_/B2 _3459_/X VGND VGND VPWR VPWR _3461_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5200_ _5200_/A _5203_/B VGND VGND VPWR VPWR _5202_/S sky130_fd_sc_hd__nand2_1
XFILLER_170_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6180_ _6180_/A _6180_/B _6180_/C _6180_/D VGND VGND VPWR VPWR _6193_/A sky130_fd_sc_hd__or4_1
X_3392_ _3392_/A _3392_/B _3392_/C _3392_/D VGND VGND VPWR VPWR _3410_/A sky130_fd_sc_hd__or4_1
XFILLER_97_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5131_ _4454_/Y _4514_/B _4815_/A _4878_/X _5008_/A VGND VGND VPWR VPWR _5132_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5062_ _5163_/B _5123_/B _5159_/A _5062_/D VGND VGND VPWR VPWR _5066_/A sky130_fd_sc_hd__nand4_1
XFILLER_97_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4013_ hold545/X _5532_/A1 _4014_/S VGND VGND VPWR VPWR _6508_/D sky130_fd_sc_hd__mux2_1
XFILLER_111_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5964_ _6329_/A1 _5964_/A2 _5964_/B1 _6324_/A1 _5963_/X VGND VGND VPWR VPWR _5967_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_52_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4915_ _4915_/A _4915_/B _4915_/C _4914_/X VGND VGND VPWR VPWR _4924_/A sky130_fd_sc_hd__or4b_1
XFILLER_178_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5895_ _6252_/B2 _5956_/A2 _5895_/B1 _5894_/X VGND VGND VPWR VPWR _5895_/X sky130_fd_sc_hd__a22o_1
X_4846_ _4846_/A _4846_/B _4846_/C _4846_/D VGND VGND VPWR VPWR _4868_/C sky130_fd_sc_hd__and4_1
X_4777_ _5094_/A _4976_/A1 _4745_/A VGND VGND VPWR VPWR _5158_/B sky130_fd_sc_hd__a21oi_2
XFILLER_21_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6516_ _7090_/CLK _6516_/D wire3945/A VGND VGND VPWR VPWR _6516_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_107_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3728_ _6010_/A1 wire915/X wire808/X _6606_/Q VGND VGND VPWR VPWR _3728_/X sky130_fd_sc_hd__a22o_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6447_ _3927_/A1 _6447_/D _6402_/X VGND VGND VPWR VPWR _6447_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3659_ _3659_/A _3659_/B _3659_/C _3659_/D VGND VGND VPWR VPWR _3660_/C sky130_fd_sc_hd__or4_1
X_6378_ _4228_/B _6378_/A2 _6378_/B1 _4228_/Y VGND VGND VPWR VPWR _6378_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5329_ hold610/X _5464_/A0 _5330_/S VGND VGND VPWR VPWR _6912_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length4020 wire4018/A VGND VGND VPWR VPWR wire4019/A sky130_fd_sc_hd__clkbuf_1
XFILLER_157_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length4053 wire4052/A VGND VGND VPWR VPWR _6499_/SET_B sky130_fd_sc_hd__clkbuf_2
Xmax_length4075 _7134_/RESET_B VGND VGND VPWR VPWR _6833_/RESET_B sky130_fd_sc_hd__buf_2
XFILLER_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length3352 _4387_/B VGND VGND VPWR VPWR _5133_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length3396 _5509_/A0 VGND VGND VPWR VPWR _5356_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_98_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length2695 _6210_/B1 VGND VGND VPWR VPWR wire2694/A sky130_fd_sc_hd__clkbuf_1
XFILLER_113_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1260 _3599_/A2 VGND VGND VPWR VPWR _3654_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_94_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1271 wire1271/A VGND VGND VPWR VPWR _3605_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1293 _3451_/A VGND VGND VPWR VPWR _3528_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4700_ _4707_/B _4704_/B _4920_/B1 _4683_/A VGND VGND VPWR VPWR _4700_/X sky130_fd_sc_hd__a31o_1
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5680_ _6962_/Q _5680_/A2 _5722_/A2 _5680_/B2 _5679_/X VGND VGND VPWR VPWR _5681_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_175_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4631_ _5083_/A _4631_/B VGND VGND VPWR VPWR _4915_/A sky130_fd_sc_hd__nand2b_1
XFILLER_175_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4562_ _4562_/A _4596_/B VGND VGND VPWR VPWR _4562_/X sky130_fd_sc_hd__or2_1
X_6301_ _6524_/Q _6301_/A2 _6301_/B1 _6764_/Q _6299_/X VGND VGND VPWR VPWR _6301_/X
+ sky130_fd_sc_hd__a221o_1
Xhold604 _7126_/Q VGND VGND VPWR VPWR hold604/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold615 _7038_/Q VGND VGND VPWR VPWR hold615/X sky130_fd_sc_hd__dlygate4sd3_1
X_3513_ _6327_/B2 _3513_/A2 _3677_/B1 _6328_/A1 VGND VGND VPWR VPWR _3513_/X sky130_fd_sc_hd__a22o_1
Xwire590 _5729_/X VGND VGND VPWR VPWR wire590/X sky130_fd_sc_hd__clkbuf_1
Xhold626 _6479_/Q VGND VGND VPWR VPWR hold626/X sky130_fd_sc_hd__dlygate4sd3_1
X_4493_ _4745_/A _4493_/B VGND VGND VPWR VPWR _4493_/X sky130_fd_sc_hd__or2_1
XFILLER_143_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold637 _6716_/Q VGND VGND VPWR VPWR hold637/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold648 _7021_/Q VGND VGND VPWR VPWR hold648/X sky130_fd_sc_hd__dlygate4sd3_1
X_6232_ _6232_/A _6232_/B _6232_/C _6232_/D VGND VGND VPWR VPWR _6232_/X sky130_fd_sc_hd__or4_1
Xhold659 _7006_/Q VGND VGND VPWR VPWR hold659/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3444_ _3444_/A1 wire943/X _5562_/A _7124_/Q _3443_/X VGND VGND VPWR VPWR _3444_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3375_ wire379/X _6789_/Q _3791_/A VGND VGND VPWR VPWR _3375_/X sky130_fd_sc_hd__mux2_1
X_6163_ _6163_/A1 _6163_/A2 _6163_/B1 _6163_/B2 VGND VGND VPWR VPWR _6163_/X sky130_fd_sc_hd__a22o_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5114_ _5114_/A _5114_/B _5114_/C _5114_/D VGND VGND VPWR VPWR _5171_/A sky130_fd_sc_hd__or4_1
XFILLER_57_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ _6119_/A _6094_/B _6094_/C _6094_/D VGND VGND VPWR VPWR _6094_/X sky130_fd_sc_hd__or4_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _5045_/A _5045_/B VGND VGND VPWR VPWR _5134_/C sky130_fd_sc_hd__or2_1
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6996_ _7076_/CLK _6996_/D fanout3976/X VGND VGND VPWR VPWR _6996_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5947_ _5969_/A1 _7172_/Q _5946_/X VGND VGND VPWR VPWR _5947_/X sky130_fd_sc_hd__a21o_1
X_5878_ _5878_/A1 _5878_/A2 _5940_/A2 _6521_/Q _5877_/X VGND VGND VPWR VPWR _5878_/X
+ sky130_fd_sc_hd__a221o_1
X_4829_ _4596_/B _4483_/A _4847_/A VGND VGND VPWR VPWR _4829_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_138_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length1202 _3320_/Y VGND VGND VPWR VPWR wire1201/A sky130_fd_sc_hd__clkbuf_1
XFILLER_119_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length1257 _5520_/A VGND VGND VPWR VPWR _3363_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_162_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length1268 _3294_/Y VGND VGND VPWR VPWR _3671_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_134_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1 hold1/A VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_94_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1090 _3450_/Y VGND VGND VPWR VPWR _5529_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6850_ _6939_/CLK _6850_/D _6407_/A VGND VGND VPWR VPWR _6850_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_35_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5801_ _5801_/A1 _5801_/A2 _5832_/B1 _5801_/B2 VGND VGND VPWR VPWR _5801_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6781_ _7196_/CLK _6781_/D wire4264/X VGND VGND VPWR VPWR _6781_/Q sky130_fd_sc_hd__dfrtp_1
X_3993_ hold577/X _4295_/A0 _4000_/S VGND VGND VPWR VPWR _6490_/D sky130_fd_sc_hd__mux2_1
XFILLER_22_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5732_ _5732_/A1 _5759_/A2 _5782_/B1 _5732_/B2 VGND VGND VPWR VPWR _5732_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5663_ _7152_/Q _5700_/C _5699_/B VGND VGND VPWR VPWR _5663_/X sky130_fd_sc_hd__and3_1
XFILLER_136_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4614_ _4614_/A _4646_/B VGND VGND VPWR VPWR _4916_/A sky130_fd_sc_hd__or2_1
XFILLER_191_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5594_ _6565_/Q _5593_/B _6564_/Q _5592_/Y VGND VGND VPWR VPWR _5604_/D sky130_fd_sc_hd__o31a_1
XFILLER_129_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold401 _6987_/Q VGND VGND VPWR VPWR hold401/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4545_ _4621_/A _4575_/B _4621_/C VGND VGND VPWR VPWR _4545_/X sky130_fd_sc_hd__or3_1
Xhold412 _7010_/Q VGND VGND VPWR VPWR hold412/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 _6603_/Q VGND VGND VPWR VPWR hold423/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold434 _6876_/Q VGND VGND VPWR VPWR hold434/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold445 _6900_/Q VGND VGND VPWR VPWR hold445/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4476_ _4476_/A _4564_/B _4588_/B _4565_/A VGND VGND VPWR VPWR _4664_/A sky130_fd_sc_hd__or4b_1
Xwire3409 _5410_/A0 VGND VGND VPWR VPWR wire3409/X sky130_fd_sc_hd__clkbuf_1
Xhold456 _6902_/Q VGND VGND VPWR VPWR hold456/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 _7136_/Q VGND VGND VPWR VPWR hold467/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 _6602_/Q VGND VGND VPWR VPWR hold478/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold489 _6661_/Q VGND VGND VPWR VPWR hold489/X sky130_fd_sc_hd__dlygate4sd3_1
X_6215_ _6215_/A1 _6215_/A2 _6215_/B1 _6215_/B2 _6214_/X VGND VGND VPWR VPWR _6216_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3427_ _6164_/A1 _5259_/A _4104_/A _3427_/B2 wire841/X VGND VGND VPWR VPWR _3431_/A
+ sky130_fd_sc_hd__a221o_1
Xwire2708 _6022_/C VGND VGND VPWR VPWR _6336_/A2 sky130_fd_sc_hd__clkbuf_2
X_7195_ _7196_/CLK _7195_/D VGND VGND VPWR VPWR _7195_/Q sky130_fd_sc_hd__dfxtp_1
Xwire2719 wire2720/X VGND VGND VPWR VPWR _6333_/B1 sky130_fd_sc_hd__clkbuf_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6146_ _7179_/Q _6145_/X _6146_/S VGND VGND VPWR VPWR _7179_/D sky130_fd_sc_hd__mux2_1
XFILLER_58_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3358_ _3358_/A1 wire941/X _3358_/B1 _6985_/Q VGND VGND VPWR VPWR _3358_/X sky130_fd_sc_hd__a22o_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6077_ _6077_/A1 _6139_/A2 _6137_/B1 _6077_/B2 _6076_/X VGND VGND VPWR VPWR _6084_/A
+ sky130_fd_sc_hd__a221o_1
X_3289_ _3313_/B _3378_/B VGND VGND VPWR VPWR _3536_/B sky130_fd_sc_hd__nand2_2
XFILLER_73_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5028_ _5074_/A2 _4781_/Y _4477_/X VGND VGND VPWR VPWR _5028_/X sky130_fd_sc_hd__a21o_1
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6979_ _6979_/CLK _6979_/D fanout4027/X VGND VGND VPWR VPWR _6979_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_80_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length979 wire981/X VGND VGND VPWR VPWR _6268_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_181_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length1043 _4252_/A VGND VGND VPWR VPWR _3513_/A2 sky130_fd_sc_hd__clkbuf_1
Xfanout3815 wire3822/X VGND VGND VPWR VPWR _4638_/A sky130_fd_sc_hd__buf_6
Xmax_length1054 _3495_/Y VGND VGND VPWR VPWR _4028_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_107_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length1076 _4318_/A VGND VGND VPWR VPWR _3652_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire3910 wire3911/X VGND VGND VPWR VPWR wire3910/X sky130_fd_sc_hd__clkbuf_1
XFILLER_150_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3921 wire3922/X VGND VGND VPWR VPWR wire3921/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3932 wire3933/X VGND VGND VPWR VPWR wire3932/X sky130_fd_sc_hd__clkbuf_1
Xwire3943 wire3943/A VGND VGND VPWR VPWR _6432_/A sky130_fd_sc_hd__clkbuf_2
Xwire3954 wire3956/X VGND VGND VPWR VPWR wire3954/X sky130_fd_sc_hd__buf_2
Xwire3965 wire3965/A VGND VGND VPWR VPWR _6440_/A sky130_fd_sc_hd__buf_2
XFILLER_103_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_588 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4330_ _4330_/A _5203_/B VGND VGND VPWR VPWR _4335_/S sky130_fd_sc_hd__nand2_2
XFILLER_126_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4261_ _6713_/Q _4273_/A1 _4263_/S VGND VGND VPWR VPWR hold71/A sky130_fd_sc_hd__mux2_1
XFILLER_5_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6000_ _6000_/A _6033_/A _6040_/B VGND VGND VPWR VPWR _6000_/X sky130_fd_sc_hd__and3_1
XFILLER_140_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3212_ _3212_/A VGND VGND VPWR VPWR _3212_/Y sky130_fd_sc_hd__inv_2
X_4192_ _6649_/Q wire364/X _4196_/S VGND VGND VPWR VPWR _6649_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6902_ _7139_/CLK _6902_/D wire4066/X VGND VGND VPWR VPWR _6902_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6833_ _7132_/CLK hold41/X _6833_/RESET_B VGND VGND VPWR VPWR hold40/A sky130_fd_sc_hd__dfrtp_1
XFILLER_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6764_ _7066_/CLK _6764_/D wire3970/X VGND VGND VPWR VPWR _6764_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3976_ hold711/X _4311_/A0 _3976_/S VGND VGND VPWR VPWR _6478_/D sky130_fd_sc_hd__mux2_1
XFILLER_10_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5715_ _7059_/Q _5715_/A2 _5715_/B1 _7075_/Q VGND VGND VPWR VPWR _5715_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6695_ _7196_/CLK _6695_/D _6780_/RESET_B VGND VGND VPWR VPWR _6695_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_148_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5646_ _5593_/Y _5609_/Y _5645_/X _6565_/Q VGND VGND VPWR VPWR _5647_/S sky130_fd_sc_hd__a22o_1
XFILLER_163_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5577_ _5577_/A0 hold393/X _5579_/S VGND VGND VPWR VPWR _7132_/D sky130_fd_sc_hd__mux2_1
Xhold220 _6899_/Q VGND VGND VPWR VPWR hold220/X sky130_fd_sc_hd__dlygate4sd3_1
X_4528_ _5126_/A _4847_/A _4882_/A _4528_/D VGND VGND VPWR VPWR _4530_/C sky130_fd_sc_hd__and4b_1
XFILLER_117_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold231 _6570_/Q VGND VGND VPWR VPWR hold231/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 _4121_/X VGND VGND VPWR VPWR _6588_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 _6724_/Q VGND VGND VPWR VPWR hold253/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 _6635_/Q VGND VGND VPWR VPWR hold264/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3206 _5105_/B2 VGND VGND VPWR VPWR _5013_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3217 _4450_/Y VGND VGND VPWR VPWR _4657_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xhold275 _6567_/Q VGND VGND VPWR VPWR hold275/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3228 _4760_/A1 VGND VGND VPWR VPWR _4748_/A sky130_fd_sc_hd__clkbuf_2
Xwire3239 _5033_/A VGND VGND VPWR VPWR _6362_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold286 _6743_/Q VGND VGND VPWR VPWR hold286/X sky130_fd_sc_hd__dlygate4sd3_1
X_4459_ _4495_/A _4459_/B VGND VGND VPWR VPWR _5035_/B sky130_fd_sc_hd__nand2_1
Xhold297 _6613_/Q VGND VGND VPWR VPWR hold297/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire2505 _6302_/B1 VGND VGND VPWR VPWR _6322_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2516 _6152_/A2 VGND VGND VPWR VPWR _6074_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7178_ _3937_/A1 _7178_/D wire4007/A VGND VGND VPWR VPWR _7178_/Q sky130_fd_sc_hd__dfrtp_1
Xwire2538 _6150_/B1 VGND VGND VPWR VPWR _6052_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire1804 wire1804/A VGND VGND VPWR VPWR wire1804/X sky130_fd_sc_hd__clkbuf_1
Xwire2549 _6175_/A2 VGND VGND VPWR VPWR _6104_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_131_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1815 wire1816/X VGND VGND VPWR VPWR _6011_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_105_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6129_ _6129_/A1 _6129_/A2 _6129_/B1 _6129_/B2 VGND VGND VPWR VPWR _6129_/X sky130_fd_sc_hd__a22o_1
Xwire1826 wire1827/X VGND VGND VPWR VPWR wire1826/X sky130_fd_sc_hd__clkbuf_1
XFILLER_85_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1837 wire1838/X VGND VGND VPWR VPWR _6031_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_86_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1848 _6104_/B2 VGND VGND VPWR VPWR _5763_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1859 wire1860/X VGND VGND VPWR VPWR _6088_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_104 _3487_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_115 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_126 _3508_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout3634 wire3662/X VGND VGND VPWR VPWR wire3642/A sky130_fd_sc_hd__buf_6
XFILLER_107_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout3678 _3235_/Y VGND VGND VPWR VPWR _5688_/A sky130_fd_sc_hd__buf_6
XFILLER_123_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3740 wire3741/X VGND VGND VPWR VPWR wire3740/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3751 wire3752/X VGND VGND VPWR VPWR _4727_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_122_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3762 wire3763/X VGND VGND VPWR VPWR wire3762/X sky130_fd_sc_hd__clkbuf_1
Xwire3773 _5593_/B VGND VGND VPWR VPWR _5859_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire3784 wire3785/X VGND VGND VPWR VPWR wire3784/X sky130_fd_sc_hd__clkbuf_1
Xwire3795 wire3796/X VGND VGND VPWR VPWR _3877_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_103_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_53_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _6956_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_45_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3830_ _3830_/A _3833_/S VGND VGND VPWR VPWR _3831_/B sky130_fd_sc_hd__nor2_1
XFILLER_177_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_68_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7074_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_60_675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3761_ _6751_/Q _4306_/A _5229_/A _6824_/Q VGND VGND VPWR VPWR _3761_/X sky130_fd_sc_hd__a22o_1
X_5500_ _5569_/A0 hold658/X _5501_/S VGND VGND VPWR VPWR _7064_/D sky130_fd_sc_hd__mux2_1
X_6480_ _7027_/CLK _6480_/D fanout3976/X VGND VGND VPWR VPWR _6480_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3692_ _6607_/Q _3692_/A2 _3691_/X _3692_/C1 VGND VGND VPWR VPWR _3722_/A sky130_fd_sc_hd__a211o_1
XFILLER_185_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5431_ _5467_/A1 hold716/X _5434_/S VGND VGND VPWR VPWR _7002_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput303 _6809_/Q VGND VGND VPWR VPWR pwr_ctrl_out[2] sky130_fd_sc_hd__buf_12
Xoutput314 wire3665/X VGND VGND VPWR VPWR spimemio_flash_io1_di sky130_fd_sc_hd__buf_12
X_5362_ _5362_/A0 hold97/X _5366_/S VGND VGND VPWR VPWR _6941_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput325 _6626_/Q VGND VGND VPWR VPWR wb_dat_o[16] sky130_fd_sc_hd__buf_12
Xoutput336 wire3718/X VGND VGND VPWR VPWR wb_dat_o[26] sky130_fd_sc_hd__buf_12
X_7101_ _7101_/CLK _7101_/D _7141_/RESET_B VGND VGND VPWR VPWR _7101_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput347 _6654_/Q VGND VGND VPWR VPWR wb_dat_o[7] sky130_fd_sc_hd__buf_12
XFILLER_113_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4313_ hold613/X _4325_/A1 _4316_/S VGND VGND VPWR VPWR _6756_/D sky130_fd_sc_hd__mux2_1
X_5293_ _5482_/A0 hold214/X _5294_/S VGND VGND VPWR VPWR _6880_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7032_ _7064_/CLK _7032_/D wire4045/X VGND VGND VPWR VPWR _7032_/Q sky130_fd_sc_hd__dfrtp_1
X_4244_ hold436/X _5533_/A1 _4245_/S VGND VGND VPWR VPWR _6689_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4175_ _4223_/A0 hold258/X _4179_/S VGND VGND VPWR VPWR _6634_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6816_ _7080_/CLK _6816_/D wire3992/X VGND VGND VPWR VPWR _6816_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6747_ _7111_/CLK _6747_/D fanout4027/X VGND VGND VPWR VPWR _6747_/Q sky130_fd_sc_hd__dfrtp_1
X_3959_ _3959_/A input1/X VGND VGND VPWR VPWR _3959_/X sky130_fd_sc_hd__and2_1
Xwire408 _4070_/X VGND VGND VPWR VPWR wire408/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire419 wire420/X VGND VGND VPWR VPWR wire419/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6678_ _7091_/CLK _6678_/D wire4029/A VGND VGND VPWR VPWR _6678_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3759 _3941_/A VGND VGND VPWR VPWR _3265_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_164_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5629_ _7154_/Q _7153_/Q VGND VGND VPWR VPWR _6040_/A sky130_fd_sc_hd__and2b_1
XFILLER_136_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3003 _5760_/A2 VGND VGND VPWR VPWR _5789_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3014 _5757_/A2 VGND VGND VPWR VPWR _5747_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3025 _5831_/B1 VGND VGND VPWR VPWR _5722_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire3036 wire3037/X VGND VGND VPWR VPWR _5918_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire2302 wire2303/X VGND VGND VPWR VPWR _3683_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire3047 _5672_/X VGND VGND VPWR VPWR _5826_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2313 _6618_/Q VGND VGND VPWR VPWR _5906_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2324 _6611_/Q VGND VGND VPWR VPWR _6225_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3069 _5670_/X VGND VGND VPWR VPWR _5826_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2335 _6604_/Q VGND VGND VPWR VPWR _3556_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2346 _6571_/Q VGND VGND VPWR VPWR _3938_/A0 sky130_fd_sc_hd__clkbuf_1
Xwire1601 _7088_/Q VGND VGND VPWR VPWR wire1601/X sky130_fd_sc_hd__clkbuf_1
Xwire2357 wire2357/A VGND VGND VPWR VPWR _3645_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire1612 _7083_/Q VGND VGND VPWR VPWR _6051_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2368 _6535_/Q VGND VGND VPWR VPWR _6336_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire1623 _5757_/B2 VGND VGND VPWR VPWR wire1623/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1634 _7069_/Q VGND VGND VPWR VPWR _6099_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire2379 _6528_/Q VGND VGND VPWR VPWR _6285_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1645 _7061_/Q VGND VGND VPWR VPWR _6101_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1656 _7056_/Q VGND VGND VPWR VPWR wire1656/X sky130_fd_sc_hd__clkbuf_1
Xwire1667 _5744_/A1 VGND VGND VPWR VPWR _3654_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire1678 wire1679/X VGND VGND VPWR VPWR _3498_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire1689 _7044_/Q VGND VGND VPWR VPWR _6078_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire920 wire920/A VGND VGND VPWR VPWR wire920/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_127_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire942 wire943/X VGND VGND VPWR VPWR wire942/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire953 _3306_/Y VGND VGND VPWR VPWR wire953/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire964 wire965/X VGND VGND VPWR VPWR _5553_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_182_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire975 _6068_/X VGND VGND VPWR VPWR _6069_/D sky130_fd_sc_hd__clkbuf_1
Xwire986 wire992/X VGND VGND VPWR VPWR _6292_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_182_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire997 wire998/X VGND VGND VPWR VPWR wire997/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4260 wire4261/X VGND VGND VPWR VPWR wire4260/X sky130_fd_sc_hd__clkbuf_4
Xwire4271 wire4272/X VGND VGND VPWR VPWR wire4271/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3570 hold22/X VGND VGND VPWR VPWR _4273_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_173_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3592 _6394_/A0 VGND VGND VPWR VPWR _5531_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2880 _5701_/A2 VGND VGND VPWR VPWR _5877_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire2891 _5698_/B1 VGND VGND VPWR VPWR _5777_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5980_ _6021_/A _6038_/B VGND VGND VPWR VPWR _5980_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4931_ _4931_/A _4931_/B VGND VGND VPWR VPWR _4932_/B sky130_fd_sc_hd__nor2_1
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4862_ _4862_/A _4862_/B _4862_/C _4862_/D VGND VGND VPWR VPWR _4864_/C sky130_fd_sc_hd__or4_1
XFILLER_177_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6601_ _7090_/CLK _6601_/D wire3945/X VGND VGND VPWR VPWR _6601_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_60_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3813_ _6468_/Q _6467_/Q _3821_/S hold60/A VGND VGND VPWR VPWR _3813_/X sky130_fd_sc_hd__a31o_1
XFILLER_177_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_15 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4793_ _4793_/A _4793_/B VGND VGND VPWR VPWR _4794_/C sky130_fd_sc_hd__or2_1
XANTENNA_26 wire813/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_37 wire1286/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 wire1353/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6532_ _7210_/CLK _6532_/D wire3950/X VGND VGND VPWR VPWR _6532_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_59 wire1586/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3744_ _5377_/A1 _3744_/A2 _4258_/A _6711_/Q wire747/X VGND VGND VPWR VPWR _3749_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6463_ _3945_/A1 _6463_/D _6418_/X VGND VGND VPWR VPWR hold81/A sky130_fd_sc_hd__dfrtp_2
X_3675_ _6799_/Q _5193_/A _5184_/A _6792_/Q VGND VGND VPWR VPWR _3675_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5414_ _5450_/A0 hold401/X _5414_/S VGND VGND VPWR VPWR _6987_/D sky130_fd_sc_hd__mux2_1
XFILLER_134_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6394_ _6394_/A0 hold540/X _6397_/S VGND VGND VPWR VPWR _7208_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5345_ _5576_/A0 hold130/X _5345_/S VGND VGND VPWR VPWR _6926_/D sky130_fd_sc_hd__mux2_1
Xoutput177 _3223_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[11] sky130_fd_sc_hd__buf_12
Xoutput188 _3213_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[21] sky130_fd_sc_hd__buf_12
XFILLER_102_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput199 _3203_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[31] sky130_fd_sc_hd__buf_12
X_5276_ _5339_/A0 hold653/X _5276_/S VGND VGND VPWR VPWR _6865_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7015_ _7017_/CLK _7015_/D fanout4077/X VGND VGND VPWR VPWR _7015_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_101_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4227_ _4263_/A1 hold355/X _4227_/S VGND VGND VPWR VPWR _6679_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4158_ _4263_/A1 hold354/X hold58/X VGND VGND VPWR VPWR _6620_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4089_ hold408/X _4088_/X _4097_/S VGND VGND VPWR VPWR _6566_/D sky130_fd_sc_hd__mux2_1
XFILLER_43_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4257 _6348_/B VGND VGND VPWR VPWR _6780_/RESET_B sky130_fd_sc_hd__buf_2
Xmax_length2800 _6022_/B VGND VGND VPWR VPWR wire2799/A sky130_fd_sc_hd__clkbuf_1
XFILLER_149_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length2822 _6125_/A2 VGND VGND VPWR VPWR _6149_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_164_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3589 _5504_/A0 VGND VGND VPWR VPWR wire3587/A sky130_fd_sc_hd__clkbuf_1
XFILLER_164_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length2866 _5702_/X VGND VGND VPWR VPWR wire2861/A sky130_fd_sc_hd__clkbuf_1
XFILLER_117_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2110 _3380_/S VGND VGND VPWR VPWR _3706_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_105_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2121 wire2122/X VGND VGND VPWR VPWR wire2121/X sky130_fd_sc_hd__clkbuf_1
Xwire2132 wire2133/X VGND VGND VPWR VPWR wire2132/X sky130_fd_sc_hd__clkbuf_1
Xwire2143 _6793_/Q VGND VGND VPWR VPWR _3772_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2165 _6751_/Q VGND VGND VPWR VPWR _6227_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1420 _5817_/X VGND VGND VPWR VPWR wire1420/X sky130_fd_sc_hd__clkbuf_1
Xwire2176 _6747_/Q VGND VGND VPWR VPWR _6259_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire1431 _4901_/X VGND VGND VPWR VPWR _4905_/A sky130_fd_sc_hd__clkbuf_1
Xwire2187 wire2188/X VGND VGND VPWR VPWR wire2187/X sky130_fd_sc_hd__clkbuf_1
Xwire1442 _4433_/X VGND VGND VPWR VPWR _4759_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1453 wire1454/X VGND VGND VPWR VPWR wire1453/X sky130_fd_sc_hd__clkbuf_2
Xwire2198 _6737_/Q VGND VGND VPWR VPWR _6250_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1464 wire1465/X VGND VGND VPWR VPWR wire1464/X sky130_fd_sc_hd__clkbuf_1
Xwire1475 wire1476/X VGND VGND VPWR VPWR wire1475/X sky130_fd_sc_hd__clkbuf_1
Xwire1486 wire1487/X VGND VGND VPWR VPWR wire1486/X sky130_fd_sc_hd__clkbuf_1
XFILLER_46_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput13 mask_rev_in[18] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput24 mask_rev_in[28] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__clkbuf_1
Xinput35 mask_rev_in[9] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__clkbuf_1
Xwire750 wire751/X VGND VGND VPWR VPWR wire750/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire761 _3702_/X VGND VGND VPWR VPWR wire761/X sky130_fd_sc_hd__clkbuf_1
Xinput46 mgmt_gpio_in[19] VGND VGND VPWR VPWR input46/X sky130_fd_sc_hd__clkbuf_1
Xinput57 mgmt_gpio_in[29] VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__clkbuf_1
Xwire772 _3657_/X VGND VGND VPWR VPWR _3658_/D sky130_fd_sc_hd__clkbuf_1
Xinput68 mgmt_gpio_in[5] VGND VGND VPWR VPWR input68/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire783 _3556_/X VGND VGND VPWR VPWR wire783/X sky130_fd_sc_hd__clkbuf_1
XFILLER_115_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput79 spi_enabled VGND VGND VPWR VPWR _3958_/B sky130_fd_sc_hd__clkbuf_2
X_3460_ _3490_/A _3460_/B VGND VGND VPWR VPWR _3460_/Y sky130_fd_sc_hd__nor2_1
XFILLER_143_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3391_ input9/X _3439_/A2 _5448_/A _7024_/Q _3385_/X VGND VGND VPWR VPWR _3391_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_184_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5130_ _5130_/A _5130_/B _5130_/C wire400/X VGND VGND VPWR VPWR _5148_/C sky130_fd_sc_hd__or4b_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire4090 wire4091/X VGND VGND VPWR VPWR wire4090/X sky130_fd_sc_hd__buf_2
XFILLER_69_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5061_ _5158_/C _5127_/C VGND VGND VPWR VPWR _5062_/D sky130_fd_sc_hd__nor2_1
XFILLER_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4012_ hold479/X _4248_/A0 _4015_/S VGND VGND VPWR VPWR _6507_/D sky130_fd_sc_hd__mux2_1
XFILLER_111_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5963_ _6321_/B2 _5963_/A2 _5963_/B1 _6334_/A1 VGND VGND VPWR VPWR _5963_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4914_ _4589_/B _4680_/B _4912_/X _4913_/X _4713_/A VGND VGND VPWR VPWR _4914_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_21_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5894_ _6712_/Q _5894_/B VGND VGND VPWR VPWR _5894_/X sky130_fd_sc_hd__or2_1
XFILLER_178_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4845_ _4745_/B _4493_/B _4745_/A VGND VGND VPWR VPWR _4930_/C sky130_fd_sc_hd__a21oi_1
XFILLER_32_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4776_ _4536_/Y _4723_/X _4775_/X _5034_/B1 _4776_/B2 VGND VGND VPWR VPWR _6776_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_165_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6515_ _7210_/CLK _6515_/D fanout3944/X VGND VGND VPWR VPWR _6515_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3727_ _5212_/A _5212_/B VGND VGND VPWR VPWR _3727_/Y sky130_fd_sc_hd__nor2_1
XFILLER_173_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6446_ _3927_/A1 _6446_/D _6401_/X VGND VGND VPWR VPWR hold35/A sky130_fd_sc_hd__dfrtp_1
X_3658_ _3658_/A _3658_/B _3658_/C _3658_/D VGND VGND VPWR VPWR _3659_/D sky130_fd_sc_hd__or4_1
XFILLER_161_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_558 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6377_ _6376_/X _7201_/Q _6386_/S VGND VGND VPWR VPWR _7201_/D sky130_fd_sc_hd__mux2_1
X_3589_ _6485_/Q _3735_/A2 _4306_/A _6754_/Q _3551_/X VGND VGND VPWR VPWR _3593_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5328_ hold528/X _5517_/A0 _5330_/S VGND VGND VPWR VPWR _6911_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5259_ _5259_/A _5571_/B VGND VGND VPWR VPWR _5267_/S sky130_fd_sc_hd__nand2_1
XFILLER_87_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length4010 fanout4005/X VGND VGND VPWR VPWR _6767_/RESET_B sky130_fd_sc_hd__clkbuf_2
XFILLER_12_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length4032 _6407_/A VGND VGND VPWR VPWR _6923_/SET_B sky130_fd_sc_hd__clkbuf_2
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length4076 fanout4073/X VGND VGND VPWR VPWR _7134_/RESET_B sky130_fd_sc_hd__buf_4
XFILLER_8_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3342 _4493_/B VGND VGND VPWR VPWR _4832_/B sky130_fd_sc_hd__clkbuf_2
Xmax_length3353 _4999_/B VGND VGND VPWR VPWR _4387_/B sky130_fd_sc_hd__clkbuf_2
Xmax_length2641 _6141_/B1 VGND VGND VPWR VPWR _6164_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_164_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length1962 _6916_/Q VGND VGND VPWR VPWR _6091_/B2 sky130_fd_sc_hd__clkbuf_1
Xmax_length1984 _6903_/Q VGND VGND VPWR VPWR wire1983/A sky130_fd_sc_hd__clkbuf_1
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1250 _3480_/A2 VGND VGND VPWR VPWR _3423_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire1261 _3296_/Y VGND VGND VPWR VPWR _3599_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1283 _3698_/A2 VGND VGND VPWR VPWR _3433_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_74_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1294 _3726_/A VGND VGND VPWR VPWR _5241_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_170_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4630_ _4630_/A _5017_/A VGND VGND VPWR VPWR _4631_/B sky130_fd_sc_hd__or2_1
XFILLER_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4561_ _4562_/A _4596_/B VGND VGND VPWR VPWR _4561_/Y sky130_fd_sc_hd__nor2_1
XFILLER_128_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6300_ _6300_/A1 _6335_/A2 _6300_/B1 _6300_/B2 _6297_/X VGND VGND VPWR VPWR _6315_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3512_ _3536_/B _3512_/B VGND VGND VPWR VPWR _3512_/Y sky130_fd_sc_hd__nor2_1
Xwire580 wire581/X VGND VGND VPWR VPWR _3355_/B sky130_fd_sc_hd__clkbuf_1
Xwire591 _5542_/S VGND VGND VPWR VPWR _5538_/S sky130_fd_sc_hd__dlymetal6s2s_1
Xhold605 _7122_/Q VGND VGND VPWR VPWR hold605/X sky130_fd_sc_hd__dlygate4sd3_1
X_4492_ _4492_/A _4721_/A _4668_/A VGND VGND VPWR VPWR _4926_/A sky130_fd_sc_hd__or3_1
Xhold616 _7032_/Q VGND VGND VPWR VPWR hold616/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold627 _7020_/Q VGND VGND VPWR VPWR hold627/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 _6718_/Q VGND VGND VPWR VPWR hold638/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6231_ _5872_/A _6333_/A2 _6306_/B1 _6231_/B2 _6230_/X VGND VGND VPWR VPWR _6232_/D
+ sky130_fd_sc_hd__a221o_1
Xhold649 _7141_/Q VGND VGND VPWR VPWR hold649/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3443_ _5800_/A1 _3443_/A2 wire870/X _6147_/B2 VGND VGND VPWR VPWR _3443_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _6162_/A1 _6162_/A2 _6162_/B1 _6887_/Q _6161_/X VGND VGND VPWR VPWR _6167_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _6456_/Q _6543_/Q VGND VGND VPWR VPWR _3917_/A sky130_fd_sc_hd__nand2_2
XFILLER_97_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _5113_/A1 _5113_/A2 _4646_/X VGND VGND VPWR VPWR _5114_/D sky130_fd_sc_hd__o21ai_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ _6093_/A1 _6093_/A2 _6090_/X _6092_/X VGND VGND VPWR VPWR _6094_/D sky130_fd_sc_hd__a211o_1
XFILLER_112_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _5136_/A _5044_/B _5130_/C _5174_/B VGND VGND VPWR VPWR _5044_/X sky130_fd_sc_hd__or4_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6995_ _7076_/CLK _6995_/D wire3981/X VGND VGND VPWR VPWR _6995_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_41_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5946_ _6317_/B2 _5946_/A2 _5935_/X _5945_/X _5946_/C1 VGND VGND VPWR VPWR _5946_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5877_ _6761_/Q _5949_/B1 _5877_/B1 _5877_/B2 VGND VGND VPWR VPWR _5877_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4828_ _4562_/A _4459_/B _4425_/B _4675_/Y VGND VGND VPWR VPWR _4828_/X sky130_fd_sc_hd__a31o_1
XFILLER_193_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4759_ _4759_/A _4759_/B VGND VGND VPWR VPWR _4759_/Y sky130_fd_sc_hd__nand2_1
XFILLER_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6429_ _6429_/A _6431_/B VGND VGND VPWR VPWR _6429_/X sky130_fd_sc_hd__and2_1
XFILLER_122_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length3150 _5824_/A2 VGND VGND VPWR VPWR wire3142/A sky130_fd_sc_hd__clkbuf_1
Xmax_length3161 _6214_/A2 VGND VGND VPWR VPWR wire3160/A sky130_fd_sc_hd__clkbuf_1
XFILLER_152_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2 hold2/A VGND VGND VPWR VPWR hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1080 _4294_/A VGND VGND VPWR VPWR _3636_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire1091 _3453_/B1 VGND VGND VPWR VPWR _3705_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_81_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5800_ _5800_/A1 _5800_/A2 _5800_/B1 _7031_/Q _5796_/X VGND VGND VPWR VPWR _5800_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6780_ _7196_/CLK _6780_/D _6780_/RESET_B VGND VGND VPWR VPWR _6780_/Q sky130_fd_sc_hd__dfrtp_1
X_3992_ _3992_/A _5229_/B VGND VGND VPWR VPWR _4000_/S sky130_fd_sc_hd__and2_2
X_5731_ _7163_/Q _5730_/X _6122_/S VGND VGND VPWR VPWR _7163_/D sky130_fd_sc_hd__mux2_1
XFILLER_188_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5662_ _6954_/Q _5712_/A2 _5735_/A2 _6032_/B2 _5657_/X VGND VGND VPWR VPWR _5681_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_175_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4613_ _4613_/A _4613_/B VGND VGND VPWR VPWR _4646_/B sky130_fd_sc_hd__or2_1
X_5593_ _6565_/Q _5593_/B VGND VGND VPWR VPWR _5593_/Y sky130_fd_sc_hd__nor2_1
XFILLER_190_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4544_ _4402_/A _4544_/B VGND VGND VPWR VPWR _4544_/X sky130_fd_sc_hd__and2b_1
Xhold402 _7019_/Q VGND VGND VPWR VPWR hold402/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 _6988_/Q VGND VGND VPWR VPWR hold413/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold424 _6791_/Q VGND VGND VPWR VPWR hold424/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 _6535_/Q VGND VGND VPWR VPWR hold435/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4475_ _4475_/A _4488_/B VGND VGND VPWR VPWR _4530_/A sky130_fd_sc_hd__nand2_1
Xhold446 _6799_/Q VGND VGND VPWR VPWR hold446/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 _6676_/Q VGND VGND VPWR VPWR hold457/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold468 _7120_/Q VGND VGND VPWR VPWR hold468/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6214_ _6214_/A1 _6214_/A2 _6214_/B1 _6937_/Q VGND VGND VPWR VPWR _6214_/X sky130_fd_sc_hd__a22o_1
XFILLER_104_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold479 _6507_/Q VGND VGND VPWR VPWR hold479/X sky130_fd_sc_hd__dlygate4sd3_1
X_3426_ _6169_/A1 _3426_/A2 _3426_/B1 _3426_/B2 VGND VGND VPWR VPWR _3426_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7194_ _7196_/CLK _7194_/D VGND VGND VPWR VPWR _7194_/Q sky130_fd_sc_hd__dfxtp_1
Xwire2709 _6014_/X VGND VGND VPWR VPWR _6022_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6145_ _7178_/Q _6144_/X _6219_/S VGND VGND VPWR VPWR _6145_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3357_ _6961_/Q _3437_/A2 _3441_/A2 _5849_/A1 wire855/X VGND VGND VPWR VPWR _3357_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ _6076_/A1 _6076_/A2 _6141_/B1 _6076_/B2 VGND VGND VPWR VPWR _6076_/X sky130_fd_sc_hd__a22o_1
X_3288_ _3288_/A hold83/X VGND VGND VPWR VPWR _3378_/B sky130_fd_sc_hd__and2_1
XFILLER_45_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5027_ _5027_/A _5027_/B VGND VGND VPWR VPWR _5109_/B sky130_fd_sc_hd__nor2_1
XFILLER_73_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6978_ _7083_/CLK _6978_/D wire4037/X VGND VGND VPWR VPWR _6978_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_179_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5929_ _6764_/Q _5949_/B1 _5929_/B1 _6313_/A1 VGND VGND VPWR VPWR _5929_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length925 _3318_/Y VGND VGND VPWR VPWR wire917/A sky130_fd_sc_hd__clkbuf_1
XFILLER_126_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout3838 wire3847/A VGND VGND VPWR VPWR _4070_/A2 sky130_fd_sc_hd__buf_6
XFILLER_122_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3900 wire3901/X VGND VGND VPWR VPWR wire3900/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3911 wire3912/X VGND VGND VPWR VPWR wire3911/X sky130_fd_sc_hd__clkbuf_1
XFILLER_150_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3922 input83/X VGND VGND VPWR VPWR wire3922/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3933 input76/X VGND VGND VPWR VPWR wire3933/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3999 wire3999/A VGND VGND VPWR VPWR wire3999/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4260_ hold639/X _6394_/A0 _4263_/S VGND VGND VPWR VPWR _6712_/D sky130_fd_sc_hd__mux2_1
XFILLER_4_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3211_ hold92/A VGND VGND VPWR VPWR _3211_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4191_ _6648_/Q wire360/X _4196_/S VGND VGND VPWR VPWR _6648_/D sky130_fd_sc_hd__mux2_1
XFILLER_140_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6901_ _7031_/CLK _6901_/D wire4044/X VGND VGND VPWR VPWR _6901_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6832_ _7132_/CLK _6832_/D _6833_/RESET_B VGND VGND VPWR VPWR _6832_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3975_ hold14/X hold119/X _3981_/S VGND VGND VPWR VPWR hold15/A sky130_fd_sc_hd__mux2_1
X_6763_ _7067_/CLK _6763_/D wire3968/X VGND VGND VPWR VPWR _6763_/Q sky130_fd_sc_hd__dfstp_1
X_5714_ _5714_/A1 _5714_/A2 _5714_/B1 _5714_/B2 _5713_/X VGND VGND VPWR VPWR _5719_/B
+ sky130_fd_sc_hd__a221o_1
X_6694_ _7206_/CLK _6694_/D _4189_/B VGND VGND VPWR VPWR _6694_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5645_ _7146_/Q _7147_/Q _5600_/Y VGND VGND VPWR VPWR _5645_/X sky130_fd_sc_hd__or3b_1
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5576_ _5576_/A0 hold137/X _5576_/S VGND VGND VPWR VPWR _7131_/D sky130_fd_sc_hd__mux2_1
XFILLER_156_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold210 _6947_/Q VGND VGND VPWR VPWR hold210/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4527_ _4527_/A1 _4872_/A _4652_/A _4940_/A _4525_/X VGND VGND VPWR VPWR _4528_/D
+ sky130_fd_sc_hd__o221a_1
Xhold221 _7088_/Q VGND VGND VPWR VPWR hold221/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 _7108_/Q VGND VGND VPWR VPWR hold232/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 _6680_/Q VGND VGND VPWR VPWR hold243/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 _6619_/Q VGND VGND VPWR VPWR hold254/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3207 _4482_/B VGND VGND VPWR VPWR _4637_/A1 sky130_fd_sc_hd__clkbuf_1
Xhold265 _7113_/Q VGND VGND VPWR VPWR hold265/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold276 _6539_/Q VGND VGND VPWR VPWR hold276/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3218 _4485_/B VGND VGND VPWR VPWR _4521_/A sky130_fd_sc_hd__clkbuf_2
X_4458_ _4846_/C _4738_/A VGND VGND VPWR VPWR _5001_/B sky130_fd_sc_hd__nor2_1
Xhold287 _4297_/X VGND VGND VPWR VPWR _6743_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2506 wire2506/A VGND VGND VPWR VPWR _6302_/B1 sky130_fd_sc_hd__clkbuf_2
Xhold298 _7068_/Q VGND VGND VPWR VPWR hold298/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3409_ _3409_/A _3409_/B _3409_/C _3409_/D VGND VGND VPWR VPWR _3409_/X sky130_fd_sc_hd__or4_1
Xwire2517 _6204_/A2 VGND VGND VPWR VPWR _6152_/A2 sky130_fd_sc_hd__clkbuf_2
X_7177_ _3937_/A1 _7177_/D wire4007/A VGND VGND VPWR VPWR _7177_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4389_ _4654_/A _4547_/A VGND VGND VPWR VPWR _4389_/Y sky130_fd_sc_hd__nor2_1
Xwire2528 _6162_/A2 VGND VGND VPWR VPWR _6139_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2539 _6127_/B1 VGND VGND VPWR VPWR _6150_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6128_ _7030_/Q _6186_/A2 _6128_/B1 _6128_/B2 VGND VGND VPWR VPWR _6128_/X sky130_fd_sc_hd__a22o_1
Xwire1816 wire1817/X VGND VGND VPWR VPWR wire1816/X sky130_fd_sc_hd__clkbuf_1
XFILLER_105_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1827 _6998_/Q VGND VGND VPWR VPWR wire1827/X sky130_fd_sc_hd__clkbuf_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1838 wire1839/X VGND VGND VPWR VPWR wire1838/X sky130_fd_sc_hd__clkbuf_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1849 wire1850/X VGND VGND VPWR VPWR _6104_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6059_ _6059_/A1 _6296_/A2 _6296_/B1 _6059_/B2 _6050_/X VGND VGND VPWR VPWR _6059_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_39_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_105 clkbuf_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_116 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 wire2819/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3730 _6779_/Q VGND VGND VPWR VPWR _5088_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire3741 _4776_/B2 VGND VGND VPWR VPWR wire3741/X sky130_fd_sc_hd__clkbuf_1
Xwire3752 wire3753/X VGND VGND VPWR VPWR wire3752/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3763 wire3764/X VGND VGND VPWR VPWR wire3763/X sky130_fd_sc_hd__clkbuf_1
Xwire3774 wire3775/X VGND VGND VPWR VPWR _6170_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire3785 wire3786/X VGND VGND VPWR VPWR wire3785/X sky130_fd_sc_hd__clkbuf_1
Xwire3796 _6458_/Q VGND VGND VPWR VPWR wire3796/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3760_ _3760_/A _3760_/B _3760_/C _3760_/D VGND VGND VPWR VPWR _3760_/X sky130_fd_sc_hd__or4_1
XFILLER_192_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3691_ _3691_/A1 wire929/A wire872/X _6059_/B2 _3690_/X VGND VGND VPWR VPWR _3691_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5430_ _5430_/A _5430_/B VGND VGND VPWR VPWR _5438_/S sky130_fd_sc_hd__nand2_2
XFILLER_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5361_ _5574_/A0 hold266/X _5361_/S VGND VGND VPWR VPWR _6940_/D sky130_fd_sc_hd__mux2_1
Xoutput304 _6810_/Q VGND VGND VPWR VPWR pwr_ctrl_out[3] sky130_fd_sc_hd__buf_12
XFILLER_161_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput315 wire3712/X VGND VGND VPWR VPWR spimemio_flash_io2_di sky130_fd_sc_hd__buf_12
Xoutput326 _6627_/Q VGND VGND VPWR VPWR wb_dat_o[17] sky130_fd_sc_hd__buf_12
Xoutput337 wire3717/X VGND VGND VPWR VPWR wb_dat_o[27] sky130_fd_sc_hd__buf_12
X_4312_ _4312_/A _4324_/B VGND VGND VPWR VPWR _4317_/S sky130_fd_sc_hd__and2_1
X_7100_ _7102_/CLK _7100_/D wire4004/A VGND VGND VPWR VPWR _7100_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput348 _6639_/Q VGND VGND VPWR VPWR wb_dat_o[8] sky130_fd_sc_hd__buf_12
XFILLER_99_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5292_ _5490_/A0 hold499/X _5294_/S VGND VGND VPWR VPWR _6879_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7031_ _7031_/CLK _7031_/D wire4048/X VGND VGND VPWR VPWR _7031_/Q sky130_fd_sc_hd__dfrtp_1
X_4243_ hold432/X _4249_/A0 _4245_/S VGND VGND VPWR VPWR _6688_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4174_ _4174_/A _4222_/B VGND VGND VPWR VPWR _4179_/S sky130_fd_sc_hd__nand2_2
XFILLER_95_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6815_ _7080_/CLK _6815_/D wire3992/A VGND VGND VPWR VPWR _6815_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6746_ _6963_/CLK _6746_/D _6401_/A VGND VGND VPWR VPWR _6746_/Q sky130_fd_sc_hd__dfrtp_1
Xmax_length3705 _3195_/Y VGND VGND VPWR VPWR wire3704/A sky130_fd_sc_hd__clkbuf_1
XFILLER_50_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3958_ _3958_/A _3958_/B VGND VGND VPWR VPWR _3958_/X sky130_fd_sc_hd__and2_1
XFILLER_50_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire409 _4082_/S VGND VGND VPWR VPWR _4078_/S sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_length3716 _7193_/Q VGND VGND VPWR VPWR wire3715/A sky130_fd_sc_hd__clkbuf_1
XFILLER_137_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3889_ _6696_/Q _3876_/X _3888_/B _6691_/Q VGND VGND VPWR VPWR _6696_/D sky130_fd_sc_hd__a22o_1
X_6677_ _7091_/CLK _6677_/D fanout4028/X VGND VGND VPWR VPWR _6677_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_137_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5628_ _6564_/Q _7154_/Q _7153_/Q VGND VGND VPWR VPWR _5637_/B sky130_fd_sc_hd__and3_1
XFILLER_191_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5559_ _5586_/A0 hold600/X _5561_/S VGND VGND VPWR VPWR _7116_/D sky130_fd_sc_hd__mux2_1
Xwire3004 _5839_/A2 VGND VGND VPWR VPWR _5760_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_144_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3026 wire3027/X VGND VGND VPWR VPWR _5831_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire3037 _5675_/X VGND VGND VPWR VPWR wire3037/X sky130_fd_sc_hd__clkbuf_1
XFILLER_78_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2303 _6261_/B2 VGND VGND VPWR VPWR wire2303/X sky130_fd_sc_hd__clkbuf_1
Xwire3048 _5951_/B1 VGND VGND VPWR VPWR _5883_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_104_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3059 wire3060/X VGND VGND VPWR VPWR _5868_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire2314 _6617_/Q VGND VGND VPWR VPWR _6246_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2325 _6610_/Q VGND VGND VPWR VPWR _3520_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire2336 _6604_/Q VGND VGND VPWR VPWR _6314_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1602 _7087_/Q VGND VGND VPWR VPWR _6149_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_76_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2347 _6569_/Q VGND VGND VPWR VPWR wire2347/X sky130_fd_sc_hd__clkbuf_2
Xwire2358 _5907_/B2 VGND VGND VPWR VPWR _6289_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire1613 wire1614/X VGND VGND VPWR VPWR _6201_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire2369 wire2370/X VGND VGND VPWR VPWR _6248_/A sky130_fd_sc_hd__clkbuf_2
Xwire1624 _7077_/Q VGND VGND VPWR VPWR _5757_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1635 _7067_/Q VGND VGND VPWR VPWR _6053_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1646 _5734_/A1 VGND VGND VPWR VPWR _6088_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire1657 _6165_/A1 VGND VGND VPWR VPWR _3426_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_100_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1668 _7052_/Q VGND VGND VPWR VPWR _5744_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1679 wire1680/X VGND VGND VPWR VPWR wire1679/X sky130_fd_sc_hd__clkbuf_1
XFILLER_74_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_1_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A VGND VGND VPWR VPWR _7187_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_27_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire910 wire911/X VGND VGND VPWR VPWR wire910/X sky130_fd_sc_hd__clkbuf_2
Xwire921 wire922/X VGND VGND VPWR VPWR wire921/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire932 _3312_/Y VGND VGND VPWR VPWR _5268_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xwire943 wire944/X VGND VGND VPWR VPWR wire943/X sky130_fd_sc_hd__clkbuf_1
Xwire954 _5304_/A VGND VGND VPWR VPWR wire954/X sky130_fd_sc_hd__clkbuf_1
XFILLER_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire965 wire966/X VGND VGND VPWR VPWR wire965/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire987 _6217_/A VGND VGND VPWR VPWR _6119_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire998 wire999/X VGND VGND VPWR VPWR wire998/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length596 _5515_/S VGND VGND VPWR VPWR _5517_/S sky130_fd_sc_hd__clkbuf_1
XFILLER_170_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4250 input18/X VGND VGND VPWR VPWR wire4250/X sky130_fd_sc_hd__clkbuf_1
Xfanout3454 wire3466/A VGND VGND VPWR VPWR _4179_/A0 sky130_fd_sc_hd__clkbuf_1
Xwire4261 wire4262/X VGND VGND VPWR VPWR wire4261/X sky130_fd_sc_hd__clkbuf_2
Xwire4272 input16/X VGND VGND VPWR VPWR wire4272/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire4283 _4476_/A VGND VGND VPWR VPWR _4588_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3560 _5352_/A0 VGND VGND VPWR VPWR _4114_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3571 wire3572/X VGND VGND VPWR VPWR wire3571/X sky130_fd_sc_hd__clkbuf_1
Xwire3582 _4206_/A1 VGND VGND VPWR VPWR _4122_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_96_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3593 _5555_/A0 VGND VGND VPWR VPWR _6394_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2870 _5700_/X VGND VGND VPWR VPWR _5701_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2881 _5699_/X VGND VGND VPWR VPWR _5701_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_77_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2892 _5697_/X VGND VGND VPWR VPWR _5698_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4930_ _4930_/A _4964_/A _4930_/C VGND VGND VPWR VPWR _5068_/B sky130_fd_sc_hd__or3_1
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4861_ _4639_/B _4707_/B _4510_/A VGND VGND VPWR VPWR _4862_/D sky130_fd_sc_hd__o21ai_1
XFILLER_60_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6600_ _7090_/CLK _6600_/D wire3948/X VGND VGND VPWR VPWR _6600_/Q sky130_fd_sc_hd__dfstp_1
X_3812_ _3828_/S _3811_/X _3810_/Y VGND VGND VPWR VPWR _6470_/D sky130_fd_sc_hd__o21ai_1
X_4792_ _4792_/A _4792_/B _4792_/C VGND VGND VPWR VPWR _4795_/B sky130_fd_sc_hd__or3_1
XANTENNA_16 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_27 wire903/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_38 _6257_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6531_ _7210_/CLK _6531_/D wire3950/X VGND VGND VPWR VPWR _6531_/Q sky130_fd_sc_hd__dfrtp_1
X_3743_ _6681_/Q _4234_/A _4222_/A _6675_/Q VGND VGND VPWR VPWR _3743_/X sky130_fd_sc_hd__a22o_1
XANTENNA_49 _6208_/C1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6462_ _6545_/CLK _6462_/D _6417_/X VGND VGND VPWR VPWR _6462_/Q sky130_fd_sc_hd__dfrtp_1
X_3674_ _5212_/A _3674_/B VGND VGND VPWR VPWR _3674_/Y sky130_fd_sc_hd__nor2_1
XFILLER_134_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5413_ _5485_/A0 hold560/X _5413_/S VGND VGND VPWR VPWR _6986_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6393_ _6393_/A0 hold373/X _6395_/S VGND VGND VPWR VPWR _7207_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5344_ _5398_/A1 _5344_/A1 _5348_/S VGND VGND VPWR VPWR _6925_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput178 _3222_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[12] sky130_fd_sc_hd__buf_12
Xoutput189 _3212_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[22] sky130_fd_sc_hd__buf_12
X_5275_ _5356_/A0 hold500/X _5275_/S VGND VGND VPWR VPWR _6864_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7014_ _7134_/CLK _7014_/D fanout4057/X VGND VGND VPWR VPWR _7014_/Q sky130_fd_sc_hd__dfrtp_1
X_4226_ _4256_/A1 _4226_/A1 _4227_/S VGND VGND VPWR VPWR _6678_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4157_ _4274_/A1 hold254/X hold58/X VGND VGND VPWR VPWR _6619_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4088_ hold330/X _5242_/A0 _4100_/S VGND VGND VPWR VPWR _4088_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4258 _4189_/B VGND VGND VPWR VPWR _6348_/B sky130_fd_sc_hd__buf_4
X_6729_ _7104_/CLK _6729_/D wire4040/X VGND VGND VPWR VPWR _6729_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_149_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length2812 _6138_/A2 VGND VGND VPWR VPWR _5985_/A2 sky130_fd_sc_hd__clkbuf_1
Xmax_length3557 _5487_/A0 VGND VGND VPWR VPWR _5523_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_192_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_52_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7142_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_191_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2100 wire2101/X VGND VGND VPWR VPWR _3783_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2111 _6818_/Q VGND VGND VPWR VPWR _3380_/S sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2122 _6810_/Q VGND VGND VPWR VPWR wire2122/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_67_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7027_/CLK sky130_fd_sc_hd__clkbuf_16
Xwire2133 wire2134/X VGND VGND VPWR VPWR wire2133/X sky130_fd_sc_hd__clkbuf_1
Xwire2144 _6791_/Q VGND VGND VPWR VPWR _3782_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_59_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2155 _6772_/Q VGND VGND VPWR VPWR _6254_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire1410 _6221_/X VGND VGND VPWR VPWR wire1410/X sky130_fd_sc_hd__clkbuf_1
Xwire2166 _3491_/B2 VGND VGND VPWR VPWR _6322_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire1421 _5746_/X VGND VGND VPWR VPWR _5747_/C1 sky130_fd_sc_hd__clkbuf_1
Xwire2177 wire2178/X VGND VGND VPWR VPWR _6234_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_59_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1432 _4982_/A VGND VGND VPWR VPWR _4634_/D sky130_fd_sc_hd__clkbuf_1
Xwire2188 _6742_/Q VGND VGND VPWR VPWR wire2188/X sky130_fd_sc_hd__clkbuf_1
XFILLER_101_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1443 _5135_/A1 VGND VGND VPWR VPWR _4858_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1454 wire1455/X VGND VGND VPWR VPWR wire1454/X sky130_fd_sc_hd__clkbuf_1
Xwire2199 wire2200/X VGND VGND VPWR VPWR _6223_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire1465 wire1466/X VGND VGND VPWR VPWR wire1465/X sky130_fd_sc_hd__clkbuf_1
Xwire1476 wire1477/X VGND VGND VPWR VPWR wire1476/X sky130_fd_sc_hd__clkbuf_1
Xwire1487 _3923_/X VGND VGND VPWR VPWR wire1487/X sky130_fd_sc_hd__clkbuf_1
XFILLER_74_554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1498 _3478_/B VGND VGND VPWR VPWR _3492_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_34_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput14 mask_rev_in[19] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__clkbuf_1
XFILLER_168_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput25 mask_rev_in[29] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__clkbuf_1
Xwire740 wire741/X VGND VGND VPWR VPWR wire740/X sky130_fd_sc_hd__clkbuf_1
Xinput36 mgmt_gpio_in[0] VGND VGND VPWR VPWR input36/X sky130_fd_sc_hd__clkbuf_1
Xwire751 _3717_/X VGND VGND VPWR VPWR wire751/X sky130_fd_sc_hd__clkbuf_1
Xinput47 mgmt_gpio_in[1] VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__clkbuf_1
Xwire762 _3693_/X VGND VGND VPWR VPWR wire762/X sky130_fd_sc_hd__clkbuf_1
Xinput58 mgmt_gpio_in[2] VGND VGND VPWR VPWR input58/X sky130_fd_sc_hd__clkbuf_2
Xwire773 _3615_/X VGND VGND VPWR VPWR wire773/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire784 _3554_/X VGND VGND VPWR VPWR wire784/X sky130_fd_sc_hd__clkbuf_1
Xinput69 mgmt_gpio_in[6] VGND VGND VPWR VPWR input69/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire795 wire795/A VGND VGND VPWR VPWR wire795/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3390_ _6904_/Q _5313_/A wire907/X input41/X _3389_/X VGND VGND VPWR VPWR _3390_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4080 wire4086/A VGND VGND VPWR VPWR wire4080/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire4091 wire4092/X VGND VGND VPWR VPWR wire4091/X sky130_fd_sc_hd__clkbuf_2
X_5060_ _5060_/A _5060_/B VGND VGND VPWR VPWR _5127_/C sky130_fd_sc_hd__and2_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3390 hold3/X VGND VGND VPWR VPWR _5240_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
X_4011_ hold551/X _5530_/A1 _4014_/S VGND VGND VPWR VPWR _6506_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5962_ _6337_/A1 _5962_/A2 _5962_/B1 _6327_/B2 _5961_/X VGND VGND VPWR VPWR _5967_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_52_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4913_ _4400_/B _5105_/B2 _4913_/B1 _5023_/B VGND VGND VPWR VPWR _4913_/X sky130_fd_sc_hd__o22a_1
X_5893_ _6666_/Q _5905_/A2 _5893_/B1 _6264_/A1 _5892_/X VGND VGND VPWR VPWR _5901_/A
+ sky130_fd_sc_hd__a221o_1
X_4844_ _4926_/A _5050_/B VGND VGND VPWR VPWR _5068_/A sky130_fd_sc_hd__nand2_1
XFILLER_138_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4775_ _4899_/B _4875_/B _4773_/X _4774_/Y _4992_/C VGND VGND VPWR VPWR _4775_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_119_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6514_ _6799_/CLK _6514_/D wire3935/X VGND VGND VPWR VPWR _6514_/Q sky130_fd_sc_hd__dfrtp_1
X_3726_ _3726_/A _3726_/B VGND VGND VPWR VPWR _5223_/A sky130_fd_sc_hd__nor2_1
XFILLER_174_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6445_ _3945_/A1 _6445_/D _6400_/X VGND VGND VPWR VPWR _6445_/Q sky130_fd_sc_hd__dfrtp_2
X_3657_ _3657_/A1_N _3525_/B _4135_/A _6603_/Q VGND VGND VPWR VPWR _3657_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_134_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6376_ _4228_/C _6376_/A2 _6376_/B1 _4228_/A _6375_/X VGND VGND VPWR VPWR _6376_/X
+ sky130_fd_sc_hd__a221o_1
X_3588_ _3588_/A _3588_/B _3588_/C _3588_/D VGND VGND VPWR VPWR _3601_/B sky130_fd_sc_hd__or4_1
X_5327_ hold289/X _5585_/A0 _5327_/S VGND VGND VPWR VPWR _6910_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5258_ hold652/X _5456_/A0 _5258_/S VGND VGND VPWR VPWR _6849_/D sky130_fd_sc_hd__mux2_1
XFILLER_57_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4209_ hold484/X _4209_/A1 _4209_/S VGND VGND VPWR VPWR _6664_/D sky130_fd_sc_hd__mux2_1
X_5189_ _5195_/A0 hold495/X _5192_/S VGND VGND VPWR VPWR _6794_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_579 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length4000 wire4001/X VGND VGND VPWR VPWR wire3999/A sky130_fd_sc_hd__buf_2
XFILLER_12_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3376 _5561_/A0 VGND VGND VPWR VPWR _5579_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_165_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length1930 _6930_/Q VGND VGND VPWR VPWR wire1927/A sky130_fd_sc_hd__clkbuf_1
XFILLER_98_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length1974 _6909_/Q VGND VGND VPWR VPWR wire1973/A sky130_fd_sc_hd__clkbuf_1
XFILLER_79_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length1996 _6895_/Q VGND VGND VPWR VPWR _3438_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_79_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1240 _3783_/A2 VGND VGND VPWR VPWR _3605_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1251 _3617_/A2 VGND VGND VPWR VPWR _3480_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1262 _3295_/Y VGND VGND VPWR VPWR _3678_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1273 _5502_/A VGND VGND VPWR VPWR _3393_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire1284 wire1285/X VGND VGND VPWR VPWR _3698_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1295 _3490_/A VGND VGND VPWR VPWR _3726_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_19_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4560_ _4560_/A _4573_/B VGND VGND VPWR VPWR _4560_/Y sky130_fd_sc_hd__nand2_1
XFILLER_190_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire570 _3458_/X VGND VGND VPWR VPWR _3468_/B sky130_fd_sc_hd__clkbuf_1
X_3511_ _3511_/A _3511_/B VGND VGND VPWR VPWR _3511_/Y sky130_fd_sc_hd__nor2_1
Xwire581 _3350_/X VGND VGND VPWR VPWR wire581/X sky130_fd_sc_hd__clkbuf_1
Xhold606 _6845_/Q VGND VGND VPWR VPWR hold606/X sky130_fd_sc_hd__dlygate4sd3_1
X_4491_ _4520_/A _4491_/B VGND VGND VPWR VPWR _4993_/B sky130_fd_sc_hd__nand2_1
Xhold617 _7040_/Q VGND VGND VPWR VPWR hold617/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire592 _5542_/S VGND VGND VPWR VPWR _5543_/S sky130_fd_sc_hd__clkbuf_2
Xhold628 _6992_/Q VGND VGND VPWR VPWR hold628/X sky130_fd_sc_hd__dlygate4sd3_1
X_6230_ _6230_/A1 _6336_/A2 _6273_/B1 _7207_/Q VGND VGND VPWR VPWR _6230_/X sky130_fd_sc_hd__a22o_1
X_3442_ _3442_/A1 _3442_/A2 _3442_/B1 _3442_/B2 _3441_/X VGND VGND VPWR VPWR _3445_/C
+ sky130_fd_sc_hd__a221o_1
Xhold639 _6712_/Q VGND VGND VPWR VPWR hold639/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3373_ _3373_/A _3373_/B _3373_/C VGND VGND VPWR VPWR _3373_/X sky130_fd_sc_hd__or3_1
XFILLER_97_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6161_ _6951_/Q _6161_/A2 _6173_/B1 _7047_/Q VGND VGND VPWR VPWR _6161_/X sky130_fd_sc_hd__a22o_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _5112_/A _5112_/B _5112_/C _5112_/D VGND VGND VPWR VPWR _5140_/B sky130_fd_sc_hd__or4_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ _7137_/Q _6092_/A2 _6092_/B1 _6092_/B2 _6091_/X VGND VGND VPWR VPWR _6092_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _5043_/A1 _4448_/B _4506_/Y _4984_/B _5007_/B VGND VGND VPWR VPWR _5174_/B
+ sky130_fd_sc_hd__a2111o_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_wbbd_sck _7205_/Q VGND VGND VPWR VPWR clkbuf_0_wbbd_sck/X sky130_fd_sc_hd__clkbuf_16
XFILLER_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6994_ _7076_/CLK _6994_/D wire3974/X VGND VGND VPWR VPWR _6994_/Q sky130_fd_sc_hd__dfstp_1
X_5945_ _5945_/A _5945_/B _5945_/C _5945_/D VGND VGND VPWR VPWR _5945_/X sky130_fd_sc_hd__or4_1
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5876_ _6238_/B2 _5936_/A2 _5920_/A2 _6222_/A _5875_/X VGND VGND VPWR VPWR _5879_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4827_ _4848_/A1 _4679_/B _4510_/C VGND VGND VPWR VPWR _5064_/B sky130_fd_sc_hd__o21ai_1
X_4758_ _4758_/A _4758_/B _4758_/C _4876_/B VGND VGND VPWR VPWR _4758_/Y sky130_fd_sc_hd__nand4_4
XFILLER_193_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3709_ _3709_/A1 _3709_/A2 wire887/X _3709_/B2 _3708_/X VGND VGND VPWR VPWR _3710_/D
+ sky130_fd_sc_hd__a221o_1
Xmax_length1204 _5394_/A VGND VGND VPWR VPWR _3570_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_162_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4689_ _4689_/A _4689_/B VGND VGND VPWR VPWR _4689_/X sky130_fd_sc_hd__or2_1
X_6428_ _6433_/A _6428_/B VGND VGND VPWR VPWR _6428_/X sky130_fd_sc_hd__and2_1
XFILLER_122_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6359_ _4228_/C _6357_/Y _6358_/Y _4228_/B VGND VGND VPWR VPWR _6362_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length3195 _4802_/A VGND VGND VPWR VPWR _4807_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_125_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length2494 _6211_/B1 VGND VGND VPWR VPWR wire2493/A sky130_fd_sc_hd__clkbuf_1
XFILLER_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3 hold3/A VGND VGND VPWR VPWR hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_94_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1070 _3596_/B1 VGND VGND VPWR VPWR _3480_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1081 _3464_/B1 VGND VGND VPWR VPWR _3664_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire1092 _3594_/B1 VGND VGND VPWR VPWR _3453_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_663 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3991_ hold705/X _3991_/A1 _3991_/S VGND VGND VPWR VPWR _6489_/D sky130_fd_sc_hd__mux2_1
X_5730_ _6121_/A1 _7162_/Q wire589/X VGND VGND VPWR VPWR _5730_/X sky130_fd_sc_hd__a21o_1
XFILLER_62_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5661_ _5683_/A _5700_/C _5703_/C VGND VGND VPWR VPWR _5661_/X sky130_fd_sc_hd__and3_1
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4612_ _4784_/B _5018_/C VGND VGND VPWR VPWR _4618_/C sky130_fd_sc_hd__or2_1
XFILLER_191_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5592_ _5593_/B _5592_/B VGND VGND VPWR VPWR _5592_/Y sky130_fd_sc_hd__nand2_1
XFILLER_129_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4543_ _4935_/A _4588_/A VGND VGND VPWR VPWR _4621_/C sky130_fd_sc_hd__nand2b_1
XFILLER_156_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold403 _7137_/Q VGND VGND VPWR VPWR hold403/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold414 _6804_/Q VGND VGND VPWR VPWR hold414/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold425 _6868_/Q VGND VGND VPWR VPWR hold425/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold436 _6689_/Q VGND VGND VPWR VPWR hold436/X sky130_fd_sc_hd__dlygate4sd3_1
X_4474_ _4474_/A _4839_/B VGND VGND VPWR VPWR _5060_/A sky130_fd_sc_hd__nor2_1
Xhold447 _6852_/Q VGND VGND VPWR VPWR hold447/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 _6800_/Q VGND VGND VPWR VPWR hold458/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold469 _7033_/Q VGND VGND VPWR VPWR hold469/X sky130_fd_sc_hd__dlygate4sd3_1
X_6213_ _6865_/Q _6213_/A2 _6213_/B1 _6213_/B2 _6212_/X VGND VGND VPWR VPWR _6216_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_116_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3425_ input17/X _3682_/A2 _3425_/B1 _3425_/B2 VGND VGND VPWR VPWR _3425_/X sky130_fd_sc_hd__a22o_1
X_7193_ _7193_/CLK _7193_/D VGND VGND VPWR VPWR _7193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3356_ _7033_/Q _5457_/A _3682_/B1 input28/X VGND VGND VPWR VPWR _3356_/X sky130_fd_sc_hd__a22o_1
X_6144_ _6144_/A1 _6133_/X wire584/X _6046_/B _6846_/Q VGND VGND VPWR VPWR _6144_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3287_ _3510_/A _3714_/A VGND VGND VPWR VPWR _3287_/Y sky130_fd_sc_hd__nor2_2
X_6075_ _6075_/A1 _6075_/A2 _6075_/B1 _6075_/B2 _6074_/X VGND VGND VPWR VPWR _6085_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5026_ _5152_/A1 _4655_/B _4679_/B _5027_/B VGND VGND VPWR VPWR _5029_/D sky130_fd_sc_hd__a31o_1
XFILLER_72_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_671 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6977_ _7031_/CLK _6977_/D wire4048/X VGND VGND VPWR VPWR _6977_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5928_ _6744_/Q _5928_/A2 _5928_/B1 _6534_/Q _5928_/C1 VGND VGND VPWR VPWR _5935_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5859_ _5859_/A1 _7168_/Q _5858_/X VGND VGND VPWR VPWR _5859_/X sky130_fd_sc_hd__a21o_1
XFILLER_139_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire3901 wire3902/X VGND VGND VPWR VPWR wire3901/X sky130_fd_sc_hd__clkbuf_1
Xwire3912 wire3913/X VGND VGND VPWR VPWR wire3912/X sky130_fd_sc_hd__clkbuf_1
Xwire3923 input82/X VGND VGND VPWR VPWR _3922_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_134_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3945 wire3945/A VGND VGND VPWR VPWR wire3945/X sky130_fd_sc_hd__clkbuf_4
Xwire3956 wire3956/A VGND VGND VPWR VPWR wire3956/X sky130_fd_sc_hd__buf_2
XFILLER_1_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3978 wire3981/A VGND VGND VPWR VPWR wire3978/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3210_ _3210_/A VGND VGND VPWR VPWR _3210_/Y sky130_fd_sc_hd__inv_2
X_4190_ _6647_/Q wire358/X _4196_/S VGND VGND VPWR VPWR _6647_/D sky130_fd_sc_hd__mux2_1
XFILLER_192_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6900_ _7084_/CLK _6900_/D wire4052/X VGND VGND VPWR VPWR _6900_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6831_ _7132_/CLK _6831_/D _6833_/RESET_B VGND VGND VPWR VPWR _6831_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6762_ _7067_/CLK _6762_/D wire3968/X VGND VGND VPWR VPWR _6762_/Q sky130_fd_sc_hd__dfrtp_1
X_3974_ hold712/X _3974_/A1 _3976_/S VGND VGND VPWR VPWR _6477_/D sky130_fd_sc_hd__mux2_1
XFILLER_149_702 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5713_ _6987_/Q _5713_/A2 _5713_/B1 _6979_/Q VGND VGND VPWR VPWR _5713_/X sky130_fd_sc_hd__a22o_1
X_6693_ _7193_/CLK _6693_/D _6348_/B VGND VGND VPWR VPWR _6693_/Q sky130_fd_sc_hd__dfrtp_1
X_5644_ _6564_/Q _5642_/X _5643_/Y _7158_/Q VGND VGND VPWR VPWR _7158_/D sky130_fd_sc_hd__a22o_1
XFILLER_136_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5575_ _5575_/A0 _3198_/A _5579_/S VGND VGND VPWR VPWR _7130_/D sky130_fd_sc_hd__mux2_1
Xhold200 _7106_/Q VGND VGND VPWR VPWR hold200/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 _6881_/Q VGND VGND VPWR VPWR hold211/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4526_ _4872_/A _4526_/B VGND VGND VPWR VPWR _4843_/A sky130_fd_sc_hd__nor2_1
Xhold222 _6931_/Q VGND VGND VPWR VPWR hold222/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 _6831_/Q VGND VGND VPWR VPWR hold233/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 _3281_/X VGND VGND VPWR VPWR hold244/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 _7060_/Q VGND VGND VPWR VPWR hold255/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3208 _4482_/B VGND VGND VPWR VPWR _4687_/B sky130_fd_sc_hd__clkbuf_2
Xhold266 _6940_/Q VGND VGND VPWR VPWR hold266/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4457_ _4460_/A _4521_/A VGND VGND VPWR VPWR _4504_/B sky130_fd_sc_hd__nand2_1
Xwire3219 _4450_/Y VGND VGND VPWR VPWR _4485_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold277 _6540_/Q VGND VGND VPWR VPWR hold277/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold288 _6625_/Q VGND VGND VPWR VPWR hold288/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold299 _6515_/Q VGND VGND VPWR VPWR hold299/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire2507 _6128_/B1 VGND VGND VPWR VPWR _6111_/A2 sky130_fd_sc_hd__clkbuf_1
X_3408_ _3408_/A _3408_/B _3408_/C _3408_/D VGND VGND VPWR VPWR _3409_/D sky130_fd_sc_hd__or4_1
XFILLER_132_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7176_ _7185_/CLK _7176_/D _7176_/RESET_B VGND VGND VPWR VPWR _7176_/Q sky130_fd_sc_hd__dfrtp_1
Xwire2518 _6176_/B1 VGND VGND VPWR VPWR _6204_/A2 sky130_fd_sc_hd__clkbuf_2
X_4388_ _4390_/A _4654_/A VGND VGND VPWR VPWR _4467_/C sky130_fd_sc_hd__nor2_1
Xwire2529 _6213_/A2 VGND VGND VPWR VPWR _6162_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_86_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1806 _5732_/A1 VGND VGND VPWR VPWR _6073_/A1 sky130_fd_sc_hd__clkbuf_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6127_ _7078_/Q _6127_/A2 _6127_/B1 _6127_/B2 _6125_/X VGND VGND VPWR VPWR _6127_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1817 wire1818/X VGND VGND VPWR VPWR wire1817/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3339_ _3466_/A _3339_/B VGND VGND VPWR VPWR _3339_/Y sky130_fd_sc_hd__nor2_1
Xwire1828 wire1829/X VGND VGND VPWR VPWR _3215_/A sky130_fd_sc_hd__clkbuf_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1839 wire1840/X VGND VGND VPWR VPWR wire1839/X sky130_fd_sc_hd__clkbuf_1
XFILLER_39_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6058_ _6058_/A _6058_/B _6058_/C _6058_/D VGND VGND VPWR VPWR _6069_/B sky130_fd_sc_hd__or4_1
XFILLER_85_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5009_ _5009_/A _5045_/B _5049_/D _5009_/D VGND VGND VPWR VPWR _5010_/D sky130_fd_sc_hd__or4_1
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_106 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_117 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_128 _4000_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout3603 hold37/X VGND VGND VPWR VPWR hold38/A sky130_fd_sc_hd__buf_6
XFILLER_146_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3720 wire3721/X VGND VGND VPWR VPWR _5881_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_123_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3731 hold140/X VGND VGND VPWR VPWR _3258_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire3742 _6776_/Q VGND VGND VPWR VPWR _4776_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3753 _6698_/Q VGND VGND VPWR VPWR wire3753/X sky130_fd_sc_hd__clkbuf_1
Xwire3764 _3963_/B VGND VGND VPWR VPWR wire3764/X sky130_fd_sc_hd__clkbuf_1
Xwire3775 _6563_/Q VGND VGND VPWR VPWR wire3775/X sky130_fd_sc_hd__clkbuf_1
XFILLER_39_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3786 wire3787/X VGND VGND VPWR VPWR wire3786/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3797 hold6/X VGND VGND VPWR VPWR _3965_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3690_ _7104_/Q wire867/X _4276_/A _6727_/Q VGND VGND VPWR VPWR _3690_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5360_ _5573_/A0 hold186/X _5361_/S VGND VGND VPWR VPWR _6939_/D sky130_fd_sc_hd__mux2_1
Xoutput305 _3730_/X VGND VGND VPWR VPWR reset sky130_fd_sc_hd__buf_12
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput316 _7215_/X VGND VGND VPWR VPWR spimemio_flash_io3_di sky130_fd_sc_hd__buf_12
Xoutput327 _6628_/Q VGND VGND VPWR VPWR wb_dat_o[18] sky130_fd_sc_hd__buf_12
X_4311_ _4311_/A0 hold360/X _4311_/S VGND VGND VPWR VPWR _6755_/D sky130_fd_sc_hd__mux2_1
Xoutput338 wire3715/X VGND VGND VPWR VPWR wb_dat_o[28] sky130_fd_sc_hd__buf_12
Xoutput349 _6640_/Q VGND VGND VPWR VPWR wb_dat_o[9] sky130_fd_sc_hd__buf_12
X_5291_ _5291_/A0 hold75/X _5291_/S VGND VGND VPWR VPWR hold76/A sky130_fd_sc_hd__mux2_1
XFILLER_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7030_ _7115_/CLK _7030_/D _7030_/RESET_B VGND VGND VPWR VPWR _7030_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4242_ hold438/X _4242_/A1 _4245_/S VGND VGND VPWR VPWR _6687_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4173_ _6633_/Q wire378/X _4173_/S VGND VGND VPWR VPWR _6633_/D sky130_fd_sc_hd__mux2_1
XFILLER_122_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6814_ _7080_/CLK _6814_/D wire3992/A VGND VGND VPWR VPWR _6814_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6745_ _6799_/CLK _6745_/D _6743_/SET_B VGND VGND VPWR VPWR _6745_/Q sky130_fd_sc_hd__dfrtp_1
X_3957_ _3957_/A _3957_/B VGND VGND VPWR VPWR _3957_/X sky130_fd_sc_hd__and2_1
XFILLER_31_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6676_ _7091_/CLK _6676_/D wire4029/A VGND VGND VPWR VPWR _6676_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3888_ _6691_/Q _3888_/B VGND VGND VPWR VPWR _3888_/Y sky130_fd_sc_hd__nand2_1
XFILLER_149_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5627_ _7154_/Q _7153_/Q VGND VGND VPWR VPWR _6033_/A sky130_fd_sc_hd__and2_2
X_5558_ _5558_/A0 hold667/X _5560_/S VGND VGND VPWR VPWR _7115_/D sky130_fd_sc_hd__mux2_1
XFILLER_191_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4509_ _4512_/B _4514_/B VGND VGND VPWR VPWR _4510_/C sky130_fd_sc_hd__nand2_1
XFILLER_132_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5489_ _5489_/A0 hold452/X _5489_/S VGND VGND VPWR VPWR _7054_/D sky130_fd_sc_hd__mux2_1
XFILLER_4_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3005 _5830_/A2 VGND VGND VPWR VPWR _5839_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3027 _5848_/B1 VGND VGND VPWR VPWR wire3027/X sky130_fd_sc_hd__clkbuf_1
Xwire3038 _5675_/X VGND VGND VPWR VPWR _5849_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3049 _5943_/A2 VGND VGND VPWR VPWR _5951_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire2304 _6635_/Q VGND VGND VPWR VPWR _6261_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2315 wire2316/X VGND VGND VPWR VPWR _5878_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2326 _6610_/Q VGND VGND VPWR VPWR _6326_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_76_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2337 _6602_/Q VGND VGND VPWR VPWR _6264_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
X_7159_ _7180_/CLK _7159_/D _7159_/RESET_B VGND VGND VPWR VPWR _7159_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2348 _6568_/Q VGND VGND VPWR VPWR _3926_/A0 sky130_fd_sc_hd__clkbuf_1
Xwire1603 _7086_/Q VGND VGND VPWR VPWR _6125_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire1614 _3345_/B2 VGND VGND VPWR VPWR wire1614/X sky130_fd_sc_hd__clkbuf_1
Xwire2359 _6538_/Q VGND VGND VPWR VPWR _5907_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1625 wire1626/X VGND VGND VPWR VPWR _6091_/A1 sky130_fd_sc_hd__clkbuf_2
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1636 wire1637/X VGND VGND VPWR VPWR _6042_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire1647 _7060_/Q VGND VGND VPWR VPWR _5734_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1658 _7055_/Q VGND VGND VPWR VPWR _6165_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1669 _7051_/Q VGND VGND VPWR VPWR _5711_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire900 wire903/X VGND VGND VPWR VPWR wire900/X sky130_fd_sc_hd__clkbuf_1
Xwire911 wire912/X VGND VGND VPWR VPWR wire911/X sky130_fd_sc_hd__dlymetal6s2s_1
Xwire922 wire924/X VGND VGND VPWR VPWR wire922/X sky130_fd_sc_hd__clkbuf_2
Xwire933 wire937/X VGND VGND VPWR VPWR wire933/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire944 _3308_/Y VGND VGND VPWR VPWR wire944/X sky130_fd_sc_hd__clkbuf_2
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire955 _3280_/Y VGND VGND VPWR VPWR _5304_/A sky130_fd_sc_hd__clkbuf_2
Xwire966 wire966/A VGND VGND VPWR VPWR wire966/X sky130_fd_sc_hd__clkbuf_1
Xwire977 _6046_/B VGND VGND VPWR VPWR wire977/X sky130_fd_sc_hd__clkbuf_2
XFILLER_127_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire988 _6168_/A VGND VGND VPWR VPWR _6069_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_170_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire999 wire999/A VGND VGND VPWR VPWR wire999/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4240 input27/X VGND VGND VPWR VPWR wire4240/X sky130_fd_sc_hd__clkbuf_1
XFILLER_123_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4251 wire4252/X VGND VGND VPWR VPWR wire4251/X sky130_fd_sc_hd__clkbuf_1
XFILLER_123_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4262 wire4263/X VGND VGND VPWR VPWR wire4262/X sky130_fd_sc_hd__clkbuf_1
XFILLER_150_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4273 wire4274/X VGND VGND VPWR VPWR _3697_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_151_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire4284 _4476_/A VGND VGND VPWR VPWR _4379_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout3488 wire3498/X VGND VGND VPWR VPWR _6396_/A0 sky130_fd_sc_hd__buf_6
Xwire4295 _4846_/B VGND VGND VPWR VPWR _4566_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_1_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3550 _5451_/A0 VGND VGND VPWR VPWR _5208_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_123_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3561 _5574_/A0 VGND VGND VPWR VPWR _5352_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3572 wire3573/X VGND VGND VPWR VPWR wire3572/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3594 _5495_/A0 VGND VGND VPWR VPWR _5555_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2860 _5782_/A2 VGND VGND VPWR VPWR _5958_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire2871 _5733_/B1 VGND VGND VPWR VPWR _5712_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire2882 _5817_/B1 VGND VGND VPWR VPWR _5783_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_64_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2893 _5803_/A2 VGND VGND VPWR VPWR _5763_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_66_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4860_ _4860_/A _4860_/B _4860_/C _4860_/D VGND VGND VPWR VPWR _4862_/C sky130_fd_sc_hd__nand4_1
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3811_ _3242_/X _3243_/Y _3811_/S VGND VGND VPWR VPWR _3811_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4791_ _4994_/A _4805_/B2 _4799_/B1 _5027_/A VGND VGND VPWR VPWR _4987_/C sky130_fd_sc_hd__o22ai_1
XANTENNA_17 input64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 _4252_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6530_ _6811_/CLK _6530_/D wire3935/X VGND VGND VPWR VPWR _6530_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_39 _6180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3742_ _6032_/B2 wire919/X wire875/X _5981_/B2 _3741_/X VGND VGND VPWR VPWR _3749_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_186_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6461_ _6545_/CLK _6461_/D _6416_/X VGND VGND VPWR VPWR _6461_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_158_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3673_ _6955_/Q _3744_/A2 _4270_/A _6256_/B2 _3672_/X VGND VGND VPWR VPWR _3673_/X
+ sky130_fd_sc_hd__a221o_1
X_5412_ _5412_/A _5535_/B VGND VGND VPWR VPWR _5417_/S sky130_fd_sc_hd__nand2_1
XFILLER_161_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6392_ _6392_/A _6392_/B VGND VGND VPWR VPWR _6396_/S sky130_fd_sc_hd__nand2_1
XFILLER_133_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5343_ _5343_/A0 hold307/X _5343_/S VGND VGND VPWR VPWR _6924_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput179 _3221_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[13] sky130_fd_sc_hd__buf_12
X_5274_ _5364_/A0 hold623/X _5274_/S VGND VGND VPWR VPWR _6863_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7013_ _7130_/CLK _7013_/D wire4061/X VGND VGND VPWR VPWR _7013_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_102_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4225_ _4255_/A1 _4225_/A1 _4227_/S VGND VGND VPWR VPWR _6677_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4156_ _4273_/A1 _6618_/Q hold58/X VGND VGND VPWR VPWR hold59/A sky130_fd_sc_hd__mux2_1
XFILLER_83_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4087_ _5241_/B _5241_/C _4052_/X _3333_/Y _5286_/B VGND VGND VPWR VPWR _4087_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_83_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4989_ _4980_/X _5119_/B _4989_/C _4989_/D VGND VGND VPWR VPWR _4990_/B sky130_fd_sc_hd__and4bb_1
X_6728_ _7104_/CLK _6728_/D wire4042/A VGND VGND VPWR VPWR _6728_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_137_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length3536 _4309_/A0 VGND VGND VPWR VPWR _5196_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_149_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6659_ _7094_/CLK _6659_/D wire3965/A VGND VGND VPWR VPWR _6659_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_137_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length2835 _5706_/X VGND VGND VPWR VPWR _5822_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_192_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length2846 _5705_/X VGND VGND VPWR VPWR wire2845/A sky130_fd_sc_hd__clkbuf_1
XFILLER_164_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2868 _5931_/B1 VGND VGND VPWR VPWR _5875_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_191_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2101 wire2101/A VGND VGND VPWR VPWR wire2101/X sky130_fd_sc_hd__clkbuf_1
XFILLER_160_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2123 wire2124/X VGND VGND VPWR VPWR _3604_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_120_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2134 _6807_/Q VGND VGND VPWR VPWR wire2134/X sky130_fd_sc_hd__clkbuf_1
Xwire1400 _3472_/A VGND VGND VPWR VPWR _3314_/A sky130_fd_sc_hd__clkbuf_2
Xwire2145 _3535_/B2 VGND VGND VPWR VPWR _6321_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2156 _6771_/Q VGND VGND VPWR VPWR _6229_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1411 _6197_/X VGND VGND VPWR VPWR _6208_/C1 sky130_fd_sc_hd__clkbuf_1
Xwire2167 _6750_/Q VGND VGND VPWR VPWR _3491_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1422 _5741_/X VGND VGND VPWR VPWR _5742_/C1 sky130_fd_sc_hd__clkbuf_1
Xwire1433 _4560_/Y VGND VGND VPWR VPWR _4794_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_19_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2178 wire2179/X VGND VGND VPWR VPWR wire2178/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1444 _4424_/Y VGND VGND VPWR VPWR _5135_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire2189 _6741_/Q VGND VGND VPWR VPWR _6234_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1455 wire1456/X VGND VGND VPWR VPWR wire1455/X sky130_fd_sc_hd__clkbuf_1
XFILLER_74_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1466 wire1467/X VGND VGND VPWR VPWR wire1466/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1477 wire1478/X VGND VGND VPWR VPWR wire1477/X sky130_fd_sc_hd__clkbuf_1
Xwire1488 wire1489/X VGND VGND VPWR VPWR wire1488/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1499 _3414_/Y VGND VGND VPWR VPWR _3478_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_74_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput15 mask_rev_in[1] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__clkbuf_1
Xwire730 _4003_/S VGND VGND VPWR VPWR _4007_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_167_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput26 mask_rev_in[2] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__clkbuf_1
Xwire741 wire742/X VGND VGND VPWR VPWR wire741/X sky130_fd_sc_hd__clkbuf_1
Xwire752 wire753/X VGND VGND VPWR VPWR wire752/X sky130_fd_sc_hd__clkbuf_1
Xinput37 mgmt_gpio_in[10] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__clkbuf_1
Xinput48 mgmt_gpio_in[20] VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__clkbuf_1
Xwire763 _3684_/X VGND VGND VPWR VPWR wire763/X sky130_fd_sc_hd__clkbuf_1
Xinput59 mgmt_gpio_in[30] VGND VGND VPWR VPWR input59/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire774 _3613_/X VGND VGND VPWR VPWR wire774/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire785 _3552_/X VGND VGND VPWR VPWR wire785/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire4081 wire4082/X VGND VGND VPWR VPWR wire4081/X sky130_fd_sc_hd__buf_2
Xwire4092 wire4092/A VGND VGND VPWR VPWR wire4092/X sky130_fd_sc_hd__clkbuf_1
Xwire3380 _5429_/A0 VGND VGND VPWR VPWR _5519_/A0 sky130_fd_sc_hd__clkbuf_2
Xwire3391 hold2/X VGND VGND VPWR VPWR hold3/A sky130_fd_sc_hd__clkbuf_2
X_4010_ _4010_/A _4135_/B VGND VGND VPWR VPWR _4014_/S sky130_fd_sc_hd__and2_1
XFILLER_38_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2690 _6016_/X VGND VGND VPWR VPWR _6024_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5961_ _6335_/A1 _5961_/A2 _5960_/X _5961_/B2 VGND VGND VPWR VPWR _5961_/X sky130_fd_sc_hd__a22o_1
X_4912_ _4912_/A1 _4680_/B _4910_/X _4911_/X _4646_/X VGND VGND VPWR VPWR _4912_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_61_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5892_ _6261_/A1 _5892_/A2 _5909_/B1 _6249_/B2 VGND VGND VPWR VPWR _5892_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4843_ _4843_/A _4843_/B VGND VGND VPWR VPWR _4866_/C sky130_fd_sc_hd__or2_1
XFILLER_166_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4774_ _5050_/B _4992_/B VGND VGND VPWR VPWR _4774_/Y sky130_fd_sc_hd__nand2_1
XFILLER_159_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6513_ _6799_/CLK _6513_/D wire3935/X VGND VGND VPWR VPWR _6513_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_186_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3725_ _3724_/X _6784_/Q _3791_/B VGND VGND VPWR VPWR _6784_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6444_ _6545_/CLK _6444_/D _6399_/X VGND VGND VPWR VPWR _6444_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3656_ _6276_/A1 _3656_/A2 _3656_/B1 _6288_/B2 _3655_/X VGND VGND VPWR VPWR _3658_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6375_ _4228_/B _6375_/A2 _6375_/B1 _4228_/Y VGND VGND VPWR VPWR _6375_/X sky130_fd_sc_hd__a22o_1
X_3587_ _3587_/A1 _3706_/B1 _3526_/Y _3587_/B2 wire786/X VGND VGND VPWR VPWR _3588_/D
+ sky130_fd_sc_hd__a221o_1
X_5326_ hold441/X _5380_/A0 _5330_/S VGND VGND VPWR VPWR _6909_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5257_ hold643/X _5509_/A0 _5258_/S VGND VGND VPWR VPWR _6848_/D sky130_fd_sc_hd__mux2_1
XFILLER_57_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4208_ hold490/X _4208_/A1 _4209_/S VGND VGND VPWR VPWR _6663_/D sky130_fd_sc_hd__mux2_1
XFILLER_180_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5188_ _5211_/A0 hold472/X _5192_/S VGND VGND VPWR VPWR _6793_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4139_ hold428/X _4139_/A1 _4139_/S VGND VGND VPWR VPWR _6604_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length4012 wire4013/X VGND VGND VPWR VPWR fanout4005/A sky130_fd_sc_hd__clkbuf_1
Xmax_length4023 wire4018/A VGND VGND VPWR VPWR wire4022/A sky130_fd_sc_hd__clkbuf_1
XFILLER_11_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4089 wire4090/X VGND VGND VPWR VPWR _7051_/SET_B sky130_fd_sc_hd__clkbuf_2
XFILLER_22_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length2610 _4742_/B VGND VGND VPWR VPWR _4758_/A sky130_fd_sc_hd__buf_2
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3366 _4369_/X VGND VGND VPWR VPWR _4497_/A sky130_fd_sc_hd__clkbuf_2
Xmax_length2621 _6212_/B1 VGND VGND VPWR VPWR _6103_/B1 sky130_fd_sc_hd__clkbuf_1
Xmax_length2632 _6148_/B VGND VGND VPWR VPWR _6099_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_125_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length3388 _5348_/A0 VGND VGND VPWR VPWR _5528_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_165_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3399 _5464_/A0 VGND VGND VPWR VPWR _5569_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_152_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1230 _3641_/A2 VGND VGND VPWR VPWR _3763_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1252 _3298_/Y VGND VGND VPWR VPWR _3617_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1263 _3439_/A2 VGND VGND VPWR VPWR _3777_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1274 _3292_/Y VGND VGND VPWR VPWR _5502_/A sky130_fd_sc_hd__clkbuf_1
Xwire1285 wire1286/X VGND VGND VPWR VPWR wire1285/X sky130_fd_sc_hd__clkbuf_1
XFILLER_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1296 _3518_/B VGND VGND VPWR VPWR _3546_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3510_ _3510_/A _3510_/B VGND VGND VPWR VPWR _4324_/A sky130_fd_sc_hd__nor2_1
Xwire560 _3565_/X VGND VGND VPWR VPWR wire560/X sky130_fd_sc_hd__clkbuf_1
Xwire571 wire572/X VGND VGND VPWR VPWR wire571/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire582 _6395_/S VGND VGND VPWR VPWR _6397_/S sky130_fd_sc_hd__clkbuf_2
X_4490_ _4872_/A _4942_/A VGND VGND VPWR VPWR _4490_/X sky130_fd_sc_hd__or2_1
XFILLER_155_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold607 _6898_/Q VGND VGND VPWR VPWR hold607/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 _6757_/Q VGND VGND VPWR VPWR hold618/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire593 _5533_/S VGND VGND VPWR VPWR _5534_/S sky130_fd_sc_hd__clkbuf_2
Xhold629 _6935_/Q VGND VGND VPWR VPWR hold629/X sky130_fd_sc_hd__dlygate4sd3_1
X_3441_ _3441_/A1 _3441_/A2 _3533_/A2 _3441_/B2 VGND VGND VPWR VPWR _3441_/X sky130_fd_sc_hd__a22o_1
XFILLER_109_590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6160_ _6927_/Q _6160_/A2 _6160_/B1 _6160_/B2 _6159_/X VGND VGND VPWR VPWR _6167_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3372_ _3372_/A _3372_/B VGND VGND VPWR VPWR _3373_/C sky130_fd_sc_hd__or2_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5111_ _5111_/A1 _5071_/A _5070_/Y _5110_/X VGND VGND VPWR VPWR _5139_/A sky130_fd_sc_hd__a22o_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _6091_/A1 _6201_/A2 _6115_/B1 _6091_/B2 VGND VGND VPWR VPWR _6091_/X sky130_fd_sc_hd__a22o_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5042_ _5042_/A _5042_/B _5042_/C VGND VGND VPWR VPWR _5130_/C sky130_fd_sc_hd__or3_1
XFILLER_69_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6993_ _7110_/CLK _6993_/D _7110_/RESET_B VGND VGND VPWR VPWR _6993_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_92_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_51_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7126_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_53_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5944_ _6304_/A1 _5944_/A2 _5944_/B1 _6298_/B2 _5943_/X VGND VGND VPWR VPWR _5945_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5875_ _6227_/A1 _5875_/A2 _5941_/B1 _6235_/B2 VGND VGND VPWR VPWR _5875_/X sky130_fd_sc_hd__a22o_1
XFILLER_33_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4826_ _4704_/A _4707_/B _4515_/B VGND VGND VPWR VPWR _5064_/A sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_66_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7056_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_147_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4757_ _4760_/A1 _5113_/A2 _5135_/A1 VGND VGND VPWR VPWR _4761_/C sky130_fd_sc_hd__a21oi_1
XFILLER_193_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3708_ _7112_/Q wire963/X _3747_/B1 _6261_/A1 VGND VGND VPWR VPWR _3708_/X sky130_fd_sc_hd__a22o_1
XFILLER_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4688_ _5021_/A _4688_/B _5021_/C VGND VGND VPWR VPWR _4713_/B sky130_fd_sc_hd__or3_1
XFILLER_161_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6427_ _6433_/A _6428_/B VGND VGND VPWR VPWR _6427_/X sky130_fd_sc_hd__and2_1
X_3639_ _3639_/A1 _3331_/Y _5221_/B _3639_/B2 _3638_/X VGND VGND VPWR VPWR _3642_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_108_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6358_ _6358_/A _6358_/B VGND VGND VPWR VPWR _6358_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5309_ _5309_/A0 hold494/X _5311_/S VGND VGND VPWR VPWR _6894_/D sky130_fd_sc_hd__mux2_1
X_6289_ _6289_/A1 _6289_/A2 _6325_/A2 _6657_/Q VGND VGND VPWR VPWR _6289_/X sky130_fd_sc_hd__a22o_1
XFILLER_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_19_csclk _6579_/CLK VGND VGND VPWR VPWR _6939_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__1134_ clkbuf_0__1134_/X VGND VGND VPWR VPWR _6353_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_138_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold4 hold4/A VGND VGND VPWR VPWR hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1060 _3486_/B1 VGND VGND VPWR VPWR _3699_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire1071 _3476_/Y VGND VGND VPWR VPWR _3596_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1082 wire1083/X VGND VGND VPWR VPWR _3464_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_35_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3990_ hold706/X _5437_/A0 _3991_/S VGND VGND VPWR VPWR _6488_/D sky130_fd_sc_hd__mux2_1
XFILLER_90_675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5660_ _7149_/Q _7148_/Q VGND VGND VPWR VPWR _5703_/C sky130_fd_sc_hd__and2b_1
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4611_ _4611_/A _4645_/B VGND VGND VPWR VPWR _4611_/X sky130_fd_sc_hd__or2_1
X_5591_ _5593_/B _6564_/Q VGND VGND VPWR VPWR _5651_/B sky130_fd_sc_hd__nor2_1
X_4542_ _4542_/A _4792_/A VGND VGND VPWR VPWR _4546_/B sky130_fd_sc_hd__nand2_1
XFILLER_116_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold404 _6668_/Q VGND VGND VPWR VPWR hold404/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire390 _3446_/X VGND VGND VPWR VPWR wire390/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold415 _6655_/Q VGND VGND VPWR VPWR hold415/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold426 _6686_/Q VGND VGND VPWR VPWR hold426/X sky130_fd_sc_hd__dlygate4sd3_1
X_4473_ _4944_/A _4947_/A VGND VGND VPWR VPWR _4839_/B sky130_fd_sc_hd__or2_1
Xhold437 _6690_/Q VGND VGND VPWR VPWR hold437/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold448 _6884_/Q VGND VGND VPWR VPWR hold448/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold459 _6675_/Q VGND VGND VPWR VPWR hold459/X sky130_fd_sc_hd__dlygate4sd3_1
X_6212_ _6212_/A1 _6212_/A2 _6212_/B1 _7049_/Q VGND VGND VPWR VPWR _6212_/X sky130_fd_sc_hd__a22o_1
X_3424_ input40/X wire907/X _5322_/A _6911_/Q VGND VGND VPWR VPWR _3424_/X sky130_fd_sc_hd__a22o_1
X_7192_ _7193_/CLK _7192_/D VGND VGND VPWR VPWR _7192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6143_ _6168_/A _6143_/B _6143_/C VGND VGND VPWR VPWR _6143_/X sky130_fd_sc_hd__or3_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3355_ _3355_/A _3355_/B _3355_/C _3355_/D VGND VGND VPWR VPWR _3373_/A sky130_fd_sc_hd__or4_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6074_ _6074_/A1 _6074_/A2 _6074_/B1 _6074_/B2 _6073_/X VGND VGND VPWR VPWR _6074_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3286_ _3714_/A VGND VGND VPWR VPWR _3286_/Y sky130_fd_sc_hd__inv_2
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5025_ _4582_/B _5108_/A _5024_/A _5027_/B VGND VGND VPWR VPWR _5029_/C sky130_fd_sc_hd__a31o_1
XFILLER_66_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6976_ _7031_/CLK _6976_/D wire4048/X VGND VGND VPWR VPWR _6976_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5927_ _6619_/Q _5927_/A2 _5927_/B1 _5927_/B2 VGND VGND VPWR VPWR _5927_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5858_ _6849_/Q _5858_/A2 _5847_/X _5857_/X _5858_/C1 VGND VGND VPWR VPWR _5858_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_22_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4809_ _5095_/B _4809_/B _4809_/C VGND VGND VPWR VPWR _4810_/B sky130_fd_sc_hd__and3b_1
XFILLER_166_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length916 _3319_/Y VGND VGND VPWR VPWR _3571_/A2 sky130_fd_sc_hd__clkbuf_1
X_5789_ _5789_/A1 _5789_/A2 _5789_/B1 _6125_/A1 _5788_/X VGND VGND VPWR VPWR _5792_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_182_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length949 wire950/X VGND VGND VPWR VPWR wire946/A sky130_fd_sc_hd__clkbuf_1
XFILLER_119_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length1046 _3511_/Y VGND VGND VPWR VPWR _3754_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_150_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3902 input87/X VGND VGND VPWR VPWR wire3902/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3913 input85/X VGND VGND VPWR VPWR wire3913/X sky130_fd_sc_hd__clkbuf_1
Xwire3924 input81/X VGND VGND VPWR VPWR _3925_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_135_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3935 wire3935/A VGND VGND VPWR VPWR wire3935/X sky130_fd_sc_hd__clkbuf_4
XFILLER_103_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3968 wire3968/A VGND VGND VPWR VPWR wire3968/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6830_ _7130_/CLK hold34/X _6833_/RESET_B VGND VGND VPWR VPWR hold33/A sky130_fd_sc_hd__dfrtp_1
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6761_ _6761_/CLK _6761_/D wire4019/X VGND VGND VPWR VPWR _6761_/Q sky130_fd_sc_hd__dfrtp_1
X_3973_ hold47/X hold722/X _3981_/S VGND VGND VPWR VPWR hold48/A sky130_fd_sc_hd__mux2_1
X_5712_ _6955_/Q _5712_/A2 _5712_/B1 _6049_/A _5711_/X VGND VGND VPWR VPWR _5719_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_149_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6692_ _7193_/CLK _6692_/D _6780_/RESET_B VGND VGND VPWR VPWR _6692_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5643_ _5643_/A _5643_/B VGND VGND VPWR VPWR _5643_/Y sky130_fd_sc_hd__nor2_1
XFILLER_176_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5574_ _5574_/A0 hold261/X _5576_/S VGND VGND VPWR VPWR _7129_/D sky130_fd_sc_hd__mux2_1
Xhold201 _6829_/Q VGND VGND VPWR VPWR hold201/X sky130_fd_sc_hd__dlygate4sd3_1
X_4525_ _4527_/A1 _4997_/A _4490_/X _4522_/X _4524_/Y VGND VGND VPWR VPWR _4525_/X
+ sky130_fd_sc_hd__o2111a_1
Xhold212 _7134_/Q VGND VGND VPWR VPWR hold212/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 _6725_/Q VGND VGND VPWR VPWR hold223/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 _6740_/Q VGND VGND VPWR VPWR hold234/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 _6396_/X VGND VGND VPWR VPWR _7210_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 _6512_/Q VGND VGND VPWR VPWR hold256/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4456_ _4456_/A _4724_/B VGND VGND VPWR VPWR _4997_/A sky130_fd_sc_hd__or2_2
Xhold267 _6514_/Q VGND VGND VPWR VPWR hold267/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold278 _6745_/Q VGND VGND VPWR VPWR hold278/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold289 _6910_/Q VGND VGND VPWR VPWR hold289/X sky130_fd_sc_hd__dlygate4sd3_1
X_3407_ _3407_/A1 _3407_/A2 wire971/X _3407_/B2 _3406_/X VGND VGND VPWR VPWR _3408_/D
+ sky130_fd_sc_hd__a221o_1
Xwire2508 _6006_/Y VGND VGND VPWR VPWR _6128_/B1 sky130_fd_sc_hd__clkbuf_1
X_7175_ _7185_/CLK _7175_/D wire4007/A VGND VGND VPWR VPWR _7175_/Q sky130_fd_sc_hd__dfrtp_1
X_4387_ _4538_/A _4387_/B VGND VGND VPWR VPWR _4387_/Y sky130_fd_sc_hd__nand2_1
XFILLER_86_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6126_ _6902_/Q _6126_/A2 _6166_/B1 _6966_/Q _6124_/X VGND VGND VPWR VPWR _6142_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1807 _3653_/B2 VGND VGND VPWR VPWR _5732_/A1 sky130_fd_sc_hd__clkbuf_1
X_3338_ _3502_/B _3338_/B VGND VGND VPWR VPWR _3338_/Y sky130_fd_sc_hd__nor2_1
XFILLER_140_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1818 _7002_/Q VGND VGND VPWR VPWR wire1818/X sky130_fd_sc_hd__clkbuf_1
XFILLER_98_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1829 _6116_/B2 VGND VGND VPWR VPWR wire1829/X sky130_fd_sc_hd__clkbuf_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6057_ _6057_/A1 _6057_/A2 _6057_/B1 _6979_/Q _6056_/X VGND VGND VPWR VPWR _6058_/D
+ sky130_fd_sc_hd__a221o_1
X_3269_ _3941_/A hold159/X hold61/X VGND VGND VPWR VPWR _3297_/A sky130_fd_sc_hd__o21ai_1
X_5008_ _5008_/A _5008_/B _5008_/C _5008_/D VGND VGND VPWR VPWR _5009_/D sky130_fd_sc_hd__or4_1
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_129 _7185_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6959_ _7031_/CLK _6959_/D wire4048/X VGND VGND VPWR VPWR _6959_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_41_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout3626 wire3642/A VGND VGND VPWR VPWR _4235_/A0 sky130_fd_sc_hd__buf_6
XFILLER_122_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout3648 wire3661/A VGND VGND VPWR VPWR wire3652/A sky130_fd_sc_hd__buf_6
XFILLER_150_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3721 _5860_/A0 VGND VGND VPWR VPWR wire3721/X sky130_fd_sc_hd__clkbuf_1
XFILLER_150_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3732 wire3733/X VGND VGND VPWR VPWR _3260_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_123_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire3743 wire3744/X VGND VGND VPWR VPWR _4228_/C sky130_fd_sc_hd__buf_4
XFILLER_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3754 wire3755/X VGND VGND VPWR VPWR wire3754/X sky130_fd_sc_hd__clkbuf_1
XFILLER_150_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3765 wire3766/X VGND VGND VPWR VPWR _3981_/S sky130_fd_sc_hd__buf_4
Xwire3776 wire3777/X VGND VGND VPWR VPWR _5969_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire3787 _6462_/Q VGND VGND VPWR VPWR wire3787/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput306 _3957_/X VGND VGND VPWR VPWR ser_rx sky130_fd_sc_hd__buf_12
XFILLER_126_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput317 wire3719/X VGND VGND VPWR VPWR wb_ack_o sky130_fd_sc_hd__buf_12
X_4310_ _4334_/A0 hold353/X _4311_/S VGND VGND VPWR VPWR _6754_/D sky130_fd_sc_hd__mux2_1
Xoutput328 _6629_/Q VGND VGND VPWR VPWR wb_dat_o[19] sky130_fd_sc_hd__buf_12
XFILLER_99_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5290_ _5479_/A0 hold96/X _5294_/S VGND VGND VPWR VPWR _6877_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput339 _7194_/Q VGND VGND VPWR VPWR wb_dat_o[29] sky130_fd_sc_hd__buf_12
XFILLER_113_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4241_ hold426/X _4247_/A0 _4245_/S VGND VGND VPWR VPWR _6686_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4172_ _6632_/Q wire375/X _4173_/S VGND VGND VPWR VPWR _6632_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6813_ _7080_/CLK _6813_/D wire3992/A VGND VGND VPWR VPWR _6813_/Q sky130_fd_sc_hd__dfrtp_1
X_6744_ _6803_/CLK _6744_/D wire3950/A VGND VGND VPWR VPWR _6744_/Q sky130_fd_sc_hd__dfrtp_1
X_3956_ _6699_/Q _3962_/B VGND VGND VPWR VPWR _6693_/D sky130_fd_sc_hd__and2_1
XFILLER_188_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6675_ _7091_/CLK _6675_/D fanout4028/X VGND VGND VPWR VPWR _6675_/Q sky130_fd_sc_hd__dfrtp_1
X_3887_ _3887_/A _3887_/B _3887_/C _3887_/D VGND VGND VPWR VPWR _3887_/Y sky130_fd_sc_hd__nor4_1
X_5626_ _5610_/X _5650_/B _7153_/Q VGND VGND VPWR VPWR _7153_/D sky130_fd_sc_hd__mux2_1
X_5557_ _5575_/A0 hold202/X _5557_/S VGND VGND VPWR VPWR _7114_/D sky130_fd_sc_hd__mux2_1
XFILLER_151_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4508_ _4871_/A _4995_/A _4447_/Y _4505_/X _4507_/X VGND VGND VPWR VPWR _4508_/X
+ sky130_fd_sc_hd__o2111a_1
X_5488_ _5575_/A0 hold208/X _5490_/S VGND VGND VPWR VPWR _7053_/D sky130_fd_sc_hd__mux2_1
XFILLER_104_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3006 _5678_/X VGND VGND VPWR VPWR _5830_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3017 _5829_/A2 VGND VGND VPWR VPWR _5856_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3028 _5676_/X VGND VGND VPWR VPWR _5848_/B1 sky130_fd_sc_hd__clkbuf_2
X_4439_ _4443_/B _4456_/A VGND VGND VPWR VPWR _4486_/A sky130_fd_sc_hd__or2_1
Xwire3039 _5955_/A2 VGND VGND VPWR VPWR _5941_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2305 wire2306/X VGND VGND VPWR VPWR _6236_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_132_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2316 _6221_/B2 VGND VGND VPWR VPWR wire2316/X sky130_fd_sc_hd__clkbuf_1
Xwire2327 wire2328/X VGND VGND VPWR VPWR _6313_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_116_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7158_ _7180_/CLK _7158_/D wire4014/X VGND VGND VPWR VPWR _7158_/Q sky130_fd_sc_hd__dfrtp_2
Xwire2338 _6601_/Q VGND VGND VPWR VPWR _5864_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1604 _7085_/Q VGND VGND VPWR VPWR _3204_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_98_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2349 wire2350/X VGND VGND VPWR VPWR _3927_/A0 sky130_fd_sc_hd__clkbuf_1
Xwire1615 _7081_/Q VGND VGND VPWR VPWR _3345_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1626 _7076_/Q VGND VGND VPWR VPWR wire1626/X sky130_fd_sc_hd__clkbuf_1
X_6109_ _6109_/A _6109_/B _6109_/C _6109_/D VGND VGND VPWR VPWR _6110_/B sky130_fd_sc_hd__or4_1
XFILLER_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1637 wire1638/X VGND VGND VPWR VPWR wire1637/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1648 wire1649/X VGND VGND VPWR VPWR _3771_/A1 sky130_fd_sc_hd__clkbuf_1
X_7089_ _7089_/CLK _7089_/D wire4071/X VGND VGND VPWR VPWR _7089_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1659 wire1660/X VGND VGND VPWR VPWR _3487_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_58_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire901 wire902/X VGND VGND VPWR VPWR wire901/X sky130_fd_sc_hd__clkbuf_2
XFILLER_167_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire912 _3319_/Y VGND VGND VPWR VPWR wire912/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire934 wire935/X VGND VGND VPWR VPWR wire934/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire956 wire957/X VGND VGND VPWR VPWR wire956/X sky130_fd_sc_hd__clkbuf_1
XFILLER_157_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire978 wire981/X VGND VGND VPWR VPWR wire978/X sky130_fd_sc_hd__clkbuf_1
Xwire989 _6217_/A VGND VGND VPWR VPWR _6168_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_157_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout3423 wire3438/A VGND VGND VPWR VPWR _4110_/A0 sky130_fd_sc_hd__clkbuf_1
Xwire4230 input36/X VGND VGND VPWR VPWR wire4230/X sky130_fd_sc_hd__clkbuf_1
Xwire4241 input26/X VGND VGND VPWR VPWR _3641_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout3445 wire3466/X VGND VGND VPWR VPWR _4033_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_151_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4252 wire4253/X VGND VGND VPWR VPWR wire4252/X sky130_fd_sc_hd__clkbuf_1
Xfanout3467 _5237_/A0 VGND VGND VPWR VPWR _4116_/A0 sky130_fd_sc_hd__clkbuf_1
Xwire4263 wire4264/X VGND VGND VPWR VPWR wire4263/X sky130_fd_sc_hd__clkbuf_1
Xwire4274 wire4275/X VGND VGND VPWR VPWR wire4274/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire4285 wire4285/A VGND VGND VPWR VPWR _4476_/A sky130_fd_sc_hd__clkbuf_2
Xwire4296 _4570_/C VGND VGND VPWR VPWR _4846_/B sky130_fd_sc_hd__buf_2
Xwire3551 _5514_/A0 VGND VGND VPWR VPWR _5451_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3573 hold21/X VGND VGND VPWR VPWR wire3573/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3584 _4248_/A0 VGND VGND VPWR VPWR _4242_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2850 _5703_/X VGND VGND VPWR VPWR wire2850/X sky130_fd_sc_hd__clkbuf_1
Xwire3595 _5495_/A0 VGND VGND VPWR VPWR _5582_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2861 wire2861/A VGND VGND VPWR VPWR _5782_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire2872 _5778_/B1 VGND VGND VPWR VPWR _5733_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2883 _5856_/B1 VGND VGND VPWR VPWR _5817_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire2894 _5854_/A2 VGND VGND VPWR VPWR _5803_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_66_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3810_ _6470_/Q _3828_/S VGND VGND VPWR VPWR _3810_/Y sky130_fd_sc_hd__nand2_1
X_4790_ _4784_/B _4675_/A _4759_/Y VGND VGND VPWR VPWR _5114_/A sky130_fd_sc_hd__o21ai_1
XFILLER_177_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_18 wire419/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_29 _3464_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3741_ _5674_/A1 _3741_/A2 _4270_/A _6721_/Q VGND VGND VPWR VPWR _3741_/X sky130_fd_sc_hd__a22o_1
XFILLER_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6460_ _6545_/CLK _6460_/D _6415_/X VGND VGND VPWR VPWR _6460_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3672_ _3672_/A1 _3747_/A2 _3672_/B1 _5890_/A1 VGND VGND VPWR VPWR _3672_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5411_ _5411_/A0 hold464/X _5411_/S VGND VGND VPWR VPWR _6985_/D sky130_fd_sc_hd__mux2_1
X_6391_ hold54/A _6697_/Q _6391_/A3 _6391_/B1 VGND VGND VPWR VPWR _7206_/D sky130_fd_sc_hd__o31a_1
X_5342_ _5342_/A0 hold148/X _5343_/S VGND VGND VPWR VPWR _6923_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5273_ hold16/X hold18/X _5273_/S VGND VGND VPWR VPWR hold19/A sky130_fd_sc_hd__mux2_1
XFILLER_114_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7012_ _7104_/CLK _7012_/D wire4040/X VGND VGND VPWR VPWR _7012_/Q sky130_fd_sc_hd__dfrtp_1
X_4224_ _5531_/A1 hold457/X _4227_/S VGND VGND VPWR VPWR _6676_/D sky130_fd_sc_hd__mux2_1
Xfanout3990 fanout3993/X VGND VGND VPWR VPWR wire3992/A sky130_fd_sc_hd__buf_6
XFILLER_68_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4155_ _6394_/A0 hold463/X hold58/X VGND VGND VPWR VPWR _6617_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4086_ hold496/X _4085_/X _4086_/S VGND VGND VPWR VPWR _6561_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4988_ _5090_/B _4988_/B _5170_/A _4988_/D VGND VGND VPWR VPWR _4988_/Y sky130_fd_sc_hd__nor4_1
X_6727_ _7136_/CLK _6727_/D wire4042/A VGND VGND VPWR VPWR _6727_/Q sky130_fd_sc_hd__dfrtp_1
X_3939_ _7159_/Q _6815_/Q _3940_/S VGND VGND VPWR VPWR _3939_/X sky130_fd_sc_hd__mux2_1
Xmax_length3526 _4274_/A1 VGND VGND VPWR VPWR _4256_/A1 sky130_fd_sc_hd__clkbuf_1
Xmax_length3537 _6395_/A0 VGND VGND VPWR VPWR _4309_/A0 sky130_fd_sc_hd__clkbuf_2
X_6658_ _7094_/CLK _6658_/D wire3965/A VGND VGND VPWR VPWR _6658_/Q sky130_fd_sc_hd__dfrtp_1
Xmax_length2825 _5977_/X VGND VGND VPWR VPWR wire2819/A sky130_fd_sc_hd__clkbuf_1
XFILLER_137_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5609_ _6562_/Q _6564_/Q VGND VGND VPWR VPWR _5609_/Y sky130_fd_sc_hd__nor2_1
XFILLER_152_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6589_ _6811_/CLK _6589_/D _3946_/B VGND VGND VPWR VPWR _6589_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2113 wire2114/X VGND VGND VPWR VPWR _3639_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_132_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2124 wire2125/X VGND VGND VPWR VPWR wire2124/X sky130_fd_sc_hd__clkbuf_1
Xwire2135 _6805_/Q VGND VGND VPWR VPWR _3712_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire2146 wire2147/X VGND VGND VPWR VPWR _3535_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire2157 _6767_/Q VGND VGND VPWR VPWR _6258_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire1412 wire1413/X VGND VGND VPWR VPWR _6191_/C1 sky130_fd_sc_hd__clkbuf_1
XFILLER_120_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2168 wire2169/X VGND VGND VPWR VPWR _6309_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire1423 wire1424/X VGND VGND VPWR VPWR _5707_/C1 sky130_fd_sc_hd__clkbuf_1
Xwire2179 _3758_/B2 VGND VGND VPWR VPWR wire2179/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1445 _4485_/A VGND VGND VPWR VPWR _4425_/B sky130_fd_sc_hd__clkbuf_2
Xwire1456 wire1457/X VGND VGND VPWR VPWR wire1456/X sky130_fd_sc_hd__clkbuf_1
XFILLER_47_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1467 wire1468/X VGND VGND VPWR VPWR wire1467/X sky130_fd_sc_hd__clkbuf_1
XFILLER_74_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1478 wire1479/X VGND VGND VPWR VPWR wire1478/X sky130_fd_sc_hd__clkbuf_1
Xwire1489 _3919_/X VGND VGND VPWR VPWR wire1489/X sky130_fd_sc_hd__clkbuf_1
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire720 _4120_/X VGND VGND VPWR VPWR wire720/X sky130_fd_sc_hd__clkbuf_1
Xinput16 mask_rev_in[20] VGND VGND VPWR VPWR input16/X sky130_fd_sc_hd__clkbuf_1
Xwire731 wire732/X VGND VGND VPWR VPWR _4003_/S sky130_fd_sc_hd__clkbuf_2
Xinput27 mask_rev_in[30] VGND VGND VPWR VPWR input27/X sky130_fd_sc_hd__clkbuf_1
Xwire742 _3779_/X VGND VGND VPWR VPWR wire742/X sky130_fd_sc_hd__clkbuf_1
Xwire753 wire754/X VGND VGND VPWR VPWR wire753/X sky130_fd_sc_hd__clkbuf_1
Xinput38 mgmt_gpio_in[11] VGND VGND VPWR VPWR input38/X sky130_fd_sc_hd__clkbuf_1
Xinput49 mgmt_gpio_in[21] VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__clkbuf_1
Xwire764 wire765/X VGND VGND VPWR VPWR wire764/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire775 _3574_/X VGND VGND VPWR VPWR wire775/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire786 wire787/X VGND VGND VPWR VPWR wire786/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire797 wire798/X VGND VGND VPWR VPWR _4204_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_155_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout3253 wire3261/X VGND VGND VPWR VPWR _4324_/B sky130_fd_sc_hd__buf_6
XFILLER_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire4071 wire4071/A VGND VGND VPWR VPWR wire4071/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_151_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout3275 hold57/X VGND VGND VPWR VPWR _4234_/B sky130_fd_sc_hd__buf_6
XFILLER_111_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire4082 wire4083/X VGND VGND VPWR VPWR wire4082/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3370 _4170_/S VGND VGND VPWR VPWR _4173_/S sky130_fd_sc_hd__buf_2
Xwire3381 _5543_/A1 VGND VGND VPWR VPWR _5429_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2680 _6299_/B1 VGND VGND VPWR VPWR _6323_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2691 _6210_/B1 VGND VGND VPWR VPWR _6113_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5960_ _5960_/A _5960_/B VGND VGND VPWR VPWR _5960_/X sky130_fd_sc_hd__or2_1
XFILLER_52_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4911_ _5013_/B _5016_/A _4477_/X VGND VGND VPWR VPWR _4911_/X sky130_fd_sc_hd__a21o_1
XFILLER_80_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5891_ _5891_/A _5891_/B _5891_/C _5891_/D VGND VGND VPWR VPWR _5891_/X sky130_fd_sc_hd__or4_1
XFILLER_33_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4842_ _4842_/A1 _4675_/B _4860_/A VGND VGND VPWR VPWR _4842_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_60_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4773_ _4376_/A _5042_/A _5042_/B _4772_/X _4897_/A VGND VGND VPWR VPWR _4773_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_193_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6512_ _6799_/CLK _6512_/D wire3935/X VGND VGND VPWR VPWR _6512_/Q sky130_fd_sc_hd__dfrtp_1
X_3724_ wire360/X _6783_/Q _3791_/A VGND VGND VPWR VPWR _3724_/X sky130_fd_sc_hd__mux2_1
XFILLER_159_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6443_ _6443_/CLK _6443_/D _3873_/X VGND VGND VPWR VPWR _6443_/Q sky130_fd_sc_hd__dfstp_1
X_3655_ _6276_/B2 _3655_/A2 _3784_/B1 _6285_/B2 VGND VGND VPWR VPWR _3655_/X sky130_fd_sc_hd__a22o_1
XFILLER_106_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6374_ _6373_/X _7200_/Q _6386_/S VGND VGND VPWR VPWR _7200_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3586_ _6534_/Q _4040_/A _3776_/B1 _7210_/Q _3553_/X VGND VGND VPWR VPWR _3588_/C
+ sky130_fd_sc_hd__a221o_1
X_5325_ hold138/X _5547_/A0 _5325_/S VGND VGND VPWR VPWR _6908_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5256_ _6169_/A1 _5256_/A1 _5256_/S VGND VGND VPWR VPWR _5256_/X sky130_fd_sc_hd__mux2_1
X_4207_ _5908_/B2 _5532_/A1 _4209_/S VGND VGND VPWR VPWR _6662_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5187_ _5187_/A _5193_/B VGND VGND VPWR VPWR _5192_/S sky130_fd_sc_hd__nand2_2
XFILLER_29_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4138_ hold423/X _5532_/A1 _4139_/S VGND VGND VPWR VPWR _6603_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4069_ hold12/X _4068_/X _4069_/S VGND VGND VPWR VPWR hold13/A sky130_fd_sc_hd__mux2_1
XFILLER_43_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3312 _4613_/B VGND VGND VPWR VPWR _4630_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length4068 wire4069/X VGND VGND VPWR VPWR _7087_/RESET_B sky130_fd_sc_hd__buf_2
XFILLER_149_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length3389 _5240_/A0 VGND VGND VPWR VPWR _5348_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_164_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length1910 _6940_/Q VGND VGND VPWR VPWR _6082_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_164_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2677 _6200_/B1 VGND VGND VPWR VPWR _6118_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_180_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length1954 _6920_/Q VGND VGND VPWR VPWR _6187_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_98_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1220 _3346_/A2 VGND VGND VPWR VPWR _3396_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire1231 _3641_/A2 VGND VGND VPWR VPWR _3394_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire1242 _3762_/A2 VGND VGND VPWR VPWR _5421_/A sky130_fd_sc_hd__buf_2
XFILLER_59_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1253 _3599_/A2 VGND VGND VPWR VPWR _3393_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_101_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1264 _3500_/A2 VGND VGND VPWR VPWR _3439_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1275 _3693_/A2 VGND VGND VPWR VPWR _3550_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire1286 _3287_/Y VGND VGND VPWR VPWR wire1286/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1297 _3490_/A VGND VGND VPWR VPWR _3518_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_170_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire550 wire551/X VGND VGND VPWR VPWR _3679_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_190_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire561 _3539_/X VGND VGND VPWR VPWR wire561/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire572 _3436_/X VGND VGND VPWR VPWR wire572/X sky130_fd_sc_hd__clkbuf_1
Xhold608 _6913_/Q VGND VGND VPWR VPWR hold608/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire594 _5525_/S VGND VGND VPWR VPWR _5523_/S sky130_fd_sc_hd__clkbuf_2
Xhold619 _6596_/Q VGND VGND VPWR VPWR hold619/X sky130_fd_sc_hd__dlygate4sd3_1
X_3440_ _3440_/A1 _3440_/A2 wire930/X _3440_/B2 wire839/X VGND VGND VPWR VPWR _3446_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_128_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3371_ _3371_/A _3371_/B _3371_/C _3371_/D VGND VGND VPWR VPWR _3372_/B sky130_fd_sc_hd__or4_1
XFILLER_112_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5110_ _5156_/C _5178_/B _5110_/C VGND VGND VPWR VPWR _5110_/X sky130_fd_sc_hd__or3_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6090_ _6090_/A1 _6090_/A2 _6090_/B1 _7068_/Q VGND VGND VPWR VPWR _6090_/X sky130_fd_sc_hd__a22o_1
XFILLER_88_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5041_ _5133_/A1 _4487_/B _4897_/A _5039_/X _5040_/X VGND VGND VPWR VPWR _5044_/B
+ sky130_fd_sc_hd__a2111o_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_wb_clk_i wb_clk_i VGND VGND VPWR VPWR clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_93_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6992_ _7064_/CLK _6992_/D wire4045/X VGND VGND VPWR VPWR _6992_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_92_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5943_ _6305_/B2 _5943_/A2 _5943_/B1 _7093_/Q VGND VGND VPWR VPWR _5943_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5874_ _6225_/A1 _5931_/A2 _5943_/B1 _7090_/Q _5873_/X VGND VGND VPWR VPWR _5879_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_139_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4825_ _5158_/B _4823_/X _4824_/Y _4549_/Y VGND VGND VPWR VPWR _4825_/X sky130_fd_sc_hd__o31a_1
XFILLER_166_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4756_ _4417_/X _4744_/X _4755_/X _4876_/B VGND VGND VPWR VPWR _4761_/B sky130_fd_sc_hd__o22a_1
XFILLER_147_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3707_ _3707_/A1 wire860/X _3707_/B1 _6252_/B2 wire758/X VGND VGND VPWR VPWR _3710_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4687_ _4739_/A _4687_/B VGND VGND VPWR VPWR _4770_/A sky130_fd_sc_hd__nor2_1
XFILLER_174_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3638_ _6768_/Q _3767_/A2 _4312_/A _6758_/Q VGND VGND VPWR VPWR _3638_/X sky130_fd_sc_hd__a22o_1
X_6426_ _6433_/A _6428_/B VGND VGND VPWR VPWR _6426_/X sky130_fd_sc_hd__and2_1
Xmax_length1239 _3605_/B1 VGND VGND VPWR VPWR wire1238/A sky130_fd_sc_hd__clkbuf_1
XFILLER_162_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6357_ _6357_/A _6358_/A VGND VGND VPWR VPWR _6357_/Y sky130_fd_sc_hd__nand2_1
XFILLER_103_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3569_ _6117_/A1 _5580_/A _5544_/A _6099_/A1 VGND VGND VPWR VPWR _3569_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5308_ _5308_/A0 hold541/X _5310_/S VGND VGND VPWR VPWR _6893_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6288_ _6603_/Q _6314_/A2 _6314_/B1 _6288_/B2 _6287_/X VGND VGND VPWR VPWR _6288_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5239_ _5365_/A0 hold104/X _5240_/S VGND VGND VPWR VPWR _6832_/D sky130_fd_sc_hd__mux2_1
XFILLER_124_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold5 hold5/A VGND VGND VPWR VPWR hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1050 _3784_/B1 VGND VGND VPWR VPWR _3686_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1061 wire1062/X VGND VGND VPWR VPWR _3486_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire1072 _3476_/Y VGND VGND VPWR VPWR _4010_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1083 _3463_/Y VGND VGND VPWR VPWR wire1083/X sky130_fd_sc_hd__clkbuf_1
XFILLER_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1094 wire1095/X VGND VGND VPWR VPWR _3442_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_90_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4610_ _4610_/A _4666_/B VGND VGND VPWR VPWR _4610_/X sky130_fd_sc_hd__or2_1
X_5590_ _5615_/A _5590_/A2 _6565_/Q _3896_/X _5589_/X VGND VGND VPWR VPWR _7143_/D
+ sky130_fd_sc_hd__o311a_1
X_4541_ _4553_/A _4553_/B VGND VGND VPWR VPWR _4780_/A sky130_fd_sc_hd__nand2_1
XFILLER_175_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold405 _6665_/Q VGND VGND VPWR VPWR hold405/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire380 wire381/X VGND VGND VPWR VPWR wire380/X sky130_fd_sc_hd__clkbuf_1
XFILLER_144_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4472_ _4570_/A _4570_/D _4570_/C _4570_/B VGND VGND VPWR VPWR _4472_/X sky130_fd_sc_hd__or4bb_1
XFILLER_7_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire391 _3409_/X VGND VGND VPWR VPWR _3410_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_144_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold416 _6970_/Q VGND VGND VPWR VPWR hold416/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold427 _6805_/Q VGND VGND VPWR VPWR hold427/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold438 _6687_/Q VGND VGND VPWR VPWR hold438/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 _6828_/Q VGND VGND VPWR VPWR hold449/X sky130_fd_sc_hd__dlygate4sd3_1
X_3423_ _3423_/A1 _3423_/A2 _3423_/B1 _3423_/B2 wire844/X VGND VGND VPWR VPWR _3445_/B
+ sky130_fd_sc_hd__a221o_1
X_6211_ _6211_/A1 _6211_/A2 _6211_/B1 _6897_/Q _6210_/X VGND VGND VPWR VPWR _6217_/C
+ sky130_fd_sc_hd__a221o_1
X_7191_ _7193_/CLK _7191_/D VGND VGND VPWR VPWR _7191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6142_ _6142_/A _6142_/B _6142_/C _6142_/D VGND VGND VPWR VPWR _6143_/C sky130_fd_sc_hd__or4_1
X_3354_ _7142_/Q _3354_/A2 _5475_/A _5483_/A1 _3353_/X VGND VGND VPWR VPWR _3355_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6073_ _6073_/A1 _6073_/A2 _6073_/B1 _7121_/Q VGND VGND VPWR VPWR _6073_/X sky130_fd_sc_hd__a22o_1
XFILLER_57_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3285_ _3313_/B hold84/X VGND VGND VPWR VPWR _3285_/Y sky130_fd_sc_hd__nand2_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _5024_/A _5027_/B VGND VGND VPWR VPWR _5155_/A sky130_fd_sc_hd__nor2_1
XFILLER_26_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6975_ _7079_/CLK _6975_/D wire4048/X VGND VGND VPWR VPWR _6975_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5926_ _7172_/Q _5925_/X _5948_/S VGND VGND VPWR VPWR _7172_/D sky130_fd_sc_hd__mux2_1
XFILLER_81_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5857_ _5857_/A _5857_/B _5857_/C _5857_/D VGND VGND VPWR VPWR _5857_/X sky130_fd_sc_hd__or4_1
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4808_ _4611_/A _4565_/X _4712_/B _4424_/Y _4981_/B VGND VGND VPWR VPWR _4809_/C
+ sky130_fd_sc_hd__o32a_1
XFILLER_186_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5788_ _5788_/A1 _5788_/A2 _5788_/B1 _5788_/B2 VGND VGND VPWR VPWR _5788_/X sky130_fd_sc_hd__a22o_1
X_4739_ _4739_/A _4739_/B VGND VGND VPWR VPWR _5042_/B sky130_fd_sc_hd__nor2_1
Xmax_length1003 _6171_/S VGND VGND VPWR VPWR _6122_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_134_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6409_ _6441_/A _6437_/B VGND VGND VPWR VPWR _6409_/X sky130_fd_sc_hd__and2_1
Xwire3903 wire3904/X VGND VGND VPWR VPWR _3947_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_122_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3914 wire3915/X VGND VGND VPWR VPWR _3943_/A0 sky130_fd_sc_hd__clkbuf_1
Xwire3925 input80/X VGND VGND VPWR VPWR _3923_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3958 wire3959/X VGND VGND VPWR VPWR wire3958/X sky130_fd_sc_hd__buf_2
XFILLER_0_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_50_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7124_/CLK sky130_fd_sc_hd__clkbuf_16
Xmax_length1592 _7096_/Q VGND VGND VPWR VPWR _3671_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_79_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_65_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7101_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_48_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6760_ _7076_/CLK _6760_/D wire3978/X VGND VGND VPWR VPWR _6760_/Q sky130_fd_sc_hd__dfrtp_1
X_3972_ hold713/X _4333_/A0 _3976_/S VGND VGND VPWR VPWR _6476_/D sky130_fd_sc_hd__mux2_1
XFILLER_62_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5711_ _5711_/A1 _5783_/B1 _5711_/B1 _5711_/B2 VGND VGND VPWR VPWR _5711_/X sky130_fd_sc_hd__a22o_1
X_6691_ _7206_/CLK _6691_/D _4189_/B VGND VGND VPWR VPWR _6691_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_148_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5642_ _6033_/A _6039_/A _6040_/B VGND VGND VPWR VPWR _5642_/X sky130_fd_sc_hd__and3_1
XFILLER_176_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5573_ _5573_/A0 hold103/X _5576_/S VGND VGND VPWR VPWR _7128_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold202 _7114_/Q VGND VGND VPWR VPWR hold202/X sky130_fd_sc_hd__dlygate4sd3_1
X_4524_ _4524_/A _4524_/B VGND VGND VPWR VPWR _4524_/Y sky130_fd_sc_hd__nand2_1
Xhold213 _6930_/Q VGND VGND VPWR VPWR hold213/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 _6705_/Q VGND VGND VPWR VPWR hold224/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_18_csclk _6579_/CLK VGND VGND VPWR VPWR _6963_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_144_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold235 _6965_/Q VGND VGND VPWR VPWR hold235/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 _6594_/Q VGND VGND VPWR VPWR hold246/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4455_ _4456_/A _4724_/B VGND VGND VPWR VPWR _4524_/B sky130_fd_sc_hd__nor2_2
Xhold257 _6637_/Q VGND VGND VPWR VPWR hold257/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold268 _6860_/Q VGND VGND VPWR VPWR hold268/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold279 _4299_/X VGND VGND VPWR VPWR _6745_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3406_ _3406_/A1 _3494_/B1 wire868/X _7109_/Q VGND VGND VPWR VPWR _3406_/X sky130_fd_sc_hd__a22o_1
X_7174_ _7180_/CLK _7174_/D wire3992/X VGND VGND VPWR VPWR _7174_/Q sky130_fd_sc_hd__dfrtp_1
X_4386_ _4451_/A _5035_/A VGND VGND VPWR VPWR _4759_/A sky130_fd_sc_hd__nor2_2
Xwire2509 _6151_/B1 VGND VGND VPWR VPWR _6073_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_131_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3337_ hold29/A _4120_/B VGND VGND VPWR VPWR _3337_/Y sky130_fd_sc_hd__nor2_1
X_6125_ _6125_/A1 _6125_/A2 _6175_/B1 _7123_/Q VGND VGND VPWR VPWR _6125_/X sky130_fd_sc_hd__a22o_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1808 wire1809/X VGND VGND VPWR VPWR _3653_/B2 sky130_fd_sc_hd__clkbuf_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1819 wire1820/X VGND VGND VPWR VPWR _6209_/B2 sky130_fd_sc_hd__clkbuf_2
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3268_ _5212_/A _3462_/A VGND VGND VPWR VPWR _3268_/Y sky130_fd_sc_hd__nor2_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ _6955_/Q _6056_/A2 _6056_/B1 _7059_/Q VGND VGND VPWR VPWR _6056_/X sky130_fd_sc_hd__a22o_1
XFILLER_105_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5007_ _5039_/A _5007_/B _5039_/B _5007_/D VGND VGND VPWR VPWR _5008_/D sky130_fd_sc_hd__or4_1
X_3199_ _3199_/A VGND VGND VPWR VPWR _3199_/Y sky130_fd_sc_hd__clkinv_2
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_108 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_119 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6958_ _7075_/CLK _6958_/D wire4041/X VGND VGND VPWR VPWR _6958_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5909_ _6613_/Q _5959_/B1 _5909_/B1 _6657_/Q VGND VGND VPWR VPWR _5909_/X sky130_fd_sc_hd__a22o_1
X_6889_ _7116_/CLK _6889_/D wire4071/A VGND VGND VPWR VPWR _6889_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_139_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3700 _3907_/A VGND VGND VPWR VPWR _5858_/C1 sky130_fd_sc_hd__clkbuf_2
XFILLER_122_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3711 _3190_/Y VGND VGND VPWR VPWR _3252_/B sky130_fd_sc_hd__clkbuf_2
Xwire3722 _7169_/Q VGND VGND VPWR VPWR _5860_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3733 wire3734/X VGND VGND VPWR VPWR wire3733/X sky130_fd_sc_hd__clkbuf_1
Xwire3744 wire3745/X VGND VGND VPWR VPWR wire3744/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3755 wire3756/X VGND VGND VPWR VPWR wire3755/X sky130_fd_sc_hd__clkbuf_1
Xwire3766 wire3767/X VGND VGND VPWR VPWR wire3766/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3777 wire3778/X VGND VGND VPWR VPWR wire3777/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3788 wire3789/X VGND VGND VPWR VPWR _3927_/S sky130_fd_sc_hd__clkbuf_1
XFILLER_131_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3799 _4589_/B VGND VGND VPWR VPWR _4675_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_64_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput307 _5592_/B VGND VGND VPWR VPWR serial_clock sky130_fd_sc_hd__buf_12
Xoutput318 _6647_/Q VGND VGND VPWR VPWR wb_dat_o[0] sky130_fd_sc_hd__buf_12
XFILLER_126_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput329 _6648_/Q VGND VGND VPWR VPWR wb_dat_o[1] sky130_fd_sc_hd__buf_12
XFILLER_126_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4240_ _4240_/A _4240_/B VGND VGND VPWR VPWR _4245_/S sky130_fd_sc_hd__and2_2
XFILLER_113_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4171_ _6631_/Q wire370/X _4173_/S VGND VGND VPWR VPWR _6631_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6812_ _6824_/CLK _6812_/D _6483_/SET_B VGND VGND VPWR VPWR _6812_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_63_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6743_ _6799_/CLK _6743_/D _6743_/SET_B VGND VGND VPWR VPWR _6743_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_149_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3955_ _6696_/Q _3962_/B VGND VGND VPWR VPWR _6694_/D sky130_fd_sc_hd__and2_1
XFILLER_189_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6674_ _6702_/CLK _6674_/D _6440_/A VGND VGND VPWR VPWR _6674_/Q sky130_fd_sc_hd__dfrtp_1
X_3886_ _4467_/A _4654_/B _3886_/C _3886_/D VGND VGND VPWR VPWR _3887_/D sky130_fd_sc_hd__or4_1
XFILLER_164_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5625_ _5624_/Y _5693_/A _5625_/S VGND VGND VPWR VPWR _7152_/D sky130_fd_sc_hd__mux2_1
XFILLER_137_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5556_ _5574_/A0 hold265/X _5557_/S VGND VGND VPWR VPWR _7113_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4507_ _4527_/A1 _4942_/A _4753_/B VGND VGND VPWR VPWR _4507_/X sky130_fd_sc_hd__a21o_1
XFILLER_132_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5487_ _5487_/A0 hold433/X _5487_/S VGND VGND VPWR VPWR _7052_/D sky130_fd_sc_hd__mux2_1
XFILLER_105_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3007 _5950_/A2 VGND VGND VPWR VPWR _5905_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3018 _5677_/X VGND VGND VPWR VPWR _5829_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_132_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4438_ _4443_/B _4456_/A VGND VGND VPWR VPWR _4448_/B sky130_fd_sc_hd__nor2_1
Xwire2306 _6634_/Q VGND VGND VPWR VPWR wire2306/X sky130_fd_sc_hd__clkbuf_1
Xwire2317 _6616_/Q VGND VGND VPWR VPWR _6221_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
X_7157_ _7187_/CLK _7157_/D wire3991/X VGND VGND VPWR VPWR _7157_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_98_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2328 _6609_/Q VGND VGND VPWR VPWR wire2328/X sky130_fd_sc_hd__clkbuf_1
X_4369_ _4596_/A _4369_/B VGND VGND VPWR VPWR _4369_/X sky130_fd_sc_hd__or2_1
Xwire2339 _6600_/Q VGND VGND VPWR VPWR _6342_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1605 _5760_/B2 VGND VGND VPWR VPWR _3599_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire1616 _3385_/A1 VGND VGND VPWR VPWR _6191_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6108_ _6108_/A1 _6150_/B1 _6151_/A2 _6108_/B2 _6107_/X VGND VGND VPWR VPWR _6109_/D
+ sky130_fd_sc_hd__a221o_1
Xwire1627 _7074_/Q VGND VGND VPWR VPWR _5995_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1638 _7066_/Q VGND VGND VPWR VPWR wire1638/X sky130_fd_sc_hd__clkbuf_1
XFILLER_74_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7088_ _7088_/CLK _7088_/D wire4069/X VGND VGND VPWR VPWR _7088_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_86_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1649 wire1650/X VGND VGND VPWR VPWR wire1649/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6039_ _6039_/A _6040_/B _6039_/C VGND VGND VPWR VPWR _6039_/X sky130_fd_sc_hd__and3_1
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire902 wire903/X VGND VGND VPWR VPWR wire902/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire913 wire914/X VGND VGND VPWR VPWR wire913/X sky130_fd_sc_hd__clkbuf_1
Xwire924 _3318_/Y VGND VGND VPWR VPWR wire924/X sky130_fd_sc_hd__clkbuf_2
Xwire935 wire936/X VGND VGND VPWR VPWR wire935/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire946 wire946/A VGND VGND VPWR VPWR wire946/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire957 wire958/X VGND VGND VPWR VPWR wire957/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire968 _4052_/B VGND VGND VPWR VPWR _5232_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_136_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire4220 wire4221/X VGND VGND VPWR VPWR _3549_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire4231 wire4232/X VGND VGND VPWR VPWR _3678_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire4242 wire4243/X VGND VGND VPWR VPWR _3494_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire4253 wire4254/X VGND VGND VPWR VPWR wire4253/X sky130_fd_sc_hd__clkbuf_1
Xwire4264 wire4264/A VGND VGND VPWR VPWR wire4264/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3530 wire3531/X VGND VGND VPWR VPWR wire3530/X sky130_fd_sc_hd__clkbuf_1
XFILLER_150_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire4275 wire4276/X VGND VGND VPWR VPWR wire4275/X sky130_fd_sc_hd__clkbuf_1
Xwire4286 _4605_/A VGND VGND VPWR VPWR _4588_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3552 _5538_/A1 VGND VGND VPWR VPWR _5514_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3563 wire3564/X VGND VGND VPWR VPWR _4092_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_104_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3574 _5565_/A0 VGND VGND VPWR VPWR _5442_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_173_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3585 _4200_/A1 VGND VGND VPWR VPWR _4248_/A0 sky130_fd_sc_hd__clkbuf_2
Xwire2851 _5786_/B1 VGND VGND VPWR VPWR _5746_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3596 _5333_/A0 VGND VGND VPWR VPWR _5495_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2862 _5808_/B1 VGND VGND VPWR VPWR _5741_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2873 _5849_/B1 VGND VGND VPWR VPWR _5778_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2884 wire2885/X VGND VGND VPWR VPWR _5856_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire2895 wire2896/X VGND VGND VPWR VPWR _5854_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_66_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_19 wire419/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3740_ _3740_/A1 wire929/X _4276_/A _6726_/Q VGND VGND VPWR VPWR _3740_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3671_ _3671_/A1 _3671_/A2 _3767_/B1 _3671_/B2 _3670_/X VGND VGND VPWR VPWR _3671_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5410_ _5410_/A0 hold703/X _5410_/S VGND VGND VPWR VPWR _6984_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_559 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6390_ _6390_/A1 _4228_/Y _6360_/X _6389_/X _6358_/A VGND VGND VPWR VPWR _6390_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_126_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5341_ _5359_/A0 hold342/X _5343_/S VGND VGND VPWR VPWR _6922_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5272_ _5308_/A0 hold547/X _5276_/S VGND VGND VPWR VPWR _6861_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7011_ _7135_/CLK _7011_/D _7051_/SET_B VGND VGND VPWR VPWR _7011_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_141_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4223_ _4223_/A0 hold459/X _4227_/S VGND VGND VPWR VPWR _6675_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4154_ _4259_/A1 hold462/X hold58/X VGND VGND VPWR VPWR _6616_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4085_ hold419/X _5552_/A0 _4085_/S VGND VGND VPWR VPWR _4085_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4987_ _4987_/A _4987_/B _4987_/C VGND VGND VPWR VPWR _4988_/D sky130_fd_sc_hd__or3_1
X_6726_ _7104_/CLK _6726_/D wire4040/X VGND VGND VPWR VPWR _6726_/Q sky130_fd_sc_hd__dfrtp_1
X_3938_ _3938_/A0 _3938_/A1 _6823_/Q VGND VGND VPWR VPWR _3938_/X sky130_fd_sc_hd__mux2_1
Xmax_length3516 _5479_/A0 VGND VGND VPWR VPWR _5584_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_177_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6657_ _6683_/CLK _6657_/D wire3965/A VGND VGND VPWR VPWR _6657_/Q sky130_fd_sc_hd__dfstp_1
X_3869_ _3184_/Y _3951_/A1 _3868_/B _3868_/Y VGND VGND VPWR VPWR _6445_/D sky130_fd_sc_hd__a31o_1
XFILLER_176_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5608_ _7147_/Q _5605_/A _5607_/Y VGND VGND VPWR VPWR _7147_/D sky130_fd_sc_hd__o21a_1
X_6588_ _6811_/CLK _6588_/D _3946_/B VGND VGND VPWR VPWR _6588_/Q sky130_fd_sc_hd__dfrtp_1
Xmax_length2859 _5958_/A2 VGND VGND VPWR VPWR _5889_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_192_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5539_ hold568/X _5539_/A1 _5542_/S VGND VGND VPWR VPWR _7098_/D sky130_fd_sc_hd__mux2_1
XFILLER_105_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7209_ _7210_/CLK _7209_/D fanout3952/X VGND VGND VPWR VPWR _7209_/Q sky130_fd_sc_hd__dfstp_1
Xwire2103 _6822_/Q VGND VGND VPWR VPWR _5227_/A0 sky130_fd_sc_hd__clkbuf_1
Xwire2114 _6815_/Q VGND VGND VPWR VPWR wire2114/X sky130_fd_sc_hd__clkbuf_1
Xwire2125 wire2126/X VGND VGND VPWR VPWR wire2125/X sky130_fd_sc_hd__clkbuf_1
XFILLER_59_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2136 wire2137/X VGND VGND VPWR VPWR _3442_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_59_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2147 _6775_/Q VGND VGND VPWR VPWR wire2147/X sky130_fd_sc_hd__clkbuf_1
Xwire1402 _3255_/X VGND VGND VPWR VPWR _3472_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_143_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2158 _6760_/Q VGND VGND VPWR VPWR _6339_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire1413 _6190_/X VGND VGND VPWR VPWR wire1413/X sky130_fd_sc_hd__clkbuf_1
Xwire2169 _3549_/B2 VGND VGND VPWR VPWR wire2169/X sky130_fd_sc_hd__clkbuf_1
Xwire1424 wire1425/X VGND VGND VPWR VPWR wire1424/X sky130_fd_sc_hd__clkbuf_1
Xwire1435 _4468_/X VGND VGND VPWR VPWR _4940_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1457 _3933_/X VGND VGND VPWR VPWR wire1457/X sky130_fd_sc_hd__clkbuf_1
XFILLER_46_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1468 wire1469/X VGND VGND VPWR VPWR wire1468/X sky130_fd_sc_hd__clkbuf_1
Xwire1479 _3924_/X VGND VGND VPWR VPWR wire1479/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire710 hold8/X VGND VGND VPWR VPWR _5249_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_52_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire721 _4128_/S VGND VGND VPWR VPWR _4125_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_168_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput17 mask_rev_in[21] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__clkbuf_1
Xwire732 wire733/X VGND VGND VPWR VPWR wire732/X sky130_fd_sc_hd__clkbuf_1
XFILLER_168_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire743 _3777_/X VGND VGND VPWR VPWR wire743/X sky130_fd_sc_hd__clkbuf_1
Xinput28 mask_rev_in[31] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__clkbuf_1
Xwire754 _3715_/X VGND VGND VPWR VPWR wire754/X sky130_fd_sc_hd__clkbuf_1
Xinput39 mgmt_gpio_in[12] VGND VGND VPWR VPWR input39/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire765 wire766/X VGND VGND VPWR VPWR wire765/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire776 wire777/X VGND VGND VPWR VPWR wire776/X sky130_fd_sc_hd__clkbuf_1
Xwire787 wire788/X VGND VGND VPWR VPWR wire787/X sky130_fd_sc_hd__clkbuf_1
Xwire798 _3531_/Y VGND VGND VPWR VPWR wire798/X sky130_fd_sc_hd__clkbuf_1
XFILLER_108_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire4061 wire4061/A VGND VGND VPWR VPWR wire4061/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire4083 wire4086/X VGND VGND VPWR VPWR wire4083/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire4094 wire4095/X VGND VGND VPWR VPWR wire4094/X sky130_fd_sc_hd__clkbuf_2
Xwire3360 _4495_/B VGND VGND VPWR VPWR _4993_/A sky130_fd_sc_hd__clkbuf_2
Xwire3382 _5456_/A0 VGND VGND VPWR VPWR _5552_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2670 _6225_/B1 VGND VGND VPWR VPWR _6327_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2681 _6022_/D VGND VGND VPWR VPWR _6299_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2692 _6159_/B1 VGND VGND VPWR VPWR _6082_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_92_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1980 _6907_/Q VGND VGND VPWR VPWR _5721_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire1991 _3740_/A1 VGND VGND VPWR VPWR _5990_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4910_ _4545_/X _4646_/A _4910_/B1 VGND VGND VPWR VPWR _4910_/X sky130_fd_sc_hd__a21o_1
XFILLER_45_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5890_ _5890_/A1 _5890_/A2 _5890_/B1 _6249_/A1 _5889_/X VGND VGND VPWR VPWR _5891_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_178_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4841_ _4940_/B _4677_/B _4520_/X VGND VGND VPWR VPWR _5162_/B sky130_fd_sc_hd__o21ai_2
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4772_ _4657_/C _5133_/A2 _4770_/X _4771_/X VGND VGND VPWR VPWR _4772_/X sky130_fd_sc_hd__a211o_1
XFILLER_21_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6511_ _7210_/CLK _6511_/D wire3935/X VGND VGND VPWR VPWR _6511_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_186_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3723_ _3723_/A _3723_/B _3723_/C VGND VGND VPWR VPWR _3723_/X sky130_fd_sc_hd__or3_1
XFILLER_186_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6442_ _6545_/CLK _6442_/D _6398_/X VGND VGND VPWR VPWR hold5/A sky130_fd_sc_hd__dfrtn_1
X_3654_ _5748_/B2 _3654_/A2 _3654_/B1 _3654_/B2 _3605_/X VGND VGND VPWR VPWR _3659_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6373_ _4228_/C _6373_/A2 _6373_/B1 _4228_/Y _6372_/X VGND VGND VPWR VPWR _6373_/X
+ sky130_fd_sc_hd__a221o_1
Xclkbuf_3_0_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A VGND VGND VPWR VPWR _7185_/CLK sky130_fd_sc_hd__clkbuf_8
X_3585_ _3585_/A1 _3585_/A2 _3547_/Y _3585_/B2 wire785/X VGND VGND VPWR VPWR _3588_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5324_ hold151/X _5522_/A0 _5325_/S VGND VGND VPWR VPWR _6907_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5255_ hold681/X _5255_/A1 _5255_/S VGND VGND VPWR VPWR _6846_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4206_ _4206_/A0 _4206_/A1 _4209_/S VGND VGND VPWR VPWR _6661_/D sky130_fd_sc_hd__mux2_1
X_5186_ _5195_/A0 hold431/X _5186_/S VGND VGND VPWR VPWR _6792_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4137_ hold478/X _4248_/A0 _4140_/S VGND VGND VPWR VPWR _6602_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4068_ _6587_/Q hold3/X _4068_/S VGND VGND VPWR VPWR _4068_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length4003 wire4004/X VGND VGND VPWR VPWR _7110_/RESET_B sky130_fd_sc_hd__clkbuf_2
Xmax_length4025 wire4026/X VGND VGND VPWR VPWR _7112_/SET_B sky130_fd_sc_hd__buf_2
XFILLER_184_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length4036 _6401_/A VGND VGND VPWR VPWR _7042_/SET_B sky130_fd_sc_hd__buf_2
Xmax_length3302 _4639_/B VGND VGND VPWR VPWR _4624_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6709_ _7091_/CLK _6709_/D wire4029/A VGND VGND VPWR VPWR _6709_/Q sky130_fd_sc_hd__dfrtp_1
Xmax_length3324 _4784_/A VGND VGND VPWR VPWR _4680_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_177_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length2656 _6205_/B1 VGND VGND VPWR VPWR wire2650/A sky130_fd_sc_hd__clkbuf_1
XFILLER_106_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1210 _3719_/A2 VGND VGND VPWR VPWR wire1210/X sky130_fd_sc_hd__clkbuf_1
XFILLER_47_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1232 _3304_/Y VGND VGND VPWR VPWR _3641_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1243 _3300_/Y VGND VGND VPWR VPWR _3762_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire1254 wire1255/X VGND VGND VPWR VPWR _3779_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_101_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1265 wire1265/A VGND VGND VPWR VPWR _3500_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_74_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1276 _3292_/Y VGND VGND VPWR VPWR _3693_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_74_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1287 _4001_/A VGND VGND VPWR VPWR _3383_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1298 hold29/X VGND VGND VPWR VPWR _3490_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire540 _3737_/X VGND VGND VPWR VPWR wire540/X sky130_fd_sc_hd__clkbuf_1
Xwire551 _3671_/X VGND VGND VPWR VPWR wire551/X sky130_fd_sc_hd__clkbuf_1
Xwire562 _3532_/X VGND VGND VPWR VPWR wire562/X sky130_fd_sc_hd__clkbuf_1
Xwire573 _3394_/X VGND VGND VPWR VPWR wire573/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold609 _6592_/Q VGND VGND VPWR VPWR hold609/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire584 wire585/X VGND VGND VPWR VPWR wire584/X sky130_fd_sc_hd__clkbuf_1
XFILLER_156_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire595 _5528_/S VGND VGND VPWR VPWR _5525_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3370_ _6206_/A1 _5394_/A wire910/X _6199_/B2 _3369_/X VGND VGND VPWR VPWR _3371_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5040_ _5133_/A1 _5133_/A2 _5130_/A VGND VGND VPWR VPWR _5040_/X sky130_fd_sc_hd__a21o_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6991_ _7110_/CLK _6991_/D _7110_/RESET_B VGND VGND VPWR VPWR _6991_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5942_ _6689_/Q _5962_/A2 _5963_/B1 _6299_/A1 _5941_/X VGND VGND VPWR VPWR _5945_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5873_ _6234_/B2 _5928_/A2 _5917_/B1 _5872_/X VGND VGND VPWR VPWR _5873_/X sky130_fd_sc_hd__a22o_1
XFILLER_178_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4824_ _4824_/A _4992_/B VGND VGND VPWR VPWR _4824_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4755_ _4759_/A _4758_/A _5001_/A _4758_/B _4495_/B VGND VGND VPWR VPWR _4755_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_119_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3706_ _3706_/A1 _3776_/A2 _3706_/B1 _6512_/Q VGND VGND VPWR VPWR _3706_/X sky130_fd_sc_hd__a22o_1
X_4686_ _4687_/B _4686_/B VGND VGND VPWR VPWR _4686_/X sky130_fd_sc_hd__or2_1
Xmax_length1207 _3316_/Y VGND VGND VPWR VPWR wire1206/A sky130_fd_sc_hd__clkbuf_1
X_6425_ _6437_/A _6437_/B VGND VGND VPWR VPWR _6425_/X sky130_fd_sc_hd__and2_1
X_3637_ input5/X _3777_/A2 _3992_/A _6492_/Q _3636_/X VGND VGND VPWR VPWR _3637_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6356_ _7196_/Q wire378/X _6356_/S VGND VGND VPWR VPWR _7196_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3568_ _3568_/A1 _3568_/A2 wire795/X _3568_/B2 wire776/X VGND VGND VPWR VPWR _3573_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5307_ _5343_/A0 hold312/X _5307_/S VGND VGND VPWR VPWR _6892_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6287_ _7092_/Q _6298_/A2 _6298_/B1 _6287_/B2 VGND VGND VPWR VPWR _6287_/X sky130_fd_sc_hd__a22o_1
X_3499_ _3499_/A _3499_/B _3499_/C _3499_/D VGND VGND VPWR VPWR _3542_/A sky130_fd_sc_hd__or4_2
XFILLER_102_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5238_ _5550_/A0 hold233/X _5240_/S VGND VGND VPWR VPWR _6831_/D sky130_fd_sc_hd__mux2_1
XFILLER_76_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5169_ _5169_/A1 _4623_/A _4728_/Y _4743_/B _4626_/Y VGND VGND VPWR VPWR _5169_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_84_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length3176 _4638_/X VGND VGND VPWR VPWR _4689_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_125_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3198 _4734_/B VGND VGND VPWR VPWR _4816_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_180_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length2475 _6182_/B1 VGND VGND VPWR VPWR wire2474/A sky130_fd_sc_hd__clkbuf_1
XFILLER_152_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length1752 _7022_/Q VGND VGND VPWR VPWR wire1751/A sky130_fd_sc_hd__clkbuf_1
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold6 hold6/A VGND VGND VPWR VPWR hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1040 _3512_/Y VGND VGND VPWR VPWR _3770_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire1051 _3507_/Y VGND VGND VPWR VPWR _3784_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1062 _3776_/B1 VGND VGND VPWR VPWR wire1062/X sky130_fd_sc_hd__clkbuf_1
XFILLER_47_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1095 _3585_/A2 VGND VGND VPWR VPWR wire1095/X sky130_fd_sc_hd__clkbuf_1
XFILLER_75_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4540_ _4553_/A _4819_/C _4819_/D VGND VGND VPWR VPWR _4792_/A sky130_fd_sc_hd__and3_1
XFILLER_156_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire370 wire371/X VGND VGND VPWR VPWR wire370/X sky130_fd_sc_hd__dlymetal6s2s_1
Xwire381 _3373_/X VGND VGND VPWR VPWR wire381/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4471_ _4495_/A _4471_/B VGND VGND VPWR VPWR _4475_/A sky130_fd_sc_hd__nor2_1
Xhold406 _6669_/Q VGND VGND VPWR VPWR hold406/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire392 wire393/X VGND VGND VPWR VPWR _3790_/D sky130_fd_sc_hd__clkbuf_1
Xhold417 _6546_/Q VGND VGND VPWR VPWR hold417/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold428 _6604_/Q VGND VGND VPWR VPWR hold428/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold439 _6533_/Q VGND VGND VPWR VPWR hold439/X sky130_fd_sc_hd__dlygate4sd3_1
X_6210_ _6921_/Q _6210_/A2 _6210_/B1 _6210_/B2 VGND VGND VPWR VPWR _6210_/X sky130_fd_sc_hd__a22o_1
X_3422_ input31/X _3763_/A2 _3983_/A _6487_/Q VGND VGND VPWR VPWR _3422_/X sky130_fd_sc_hd__a22o_1
XFILLER_99_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7190_ _7196_/CLK _7190_/D VGND VGND VPWR VPWR _7190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6141_ _6141_/A1 _6141_/A2 _6141_/B1 _6141_/B2 _6140_/X VGND VGND VPWR VPWR _6142_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _7073_/Q _3550_/A2 wire892/X _6198_/B2 VGND VGND VPWR VPWR _3353_/X sky130_fd_sc_hd__a22o_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ _7176_/Q _6071_/X _6122_/S VGND VGND VPWR VPWR _7176_/D sky130_fd_sc_hd__mux2_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ _3284_/A hold83/X VGND VGND VPWR VPWR hold84/A sky130_fd_sc_hd__nor2_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5023_ _5023_/A _5023_/B _5023_/C VGND VGND VPWR VPWR _5027_/B sky130_fd_sc_hd__and3_2
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6974_ _7121_/CLK _6974_/D fanout4047/A VGND VGND VPWR VPWR _6974_/Q sky130_fd_sc_hd__dfrtp_1
X_5925_ _5969_/A1 _7171_/Q wire460/X VGND VGND VPWR VPWR _5925_/X sky130_fd_sc_hd__a21o_1
XFILLER_41_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5856_ _6921_/Q _5856_/A2 _5856_/B1 _7057_/Q _5855_/X VGND VGND VPWR VPWR _5857_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_166_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4807_ _4794_/A _4562_/X _4610_/X _5094_/B _4807_/B2 VGND VGND VPWR VPWR _4809_/B
+ sky130_fd_sc_hd__o32a_1
X_5787_ _5787_/A1 _5787_/A2 _5775_/X _5786_/X VGND VGND VPWR VPWR _5792_/A sky130_fd_sc_hd__a211o_1
XFILLER_119_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4738_ _4738_/A _4739_/B VGND VGND VPWR VPWR _5042_/A sky130_fd_sc_hd__nor2_1
XFILLER_119_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4669_ _4663_/Y _4666_/Y _4667_/X _4665_/Y _4669_/B2 VGND VGND VPWR VPWR _4669_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_107_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length1048 _4324_/A VGND VGND VPWR VPWR _3767_/A2 sky130_fd_sc_hd__clkbuf_2
X_6408_ _6441_/A _6431_/B VGND VGND VPWR VPWR _6408_/X sky130_fd_sc_hd__and2_1
XFILLER_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3904 wire3905/X VGND VGND VPWR VPWR wire3904/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3915 wire3916/X VGND VGND VPWR VPWR wire3915/X sky130_fd_sc_hd__clkbuf_1
Xwire3926 input78/X VGND VGND VPWR VPWR _3924_/A1 sky130_fd_sc_hd__clkbuf_1
X_6339_ _6339_/A1 _6339_/A2 _6339_/B1 _6339_/B2 _6338_/X VGND VGND VPWR VPWR _6339_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3948 wire3948/A VGND VGND VPWR VPWR wire3948/X sky130_fd_sc_hd__buf_2
Xwire3959 wire3959/A VGND VGND VPWR VPWR wire3959/X sky130_fd_sc_hd__buf_2
XFILLER_103_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2261 _6679_/Q VGND VGND VPWR VPWR wire2259/A sky130_fd_sc_hd__clkbuf_1
XFILLER_125_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length2294 hold415/X VGND VGND VPWR VPWR _4199_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_180_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length1582 _7099_/Q VGND VGND VPWR VPWR wire1581/A sky130_fd_sc_hd__clkbuf_1
XFILLER_192_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3971_ hold20/X hold77/X _3981_/S VGND VGND VPWR VPWR hold21/A sky130_fd_sc_hd__mux2_1
XFILLER_63_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5710_ _7162_/Q _5652_/Y _5709_/X VGND VGND VPWR VPWR _7162_/D sky130_fd_sc_hd__a21o_1
XFILLER_188_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6690_ _7093_/CLK _6690_/D wire3959/X VGND VGND VPWR VPWR _6690_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5641_ _7158_/Q _7157_/Q VGND VGND VPWR VPWR _6038_/A sky130_fd_sc_hd__nand2b_1
XFILLER_188_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5572_ _5572_/A0 hold205/X _5576_/S VGND VGND VPWR VPWR _7127_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_1_csclk clkbuf_1_0_1_csclk/A VGND VGND VPWR VPWR clkbuf_2_1_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_117_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4523_ _4997_/A _4526_/B VGND VGND VPWR VPWR _5049_/A sky130_fd_sc_hd__nor2_1
XFILLER_144_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold203 _6925_/Q VGND VGND VPWR VPWR hold203/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold214 _6880_/Q VGND VGND VPWR VPWR hold214/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 _6703_/Q VGND VGND VPWR VPWR hold225/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4454_ _5002_/A VGND VGND VPWR VPWR _4454_/Y sky130_fd_sc_hd__clkinv_2
Xhold236 _6750_/Q VGND VGND VPWR VPWR hold236/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 _6609_/Q VGND VGND VPWR VPWR hold247/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 _6634_/Q VGND VGND VPWR VPWR hold258/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 _6963_/Q VGND VGND VPWR VPWR hold269/X sky130_fd_sc_hd__dlygate4sd3_1
X_3405_ _6183_/A1 wire898/X wire885/X input69/X _3384_/X VGND VGND VPWR VPWR _3408_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_171_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7173_ _7185_/CLK _7173_/D wire3950/X VGND VGND VPWR VPWR _7173_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4385_ _4495_/A _4385_/B VGND VGND VPWR VPWR _5035_/A sky130_fd_sc_hd__or2_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6124_ _6124_/A1 _6124_/A2 _6166_/A2 _6870_/Q VGND VGND VPWR VPWR _6124_/X sky130_fd_sc_hd__a22o_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3336_ _3518_/B hold85/X VGND VGND VPWR VPWR _3336_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1809 _7004_/Q VGND VGND VPWR VPWR wire1809/X sky130_fd_sc_hd__clkbuf_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__1134_ _3543_/X VGND VGND VPWR VPWR clkbuf_0__1134_/X sky130_fd_sc_hd__clkbuf_16
X_6055_ _6055_/A1 _6074_/A2 _6055_/B1 _7104_/Q _6054_/X VGND VGND VPWR VPWR _6058_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_39_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ _3303_/A _3416_/A VGND VGND VPWR VPWR _3267_/Y sky130_fd_sc_hd__nand2_1
XFILLER_100_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5006_ _4418_/B _4485_/A _4744_/X _4993_/B _4495_/B VGND VGND VPWR VPWR _5007_/D
+ sky130_fd_sc_hd__o32a_1
X_3198_ _3198_/A VGND VGND VPWR VPWR _3198_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_54_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_109 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6957_ _7031_/CLK _6957_/D wire4048/X VGND VGND VPWR VPWR _6957_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_54_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5908_ _5908_/A1 _5963_/B1 _5934_/A2 _5908_/B2 _5907_/X VGND VGND VPWR VPWR _5913_/B
+ sky130_fd_sc_hd__a221o_1
X_6888_ _7116_/CLK _6888_/D wire4071/A VGND VGND VPWR VPWR _6888_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5839_ _7073_/Q _5839_/A2 _5839_/B1 _6201_/B2 VGND VGND VPWR VPWR _5839_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length704 _5331_/Y VGND VGND VPWR VPWR wire703/A sky130_fd_sc_hd__clkbuf_1
XFILLER_167_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3701 _6095_/C1 VGND VGND VPWR VPWR _5729_/C1 sky130_fd_sc_hd__clkbuf_1
Xwire3712 wire3713/X VGND VGND VPWR VPWR wire3712/X sky130_fd_sc_hd__clkbuf_2
XFILLER_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3723 wire3724/X VGND VGND VPWR VPWR _3776_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_89_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3734 _6778_/Q VGND VGND VPWR VPWR wire3734/X sky130_fd_sc_hd__clkbuf_1
Xwire3745 _6700_/Q VGND VGND VPWR VPWR wire3745/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3756 wire3757/X VGND VGND VPWR VPWR wire3756/X sky130_fd_sc_hd__clkbuf_1
Xwire3767 _6680_/Q VGND VGND VPWR VPWR wire3767/X sky130_fd_sc_hd__clkbuf_1
X_3234__1 _6545_/CLK VGND VGND VPWR VPWR _6443_/CLK sky130_fd_sc_hd__inv_2
Xwire3778 _6563_/Q VGND VGND VPWR VPWR wire3778/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3789 wire3790/X VGND VGND VPWR VPWR wire3789/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput308 _3413_/X VGND VGND VPWR VPWR serial_data_1 sky130_fd_sc_hd__buf_12
Xoutput319 _6641_/Q VGND VGND VPWR VPWR wb_dat_o[10] sky130_fd_sc_hd__buf_12
XFILLER_114_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4170_ _6630_/Q _6353_/A1 _4170_/S VGND VGND VPWR VPWR _6630_/D sky130_fd_sc_hd__mux2_1
XFILLER_36_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6811_ _6811_/CLK _6811_/D _3946_/B VGND VGND VPWR VPWR _6811_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_51_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6742_ _6799_/CLK _6742_/D fanout3952/X VGND VGND VPWR VPWR _6742_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_51_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3954_ _6698_/Q _3962_/B VGND VGND VPWR VPWR _6695_/D sky130_fd_sc_hd__and2_1
XFILLER_50_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6673_ _6702_/CLK _6673_/D wire3961/X VGND VGND VPWR VPWR _6673_/Q sky130_fd_sc_hd__dfrtp_1
X_3885_ _3885_/A _3885_/B input120/X input117/X VGND VGND VPWR VPWR _3886_/D sky130_fd_sc_hd__or4bb_1
XFILLER_176_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5624_ _5693_/A _5624_/B VGND VGND VPWR VPWR _5624_/Y sky130_fd_sc_hd__nand2_1
XFILLER_176_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5555_ _5555_/A0 hold481/X _5555_/S VGND VGND VPWR VPWR _7112_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4506_ _4996_/A _4506_/B VGND VGND VPWR VPWR _4506_/Y sky130_fd_sc_hd__nor2_2
XFILLER_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5486_ _5573_/A0 hold181/X _5487_/S VGND VGND VPWR VPWR _7051_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3008 _5865_/A2 VGND VGND VPWR VPWR _5950_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4437_ _4758_/A _4744_/C VGND VGND VPWR VPWR _4456_/A sky130_fd_sc_hd__nand2_1
Xwire3019 _5952_/A2 VGND VGND VPWR VPWR _5883_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_132_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7156_ _7187_/CLK _7156_/D wire4014/X VGND VGND VPWR VPWR _7156_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2318 _6615_/Q VGND VGND VPWR VPWR _5959_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
X_4368_ _4596_/A _4369_/B VGND VGND VPWR VPWR _4397_/A sky130_fd_sc_hd__nor2_1
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1606 _6112_/A1 VGND VGND VPWR VPWR _5760_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_112_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6107_ _7077_/Q _6150_/A2 _6152_/A2 _6107_/B2 VGND VGND VPWR VPWR _6107_/X sky130_fd_sc_hd__a22o_1
Xwire1617 _7080_/Q VGND VGND VPWR VPWR _3385_/A1 sky130_fd_sc_hd__clkbuf_1
X_3319_ _3466_/A hold85/A VGND VGND VPWR VPWR _3319_/Y sky130_fd_sc_hd__nor2_1
X_7087_ _7089_/CLK _7087_/D _7087_/RESET_B VGND VGND VPWR VPWR _7087_/Q sky130_fd_sc_hd__dfrtp_1
Xwire1628 _3438_/B2 VGND VGND VPWR VPWR _6148_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_100_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4299_ _5198_/A0 hold278/X _4299_/S VGND VGND VPWR VPWR _4299_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1639 _7065_/Q VGND VGND VPWR VPWR _6205_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6038_ _6038_/A _6038_/B VGND VGND VPWR VPWR _6038_/Y sky130_fd_sc_hd__nor2_1
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire903 wire904/A VGND VGND VPWR VPWR wire903/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire914 wire915/X VGND VGND VPWR VPWR wire914/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_64_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7001_/CLK sky130_fd_sc_hd__clkbuf_16
Xwire936 wire937/X VGND VGND VPWR VPWR wire936/X sky130_fd_sc_hd__clkbuf_1
XFILLER_127_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire947 wire948/X VGND VGND VPWR VPWR _5580_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_155_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire958 _3280_/Y VGND VGND VPWR VPWR wire958/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire969 wire970/X VGND VGND VPWR VPWR _4052_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_41_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire4210 wire4211/X VGND VGND VPWR VPWR wire4210/X sky130_fd_sc_hd__clkbuf_1
Xwire4221 wire4222/X VGND VGND VPWR VPWR wire4221/X sky130_fd_sc_hd__clkbuf_1
Xwire4232 wire4233/X VGND VGND VPWR VPWR wire4232/X sky130_fd_sc_hd__clkbuf_1
XFILLER_150_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_79_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6825_/CLK sky130_fd_sc_hd__clkbuf_16
Xwire4243 wire4244/X VGND VGND VPWR VPWR wire4243/X sky130_fd_sc_hd__clkbuf_1
Xfanout3458 wire3484/X VGND VGND VPWR VPWR wire3466/A sky130_fd_sc_hd__clkbuf_1
Xwire4254 wire4255/X VGND VGND VPWR VPWR wire4254/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire4265 wire4266/X VGND VGND VPWR VPWR wire4265/X sky130_fd_sc_hd__clkbuf_1
Xwire3520 _5380_/A0 VGND VGND VPWR VPWR _5353_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire4276 input15/X VGND VGND VPWR VPWR wire4276/X sky130_fd_sc_hd__clkbuf_1
Xwire3531 wire3532/X VGND VGND VPWR VPWR wire3531/X sky130_fd_sc_hd__clkbuf_1
XFILLER_173_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3553 _5505_/A0 VGND VGND VPWR VPWR _5538_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4298 _4398_/C VGND VGND VPWR VPWR _4562_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3564 _5406_/A0 VGND VGND VPWR VPWR wire3564/X sky130_fd_sc_hd__clkbuf_1
Xwire2830 _5755_/B1 VGND VGND VPWR VPWR _5711_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire3575 wire3575/A VGND VGND VPWR VPWR _5565_/A0 sky130_fd_sc_hd__clkbuf_1
Xwire3586 _4314_/A1 VGND VGND VPWR VPWR _4284_/A0 sky130_fd_sc_hd__clkbuf_1
Xwire2841 _5705_/X VGND VGND VPWR VPWR _5707_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2852 _5754_/B1 VGND VGND VPWR VPWR _5786_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2863 wire2864/X VGND VGND VPWR VPWR _5808_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_65_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2874 _5800_/B1 VGND VGND VPWR VPWR _5764_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire2885 _5699_/X VGND VGND VPWR VPWR wire2885/X sky130_fd_sc_hd__clkbuf_1
Xwire2896 _5697_/X VGND VGND VPWR VPWR wire2896/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3670_ _3670_/A1 _3496_/Y _3774_/B1 _6757_/Q VGND VGND VPWR VPWR _3670_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5340_ _5340_/A _5571_/B VGND VGND VPWR VPWR _5348_/S sky130_fd_sc_hd__nand2_2
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5271_ _5574_/A0 hold268/X _5273_/S VGND VGND VPWR VPWR _6860_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7010_ _7046_/CLK _7010_/D wire4052/A VGND VGND VPWR VPWR _7010_/Q sky130_fd_sc_hd__dfstp_1
X_4222_ _4222_/A _4222_/B VGND VGND VPWR VPWR _4227_/S sky130_fd_sc_hd__nand2_2
XFILLER_102_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4153_ _4153_/A _4222_/B VGND VGND VPWR VPWR hold58/A sky130_fd_sc_hd__nand2_2
XFILLER_56_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4084_ hold493/X _4083_/X _4084_/S VGND VGND VPWR VPWR _6560_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4986_ _4986_/A _4986_/B _4799_/X VGND VGND VPWR VPWR _5170_/A sky130_fd_sc_hd__or3b_1
XFILLER_23_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6725_ _6979_/CLK _6725_/D fanout4027/X VGND VGND VPWR VPWR _6725_/Q sky130_fd_sc_hd__dfrtp_1
X_3937_ _6572_/Q _3937_/A1 _3937_/S VGND VGND VPWR VPWR _3937_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6656_ _6683_/CLK _6656_/D _6672_/SET_B VGND VGND VPWR VPWR _6656_/Q sky130_fd_sc_hd__dfrtp_1
X_3868_ _3868_/A _3868_/B VGND VGND VPWR VPWR _3868_/Y sky130_fd_sc_hd__nor2_1
XFILLER_109_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5607_ _7147_/Q _5605_/A _5606_/A VGND VGND VPWR VPWR _5607_/Y sky130_fd_sc_hd__a21boi_1
X_6587_ _7130_/CLK hold4/X wire4058/X VGND VGND VPWR VPWR _6587_/Q sky130_fd_sc_hd__dfrtp_1
X_3799_ _6471_/Q _3801_/B _6472_/Q VGND VGND VPWR VPWR _3800_/B sky130_fd_sc_hd__a21oi_1
XFILLER_152_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5538_ hold410/X _5538_/A1 _5538_/S VGND VGND VPWR VPWR _7097_/D sky130_fd_sc_hd__mux2_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5469_ hold666/X _5469_/A1 _5469_/S VGND VGND VPWR VPWR _7036_/D sky130_fd_sc_hd__mux2_1
XFILLER_105_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7208_ _7208_/CLK _7208_/D wire4026/X VGND VGND VPWR VPWR _7208_/Q sky130_fd_sc_hd__dfrtp_1
Xwire2104 _6821_/Q VGND VGND VPWR VPWR _3937_/S sky130_fd_sc_hd__clkbuf_1
Xwire2115 hold521/X VGND VGND VPWR VPWR _5216_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_120_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2126 _6809_/Q VGND VGND VPWR VPWR wire2126/X sky130_fd_sc_hd__clkbuf_1
Xwire2137 wire2138/X VGND VGND VPWR VPWR wire2137/X sky130_fd_sc_hd__clkbuf_1
Xwire2148 wire2148/A VGND VGND VPWR VPWR _3599_/B2 sky130_fd_sc_hd__clkbuf_1
X_7139_ _7139_/CLK _7139_/D wire4065/X VGND VGND VPWR VPWR _7139_/Q sky130_fd_sc_hd__dfrtp_1
Xwire2159 wire2160/X VGND VGND VPWR VPWR _6322_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire1414 _6131_/X VGND VGND VPWR VPWR _6132_/C1 sky130_fd_sc_hd__clkbuf_1
Xwire1425 wire1426/X VGND VGND VPWR VPWR wire1425/X sky130_fd_sc_hd__clkbuf_1
Xwire1458 wire1459/X VGND VGND VPWR VPWR wire1458/X sky130_fd_sc_hd__clkbuf_2
XFILLER_101_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1469 wire1470/X VGND VGND VPWR VPWR wire1469/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire700 _5331_/Y VGND VGND VPWR VPWR _5334_/S sky130_fd_sc_hd__clkbuf_1
Xwire711 _5059_/Y VGND VGND VPWR VPWR _5159_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire722 wire723/X VGND VGND VPWR VPWR _4128_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_128_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput18 mask_rev_in[22] VGND VGND VPWR VPWR input18/X sky130_fd_sc_hd__clkbuf_1
Xwire733 wire734/X VGND VGND VPWR VPWR wire733/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire744 _3768_/X VGND VGND VPWR VPWR wire744/X sky130_fd_sc_hd__clkbuf_1
Xinput29 mask_rev_in[3] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__clkbuf_1
Xwire755 wire756/X VGND VGND VPWR VPWR wire755/X sky130_fd_sc_hd__clkbuf_1
XFILLER_182_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire766 _3682_/X VGND VGND VPWR VPWR wire766/X sky130_fd_sc_hd__clkbuf_1
Xwire777 wire778/X VGND VGND VPWR VPWR wire777/X sky130_fd_sc_hd__clkbuf_1
Xwire788 wire789/X VGND VGND VPWR VPWR wire788/X sky130_fd_sc_hd__clkbuf_1
XFILLER_170_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire799 wire802/X VGND VGND VPWR VPWR wire799/X sky130_fd_sc_hd__clkbuf_1
XFILLER_182_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire4040 wire4042/A VGND VGND VPWR VPWR wire4040/X sky130_fd_sc_hd__buf_2
XFILLER_151_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4095 wire4096/X VGND VGND VPWR VPWR wire4095/X sky130_fd_sc_hd__clkbuf_1
Xwire3361 _4778_/A VGND VGND VPWR VPWR _4495_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3372 _5501_/A0 VGND VGND VPWR VPWR _5588_/A0 sky130_fd_sc_hd__clkbuf_2
Xwire3383 _5543_/A1 VGND VGND VPWR VPWR _5456_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3394 _5491_/A0 VGND VGND VPWR VPWR _5518_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2660 _6282_/B1 VGND VGND VPWR VPWR _6321_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2671 wire2672/X VGND VGND VPWR VPWR _6225_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire2682 _6017_/X VGND VGND VPWR VPWR _6022_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2693 _6172_/B1 VGND VGND VPWR VPWR _6159_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1970 _6910_/Q VGND VGND VPWR VPWR _5779_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1981 _6906_/Q VGND VGND VPWR VPWR _6031_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_18_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1992 _6898_/Q VGND VGND VPWR VPWR _3740_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_80_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4840_ _4940_/B _4659_/B _4447_/Y VGND VGND VPWR VPWR _5065_/C sky130_fd_sc_hd__o21ai_1
XFILLER_178_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4771_ _4657_/C _4846_/D _4771_/B1 VGND VGND VPWR VPWR _4771_/X sky130_fd_sc_hd__a21o_1
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6510_ _6705_/CLK _6510_/D wire3958/X VGND VGND VPWR VPWR _6510_/Q sky130_fd_sc_hd__dfrtp_1
X_3722_ _3722_/A _3722_/B _3722_/C _3722_/D VGND VGND VPWR VPWR _3723_/C sky130_fd_sc_hd__or4_1
XFILLER_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6441_ _6441_/A _6441_/B VGND VGND VPWR VPWR _6441_/X sky130_fd_sc_hd__and2_1
X_3653_ _6086_/B2 _3653_/A2 _3332_/Y _3653_/B2 _3652_/X VGND VGND VPWR VPWR _3659_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6372_ _4228_/B _6372_/A2 _6372_/B1 _4228_/A VGND VGND VPWR VPWR _6372_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3584_ _7021_/Q _3736_/B1 _3777_/B1 _3584_/B2 _3559_/X VGND VGND VPWR VPWR _3588_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5323_ hold195/X _5476_/A0 _5325_/S VGND VGND VPWR VPWR _6906_/D sky130_fd_sc_hd__mux2_1
X_5254_ hold606/X _5254_/A1 _5254_/S VGND VGND VPWR VPWR _6845_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4205_ hold524/X _5530_/A1 _4209_/S VGND VGND VPWR VPWR _6660_/D sky130_fd_sc_hd__mux2_1
X_5185_ _5211_/A0 hold424/X _5186_/S VGND VGND VPWR VPWR _6791_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_3_6_0_csclk clkbuf_3_7_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_6_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_68_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4136_ hold420/X _5530_/A1 _4139_/S VGND VGND VPWR VPWR _6601_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4067_ hold87/X _4066_/X _4069_/S VGND VGND VPWR VPWR hold88/A sky130_fd_sc_hd__mux2_1
XFILLER_83_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4969_ _4969_/A _4969_/B VGND VGND VPWR VPWR _5114_/B sky130_fd_sc_hd__nand2_1
XFILLER_11_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length4059 fanout4057/X VGND VGND VPWR VPWR wire4058/A sky130_fd_sc_hd__buf_2
X_6708_ _7091_/CLK _6708_/D wire4029/X VGND VGND VPWR VPWR _6708_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_177_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length2624 _6040_/X VGND VGND VPWR VPWR wire2617/A sky130_fd_sc_hd__clkbuf_1
X_6639_ _7206_/CLK _6639_/D VGND VGND VPWR VPWR _6639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1200 _3320_/Y VGND VGND VPWR VPWR _3615_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_87_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1211 wire1212/X VGND VGND VPWR VPWR _3719_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire1222 _3615_/A2 VGND VGND VPWR VPWR _3346_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1233 _3540_/A2 VGND VGND VPWR VPWR _3697_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_170_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1244 _3653_/A2 VGND VGND VPWR VPWR _3440_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_47_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1255 _3681_/A2 VGND VGND VPWR VPWR wire1255/X sky130_fd_sc_hd__clkbuf_1
Xwire1277 wire1277/A VGND VGND VPWR VPWR _3361_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire1288 _3287_/Y VGND VGND VPWR VPWR _4001_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1299 hold28/X VGND VGND VPWR VPWR hold29/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire530 wire531/X VGND VGND VPWR VPWR wire530/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire541 wire542/X VGND VGND VPWR VPWR wire541/X sky130_fd_sc_hd__clkbuf_1
Xwire552 _3644_/X VGND VGND VPWR VPWR _3651_/A sky130_fd_sc_hd__clkbuf_1
Xwire563 _3520_/X VGND VGND VPWR VPWR _3524_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_171_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire574 wire575/X VGND VGND VPWR VPWR _3392_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire585 _6143_/X VGND VGND VPWR VPWR wire585/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3180 _4595_/Y VGND VGND VPWR VPWR _4655_/B sky130_fd_sc_hd__buf_2
Xwire3191 _5076_/B VGND VGND VPWR VPWR _4799_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_78_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2490 _6018_/Y VGND VGND VPWR VPWR _6023_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6990_ _7115_/CLK _6990_/D _7030_/RESET_B VGND VGND VPWR VPWR _6990_/Q sky130_fd_sc_hd__dfrtp_1
X_5941_ _6311_/A1 _5941_/A2 _5941_/B1 _6684_/Q VGND VGND VPWR VPWR _5941_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5872_ _5872_/A _5872_/B VGND VGND VPWR VPWR _5872_/X sky130_fd_sc_hd__or2_1
XFILLER_61_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4823_ _4823_/A _5158_/A _4823_/C _4778_/Y VGND VGND VPWR VPWR _4823_/X sky130_fd_sc_hd__or4b_1
XFILLER_178_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4754_ _4995_/A _4754_/B VGND VGND VPWR VPWR _4984_/B sky130_fd_sc_hd__nor2_1
XFILLER_193_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3705_ _7091_/Q _3705_/A2 _3460_/Y _6250_/B2 _3704_/X VGND VGND VPWR VPWR _3710_/B
+ sky130_fd_sc_hd__a221o_1
X_4685_ _4687_/B _4685_/A2 _4672_/X VGND VGND VPWR VPWR _4714_/A sky130_fd_sc_hd__o21ai_1
XFILLER_146_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3636_ _3636_/A1 _3636_/A2 _3636_/B1 _3636_/B2 VGND VGND VPWR VPWR _3636_/X sky130_fd_sc_hd__a22o_1
X_6424_ _6437_/A _6441_/B VGND VGND VPWR VPWR _6424_/X sky130_fd_sc_hd__and2_1
XFILLER_174_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6355_ _7195_/Q wire375/X _6356_/S VGND VGND VPWR VPWR _7195_/D sky130_fd_sc_hd__mux2_1
X_3567_ _6689_/Q _4240_/A _3567_/B1 _6311_/A1 VGND VGND VPWR VPWR _3567_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5306_ _5342_/A0 hold156/X _5307_/S VGND VGND VPWR VPWR _6891_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6286_ _6286_/A1 _6286_/A2 _6286_/B1 _6623_/Q _6286_/C1 VGND VGND VPWR VPWR _6291_/B
+ sky130_fd_sc_hd__a221o_1
X_3498_ _3498_/A1 _3498_/A2 _3681_/B1 _6525_/Q wire817/X VGND VGND VPWR VPWR _3499_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5237_ _5237_/A0 hold33/X _5240_/S VGND VGND VPWR VPWR hold34/A sky130_fd_sc_hd__mux2_1
XFILLER_130_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5168_ _6781_/Q _5182_/A2 wire382/X wire353/X VGND VGND VPWR VPWR _6781_/D sky130_fd_sc_hd__a211o_1
XFILLER_124_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4119_ hold3/X _6587_/Q _4119_/S VGND VGND VPWR VPWR hold4/A sky130_fd_sc_hd__mux2_1
XFILLER_84_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5099_ _4657_/A _4667_/B _4488_/A _4607_/X _4829_/Y VGND VGND VPWR VPWR _5100_/D
+ sky130_fd_sc_hd__a311o_1
XFILLER_44_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length3166 _4692_/B VGND VGND VPWR VPWR _4920_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_153_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold7 hold7/A VGND VGND VPWR VPWR hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_181_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1041 _3512_/Y VGND VGND VPWR VPWR _4135_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_59_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1052 _3496_/Y VGND VGND VPWR VPWR _4129_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1063 _6392_/A VGND VGND VPWR VPWR _3776_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1074 _3652_/B1 VGND VGND VPWR VPWR _3719_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire1085 _3655_/A2 VGND VGND VPWR VPWR _3707_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1096 _3417_/Y VGND VGND VPWR VPWR _3585_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire360 wire361/X VGND VGND VPWR VPWR wire360/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4470_ _4512_/B _4521_/A VGND VGND VPWR VPWR _4510_/B sky130_fd_sc_hd__nand2_1
Xwire371 wire372/X VGND VGND VPWR VPWR wire371/X sky130_fd_sc_hd__clkbuf_1
XFILLER_156_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold407 _6666_/Q VGND VGND VPWR VPWR hold407/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire382 _5157_/X VGND VGND VPWR VPWR wire382/X sky130_fd_sc_hd__clkbuf_1
Xhold418 _6806_/Q VGND VGND VPWR VPWR hold418/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire393 wire394/X VGND VGND VPWR VPWR wire393/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3421_ _7100_/Q _3421_/A2 _3550_/B1 _3421_/B2 wire847/X VGND VGND VPWR VPWR _3445_/A
+ sky130_fd_sc_hd__a221o_1
Xhold429 _6968_/Q VGND VGND VPWR VPWR hold429/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6140_ _6502_/Q _6140_/A2 _6163_/B1 _6140_/B2 VGND VGND VPWR VPWR _6140_/X sky130_fd_sc_hd__a22o_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3352_ _3352_/A1 _5232_/A wire894/X _6197_/A1 _3351_/X VGND VGND VPWR VPWR _3352_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _6121_/A1 _7175_/Q wire454/X VGND VGND VPWR VPWR _6071_/X sky130_fd_sc_hd__a21o_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ hold69/X VGND VGND VPWR VPWR _3313_/B sky130_fd_sc_hd__inv_2
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _4638_/X _5017_/B _5021_/X VGND VGND VPWR VPWR _5079_/B sky130_fd_sc_hd__o21ai_1
XFILLER_38_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6973_ _6973_/CLK _6973_/D wire4069/X VGND VGND VPWR VPWR _6973_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_81_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5924_ _5924_/A1 _5946_/A2 _5913_/X _5923_/X _5946_/C1 VGND VGND VPWR VPWR _5924_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_34_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5855_ _6897_/Q _5855_/A2 _5855_/B1 _6214_/A1 VGND VGND VPWR VPWR _5855_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4806_ _4971_/A _4749_/C _4607_/D _4574_/Y VGND VGND VPWR VPWR _4806_/X sky130_fd_sc_hd__a31o_1
X_5786_ _5786_/A1 _5786_/A2 _5786_/B1 _5786_/B2 _5776_/X VGND VGND VPWR VPWR _5786_/X
+ sky130_fd_sc_hd__a221o_1
Xmax_length908 _3333_/Y VGND VGND VPWR VPWR wire904/A sky130_fd_sc_hd__clkbuf_1
XFILLER_119_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4737_ _4758_/C _5001_/C VGND VGND VPWR VPWR _4739_/B sky130_fd_sc_hd__nand2_1
XFILLER_119_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4668_ _4668_/A _4739_/A VGND VGND VPWR VPWR _4668_/X sky130_fd_sc_hd__or2_1
XFILLER_79_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length1038 _3767_/B1 VGND VGND VPWR VPWR _3555_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_107_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6407_ _6407_/A _6407_/B VGND VGND VPWR VPWR _6407_/X sky130_fd_sc_hd__and2_1
X_3619_ _3619_/A1 _3308_/Y wire926/X _6900_/Q _3618_/X VGND VGND VPWR VPWR _3619_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_190_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4599_ _5115_/A _4599_/B _4984_/A _4584_/X VGND VGND VPWR VPWR _4599_/X sky130_fd_sc_hd__or4b_1
XFILLER_162_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3905 wire3906/X VGND VGND VPWR VPWR wire3905/X sky130_fd_sc_hd__clkbuf_1
Xwire3916 wire3917/X VGND VGND VPWR VPWR wire3916/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3927 _3918_/S VGND VGND VPWR VPWR _3921_/S sky130_fd_sc_hd__clkbuf_2
X_6338_ _6720_/Q _6338_/A2 _6338_/B1 _6770_/Q VGND VGND VPWR VPWR _6338_/X sky130_fd_sc_hd__a22o_1
Xwire3938 _6430_/A VGND VGND VPWR VPWR _6433_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_115_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6269_ _7183_/Q _6343_/A2 _5650_/Y VGND VGND VPWR VPWR _6269_/X sky130_fd_sc_hd__o21ba_1
XFILLER_130_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_3_0_csclk clkbuf_2_3_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_7_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_151_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3970_ hold715/X _5231_/A0 _3976_/S VGND VGND VPWR VPWR _6475_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5640_ _7158_/Q _7157_/Q VGND VGND VPWR VPWR _6040_/B sky130_fd_sc_hd__and2b_2
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5571_ _5571_/A _5571_/B VGND VGND VPWR VPWR _5579_/S sky130_fd_sc_hd__nand2_2
XFILLER_191_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4522_ _4527_/A1 _4520_/B _4519_/X _4520_/X _5054_/A VGND VGND VPWR VPWR _4522_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_172_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold204 _6973_/Q VGND VGND VPWR VPWR hold204/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 _6889_/Q VGND VGND VPWR VPWR hold215/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 _6704_/Q VGND VGND VPWR VPWR hold226/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4453_ _4453_/A _4724_/A _4453_/C VGND VGND VPWR VPWR _4453_/X sky130_fd_sc_hd__or3_1
XFILLER_172_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold237 _6606_/Q VGND VGND VPWR VPWR hold237/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold248 _6589_/Q VGND VGND VPWR VPWR hold248/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold259 _6502_/Q VGND VGND VPWR VPWR hold259/X sky130_fd_sc_hd__dlygate4sd3_1
X_3404_ _6188_/A1 _3437_/A2 _3442_/A2 _6187_/B2 _3403_/X VGND VGND VPWR VPWR _3408_/B
+ sky130_fd_sc_hd__a221o_1
X_7172_ _7185_/CLK _7172_/D wire3950/A VGND VGND VPWR VPWR _7172_/Q sky130_fd_sc_hd__dfrtp_1
X_4384_ _4495_/A _4385_/B VGND VGND VPWR VPWR _4999_/B sky130_fd_sc_hd__nor2_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6123_ _6123_/A1 _6197_/A2 _6197_/B1 _6123_/B2 VGND VGND VPWR VPWR _6123_/X sky130_fd_sc_hd__a22o_1
X_3335_ _3546_/A _3339_/B VGND VGND VPWR VPWR _3335_/Y sky130_fd_sc_hd__nor2_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6054_ _6987_/Q _6054_/A2 _6054_/B1 _6054_/B2 VGND VGND VPWR VPWR _6054_/X sky130_fd_sc_hd__a22o_1
X_3266_ _3288_/A hold83/X VGND VGND VPWR VPWR _3416_/A sky130_fd_sc_hd__and2b_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _4931_/B _4744_/C _5001_/C _4896_/B _4770_/A VGND VGND VPWR VPWR _5134_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_100_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3197_ _7138_/Q VGND VGND VPWR VPWR _3197_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6956_ _6956_/CLK _6956_/D wire4040/X VGND VGND VPWR VPWR _6956_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_41_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5907_ _6288_/B2 _5934_/B1 _5961_/A2 _5907_/B2 VGND VGND VPWR VPWR _5907_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6887_ _7116_/CLK _6887_/D wire4071/A VGND VGND VPWR VPWR _6887_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_179_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5838_ _7168_/Q _5837_/X _5838_/S VGND VGND VPWR VPWR _7168_/D sky130_fd_sc_hd__mux2_1
XFILLER_22_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5769_ _6100_/B2 _5807_/A2 _5807_/B1 _5769_/B2 _5768_/X VGND VGND VPWR VPWR _5770_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_6_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3702 _6120_/C1 VGND VGND VPWR VPWR _6095_/C1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3713 _7214_/X VGND VGND VPWR VPWR wire3713/X sky130_fd_sc_hd__clkbuf_1
Xwire3724 _7143_/Q VGND VGND VPWR VPWR wire3724/X sky130_fd_sc_hd__clkbuf_1
Xwire3735 wire3736/X VGND VGND VPWR VPWR _3263_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire3746 _4548_/B1 VGND VGND VPWR VPWR _4228_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_89_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3757 _6696_/Q VGND VGND VPWR VPWR wire3757/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3768 _6630_/Q VGND VGND VPWR VPWR wire3768/X sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3779 _3850_/A VGND VGND VPWR VPWR _3820_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_103_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput309 _3380_/X VGND VGND VPWR VPWR serial_data_2 sky130_fd_sc_hd__buf_12
XFILLER_181_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6810_ _7081_/CLK _6810_/D _7159_/RESET_B VGND VGND VPWR VPWR _6810_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6741_ _6799_/CLK _6741_/D fanout3952/X VGND VGND VPWR VPWR _6741_/Q sky130_fd_sc_hd__dfrtp_1
X_3953_ _6459_/Q _3953_/B VGND VGND VPWR VPWR _3953_/X sky130_fd_sc_hd__and2b_1
XFILLER_16_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3884_ _3884_/A _3884_/B wire4278/X wire4251/X VGND VGND VPWR VPWR _3886_/C sky130_fd_sc_hd__or4bb_1
XFILLER_176_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6672_ _6683_/CLK _6672_/D _6672_/SET_B VGND VGND VPWR VPWR _6672_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_31_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5623_ _7151_/Q _5624_/B _5622_/B _5625_/S VGND VGND VPWR VPWR _7151_/D sky130_fd_sc_hd__a31o_1
XFILLER_149_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5554_ _5554_/A0 hold337/X _5555_/S VGND VGND VPWR VPWR _7111_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4505_ _4527_/A1 _4858_/A1 _4503_/X _4504_/X VGND VGND VPWR VPWR _4505_/X sky130_fd_sc_hd__o211a_1
X_5485_ _5485_/A0 _5990_/A1 _5491_/S VGND VGND VPWR VPWR _7050_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4436_ _4436_/A _4436_/B VGND VGND VPWR VPWR _4744_/C sky130_fd_sc_hd__nor2_1
Xwire3009 wire3010/X VGND VGND VPWR VPWR _5865_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_104_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4367_ _4846_/B _4367_/B VGND VGND VPWR VPWR _4367_/Y sky130_fd_sc_hd__nand2_1
X_7155_ _7180_/CLK _7155_/D wire3996/X VGND VGND VPWR VPWR _7155_/Q sky130_fd_sc_hd__dfrtp_1
Xwire2308 _6623_/Q VGND VGND VPWR VPWR _5922_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2319 _5931_/A1 VGND VGND VPWR VPWR _3572_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_116_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3318_ _3466_/A _3318_/B VGND VGND VPWR VPWR _3318_/Y sky130_fd_sc_hd__nor2_1
Xwire1607 wire1608/X VGND VGND VPWR VPWR _6112_/A1 sky130_fd_sc_hd__clkbuf_1
X_6106_ _6106_/A1 _6166_/A2 _6139_/B1 _6885_/Q _6105_/X VGND VGND VPWR VPWR _6109_/C
+ sky130_fd_sc_hd__a221o_1
X_7086_ _7140_/CLK _7086_/D wire4065/X VGND VGND VPWR VPWR _7086_/Q sky130_fd_sc_hd__dfrtp_1
X_4298_ _4298_/A0 hold302/X _4299_/S VGND VGND VPWR VPWR _4298_/X sky130_fd_sc_hd__mux2_1
Xwire1618 _7078_/Q VGND VGND VPWR VPWR _3469_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire1629 _7071_/Q VGND VGND VPWR VPWR _3438_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3249_ hold24/X _3820_/A _3248_/Y VGND VGND VPWR VPWR hold25/A sky130_fd_sc_hd__a21bo_1
X_6037_ _7119_/Q _6073_/B1 _6065_/B1 _6037_/B2 VGND VGND VPWR VPWR _6037_/X sky130_fd_sc_hd__a22o_1
XFILLER_39_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6939_ _6939_/CLK _6939_/D wire4090/X VGND VGND VPWR VPWR _6939_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_25_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire904 wire904/A VGND VGND VPWR VPWR _4102_/S sky130_fd_sc_hd__dlymetal6s2s_1
Xwire915 _3319_/Y VGND VGND VPWR VPWR wire915/X sky130_fd_sc_hd__clkbuf_2
XFILLER_167_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire926 wire929/A VGND VGND VPWR VPWR wire926/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire937 _3312_/Y VGND VGND VPWR VPWR wire937/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire948 wire950/X VGND VGND VPWR VPWR wire948/X sky130_fd_sc_hd__clkbuf_1
XFILLER_157_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire959 wire960/X VGND VGND VPWR VPWR wire959/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_csclk _3942_/X VGND VGND VPWR VPWR clkbuf_0_csclk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_163_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire4200 wire4201/X VGND VGND VPWR VPWR wire4200/X sky130_fd_sc_hd__clkbuf_1
XFILLER_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4211 input42/X VGND VGND VPWR VPWR wire4211/X sky130_fd_sc_hd__clkbuf_1
Xwire4222 wire4223/X VGND VGND VPWR VPWR wire4222/X sky130_fd_sc_hd__clkbuf_1
Xwire4233 wire4234/X VGND VGND VPWR VPWR wire4233/X sky130_fd_sc_hd__clkbuf_1
Xwire4244 input24/X VGND VGND VPWR VPWR wire4244/X sky130_fd_sc_hd__clkbuf_1
XFILLER_150_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire4255 wire4255/A VGND VGND VPWR VPWR wire4255/X sky130_fd_sc_hd__clkbuf_1
Xwire3510 wire3511/X VGND VGND VPWR VPWR _5506_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_123_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire4266 wire4267/X VGND VGND VPWR VPWR wire4266/X sky130_fd_sc_hd__clkbuf_1
Xhold590 _6591_/Q VGND VGND VPWR VPWR hold590/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire4277 input14/X VGND VGND VPWR VPWR _3595_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3532 wire3532/A VGND VGND VPWR VPWR wire3532/X sky130_fd_sc_hd__clkbuf_1
Xwire4288 _4379_/C VGND VGND VPWR VPWR _4591_/A sky130_fd_sc_hd__buf_2
Xwire3543 wire3543/A VGND VGND VPWR VPWR _4285_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_104_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire4299 _4376_/A VGND VGND VPWR VPWR _4495_/A sky130_fd_sc_hd__clkbuf_2
Xwire3565 _5547_/A0 VGND VGND VPWR VPWR _5343_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2820 _6051_/A2 VGND VGND VPWR VPWR _6076_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2831 _5806_/B1 VGND VGND VPWR VPWR _5755_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3587 wire3587/A VGND VGND VPWR VPWR _4314_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2842 _5780_/B1 VGND VGND VPWR VPWR _5717_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire2853 _5845_/B1 VGND VGND VPWR VPWR _5810_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire3598 _5522_/A0 VGND VGND VPWR VPWR _5387_/A0 sky130_fd_sc_hd__clkbuf_1
Xwire2864 _5854_/B1 VGND VGND VPWR VPWR wire2864/X sky130_fd_sc_hd__clkbuf_1
Xwire2875 _5834_/B1 VGND VGND VPWR VPWR _5800_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire2886 _5954_/A2 VGND VGND VPWR VPWR _5886_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2897 _5966_/B1 VGND VGND VPWR VPWR _5888_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_18_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_1_0_1_csclk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_18_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5270_ _5342_/A0 hold162/X _5273_/S VGND VGND VPWR VPWR _6859_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4221_ _5534_/A1 hold309/X _4221_/S VGND VGND VPWR VPWR _6674_/D sky130_fd_sc_hd__mux2_1
Xfanout3960 wire3970/A VGND VGND VPWR VPWR wire3963/A sky130_fd_sc_hd__clkbuf_1
XFILLER_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout3982 wire4016/A VGND VGND VPWR VPWR wire3985/A sky130_fd_sc_hd__buf_6
Xfanout3993 wire4016/X VGND VGND VPWR VPWR fanout3993/X sky130_fd_sc_hd__clkbuf_1
X_4152_ _4251_/A0 hold295/X _4152_/S VGND VGND VPWR VPWR _6615_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4083_ hold246/X _4127_/A0 _4083_/S VGND VGND VPWR VPWR _4083_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4985_ _4985_/A _4985_/B _4985_/C VGND VGND VPWR VPWR _4988_/B sky130_fd_sc_hd__or3_1
XFILLER_189_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6724_ _6979_/CLK _6724_/D fanout4027/X VGND VGND VPWR VPWR _6724_/Q sky130_fd_sc_hd__dfrtp_1
X_3936_ hold10/A user_clock _6822_/Q VGND VGND VPWR VPWR _3936_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_2_0_csclk clkbuf_3_3_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_2_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_176_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6655_ _6683_/CLK _6655_/D _6672_/SET_B VGND VGND VPWR VPWR _6655_/Q sky130_fd_sc_hd__dfrtp_1
Xmax_length3529 hold49/X VGND VGND VPWR VPWR _5281_/A0 sky130_fd_sc_hd__clkbuf_1
X_3867_ _6473_/Q _6471_/Q _6541_/Q VGND VGND VPWR VPWR _3868_/B sky130_fd_sc_hd__and3_1
XFILLER_176_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5606_ _5606_/A _5606_/B _5606_/C VGND VGND VPWR VPWR _7146_/D sky130_fd_sc_hd__and3_1
Xmax_length2817 _5982_/X VGND VGND VPWR VPWR _6024_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_192_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6586_ _7131_/CLK hold46/X wire4058/X VGND VGND VPWR VPWR _6586_/Q sky130_fd_sc_hd__dfrtp_1
X_3798_ _6473_/Q _3800_/A VGND VGND VPWR VPWR _6473_/D sky130_fd_sc_hd__xor2_1
XFILLER_191_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5537_ hold621/X _5537_/A1 _5538_/S VGND VGND VPWR VPWR _7096_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5468_ hold72/X _5468_/A1 _5468_/S VGND VGND VPWR VPWR hold73/A sky130_fd_sc_hd__mux2_1
X_7207_ _7210_/CLK _7207_/D wire4019/A VGND VGND VPWR VPWR _7207_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4419_ _4566_/A _4419_/B _4451_/A VGND VGND VPWR VPWR _4459_/B sky130_fd_sc_hd__and3b_1
Xwire2105 wire2106/X VGND VGND VPWR VPWR _3647_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_59_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2116 _6813_/Q VGND VGND VPWR VPWR _3501_/B2 sky130_fd_sc_hd__clkbuf_1
X_5399_ hold122/X _5498_/A0 _5399_/S VGND VGND VPWR VPWR _5399_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2127 wire2128/X VGND VGND VPWR VPWR _3695_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_132_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7138_ _7140_/CLK _7138_/D _7138_/RESET_B VGND VGND VPWR VPWR _7138_/Q sky130_fd_sc_hd__dfrtp_1
Xwire2138 wire2139/X VGND VGND VPWR VPWR wire2138/X sky130_fd_sc_hd__clkbuf_1
Xwire2149 _6774_/Q VGND VGND VPWR VPWR _6304_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire1404 _6320_/X VGND VGND VPWR VPWR _6332_/A sky130_fd_sc_hd__clkbuf_1
Xwire1415 wire1416/X VGND VGND VPWR VPWR _5928_/C1 sky130_fd_sc_hd__clkbuf_1
XFILLER_59_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1426 _5704_/X VGND VGND VPWR VPWR wire1426/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1448 wire1449/X VGND VGND VPWR VPWR wire1448/X sky130_fd_sc_hd__clkbuf_2
XFILLER_47_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7069_ _7137_/CLK _7069_/D _7137_/RESET_B VGND VGND VPWR VPWR _7069_/Q sky130_fd_sc_hd__dfrtp_1
Xwire1459 wire1460/X VGND VGND VPWR VPWR wire1459/X sky130_fd_sc_hd__clkbuf_1
XFILLER_46_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire701 _5336_/S VGND VGND VPWR VPWR _5337_/S sky130_fd_sc_hd__clkbuf_1
Xwire712 _5031_/X VGND VGND VPWR VPWR _5071_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_10_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire723 wire724/X VGND VGND VPWR VPWR wire723/X sky130_fd_sc_hd__clkbuf_1
Xwire734 _4004_/S VGND VGND VPWR VPWR wire734/X sky130_fd_sc_hd__clkbuf_1
Xinput19 mask_rev_in[23] VGND VGND VPWR VPWR input19/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire745 wire746/X VGND VGND VPWR VPWR wire745/X sky130_fd_sc_hd__clkbuf_1
XFILLER_168_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire756 wire757/X VGND VGND VPWR VPWR wire756/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire767 wire768/X VGND VGND VPWR VPWR wire767/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire778 _3567_/X VGND VGND VPWR VPWR wire778/X sky130_fd_sc_hd__clkbuf_1
Xwire789 _3550_/X VGND VGND VPWR VPWR wire789/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire4041 wire4042/X VGND VGND VPWR VPWR wire4041/X sky130_fd_sc_hd__clkbuf_2
XFILLER_151_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4052 wire4052/A VGND VGND VPWR VPWR wire4052/X sky130_fd_sc_hd__buf_2
XFILLER_96_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3340 _4652_/A VGND VGND VPWR VPWR _4958_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire4096 input75/X VGND VGND VPWR VPWR wire4096/X sky130_fd_sc_hd__clkbuf_1
Xwire3351 _4387_/B VGND VGND VPWR VPWR _4451_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3362 _4372_/Y VGND VGND VPWR VPWR _4778_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3373 _5501_/A0 VGND VGND VPWR VPWR _5339_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3384 _5411_/A0 VGND VGND VPWR VPWR _5543_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3395 _5587_/A0 VGND VGND VPWR VPWR _5491_/A0 sky130_fd_sc_hd__clkbuf_2
Xwire2650 wire2650/A VGND VGND VPWR VPWR _6088_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire2661 _6191_/B1 VGND VGND VPWR VPWR _6282_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire2672 _6025_/D VGND VGND VPWR VPWR wire2672/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2683 _6175_/B1 VGND VGND VPWR VPWR _6073_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire2694 wire2694/A VGND VGND VPWR VPWR _6172_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire1960 _6917_/Q VGND VGND VPWR VPWR _6115_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1971 _6909_/Q VGND VGND VPWR VPWR _5766_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire1982 wire1983/X VGND VGND VPWR VPWR _3440_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_80_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4770_ _4770_/A _4770_/B _4770_/C _4882_/B VGND VGND VPWR VPWR _4770_/X sky130_fd_sc_hd__or4b_1
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3721_ _3721_/A _3721_/B _3721_/C _3721_/D VGND VGND VPWR VPWR _3722_/D sky130_fd_sc_hd__or4_1
XFILLER_158_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6440_ _6440_/A _6440_/B VGND VGND VPWR VPWR _6440_/X sky130_fd_sc_hd__and2_1
XFILLER_174_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3652_ _6088_/B2 _3652_/A2 _3652_/B1 _6763_/Q VGND VGND VPWR VPWR _3652_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6371_ _6370_/X hold77/A _6386_/S VGND VGND VPWR VPWR _7199_/D sky130_fd_sc_hd__mux2_1
X_3583_ _3583_/A _3583_/B _3583_/C _3583_/D VGND VGND VPWR VPWR _3583_/X sky130_fd_sc_hd__or4_1
XFILLER_127_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5322_ _5322_/A _5475_/B VGND VGND VPWR VPWR _5322_/X sky130_fd_sc_hd__and2_1
XFILLER_114_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5253_ hold398/X _5583_/A0 _5253_/S VGND VGND VPWR VPWR _6844_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4204_ _4204_/A _5529_/B VGND VGND VPWR VPWR _4209_/S sky130_fd_sc_hd__and2_2
XFILLER_87_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5184_ _5184_/A _5210_/B VGND VGND VPWR VPWR _5186_/S sky130_fd_sc_hd__nand2_1
XFILLER_68_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4135_ _4135_/A _4135_/B VGND VGND VPWR VPWR _4139_/S sky130_fd_sc_hd__and2_1
XFILLER_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_63_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7080_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_28_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4066_ _6586_/Q _4118_/A0 _4068_/S VGND VGND VPWR VPWR _4066_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_78_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6824_/CLK sky130_fd_sc_hd__clkbuf_16
X_4968_ _4969_/B VGND VGND VPWR VPWR _5100_/A sky130_fd_sc_hd__clkinv_2
XFILLER_51_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6707_ _7091_/CLK _6707_/D wire4029/A VGND VGND VPWR VPWR _6707_/Q sky130_fd_sc_hd__dfrtp_1
X_3919_ _6578_/Q _3919_/A1 _3921_/S VGND VGND VPWR VPWR _3919_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4899_ _5059_/A _4899_/B VGND VGND VPWR VPWR _5130_/B sky130_fd_sc_hd__or2_1
XFILLER_20_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3348 _4662_/B VGND VGND VPWR VPWR _4669_/B2 sky130_fd_sc_hd__clkbuf_1
X_6638_ _6683_/CLK _6638_/D wire3965/A VGND VGND VPWR VPWR _6638_/Q sky130_fd_sc_hd__dfrtp_1
Xmax_length3359 _4993_/A VGND VGND VPWR VPWR _4763_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_192_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6569_ _6973_/CLK _6569_/D wire4069/X VGND VGND VPWR VPWR _6569_/Q sky130_fd_sc_hd__dfrtp_1
Xmax_length2669 _6327_/B1 VGND VGND VPWR VPWR _6265_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_106_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_16_csclk _7059_/CLK VGND VGND VPWR VPWR _6671_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_121_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1201 wire1201/A VGND VGND VPWR VPWR _3437_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire1212 _3596_/A2 VGND VGND VPWR VPWR wire1212/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1223 _3311_/Y VGND VGND VPWR VPWR _3615_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1234 _3304_/Y VGND VGND VPWR VPWR _3540_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1256 _3654_/A2 VGND VGND VPWR VPWR _3681_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire1267 _3294_/Y VGND VGND VPWR VPWR _5535_/A sky130_fd_sc_hd__clkbuf_2
Xwire1289 _3504_/A VGND VGND VPWR VPWR _3466_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_43_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire520 _5091_/X VGND VGND VPWR VPWR _5092_/D sky130_fd_sc_hd__clkbuf_1
Xwire531 wire532/X VGND VGND VPWR VPWR wire531/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire542 _3732_/X VGND VGND VPWR VPWR wire542/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire553 _3637_/X VGND VGND VPWR VPWR _3642_/B sky130_fd_sc_hd__clkbuf_1
Xwire564 _3505_/X VGND VGND VPWR VPWR wire564/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire575 wire576/X VGND VGND VPWR VPWR wire575/X sky130_fd_sc_hd__clkbuf_1
Xwire586 _6110_/X VGND VGND VPWR VPWR wire586/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire597 _5516_/S VGND VGND VPWR VPWR _5515_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_171_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3170 _4704_/B VGND VGND VPWR VPWR _5161_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3192 _5076_/B VGND VGND VPWR VPWR _4590_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2480 _6025_/C VGND VGND VPWR VPWR _6282_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2491 _6137_/B1 VGND VGND VPWR VPWR _6062_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_19_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1790 _7008_/Q VGND VGND VPWR VPWR _6177_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_92_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5940_ _6524_/Q _5940_/A2 _5952_/B1 _6314_/A1 _5939_/X VGND VGND VPWR VPWR _5945_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5871_ _6236_/B2 _5953_/A2 _5915_/A2 _6686_/Q _5870_/X VGND VGND VPWR VPWR _5879_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_179_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4822_ _4822_/A _4822_/B _4822_/C _4882_/A VGND VGND VPWR VPWR _4823_/C sky130_fd_sc_hd__or4b_1
XFILLER_61_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4753_ _4753_/A _4753_/B VGND VGND VPWR VPWR _4753_/Y sky130_fd_sc_hd__nor2_1
X_3704_ _6712_/Q _3489_/Y wire804/X _6622_/Q VGND VGND VPWR VPWR _3704_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4684_ _4684_/A _4684_/B VGND VGND VPWR VPWR _4860_/B sky130_fd_sc_hd__nand2_1
XFILLER_147_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6423_ _6438_/A _6435_/B VGND VGND VPWR VPWR _6423_/X sky130_fd_sc_hd__and2_1
X_3635_ _7068_/Q _3693_/A2 _3635_/B1 _5739_/B2 _3634_/X VGND VGND VPWR VPWR _3635_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6354_ _7194_/Q wire371/X _6356_/S VGND VGND VPWR VPWR _7194_/D sky130_fd_sc_hd__mux2_1
X_3566_ _3566_/A1 wire944/X _3566_/B1 _7122_/Q wire560/X VGND VGND VPWR VPWR _3573_/A
+ sky130_fd_sc_hd__a221o_1
X_5305_ _5581_/A0 hold340/X _5307_/S VGND VGND VPWR VPWR _6890_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3497_ _6802_/Q _3417_/Y _4129_/A _6600_/Q VGND VGND VPWR VPWR _3497_/X sky130_fd_sc_hd__a22o_1
X_6285_ _6688_/Q _6337_/A2 _6312_/B1 _6285_/B2 VGND VGND VPWR VPWR _6285_/X sky130_fd_sc_hd__a22o_1
XFILLER_88_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5236_ _5575_/A0 hold201/X _5240_/S VGND VGND VPWR VPWR _6829_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5167_ _5148_/Y _5151_/X _5166_/Y _5147_/X VGND VGND VPWR VPWR _5167_/X sky130_fd_sc_hd__a211o_1
XFILLER_96_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4118_ _4118_/A0 _6586_/Q _4119_/S VGND VGND VPWR VPWR hold46/A sky130_fd_sc_hd__mux2_1
XFILLER_68_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5098_ _4997_/A _4728_/Y _4983_/Y _4618_/D VGND VGND VPWR VPWR _5142_/B sky130_fd_sc_hd__o211ai_2
XFILLER_140_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4049_ _4049_/A0 hold291/X _4051_/S VGND VGND VPWR VPWR _6538_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3178 _4611_/X VGND VGND VPWR VPWR _4976_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_153_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length3189 _4567_/X VGND VGND VPWR VPWR _4688_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1020 wire1021/X VGND VGND VPWR VPWR wire1020/X sky130_fd_sc_hd__clkbuf_1
XFILLER_47_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold8 hold8/A VGND VGND VPWR VPWR hold8/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire1031 _3774_/B1 VGND VGND VPWR VPWR _4312_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1042 _3512_/Y VGND VGND VPWR VPWR _3677_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1053 _3495_/Y VGND VGND VPWR VPWR _3681_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_181_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1064 _4022_/A VGND VGND VPWR VPWR _3687_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1075 _4318_/A VGND VGND VPWR VPWR _3786_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_75_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1086 _4306_/A VGND VGND VPWR VPWR _3655_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_47_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire350 _4818_/X VGND VGND VPWR VPWR _4821_/B sky130_fd_sc_hd__clkbuf_1
Xwire361 wire362/X VGND VGND VPWR VPWR wire361/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire372 wire373/X VGND VGND VPWR VPWR wire372/X sky130_fd_sc_hd__clkbuf_1
Xwire383 _5140_/X VGND VGND VPWR VPWR _5172_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_144_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold408 _6566_/Q VGND VGND VPWR VPWR hold408/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_156_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire394 _3789_/X VGND VGND VPWR VPWR wire394/X sky130_fd_sc_hd__clkbuf_1
Xhold419 _6595_/Q VGND VGND VPWR VPWR hold419/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3420_ _6479_/Q _3420_/A2 _5448_/A _7023_/Q VGND VGND VPWR VPWR _3420_/X sky130_fd_sc_hd__a22o_1
XFILLER_7_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3351_ _3351_/A1 _5553_/A _5439_/A _3351_/B2 VGND VGND VPWR VPWR _3351_/X sky130_fd_sc_hd__a22o_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3282_ _3282_/A hold68/X VGND VGND VPWR VPWR hold69/A sky130_fd_sc_hd__nand2_1
XFILLER_98_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6070_ _6070_/A1 wire978/X _6069_/X _6070_/C1 VGND VGND VPWR VPWR _6070_/X sky130_fd_sc_hd__o211a_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _5021_/A _5021_/B _5021_/C VGND VGND VPWR VPWR _5021_/X sky130_fd_sc_hd__or3_1
XFILLER_85_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6972_ _7046_/CLK _6972_/D wire4052/X VGND VGND VPWR VPWR _6972_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5923_ _5923_/A _5923_/B _5923_/C _5923_/D VGND VGND VPWR VPWR _5923_/X sky130_fd_sc_hd__or4_1
XFILLER_81_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5854_ _6993_/Q _5854_/A2 _5854_/B1 _6985_/Q _5853_/X VGND VGND VPWR VPWR _5857_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4805_ _4814_/A _5169_/A1 _4590_/A _4753_/B _4805_/B2 VGND VGND VPWR VPWR _4805_/X
+ sky130_fd_sc_hd__o32a_1
X_5785_ _5785_/A _5785_/B _5785_/C _5785_/D VGND VGND VPWR VPWR _5785_/X sky130_fd_sc_hd__or4_1
XFILLER_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4736_ _4748_/A _4997_/A VGND VGND VPWR VPWR _5049_/B sky130_fd_sc_hd__nor2_1
XFILLER_175_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4667_ _4596_/A _4667_/B _4667_/C VGND VGND VPWR VPWR _4667_/X sky130_fd_sc_hd__and3b_1
XFILLER_147_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6406_ _6407_/A _6407_/B VGND VGND VPWR VPWR _6406_/X sky130_fd_sc_hd__and2_1
XFILLER_134_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3618_ _6075_/A1 wire895/X _4288_/A _3618_/B2 VGND VGND VPWR VPWR _3618_/X sky130_fd_sc_hd__a22o_1
X_4598_ _4965_/A _4598_/B _4983_/A _4598_/D VGND VGND VPWR VPWR _4599_/B sky130_fd_sc_hd__or4_1
XFILLER_122_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6337_ _6337_/A1 _6337_/A2 _6337_/B1 _6337_/B2 VGND VGND VPWR VPWR _6337_/X sky130_fd_sc_hd__a22o_1
Xwire3906 wire3907/X VGND VGND VPWR VPWR wire3906/X sky130_fd_sc_hd__clkbuf_1
X_3549_ _3549_/A1 wire900/X hold30/A _3549_/B2 VGND VGND VPWR VPWR _3549_/X sky130_fd_sc_hd__a22o_1
Xwire3917 input84/X VGND VGND VPWR VPWR wire3917/X sky130_fd_sc_hd__clkbuf_1
Xwire3928 wire3929/X VGND VGND VPWR VPWR _3918_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_143_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3939 _3946_/B VGND VGND VPWR VPWR _6430_/A sky130_fd_sc_hd__buf_2
XFILLER_115_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6268_ _6268_/A1 _6268_/A2 _6257_/X _6267_/X _6268_/C1 VGND VGND VPWR VPWR _6268_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_76_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5219_ _5518_/A0 hold514/X _5220_/S VGND VGND VPWR VPWR _6817_/D sky130_fd_sc_hd__mux2_1
X_6199_ _7057_/Q _6199_/A2 _6199_/B1 _6199_/B2 VGND VGND VPWR VPWR _6216_/A sky130_fd_sc_hd__a22o_1
XFILLER_84_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length2263 hold400/X VGND VGND VPWR VPWR _4226_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_180_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5570_ _5588_/A0 _6198_/B2 _5570_/S VGND VGND VPWR VPWR _7126_/D sky130_fd_sc_hd__mux2_1
XFILLER_157_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4521_ _4521_/A _4524_/B VGND VGND VPWR VPWR _5054_/A sky130_fd_sc_hd__nand2_1
XFILLER_144_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold205 _7127_/Q VGND VGND VPWR VPWR hold205/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold216 _7119_/Q VGND VGND VPWR VPWR hold216/X sky130_fd_sc_hd__dlygate4sd3_1
X_4452_ _4758_/A _5001_/A _4758_/B _4485_/B VGND VGND VPWR VPWR _5165_/D sky130_fd_sc_hd__nand4_1
Xhold227 _6949_/Q VGND VGND VPWR VPWR hold227/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 _6610_/Q VGND VGND VPWR VPWR hold238/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 _6623_/Q VGND VGND VPWR VPWR hold249/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3403_ _6182_/B2 wire917/X _3403_/B1 _3403_/B2 VGND VGND VPWR VPWR _3403_/X sky130_fd_sc_hd__a22o_1
X_7171_ _7185_/CLK _7171_/D fanout3952/X VGND VGND VPWR VPWR _7171_/Q sky130_fd_sc_hd__dfrtp_1
X_4383_ _4419_/B _4566_/A VGND VGND VPWR VPWR _4385_/B sky130_fd_sc_hd__nand2_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6122_ _7178_/Q _6121_/X _6122_/S VGND VGND VPWR VPWR _7178_/D sky130_fd_sc_hd__mux2_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3334_ _3511_/B _3338_/B VGND VGND VPWR VPWR _3334_/Y sky130_fd_sc_hd__nor2_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _6053_/A1 _6073_/A2 _6053_/B1 _6053_/B2 _6049_/X VGND VGND VPWR VPWR _6058_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3265_ hold82/X _3265_/A1 _3265_/S VGND VGND VPWR VPWR hold83/A sky130_fd_sc_hd__mux2_1
XFILLER_86_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _5133_/A1 _4487_/B _4897_/A VGND VGND VPWR VPWR _5148_/B sky130_fd_sc_hd__a21o_1
X_3196_ _6564_/Q VGND VGND VPWR VPWR _5650_/B sky130_fd_sc_hd__clkinv_2
XFILLER_93_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6955_ _6979_/CLK _6955_/D fanout4027/X VGND VGND VPWR VPWR _6955_/Q sky130_fd_sc_hd__dfstp_1
X_5906_ _5906_/A1 _5906_/A2 _5959_/A2 _5906_/B2 _5905_/X VGND VGND VPWR VPWR _5906_/X
+ sky130_fd_sc_hd__a221o_1
X_6886_ _7139_/CLK _6886_/D wire4065/X VGND VGND VPWR VPWR _6886_/Q sky130_fd_sc_hd__dfrtp_1
X_5837_ _5859_/A1 _7167_/Q _5836_/X VGND VGND VPWR VPWR _5837_/X sky130_fd_sc_hd__a21o_1
XFILLER_167_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5768_ _6116_/A1 _5768_/A2 _5817_/B1 _6105_/B2 _5768_/C1 VGND VGND VPWR VPWR _5768_/X
+ sky130_fd_sc_hd__a221o_1
X_4719_ _4719_/A _4721_/C VGND VGND VPWR VPWR _4720_/C sky130_fd_sc_hd__nor2_1
X_5699_ _7152_/Q _5699_/B _5699_/C VGND VGND VPWR VPWR _5699_/X sky130_fd_sc_hd__and3_1
XFILLER_30_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3703 wire3704/X VGND VGND VPWR VPWR _6120_/C1 sky130_fd_sc_hd__clkbuf_2
XFILLER_150_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3714 _7196_/Q VGND VGND VPWR VPWR wire3714/X sky130_fd_sc_hd__clkbuf_2
Xwire3725 _6782_/Q VGND VGND VPWR VPWR _5182_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire3736 wire3737/X VGND VGND VPWR VPWR wire3736/X sky130_fd_sc_hd__clkbuf_1
Xwire3747 wire3748/X VGND VGND VPWR VPWR _4548_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_131_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length1392 _3322_/A VGND VGND VPWR VPWR wire1391/A sky130_fd_sc_hd__clkbuf_1
XFILLER_95_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6740_ _6740_/CLK _6740_/D fanout4027/X VGND VGND VPWR VPWR _6740_/Q sky130_fd_sc_hd__dfrtp_1
X_3952_ _6460_/Q _3952_/B VGND VGND VPWR VPWR _3952_/X sky130_fd_sc_hd__and2b_1
XFILLER_189_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6671_ _6671_/CLK _6671_/D fanout4028/X VGND VGND VPWR VPWR _6671_/Q sky130_fd_sc_hd__dfrtp_1
X_3883_ _4390_/C _4390_/D VGND VGND VPWR VPWR _4654_/B sky130_fd_sc_hd__or2_1
XFILLER_188_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5622_ _7151_/Q _5622_/B VGND VGND VPWR VPWR _5625_/S sky130_fd_sc_hd__nor2_1
XFILLER_136_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5553_ _5553_/A _5553_/B VGND VGND VPWR VPWR _5553_/Y sky130_fd_sc_hd__nand2_1
XFILLER_191_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4504_ _4504_/A _4504_/B _4860_/A VGND VGND VPWR VPWR _4504_/X sky130_fd_sc_hd__and3_1
X_5484_ _5484_/A _5535_/B VGND VGND VPWR VPWR _5484_/Y sky130_fd_sc_hd__nand2_1
XFILLER_144_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4435_ _4435_/A _4435_/B VGND VGND VPWR VPWR _4453_/C sky130_fd_sc_hd__nand2_1
XFILLER_132_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7154_ _7187_/CLK _7154_/D wire3991/X VGND VGND VPWR VPWR _7154_/Q sky130_fd_sc_hd__dfstp_1
X_4366_ _4369_/B VGND VGND VPWR VPWR _4367_/B sky130_fd_sc_hd__inv_2
Xwire2309 _6621_/Q VGND VGND VPWR VPWR _6238_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_86_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6105_ _6105_/A1 _6141_/A2 _6172_/A2 _6105_/B2 VGND VGND VPWR VPWR _6105_/X sky130_fd_sc_hd__a22o_1
X_3317_ _3502_/B _3322_/A VGND VGND VPWR VPWR _3317_/Y sky130_fd_sc_hd__nor2_1
X_7085_ _7140_/CLK _7085_/D wire4065/X VGND VGND VPWR VPWR _7085_/Q sky130_fd_sc_hd__dfrtp_1
Xwire1608 _7085_/Q VGND VGND VPWR VPWR wire1608/X sky130_fd_sc_hd__clkbuf_1
X_4297_ _4309_/A0 hold286/X _4299_/S VGND VGND VPWR VPWR _4297_/X sky130_fd_sc_hd__mux2_1
Xwire1619 wire1620/X VGND VGND VPWR VPWR _3205_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_112_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6036_ _6040_/B _6039_/C _6040_/C VGND VGND VPWR VPWR _6036_/X sky130_fd_sc_hd__and3_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3248_ _6467_/Q _3252_/B VGND VGND VPWR VPWR _3248_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6938_ _6939_/CLK _6938_/D wire4090/X VGND VGND VPWR VPWR _6938_/Q sky130_fd_sc_hd__dfstp_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6869_ _6939_/CLK hold50/X _6404_/A VGND VGND VPWR VPWR _6869_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire905 wire907/X VGND VGND VPWR VPWR wire905/X sky130_fd_sc_hd__clkbuf_1
Xwire927 wire928/X VGND VGND VPWR VPWR _5313_/A sky130_fd_sc_hd__clkbuf_1
Xwire938 _4068_/S VGND VGND VPWR VPWR _4060_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_127_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4201 input45/X VGND VGND VPWR VPWR wire4201/X sky130_fd_sc_hd__clkbuf_1
Xfanout3405 hold44/X VGND VGND VPWR VPWR hold45/A sky130_fd_sc_hd__clkbuf_1
Xwire4212 wire4213/X VGND VGND VPWR VPWR _3961_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_2_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4223 input38/X VGND VGND VPWR VPWR wire4223/X sky130_fd_sc_hd__clkbuf_1
Xfanout3427 hold108/X VGND VGND VPWR VPWR wire3438/A sky130_fd_sc_hd__clkbuf_1
XFILLER_173_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire4234 input35/X VGND VGND VPWR VPWR wire4234/X sky130_fd_sc_hd__clkbuf_1
Xwire4245 input23/X VGND VGND VPWR VPWR _3584_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3500 _4250_/A0 VGND VGND VPWR VPWR _5533_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_151_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3511 wire3511/A VGND VGND VPWR VPWR wire3511/X sky130_fd_sc_hd__clkbuf_1
XFILLER_150_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3522 _5362_/A0 VGND VGND VPWR VPWR _5389_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_173_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire4267 wire4268/X VGND VGND VPWR VPWR wire4267/X sky130_fd_sc_hd__clkbuf_1
Xwire4278 wire4278/A VGND VGND VPWR VPWR wire4278/X sky130_fd_sc_hd__clkbuf_1
Xhold580 _6976_/Q VGND VGND VPWR VPWR hold580/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold591 _7102_/Q VGND VGND VPWR VPWR hold591/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire2810 wire2811/X VGND VGND VPWR VPWR _6237_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_77_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3555 wire3555/A VGND VGND VPWR VPWR _5505_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_103_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2821 _6125_/A2 VGND VGND VPWR VPWR _6051_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_173_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2832 _5855_/B1 VGND VGND VPWR VPWR _5806_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire3588 _5504_/A0 VGND VGND VPWR VPWR _4326_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2843 _5832_/B1 VGND VGND VPWR VPWR _5780_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2854 _5754_/B1 VGND VGND VPWR VPWR _5845_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire3599 _5477_/A0 VGND VGND VPWR VPWR _5396_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2865 _5702_/X VGND VGND VPWR VPWR _5854_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2876 _5849_/B1 VGND VGND VPWR VPWR _5834_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire2898 _5934_/B1 VGND VGND VPWR VPWR _5966_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_66_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_551 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4220_ _4250_/A0 hold308/X _4221_/S VGND VGND VPWR VPWR _6673_/D sky130_fd_sc_hd__mux2_1
X_4151_ _4250_/A0 hold311/X _4152_/S VGND VGND VPWR VPWR _6614_/D sky130_fd_sc_hd__mux2_1
XFILLER_122_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4082_ hold679/X _4081_/X _4082_/S VGND VGND VPWR VPWR _6559_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4984_ _4984_/A _4984_/B _4984_/C VGND VGND VPWR VPWR _5090_/B sky130_fd_sc_hd__or3_1
XFILLER_51_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6723_ _6979_/CLK hold65/X fanout4027/X VGND VGND VPWR VPWR _6723_/Q sky130_fd_sc_hd__dfstp_1
X_3935_ _3233_/Y input2/X input1/X VGND VGND VPWR VPWR _3935_/X sky130_fd_sc_hd__mux2_1
X_6654_ _7206_/CLK _6654_/D VGND VGND VPWR VPWR _6654_/Q sky130_fd_sc_hd__dfxtp_1
X_3866_ _3967_/A0 hold35/A _3866_/S VGND VGND VPWR VPWR _6446_/D sky130_fd_sc_hd__mux2_1
XFILLER_31_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3519 _5353_/A0 VGND VGND VPWR VPWR _5515_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_164_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5605_ _5605_/A VGND VGND VPWR VPWR _5606_/C sky130_fd_sc_hd__clkinv_2
X_6585_ _7129_/CLK _6585_/D wire4055/X VGND VGND VPWR VPWR _6585_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3797_ _6473_/Q _6472_/Q VGND VGND VPWR VPWR _3838_/B sky130_fd_sc_hd__and2_1
XFILLER_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5536_ hold704/X _5536_/A1 _5538_/S VGND VGND VPWR VPWR _7095_/D sky130_fd_sc_hd__mux2_1
XFILLER_105_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5467_ hold710/X _5467_/A1 _5469_/S VGND VGND VPWR VPWR _7034_/D sky130_fd_sc_hd__mux2_1
X_7206_ _7206_/CLK _7206_/D _6348_/B VGND VGND VPWR VPWR hold54/A sky130_fd_sc_hd__dfrtp_1
X_4418_ _4524_/A _4418_/B VGND VGND VPWR VPWR _4503_/C sky130_fd_sc_hd__nand2_1
X_5398_ hold204/X _5398_/A1 _5400_/S VGND VGND VPWR VPWR _6973_/D sky130_fd_sc_hd__mux2_1
Xwire2106 wire2107/X VGND VGND VPWR VPWR wire2106/X sky130_fd_sc_hd__clkbuf_1
XFILLER_99_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2117 wire2118/X VGND VGND VPWR VPWR wire2117/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2128 wire2129/X VGND VGND VPWR VPWR wire2128/X sky130_fd_sc_hd__clkbuf_1
X_7137_ _7137_/CLK _7137_/D _7137_/RESET_B VGND VGND VPWR VPWR _7137_/Q sky130_fd_sc_hd__dfrtp_1
X_4349_ _4404_/B _4350_/B _4654_/A VGND VGND VPWR VPWR _4351_/A sky130_fd_sc_hd__a21o_1
Xwire2139 _6803_/Q VGND VGND VPWR VPWR wire2139/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1405 wire1406/X VGND VGND VPWR VPWR _6308_/C1 sky130_fd_sc_hd__clkbuf_1
Xwire1416 _5927_/X VGND VGND VPWR VPWR wire1416/X sky130_fd_sc_hd__clkbuf_1
XFILLER_47_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1427 wire1428/X VGND VGND VPWR VPWR _5695_/C1 sky130_fd_sc_hd__clkbuf_1
XFILLER_100_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7068_ _7068_/CLK _7068_/D wire4007/X VGND VGND VPWR VPWR _7068_/Q sky130_fd_sc_hd__dfrtp_1
Xwire1438 _4453_/X VGND VGND VPWR VPWR _5002_/A sky130_fd_sc_hd__buf_2
Xwire1449 _3961_/X VGND VGND VPWR VPWR wire1449/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6019_ _6019_/A _6019_/B VGND VGND VPWR VPWR _6025_/C sky130_fd_sc_hd__nor2_1
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire702 _5336_/S VGND VGND VPWR VPWR _5333_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_168_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire713 _5142_/A VGND VGND VPWR VPWR _4979_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_155_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire724 wire725/X VGND VGND VPWR VPWR wire724/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire735 _4009_/S VGND VGND VPWR VPWR _4004_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire746 _3745_/X VGND VGND VPWR VPWR wire746/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire757 _3712_/X VGND VGND VPWR VPWR wire757/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire768 wire769/X VGND VGND VPWR VPWR wire768/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire779 _3560_/X VGND VGND VPWR VPWR wire779/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_551 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire4042 wire4042/A VGND VGND VPWR VPWR wire4042/X sky130_fd_sc_hd__buf_2
XFILLER_184_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3330 wire3331/X VGND VGND VPWR VPWR _4595_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_96_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4086 wire4086/A VGND VGND VPWR VPWR wire4086/X sky130_fd_sc_hd__clkbuf_2
Xwire3341 _4832_/B VGND VGND VPWR VPWR _4652_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire4097 input74/X VGND VGND VPWR VPWR _3953_/B sky130_fd_sc_hd__clkbuf_1
Xwire3363 _4710_/B2 VGND VGND VPWR VPWR _5076_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_77_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3374 _5375_/A0 VGND VGND VPWR VPWR _5501_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3385 wire3386/X VGND VGND VPWR VPWR _5411_/A0 sky130_fd_sc_hd__clkbuf_1
Xwire2640 _6141_/B1 VGND VGND VPWR VPWR _6065_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2651 _6131_/B1 VGND VGND VPWR VPWR _6056_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire2662 _6060_/B1 VGND VGND VPWR VPWR _6031_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire2673 _6020_/X VGND VGND VPWR VPWR _6025_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2684 _6175_/B1 VGND VGND VPWR VPWR _6149_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire1950 _6062_/A1 VGND VGND VPWR VPWR _3667_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_18_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1961 _6091_/B2 VGND VGND VPWR VPWR _3609_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1972 _3226_/A VGND VGND VPWR VPWR _6111_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1983 wire1983/A VGND VGND VPWR VPWR wire1983/X sky130_fd_sc_hd__clkbuf_1
Xwire1994 wire1995/X VGND VGND VPWR VPWR _6160_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_133_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3720_ _5714_/B2 wire915/X _3720_/B1 _3720_/B2 _3719_/X VGND VGND VPWR VPWR _3721_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_159_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3651_ _3651_/A _3651_/B _3651_/C _3651_/D VGND VGND VPWR VPWR _3651_/X sky130_fd_sc_hd__or4_1
XFILLER_9_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6370_ _4228_/C _6370_/A2 _6370_/B1 _4228_/Y _6369_/X VGND VGND VPWR VPWR _6370_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3582_ _3582_/A _3582_/B _3582_/C _3582_/D VGND VGND VPWR VPWR _3583_/D sky130_fd_sc_hd__or4_1
X_5321_ _5339_/A0 hold672/X _5321_/S VGND VGND VPWR VPWR _6905_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5252_ hold395/X _5450_/A0 _5253_/S VGND VGND VPWR VPWR _6843_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4203_ hold466/X _5534_/A1 _4203_/S VGND VGND VPWR VPWR _6659_/D sky130_fd_sc_hd__mux2_1
X_5183_ _5183_/A _5183_/B _5183_/C VGND VGND VPWR VPWR _5183_/X sky130_fd_sc_hd__or3_1
XFILLER_68_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4134_ hold695/X _4134_/A1 _4134_/S VGND VGND VPWR VPWR _6600_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_663 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4065_ hold174/X _4064_/X _4069_/S VGND VGND VPWR VPWR _4065_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4967_ _4794_/A _4565_/X _4688_/B _4810_/D _4887_/D VGND VGND VPWR VPWR _4969_/B
+ sky130_fd_sc_hd__o311a_1
Xmax_length4006 wire4007/X VGND VGND VPWR VPWR _7137_/RESET_B sky130_fd_sc_hd__clkbuf_2
XFILLER_51_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3918_ _6579_/Q _3918_/A1 _3918_/S VGND VGND VPWR VPWR _3918_/X sky130_fd_sc_hd__mux2_1
X_6706_ _7091_/CLK _6706_/D wire4029/X VGND VGND VPWR VPWR _6706_/Q sky130_fd_sc_hd__dfrtp_1
X_4898_ _5042_/A _4873_/Y _4875_/X _4897_/X _4992_/C VGND VGND VPWR VPWR _4928_/C
+ sky130_fd_sc_hd__o41a_1
XFILLER_137_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6637_ _6683_/CLK _6637_/D _6672_/SET_B VGND VGND VPWR VPWR _6637_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3849_ _6473_/Q _6472_/Q _6541_/Q _3848_/Y VGND VGND VPWR VPWR _3856_/B sky130_fd_sc_hd__o211a_1
XFILLER_20_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length2615 _6312_/B1 VGND VGND VPWR VPWR wire2614/A sky130_fd_sc_hd__clkbuf_1
XFILLER_137_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6568_ _7031_/CLK _6568_/D wire4044/X VGND VGND VPWR VPWR _6568_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5519_ _5519_/A0 hold584/X _5519_/S VGND VGND VPWR VPWR _7081_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6499_ _7139_/CLK _6499_/D _6499_/SET_B VGND VGND VPWR VPWR _6499_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_106_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1213 _3315_/Y VGND VGND VPWR VPWR _3596_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1224 _3666_/A2 VGND VGND VPWR VPWR _3459_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_170_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1235 wire1236/X VGND VGND VPWR VPWR _3703_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_87_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1246 _3298_/Y VGND VGND VPWR VPWR _5412_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_170_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1279 _3646_/A2 VGND VGND VPWR VPWR _3782_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire510 wire511/X VGND VGND VPWR VPWR _5273_/S sky130_fd_sc_hd__clkbuf_2
Xwire521 _5170_/B VGND VGND VPWR VPWR _5092_/C sky130_fd_sc_hd__clkbuf_1
Xwire532 _4110_/S VGND VGND VPWR VPWR wire532/X sky130_fd_sc_hd__clkbuf_1
Xwire543 wire544/X VGND VGND VPWR VPWR _3688_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire554 _3635_/X VGND VGND VPWR VPWR _3642_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_183_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire565 _3501_/X VGND VGND VPWR VPWR _3515_/A sky130_fd_sc_hd__clkbuf_1
Xwire576 _3391_/X VGND VGND VPWR VPWR wire576/X sky130_fd_sc_hd__clkbuf_1
Xwire587 _6085_/X VGND VGND VPWR VPWR wire587/X sky130_fd_sc_hd__clkbuf_1
Xwire598 wire599/X VGND VGND VPWR VPWR _5516_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_12_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3160 wire3160/A VGND VGND VPWR VPWR _6163_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire3171 _4660_/X VGND VGND VPWR VPWR _5016_/B sky130_fd_sc_hd__clkbuf_1
Xwire3182 _4620_/A VGND VGND VPWR VPWR _5108_/A sky130_fd_sc_hd__buf_2
XFILLER_77_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3193 _5013_/B VGND VGND VPWR VPWR _5076_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2470 _6082_/B1 VGND VGND VPWR VPWR _6032_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_38_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2481 _6060_/A2 VGND VGND VPWR VPWR _6032_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_93_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2492 _6160_/B1 VGND VGND VPWR VPWR _6137_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_65_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1780 _7012_/Q VGND VGND VPWR VPWR _6089_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1791 wire1792/X VGND VGND VPWR VPWR _6151_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_46_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5870_ _6229_/A1 _5944_/A2 _5930_/A2 _6227_/B2 VGND VGND VPWR VPWR _5870_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4821_ _4982_/B _4821_/B _4821_/C _4821_/D VGND VGND VPWR VPWR _4822_/B sky130_fd_sc_hd__or4_1
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4752_ _4753_/B _4752_/B VGND VGND VPWR VPWR _4986_/B sky130_fd_sc_hd__nor2_1
XFILLER_159_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3703_ _6070_/A1 _3703_/A2 _3503_/Y _6249_/B2 wire760/X VGND VGND VPWR VPWR _3710_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4683_ _4683_/A _4683_/B VGND VGND VPWR VPWR _4699_/B sky130_fd_sc_hd__or2_1
XFILLER_119_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6422_ _6438_/A _6435_/B VGND VGND VPWR VPWR _6422_/X sky130_fd_sc_hd__and2_1
XFILLER_147_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3634_ _6088_/A1 _3634_/A2 _3495_/Y _6523_/Q VGND VGND VPWR VPWR _3634_/X sky130_fd_sc_hd__a22o_1
XFILLER_134_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6353_ _7193_/Q _6353_/A1 _6353_/S VGND VGND VPWR VPWR _7193_/D sky130_fd_sc_hd__mux2_1
X_3565_ _6739_/Q wire830/X _4270_/A _6724_/Q VGND VGND VPWR VPWR _3565_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5304_ _5304_/A _5502_/B VGND VGND VPWR VPWR _5304_/Y sky130_fd_sc_hd__nand2_1
X_6284_ _6672_/Q _6284_/A2 _6284_/B1 _6284_/B2 _6283_/X VGND VGND VPWR VPWR _6291_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3496_ _3714_/B _3510_/B VGND VGND VPWR VPWR _3496_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5235_ _5352_/A0 hold449/X _5240_/S VGND VGND VPWR VPWR _6828_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5166_ _5128_/C _5163_/X _5180_/C _5160_/X VGND VGND VPWR VPWR _5166_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_29_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4117_ _5247_/A0 _6585_/Q _4119_/S VGND VGND VPWR VPWR _4117_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5097_ _4494_/Y _4783_/Y _5096_/X VGND VGND VPWR VPWR _5112_/D sky130_fd_sc_hd__a21o_1
X_4048_ _4122_/A0 hold283/X _4051_/S VGND VGND VPWR VPWR _6537_/D sky130_fd_sc_hd__mux2_1
XFILLER_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5999_ _5999_/A1 _5999_/A2 _5999_/B1 _5999_/B2 _5995_/X VGND VGND VPWR VPWR _5999_/X
+ sky130_fd_sc_hd__a221o_1
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3157 _5995_/A2 VGND VGND VPWR VPWR wire3153/A sky130_fd_sc_hd__clkbuf_1
XFILLER_137_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput290 _6481_/Q VGND VGND VPWR VPWR pll_trim[23] sky130_fd_sc_hd__buf_12
XFILLER_160_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1010 wire1011/X VGND VGND VPWR VPWR _6146_/S sky130_fd_sc_hd__clkbuf_1
Xhold9 hold9/A VGND VGND VPWR VPWR hold9/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire1021 _3932_/X VGND VGND VPWR VPWR wire1021/X sky130_fd_sc_hd__clkbuf_1
XFILLER_47_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1032 _3536_/Y VGND VGND VPWR VPWR _3774_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1065 _4022_/A VGND VGND VPWR VPWR _3656_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1087 _4040_/A VGND VGND VPWR VPWR _3771_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1098 _5221_/B VGND VGND VPWR VPWR _3776_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire351 _4713_/Y VGND VGND VPWR VPWR _4714_/B sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_62_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7081_/CLK sky130_fd_sc_hd__clkbuf_16
Xwire362 _3723_/X VGND VGND VPWR VPWR wire362/X sky130_fd_sc_hd__clkbuf_1
Xwire373 _3447_/X VGND VGND VPWR VPWR wire373/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold409 _6621_/Q VGND VGND VPWR VPWR hold409/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire384 _4961_/Y VGND VGND VPWR VPWR _4962_/B sky130_fd_sc_hd__clkbuf_1
Xwire395 wire396/X VGND VGND VPWR VPWR wire395/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3350_ _3350_/A1 _3500_/A2 wire901/X _3350_/B2 _3349_/X VGND VGND VPWR VPWR _3350_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_98_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_77_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6775_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ hold26/X _3301_/C _3297_/A VGND VGND VPWR VPWR _3281_/X sky130_fd_sc_hd__or3_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5020_ _4638_/A _4396_/X _4919_/X VGND VGND VPWR VPWR _5073_/B sky130_fd_sc_hd__o21ai_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6971_ _7046_/CLK _6971_/D wire4052/A VGND VGND VPWR VPWR _6971_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_19_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5922_ _5922_/A1 _5922_/A2 _5955_/A2 _5922_/B2 _5921_/X VGND VGND VPWR VPWR _5922_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5853_ _6209_/B2 _5853_/A2 _5853_/B1 _6937_/Q VGND VGND VPWR VPWR _5853_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_15_csclk _7059_/CLK VGND VGND VPWR VPWR _7091_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4804_ _4674_/A _4804_/A2 _4622_/Y _4746_/Y VGND VGND VPWR VPWR _4813_/C sky130_fd_sc_hd__a31o_1
X_5784_ _6123_/B2 _5784_/A2 _5784_/B1 _6966_/Q _5783_/X VGND VGND VPWR VPWR _5784_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_166_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4735_ _4735_/A _4876_/A VGND VGND VPWR VPWR _4810_/C sky130_fd_sc_hd__nand2_1
XFILLER_159_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4666_ _4689_/A _4666_/B VGND VGND VPWR VPWR _4666_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6405_ _6405_/A _6407_/B VGND VGND VPWR VPWR _6405_/X sky130_fd_sc_hd__and2_1
XFILLER_135_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3617_ _6988_/Q _3617_/A2 _3617_/B1 _6278_/A1 VGND VGND VPWR VPWR _3658_/B sky130_fd_sc_hd__a22o_1
XFILLER_134_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4597_ _4569_/B _5089_/B2 _4659_/B VGND VGND VPWR VPWR _4598_/D sky130_fd_sc_hd__a21oi_1
XFILLER_134_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6336_ _6705_/Q _6336_/A2 _6272_/B _6336_/B2 _6335_/X VGND VGND VPWR VPWR _6341_/C
+ sky130_fd_sc_hd__a221o_1
X_3548_ _6104_/A1 _3548_/A2 _3548_/B1 _6113_/A1 VGND VGND VPWR VPWR _3548_/X sky130_fd_sc_hd__a22o_1
Xwire3907 wire3908/X VGND VGND VPWR VPWR wire3907/X sky130_fd_sc_hd__clkbuf_1
Xwire3918 wire3919/X VGND VGND VPWR VPWR _3945_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3929 wire3930/X VGND VGND VPWR VPWR wire3929/X sky130_fd_sc_hd__clkbuf_1
XFILLER_142_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6267_ _6267_/A _6267_/B _6267_/C VGND VGND VPWR VPWR _6267_/X sky130_fd_sc_hd__or3_1
X_3479_ _6340_/A1 _3567_/B1 _4246_/A _6705_/Q VGND VGND VPWR VPWR _3479_/X sky130_fd_sc_hd__a22o_1
XFILLER_95_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5218_ _5454_/A0 hold523/X _5220_/S VGND VGND VPWR VPWR _6816_/D sky130_fd_sc_hd__mux2_1
XFILLER_103_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6198_ _6198_/A1 _6198_/A2 _6198_/B1 _6198_/B2 VGND VGND VPWR VPWR _6198_/X sky130_fd_sc_hd__a22o_1
XFILLER_57_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5149_ _4451_/B _4446_/Y _4843_/A _4894_/A _5009_/A VGND VGND VPWR VPWR _5151_/C
+ sky130_fd_sc_hd__a2111o_1
XFILLER_28_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_690 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length2286 hold492/X VGND VGND VPWR VPWR _5908_/B2 sky130_fd_sc_hd__clkbuf_1
Xmax_length1574 hold200/X VGND VGND VPWR VPWR _5548_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_106_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length1596 _7092_/Q VGND VGND VPWR VPWR _5914_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_69_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4520_ _4520_/A _4520_/B VGND VGND VPWR VPWR _4520_/X sky130_fd_sc_hd__or2_1
XFILLER_156_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold206 _7048_/Q VGND VGND VPWR VPWR hold206/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4451_ _4451_/A _4451_/B VGND VGND VPWR VPWR _4942_/A sky130_fd_sc_hd__nand2_2
XFILLER_156_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold217 _6835_/Q VGND VGND VPWR VPWR hold217/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 _6837_/Q VGND VGND VPWR VPWR hold228/X sky130_fd_sc_hd__dlygate4sd3_1
X_3402_ _6194_/A1 _5250_/A wire940/X _3402_/B2 _3401_/X VGND VGND VPWR VPWR _3408_/A
+ sky130_fd_sc_hd__a221o_1
Xhold239 _6607_/Q VGND VGND VPWR VPWR hold239/X sky130_fd_sc_hd__dlygate4sd3_1
X_7170_ _7185_/CLK _7170_/D fanout3952/X VGND VGND VPWR VPWR _7170_/Q sky130_fd_sc_hd__dfrtp_1
X_4382_ _4492_/A _4719_/A VGND VGND VPWR VPWR _4952_/A sky130_fd_sc_hd__nor2_1
XFILLER_171_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6121_ _6121_/A1 _7177_/Q wire452/X VGND VGND VPWR VPWR _6121_/X sky130_fd_sc_hd__a21o_1
XFILLER_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ _5241_/A _5241_/B VGND VGND VPWR VPWR _3333_/Y sky130_fd_sc_hd__nor2_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6052_ _7075_/Q _6052_/A2 _6052_/B1 _6052_/B2 _6051_/X VGND VGND VPWR VPWR _6058_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3264_ hold81/X _3832_/A1 _3820_/A VGND VGND VPWR VPWR hold82/A sky130_fd_sc_hd__mux2_1
XFILLER_39_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5003_ _5003_/A _5003_/B VGND VGND VPWR VPWR _5008_/C sky130_fd_sc_hd__nor2_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3195_ _5593_/B VGND VGND VPWR VPWR _3195_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_66_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6954_ _7111_/CLK _6954_/D fanout4027/X VGND VGND VPWR VPWR _6954_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_81_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5905_ _6667_/Q _5905_/A2 _5964_/B1 _6523_/Q VGND VGND VPWR VPWR _5905_/X sky130_fd_sc_hd__a22o_1
X_6885_ _7140_/CLK _6885_/D _7138_/RESET_B VGND VGND VPWR VPWR _6885_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_62_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5836_ _6848_/Q _5836_/A2 _5825_/X _5835_/X _5858_/C1 VGND VGND VPWR VPWR _5836_/X
+ sky130_fd_sc_hd__o221a_1
X_5767_ _5767_/A1 _5805_/A2 _5806_/A2 _6106_/A1 _5755_/X VGND VGND VPWR VPWR _5770_/C
+ sky130_fd_sc_hd__a221o_1
X_4718_ _4745_/A _4718_/B VGND VGND VPWR VPWR _4899_/B sky130_fd_sc_hd__nor2_1
XFILLER_147_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5698_ _5698_/A1 _5698_/A2 _5698_/B1 _5999_/A1 VGND VGND VPWR VPWR _5698_/X sky130_fd_sc_hd__a22o_1
XFILLER_30_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4649_ _4719_/A _4685_/A2 _4228_/Y VGND VGND VPWR VPWR _5031_/A sky130_fd_sc_hd__o21ai_1
XFILLER_162_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3704 wire3704/A VGND VGND VPWR VPWR wire3704/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3715 wire3715/A VGND VGND VPWR VPWR wire3715/X sky130_fd_sc_hd__clkbuf_2
Xwire3726 _6782_/Q VGND VGND VPWR VPWR wire3726/X sky130_fd_sc_hd__clkbuf_1
X_6319_ _7186_/Q _6318_/X _6319_/S VGND VGND VPWR VPWR _7186_/D sky130_fd_sc_hd__mux2_1
Xwire3737 _4929_/A1 VGND VGND VPWR VPWR wire3737/X sky130_fd_sc_hd__clkbuf_1
XFILLER_115_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3748 wire3749/X VGND VGND VPWR VPWR wire3748/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_606 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3951_ _3951_/A0 _3951_/A1 _3951_/S VGND VGND VPWR VPWR _3951_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6670_ _6671_/CLK _6670_/D fanout4028/X VGND VGND VPWR VPWR _6670_/Q sky130_fd_sc_hd__dfrtp_1
X_3882_ _4390_/A _4654_/A VGND VGND VPWR VPWR _4467_/A sky130_fd_sc_hd__and2_1
XFILLER_149_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5621_ _7151_/Q _7150_/Q VGND VGND VPWR VPWR _5703_/B sky130_fd_sc_hd__nor2_2
XFILLER_164_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5552_ _5552_/A0 hold665/X _5552_/S VGND VGND VPWR VPWR _7110_/D sky130_fd_sc_hd__mux2_1
XFILLER_191_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4503_ _4502_/X _4887_/C _4503_/C _4503_/D VGND VGND VPWR VPWR _4503_/X sky130_fd_sc_hd__and4b_1
XFILLER_145_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5483_ _5588_/A0 _5483_/A1 _5483_/S VGND VGND VPWR VPWR _7049_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4434_ _4453_/A _4434_/B _4444_/B _4724_/A VGND VGND VPWR VPWR _4434_/X sky130_fd_sc_hd__or4_1
XFILLER_6_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7153_ _7180_/CLK _7153_/D wire3991/X VGND VGND VPWR VPWR _7153_/Q sky130_fd_sc_hd__dfstp_1
X_4365_ _4846_/A _4538_/A VGND VGND VPWR VPWR _4369_/B sky130_fd_sc_hd__nand2b_2
XFILLER_160_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6104_ _6104_/A1 _6104_/A2 _6104_/B1 _6104_/B2 _6103_/X VGND VGND VPWR VPWR _6109_/B
+ sky130_fd_sc_hd__a221o_1
X_3316_ _3316_/A _3465_/B VGND VGND VPWR VPWR _3316_/Y sky130_fd_sc_hd__nor2_1
XFILLER_86_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7084_ _7084_/CLK _7084_/D _7035_/SET_B VGND VGND VPWR VPWR _7084_/Q sky130_fd_sc_hd__dfrtp_1
X_4296_ _4308_/A0 hold272/X _4299_/S VGND VGND VPWR VPWR _4296_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1609 _6076_/A1 VGND VGND VPWR VPWR _5748_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_100_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6035_ _6035_/A1 _6082_/A2 _6062_/B1 _6035_/B2 _6034_/X VGND VGND VPWR VPWR _6044_/C
+ sky130_fd_sc_hd__a221o_1
X_3247_ _3941_/A hold159/X hold61/X VGND VGND VPWR VPWR hold62/A sky130_fd_sc_hd__o21bai_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_606 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6937_ _7125_/CLK _6937_/D wire4046/X VGND VGND VPWR VPWR _6937_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6868_ _7129_/CLK _6868_/D wire4056/A VGND VGND VPWR VPWR _6868_/Q sky130_fd_sc_hd__dfrtp_1
X_5819_ _6188_/A1 _5659_/X _5819_/B1 _6176_/B2 VGND VGND VPWR VPWR _5819_/X sky130_fd_sc_hd__a22o_1
Xwire906 wire907/X VGND VGND VPWR VPWR _4100_/S sky130_fd_sc_hd__buf_2
Xwire917 wire917/A VGND VGND VPWR VPWR wire917/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6799_ _6799_/CLK _6799_/D wire3935/A VGND VGND VPWR VPWR _6799_/Q sky130_fd_sc_hd__dfstp_1
Xwire928 wire929/X VGND VGND VPWR VPWR wire928/X sky130_fd_sc_hd__clkbuf_1
XFILLER_182_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire939 wire939/A VGND VGND VPWR VPWR _4068_/S sky130_fd_sc_hd__buf_2
Xmax_length515 _5268_/Y VGND VGND VPWR VPWR _5275_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length526 _4164_/S VGND VGND VPWR VPWR _4162_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_6_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length537 _4052_/X VGND VGND VPWR VPWR wire536/A sky130_fd_sc_hd__clkbuf_1
XFILLER_41_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4202 wire4203/X VGND VGND VPWR VPWR _3696_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire4213 _3540_/B2 VGND VGND VPWR VPWR wire4213/X sky130_fd_sc_hd__clkbuf_1
Xwire4224 wire4225/X VGND VGND VPWR VPWR _3629_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_150_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4235 input33/X VGND VGND VPWR VPWR _3349_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire4246 input22/X VGND VGND VPWR VPWR _3636_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire3501 _4214_/A1 VGND VGND VPWR VPWR _4250_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold570 _6491_/Q VGND VGND VPWR VPWR hold570/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3523 wire3523/A VGND VGND VPWR VPWR _5362_/A0 sky130_fd_sc_hd__clkbuf_1
Xwire4268 wire4269/X VGND VGND VPWR VPWR wire4268/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold581 _6897_/Q VGND VGND VPWR VPWR hold581/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_173_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4279 input13/X VGND VGND VPWR VPWR _3647_/A1 sky130_fd_sc_hd__clkbuf_1
Xhold592 _6605_/Q VGND VGND VPWR VPWR hold592/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3545 _4237_/A0 VGND VGND VPWR VPWR _4249_/A0 sky130_fd_sc_hd__clkbuf_2
Xwire2811 _6024_/A VGND VGND VPWR VPWR wire2811/X sky130_fd_sc_hd__clkbuf_1
Xwire3567 hold22/X VGND VGND VPWR VPWR _5406_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3578 _4122_/A0 VGND VGND VPWR VPWR _5195_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2833 wire2834/X VGND VGND VPWR VPWR _5855_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_104_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2844 _5841_/B1 VGND VGND VPWR VPWR _5832_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire2855 _5830_/B1 VGND VGND VPWR VPWR _5754_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2877 _5700_/X VGND VGND VPWR VPWR _5849_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2888 _5698_/B1 VGND VGND VPWR VPWR _5932_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire2899 _5698_/A2 VGND VGND VPWR VPWR _5934_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_64_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout3940 wire3945/A VGND VGND VPWR VPWR wire3943/A sky130_fd_sc_hd__clkbuf_1
XFILLER_142_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout3973 wire3985/A VGND VGND VPWR VPWR fanout3973/X sky130_fd_sc_hd__buf_6
X_4150_ _4237_/A0 hold297/X _4152_/S VGND VGND VPWR VPWR _6613_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4081_ hold512/X _5508_/A0 _4085_/S VGND VGND VPWR VPWR _4081_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4983_ _4983_/A _4983_/B _4983_/C VGND VGND VPWR VPWR _4983_/Y sky130_fd_sc_hd__nor3_1
XFILLER_23_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6722_ _6979_/CLK _6722_/D fanout4027/X VGND VGND VPWR VPWR _6722_/Q sky130_fd_sc_hd__dfrtp_1
X_3934_ _3232_/Y _3934_/A1 _3934_/S VGND VGND VPWR VPWR _3934_/X sky130_fd_sc_hd__mux2_1
XFILLER_189_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3865_ hold35/A _6447_/Q _3866_/S VGND VGND VPWR VPWR _6447_/D sky130_fd_sc_hd__mux2_1
X_6653_ _7206_/CLK _6653_/D VGND VGND VPWR VPWR _6653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5604_ _7144_/Q _7145_/Q _7146_/Q _5604_/D VGND VGND VPWR VPWR _5605_/A sky130_fd_sc_hd__and4_1
XFILLER_177_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6584_ _7129_/CLK _6584_/D wire4055/X VGND VGND VPWR VPWR hold74/A sky130_fd_sc_hd__dfrtp_1
X_3796_ _6472_/Q _6471_/Q _3801_/B VGND VGND VPWR VPWR _3800_/A sky130_fd_sc_hd__and3_1
XFILLER_191_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5535_ _5535_/A _5535_/B VGND VGND VPWR VPWR _5542_/S sky130_fd_sc_hd__and2_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5466_ _5466_/A _5535_/B VGND VGND VPWR VPWR _5474_/S sky130_fd_sc_hd__and2_1
XFILLER_145_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7205_ _7206_/CLK _7205_/D _4189_/B VGND VGND VPWR VPWR _7205_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4417_ _4742_/B _5001_/A _4758_/B VGND VGND VPWR VPWR _4417_/X sky130_fd_sc_hd__and3_1
XFILLER_132_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5397_ hold161/X _5547_/A0 _5397_/S VGND VGND VPWR VPWR _6972_/D sky130_fd_sc_hd__mux2_1
Xwire2107 wire2108/X VGND VGND VPWR VPWR wire2107/X sky130_fd_sc_hd__clkbuf_1
X_4348_ _4348_/A _4348_/B _4348_/C VGND VGND VPWR VPWR _4542_/A sky130_fd_sc_hd__and3_1
Xwire2118 _6812_/Q VGND VGND VPWR VPWR wire2118/X sky130_fd_sc_hd__clkbuf_1
X_7136_ _7136_/CLK _7136_/D wire4042/X VGND VGND VPWR VPWR _7136_/Q sky130_fd_sc_hd__dfstp_1
Xwire2129 _6808_/Q VGND VGND VPWR VPWR wire2129/X sky130_fd_sc_hd__clkbuf_1
XFILLER_59_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1406 _6296_/X VGND VGND VPWR VPWR wire1406/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1417 _5828_/X VGND VGND VPWR VPWR _5829_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_98_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7067_ _7067_/CLK _7067_/D wire3968/X VGND VGND VPWR VPWR _7067_/Q sky130_fd_sc_hd__dfstp_1
X_4279_ _4279_/A0 _6728_/Q _4281_/S VGND VGND VPWR VPWR _4279_/X sky130_fd_sc_hd__mux2_1
Xwire1428 _5692_/X VGND VGND VPWR VPWR wire1428/X sky130_fd_sc_hd__clkbuf_1
Xwire1439 _5113_/A1 VGND VGND VPWR VPWR _4995_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6018_ _6018_/A _6021_/A VGND VGND VPWR VPWR _6018_/Y sky130_fd_sc_hd__nor2_1
XFILLER_39_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire703 wire703/A VGND VGND VPWR VPWR _5336_/S sky130_fd_sc_hd__clkbuf_2
Xwire714 _4857_/X VGND VGND VPWR VPWR wire714/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire725 _4120_/X VGND VGND VPWR VPWR wire725/X sky130_fd_sc_hd__clkbuf_1
XFILLER_168_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire736 _3991_/S VGND VGND VPWR VPWR _3988_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_155_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire747 _3743_/X VGND VGND VPWR VPWR wire747/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire758 wire759/X VGND VGND VPWR VPWR wire758/X sky130_fd_sc_hd__clkbuf_1
Xwire769 _3675_/X VGND VGND VPWR VPWR wire769/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4021 wire4022/X VGND VGND VPWR VPWR wire4021/X sky130_fd_sc_hd__clkbuf_1
XFILLER_151_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout3247 _4246_/B VGND VGND VPWR VPWR _4135_/B sky130_fd_sc_hd__buf_6
XFILLER_124_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout3258 hold56/X VGND VGND VPWR VPWR _4159_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_97_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3320 _4814_/C VGND VGND VPWR VPWR _4704_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_151_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4065 wire4066/X VGND VGND VPWR VPWR wire4065/X sky130_fd_sc_hd__buf_2
Xwire3331 _4544_/X VGND VGND VPWR VPWR wire3331/X sky130_fd_sc_hd__clkbuf_1
Xfanout3269 wire3280/X VGND VGND VPWR VPWR _5225_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_151_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4098 wire4099/X VGND VGND VPWR VPWR _3751_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_104_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3364 _4461_/A VGND VGND VPWR VPWR _4710_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire3375 _5579_/A0 VGND VGND VPWR VPWR _5375_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2630 _6053_/B1 VGND VGND VPWR VPWR _6042_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire3386 wire3387/X VGND VGND VPWR VPWR wire3386/X sky130_fd_sc_hd__clkbuf_1
Xwire2652 _6154_/B1 VGND VGND VPWR VPWR _6131_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3397 _5587_/A0 VGND VGND VPWR VPWR _5509_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2663 _6086_/B1 VGND VGND VPWR VPWR _6060_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire2674 _6166_/B1 VGND VGND VPWR VPWR _6078_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1940 _6926_/Q VGND VGND VPWR VPWR _6137_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2685 _6198_/B1 VGND VGND VPWR VPWR _6175_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire1951 _6923_/Q VGND VGND VPWR VPWR _6062_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire2696 wire2697/X VGND VGND VPWR VPWR _6210_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire1973 wire1973/A VGND VGND VPWR VPWR _3226_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_93_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1995 _6895_/Q VGND VGND VPWR VPWR wire1995/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3650_ _7076_/Q _3736_/A2 _3650_/B1 _6484_/Q _3649_/X VGND VGND VPWR VPWR _3651_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3581_ _6118_/A1 _3581_/A2 wire849/X _3581_/B2 wire558/X VGND VGND VPWR VPWR _3582_/D
+ sky130_fd_sc_hd__a221o_1
X_5320_ _5392_/A0 hold460/X _5320_/S VGND VGND VPWR VPWR _6904_/D sky130_fd_sc_hd__mux2_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length890 _5562_/A VGND VGND VPWR VPWR _3566_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_115_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5251_ hold583/X _5251_/A1 _5254_/S VGND VGND VPWR VPWR _6842_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4202_ hold465/X _4214_/A1 _4203_/S VGND VGND VPWR VPWR _6658_/D sky130_fd_sc_hd__mux2_1
X_5182_ _5182_/A1 _5182_/A2 _5156_/Y _5178_/X _5181_/Y VGND VGND VPWR VPWR _5183_/C
+ sky130_fd_sc_hd__a221o_1
X_4133_ hold692/X _4208_/A1 _4134_/S VGND VGND VPWR VPWR _6599_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4064_ _6585_/Q _5247_/A0 _4068_/S VGND VGND VPWR VPWR _4064_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4966_ _4567_/X _4673_/A _4758_/Y _4786_/Y VGND VGND VPWR VPWR _4969_/A sky130_fd_sc_hd__o211a_1
XFILLER_51_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6705_ _6705_/CLK _6705_/D wire3958/X VGND VGND VPWR VPWR _6705_/Q sky130_fd_sc_hd__dfrtp_1
X_3917_ _3917_/A _3917_/B VGND VGND VPWR VPWR _6443_/D sky130_fd_sc_hd__and2_1
X_4897_ _4897_/A _4897_/B _4897_/C _4530_/B VGND VGND VPWR VPWR _4897_/X sky130_fd_sc_hd__or4b_1
XFILLER_192_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6636_ _6671_/CLK _6636_/D fanout4028/X VGND VGND VPWR VPWR _6636_/Q sky130_fd_sc_hd__dfstp_1
X_3848_ _6472_/Q _6471_/Q _6473_/Q VGND VGND VPWR VPWR _3848_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_137_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6567_ _6945_/CLK _6567_/D fanout4078/X VGND VGND VPWR VPWR _6567_/Q sky130_fd_sc_hd__dfrtp_1
X_3779_ _7082_/Q _3779_/A2 _5403_/A _6978_/Q VGND VGND VPWR VPWR _3779_/X sky130_fd_sc_hd__a22o_1
XFILLER_192_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5518_ _5518_/A0 hold575/X _5519_/S VGND VGND VPWR VPWR _7080_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6498_ _7076_/CLK _6498_/D wire3981/X VGND VGND VPWR VPWR _6498_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_145_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5449_ _5467_/A1 hold709/X _5453_/S VGND VGND VPWR VPWR _7018_/D sky130_fd_sc_hd__mux2_1
XFILLER_120_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1203 _3625_/A2 VGND VGND VPWR VPWR _3733_/A2 sky130_fd_sc_hd__clkbuf_1
X_7119_ _7136_/CLK _7119_/D wire4086/X VGND VGND VPWR VPWR _7119_/Q sky130_fd_sc_hd__dfstp_1
Xwire1214 _3314_/Y VGND VGND VPWR VPWR _3992_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1225 _3666_/A2 VGND VGND VPWR VPWR _5367_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1236 _3302_/Y VGND VGND VPWR VPWR wire1236/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1247 wire1248/X VGND VGND VPWR VPWR _3663_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_74_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1258 _3522_/A2 VGND VGND VPWR VPWR _5520_/A sky130_fd_sc_hd__clkbuf_2
Xwire1269 wire1271/A VGND VGND VPWR VPWR _3399_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_101_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_wbbd_sck clkbuf_0_wbbd_sck/X VGND VGND VPWR VPWR _6387_/A1 sky130_fd_sc_hd__clkbuf_16
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire500 _5304_/Y VGND VGND VPWR VPWR wire500/X sky130_fd_sc_hd__clkbuf_1
XFILLER_168_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire511 _5269_/S VGND VGND VPWR VPWR wire511/X sky130_fd_sc_hd__clkbuf_1
Xwire522 _5068_/X VGND VGND VPWR VPWR _5160_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire533 _4109_/S VGND VGND VPWR VPWR _4110_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire544 _3687_/X VGND VGND VPWR VPWR wire544/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3851 _4793_/A VGND VGND VPWR VPWR _4436_/A sky130_fd_sc_hd__clkbuf_2
Xwire555 _3606_/X VGND VGND VPWR VPWR wire555/X sky130_fd_sc_hd__clkbuf_1
XFILLER_156_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire566 wire567/X VGND VGND VPWR VPWR wire566/X sky130_fd_sc_hd__clkbuf_1
Xwire577 _3390_/X VGND VGND VPWR VPWR _3392_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_171_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire588 _5792_/X VGND VGND VPWR VPWR wire588/X sky130_fd_sc_hd__clkbuf_1
Xwire599 wire600/X VGND VGND VPWR VPWR wire599/X sky130_fd_sc_hd__clkbuf_1
XFILLER_171_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3172 _4660_/X VGND VGND VPWR VPWR _5164_/A3 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3183 _4587_/B VGND VGND VPWR VPWR _5152_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire3194 _4976_/A1 VGND VGND VPWR VPWR _5013_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2460 _6328_/B1 VGND VGND VPWR VPWR _6256_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_93_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2471 _6139_/B1 VGND VGND VPWR VPWR _6082_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2482 _6209_/A2 VGND VGND VPWR VPWR _6060_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire2493 wire2493/A VGND VGND VPWR VPWR _6160_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire1770 hold112/X VGND VGND VPWR VPWR _5447_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire1781 _5723_/A1 VGND VGND VPWR VPWR _6052_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1792 _3441_/B2 VGND VGND VPWR VPWR wire1792/X sky130_fd_sc_hd__clkbuf_1
XFILLER_93_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4820_ _4553_/A _4819_/C _4819_/D _4797_/A _4607_/X VGND VGND VPWR VPWR _4821_/D
+ sky130_fd_sc_hd__a41o_1
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751_ _4994_/A _4754_/B VGND VGND VPWR VPWR _4987_/B sky130_fd_sc_hd__nor2_1
XFILLER_193_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3702_ _6491_/Q _3314_/Y _4040_/A _6532_/Q VGND VGND VPWR VPWR _3702_/X sky130_fd_sc_hd__a22o_1
XFILLER_147_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4682_ _4677_/A _4660_/B _4581_/X VGND VGND VPWR VPWR _4699_/A sky130_fd_sc_hd__a21o_1
XFILLER_119_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6421_ _6438_/A _6440_/B VGND VGND VPWR VPWR _6421_/X sky130_fd_sc_hd__and2_1
X_3633_ _3633_/A _3633_/B _3633_/C _3633_/D VGND VGND VPWR VPWR _3633_/X sky130_fd_sc_hd__or4_1
XFILLER_174_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6352_ _7192_/Q wire366/X _6353_/S VGND VGND VPWR VPWR _7192_/D sky130_fd_sc_hd__mux2_1
X_3564_ _6115_/B2 _3564_/A2 _3562_/X wire432/X VGND VGND VPWR VPWR _3583_/B sky130_fd_sc_hd__a211o_1
XFILLER_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5303_ _5579_/A0 hold215/X _5303_/S VGND VGND VPWR VPWR _6889_/D sky130_fd_sc_hd__mux2_1
XFILLER_170_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6283_ _6667_/Q _6283_/A2 _6325_/B1 _6683_/Q VGND VGND VPWR VPWR _6283_/X sky130_fd_sc_hd__a22o_1
X_3495_ _3536_/A _3528_/B VGND VGND VPWR VPWR _3495_/Y sky130_fd_sc_hd__nor2_1
XFILLER_88_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5234_ _5234_/A0 _6827_/Q _5240_/S VGND VGND VPWR VPWR hold39/A sky130_fd_sc_hd__mux2_1
XFILLER_88_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5165_ _4502_/A _5067_/A _5165_/C _5165_/D VGND VGND VPWR VPWR _5180_/C sky130_fd_sc_hd__and4bb_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4116_ _4116_/A0 hold74/X _4119_/S VGND VGND VPWR VPWR _6584_/D sky130_fd_sc_hd__mux2_1
XFILLER_69_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5096_ _4372_/Y _4494_/Y _4749_/B _4778_/B VGND VGND VPWR VPWR _5096_/X sky130_fd_sc_hd__o31a_1
XFILLER_96_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4047_ _5530_/A1 hold274/X _4051_/S VGND VGND VPWR VPWR _6536_/D sky130_fd_sc_hd__mux2_1
XFILLER_37_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5998_ _6038_/A _6021_/B VGND VGND VPWR VPWR _5998_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4949_ _4932_/A _4933_/A _4944_/B _4932_/B _4837_/X VGND VGND VPWR VPWR _4950_/C
+ sky130_fd_sc_hd__o41a_1
XFILLER_138_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6619_ _7112_/CLK _6619_/D wire4026/X VGND VGND VPWR VPWR _6619_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_193_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length2446 _6488_/Q VGND VGND VPWR VPWR wire2444/A sky130_fd_sc_hd__clkbuf_1
XFILLER_137_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length2479 _6282_/A2 VGND VGND VPWR VPWR wire2478/A sky130_fd_sc_hd__clkbuf_1
XFILLER_106_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput280 wire2445/X VGND VGND VPWR VPWR pll_trim[14] sky130_fd_sc_hd__buf_12
XFILLER_121_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput291 _6804_/Q VGND VGND VPWR VPWR pll_trim[24] sky130_fd_sc_hd__buf_12
Xwire1000 _5681_/X VGND VGND VPWR VPWR wire999/A sky130_fd_sc_hd__clkbuf_1
Xwire1011 _5651_/Y VGND VGND VPWR VPWR wire1011/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1022 _3731_/Y VGND VGND VPWR VPWR _5210_/A sky130_fd_sc_hd__clkbuf_1
Xwire1033 _3617_/B1 VGND VGND VPWR VPWR _3665_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_59_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1044 _3511_/Y VGND VGND VPWR VPWR _4252_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1055 _3766_/B1 VGND VGND VPWR VPWR _3493_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_47_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1066 _4246_/A VGND VGND VPWR VPWR _3676_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1077 _3465_/Y VGND VGND VPWR VPWR _3574_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1088 _3454_/Y VGND VGND VPWR VPWR _3672_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_114_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1099 _3403_/B1 VGND VGND VPWR VPWR _3432_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_90_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire352 _5183_/X VGND VGND VPWR VPWR _6782_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire363 wire364/X VGND VGND VPWR VPWR wire363/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire374 wire375/X VGND VGND VPWR VPWR wire374/X sky130_fd_sc_hd__clkbuf_2
XFILLER_156_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire385 _3765_/X VGND VGND VPWR VPWR _3790_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_183_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire396 _3760_/X VGND VGND VPWR VPWR wire396/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3280_ _3320_/A _3528_/A VGND VGND VPWR VPWR _3280_/Y sky130_fd_sc_hd__nor2_1
XFILLER_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2290 _6658_/Q VGND VGND VPWR VPWR _6300_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6970_ _7046_/CLK _6970_/D wire4052/A VGND VGND VPWR VPWR _6970_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5921_ _6763_/Q _5921_/A2 _5921_/B1 _5921_/B2 VGND VGND VPWR VPWR _5921_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5852_ _6205_/B2 _5852_/A2 _5852_/B1 _6905_/Q _5851_/X VGND VGND VPWR VPWR _5857_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4803_ _4662_/B _4804_/A2 _4592_/Y _5049_/B VGND VGND VPWR VPWR _4817_/B sky130_fd_sc_hd__a31o_1
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5783_ _6974_/Q _5783_/A2 _5783_/B1 _6124_/A1 _5783_/C1 VGND VGND VPWR VPWR _5783_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4734_ _4872_/A _4734_/B VGND VGND VPWR VPWR _4734_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4665_ _5021_/C _4665_/B VGND VGND VPWR VPWR _4665_/Y sky130_fd_sc_hd__nor2_1
XFILLER_135_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6404_ _6404_/A _6407_/B VGND VGND VPWR VPWR _6404_/X sky130_fd_sc_hd__and2_1
X_3616_ _3616_/A1 wire887/X wire867/X _3616_/B2 VGND VGND VPWR VPWR _3616_/X sky130_fd_sc_hd__a22o_1
X_4596_ _4596_/A _4596_/B VGND VGND VPWR VPWR _5021_/B sky130_fd_sc_hd__or2_2
XFILLER_134_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6335_ _6335_/A1 _6335_/A2 _6335_/B1 _6615_/Q VGND VGND VPWR VPWR _6335_/X sky130_fd_sc_hd__a22o_1
XFILLER_89_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3547_ _5212_/B _3714_/B VGND VGND VPWR VPWR _3547_/Y sky130_fd_sc_hd__nor2_2
XFILLER_89_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3908 input86/X VGND VGND VPWR VPWR wire3908/X sky130_fd_sc_hd__clkbuf_1
Xwire3919 wire3920/X VGND VGND VPWR VPWR wire3919/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3478_ hold63/X _3478_/B VGND VGND VPWR VPWR _4246_/A sky130_fd_sc_hd__nor2_1
X_6266_ _6266_/A _6266_/B _6266_/C _6266_/D VGND VGND VPWR VPWR _6267_/C sky130_fd_sc_hd__or4_1
XFILLER_142_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5217_ _5451_/A0 hold517/X _5220_/S VGND VGND VPWR VPWR _6815_/D sky130_fd_sc_hd__mux2_1
XFILLER_130_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6197_ _6197_/A1 _6197_/A2 _6197_/B1 _6197_/B2 VGND VGND VPWR VPWR _6197_/X sky130_fd_sc_hd__a22o_1
XFILLER_28_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5148_ _5148_/A _5148_/B _5148_/C _5148_/D VGND VGND VPWR VPWR _5148_/Y sky130_fd_sc_hd__nor4_2
XFILLER_28_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5079_ _5079_/A _5079_/B VGND VGND VPWR VPWR _5106_/C sky130_fd_sc_hd__or2_1
XFILLER_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length2265 hold147/X VGND VGND VPWR VPWR _4225_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_69_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4450_ _4450_/A _5035_/A VGND VGND VPWR VPWR _4450_/Y sky130_fd_sc_hd__nor2_1
Xhold207 _6883_/Q VGND VGND VPWR VPWR hold207/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 _6702_/Q VGND VGND VPWR VPWR hold218/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold229 _7075_/Q VGND VGND VPWR VPWR hold229/X sky130_fd_sc_hd__dlygate4sd3_1
X_3401_ _6188_/B2 _3401_/A2 wire864/X _6184_/B2 VGND VGND VPWR VPWR _3401_/X sky130_fd_sc_hd__a22o_1
X_4381_ _4657_/A _4667_/B VGND VGND VPWR VPWR _4719_/A sky130_fd_sc_hd__nand2_1
XFILLER_125_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3332_ _3339_/B _3507_/B VGND VGND VPWR VPWR _3332_/Y sky130_fd_sc_hd__nor2_1
X_6120_ _6120_/A1 wire981/X wire586/X _6119_/X _6120_/C1 VGND VGND VPWR VPWR _6120_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_124_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ hold115/X _3263_/A1 _3265_/S VGND VGND VPWR VPWR _3284_/A sky130_fd_sc_hd__mux2_1
X_6051_ _6051_/A1 _6051_/A2 _6073_/B1 _7120_/Q VGND VGND VPWR VPWR _6051_/X sky130_fd_sc_hd__a22o_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _5002_/A _5036_/B VGND VGND VPWR VPWR _5049_/D sky130_fd_sc_hd__nor2_1
X_3194_ _6565_/Q VGND VGND VPWR VPWR _5648_/C sky130_fd_sc_hd__inv_2
XFILLER_39_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6953_ _7133_/CLK _6953_/D _7087_/RESET_B VGND VGND VPWR VPWR _6953_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5904_ _7171_/Q _5903_/X _5948_/S VGND VGND VPWR VPWR _7171_/D sky130_fd_sc_hd__mux2_1
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6884_ _7084_/CLK _6884_/D _7035_/SET_B VGND VGND VPWR VPWR _6884_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5835_ _5835_/A _5835_/B _5835_/C _5835_/D VGND VGND VPWR VPWR _5835_/X sky130_fd_sc_hd__or4_1
XFILLER_179_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5766_ _5766_/A1 _5805_/B1 _5779_/B1 _5766_/B2 _5765_/X VGND VGND VPWR VPWR _5770_/B
+ sky130_fd_sc_hd__a221o_1
Xmax_length708 _5254_/S VGND VGND VPWR VPWR _5255_/S sky130_fd_sc_hd__clkbuf_1
X_4717_ _4745_/A _4717_/B VGND VGND VPWR VPWR _5050_/B sky130_fd_sc_hd__or2_1
XFILLER_147_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5697_ _7152_/Q _5703_/B _5699_/B VGND VGND VPWR VPWR _5697_/X sky130_fd_sc_hd__and3_1
XFILLER_163_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4648_ _4963_/A _4648_/B VGND VGND VPWR VPWR _4648_/Y sky130_fd_sc_hd__nor2_1
XFILLER_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4579_ _4693_/A _4632_/A VGND VGND VPWR VPWR _4639_/A sky130_fd_sc_hd__or2_1
X_6318_ _7185_/Q wire443/X _6318_/S VGND VGND VPWR VPWR _6318_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3727 hold723/X VGND VGND VPWR VPWR _3254_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire3738 _6777_/Q VGND VGND VPWR VPWR _4929_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3749 _6699_/Q VGND VGND VPWR VPWR wire3749/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6249_ _6249_/A1 _6289_/A2 _6325_/A2 _6249_/B2 VGND VGND VPWR VPWR _6249_/X sky130_fd_sc_hd__a22o_1
XFILLER_39_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_61_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _6989_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_76_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6761_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length1383 _3301_/X VGND VGND VPWR VPWR wire1379/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_14_csclk _7059_/CLK VGND VGND VPWR VPWR _7208_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_122_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_29_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7075_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold90 hold90/A VGND VGND VPWR VPWR hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_36_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3950_ _3950_/A VGND VGND VPWR VPWR _3950_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3881_ _4338_/C _4338_/D _4337_/A _4337_/B VGND VGND VPWR VPWR _3887_/C sky130_fd_sc_hd__or4_1
XFILLER_149_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5620_ _7150_/Q _5618_/B _5624_/B _5619_/Y VGND VGND VPWR VPWR _7150_/D sky130_fd_sc_hd__a31o_1
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5551_ _5551_/A0 hold574/X _5552_/S VGND VGND VPWR VPWR _7109_/D sky130_fd_sc_hd__mux2_1
XFILLER_157_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4502_ _4502_/A _5053_/A _5165_/D VGND VGND VPWR VPWR _4502_/X sky130_fd_sc_hd__or3b_1
XFILLER_184_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5482_ _5482_/A0 hold206/X _5482_/S VGND VGND VPWR VPWR _7048_/D sky130_fd_sc_hd__mux2_1
XFILLER_6_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4433_ _4742_/B _4436_/B _4433_/C _4758_/B VGND VGND VPWR VPWR _4433_/X sky130_fd_sc_hd__and4_1
XFILLER_172_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7152_ _7180_/CLK _7152_/D wire4014/X VGND VGND VPWR VPWR _7152_/Q sky130_fd_sc_hd__dfstp_4
X_4364_ _4474_/A _4489_/A VGND VGND VPWR VPWR _4745_/A sky130_fd_sc_hd__or2_4
XFILLER_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6103_ _6103_/A1 _6103_/A2 _6103_/B1 _6103_/B2 VGND VGND VPWR VPWR _6103_/X sky130_fd_sc_hd__a22o_1
X_3315_ _3534_/A _3674_/B VGND VGND VPWR VPWR _3315_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4295_ _4295_/A0 hold270/X _4299_/S VGND VGND VPWR VPWR _4295_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7083_ _7083_/CLK _7083_/D wire4037/X VGND VGND VPWR VPWR _7083_/Q sky130_fd_sc_hd__dfstp_1
X_3246_ hold60/X _3941_/A _3244_/X _3245_/Y VGND VGND VPWR VPWR hold61/A sky130_fd_sc_hd__o31a_1
X_6034_ _6914_/Q _6061_/A2 _6034_/B1 _7058_/Q VGND VGND VPWR VPWR _6034_/X sky130_fd_sc_hd__a22o_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6936_ _7109_/CLK _6936_/D wire3999/A VGND VGND VPWR VPWR _6936_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6867_ _6939_/CLK _6867_/D _6404_/A VGND VGND VPWR VPWR _6867_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5818_ _6183_/B2 _5844_/A2 _5682_/X _6189_/A1 _5818_/C1 VGND VGND VPWR VPWR _5825_/A
+ sky130_fd_sc_hd__a221o_1
X_6798_ _6799_/CLK _6798_/D wire3935/A VGND VGND VPWR VPWR _6798_/Q sky130_fd_sc_hd__dfrtp_2
Xwire907 _3333_/Y VGND VGND VPWR VPWR wire907/X sky130_fd_sc_hd__clkbuf_2
Xwire918 wire920/X VGND VGND VPWR VPWR _5295_/A sky130_fd_sc_hd__clkbuf_1
Xwire929 wire929/A VGND VGND VPWR VPWR wire929/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5749_ _6086_/B2 _5749_/A2 _5896_/B1 _6091_/A1 _5748_/X VGND VGND VPWR VPWR _5750_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_136_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4203 input44/X VGND VGND VPWR VPWR wire4203/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire4214 wire4215/X VGND VGND VPWR VPWR _3540_/B2 sky130_fd_sc_hd__clkbuf_2
Xfanout3418 _5577_/A0 VGND VGND VPWR VPWR _5490_/A0 sky130_fd_sc_hd__clkbuf_2
Xwire4225 input37/X VGND VGND VPWR VPWR wire4225/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4236 input32/X VGND VGND VPWR VPWR _3394_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire4247 wire4248/X VGND VGND VPWR VPWR _3347_/A1 sky130_fd_sc_hd__clkbuf_1
Xhold560 _6986_/Q VGND VGND VPWR VPWR hold560/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3502 _4178_/A0 VGND VGND VPWR VPWR _4214_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_135_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3513 _5575_/A0 VGND VGND VPWR VPWR _4115_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_173_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold571 _6496_/Q VGND VGND VPWR VPWR hold571/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire4269 wire4269/A VGND VGND VPWR VPWR wire4269/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3535 _4309_/A0 VGND VGND VPWR VPWR _4333_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold582 _6767_/Q VGND VGND VPWR VPWR hold582/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_173_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold593 _7030_/Q VGND VGND VPWR VPWR hold593/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire2801 _6335_/A2 VGND VGND VPWR VPWR _6289_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3546 _4162_/A1 VGND VGND VPWR VPWR _4237_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_103_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2823 _6198_/A2 VGND VGND VPWR VPWR _6125_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3568 _4273_/A1 VGND VGND VPWR VPWR _4279_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_131_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3579 _4308_/A0 VGND VGND VPWR VPWR _5231_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2834 _5706_/X VGND VGND VPWR VPWR wire2834/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2845 wire2845/A VGND VGND VPWR VPWR _5841_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire2856 _5703_/X VGND VGND VPWR VPWR _5830_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2867 _5931_/B1 VGND VGND VPWR VPWR _5965_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2878 _5961_/A2 VGND VGND VPWR VPWR _5890_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire2889 _5738_/A2 VGND VGND VPWR VPWR _5713_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_18_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout3952 wire3956/A VGND VGND VPWR VPWR fanout3952/X sky130_fd_sc_hd__clkbuf_4
XFILLER_122_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4080_ hold682/X _4079_/X _4082_/S VGND VGND VPWR VPWR _6558_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4982_ _4982_/A _4982_/B _4982_/C VGND VGND VPWR VPWR _5119_/B sky130_fd_sc_hd__or3_1
XFILLER_63_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6721_ _6979_/CLK _6721_/D fanout4027/X VGND VGND VPWR VPWR _6721_/Q sky130_fd_sc_hd__dfrtp_1
X_3933_ _6554_/Q input3/X input1/X VGND VGND VPWR VPWR _3933_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6652_ _7206_/CLK _6652_/D VGND VGND VPWR VPWR _6652_/Q sky130_fd_sc_hd__dfxtp_1
X_3864_ _6447_/Q hold47/A _3866_/S VGND VGND VPWR VPWR _6448_/D sky130_fd_sc_hd__mux2_1
X_5603_ _7144_/Q _7145_/Q _5604_/D _7146_/Q VGND VGND VPWR VPWR _5606_/B sky130_fd_sc_hd__a31o_1
XFILLER_164_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6583_ _6945_/CLK _6583_/D fanout4078/X VGND VGND VPWR VPWR _6583_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3795_ _3801_/B VGND VGND VPWR VPWR _3795_/Y sky130_fd_sc_hd__inv_2
X_5534_ hold516/X _5534_/A1 _5534_/S VGND VGND VPWR VPWR _7094_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5465_ _5519_/A0 hold469/X _5465_/S VGND VGND VPWR VPWR _7033_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7204_ _7204_/CLK _7204_/D wire4260/X VGND VGND VPWR VPWR _7204_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_105_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4416_ _4434_/B _4444_/B VGND VGND VPWR VPWR _4758_/B sky130_fd_sc_hd__nor2_2
XFILLER_132_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5396_ hold219/X _5396_/A1 _5397_/S VGND VGND VPWR VPWR _6971_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2108 _6821_/Q VGND VGND VPWR VPWR wire2108/X sky130_fd_sc_hd__clkbuf_1
X_7135_ _7135_/CLK _7135_/D wire4052/X VGND VGND VPWR VPWR _7135_/Q sky130_fd_sc_hd__dfstp_1
X_4347_ _4402_/A _4544_/B _4359_/B VGND VGND VPWR VPWR _4350_/B sky130_fd_sc_hd__and3_1
Xwire2119 wire2120/X VGND VGND VPWR VPWR _3568_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_113_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1407 _6285_/X VGND VGND VPWR VPWR _6286_/C1 sky130_fd_sc_hd__clkbuf_1
X_7066_ _7066_/CLK _7066_/D wire3970/X VGND VGND VPWR VPWR _7066_/Q sky130_fd_sc_hd__dfstp_1
Xwire1418 wire1419/X VGND VGND VPWR VPWR _5818_/C1 sky130_fd_sc_hd__clkbuf_1
XFILLER_143_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4278_ _5582_/A0 hold368/X _4281_/S VGND VGND VPWR VPWR _6727_/D sky130_fd_sc_hd__mux2_1
Xwire1429 _5036_/B VGND VGND VPWR VPWR _5003_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_86_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6017_ _6019_/A _6033_/A _6030_/C VGND VGND VPWR VPWR _6017_/X sky130_fd_sc_hd__and3b_1
XFILLER_46_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3229_ _3229_/A VGND VGND VPWR VPWR _3229_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_wbbd_sck clkbuf_0_wbbd_sck/X VGND VGND VPWR VPWR _3942_/A2 sky130_fd_sc_hd__clkbuf_16
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6919_ _6973_/CLK _6919_/D _7087_/RESET_B VGND VGND VPWR VPWR _6919_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire715 _4328_/S VGND VGND VPWR VPWR _4329_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire726 _4119_/S VGND VGND VPWR VPWR _4115_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_109_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire737 _3982_/S VGND VGND VPWR VPWR _3976_/S sky130_fd_sc_hd__clkbuf_2
Xwire748 wire749/X VGND VGND VPWR VPWR wire748/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire759 _3706_/X VGND VGND VPWR VPWR wire759/X sky130_fd_sc_hd__clkbuf_1
XFILLER_184_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire4022 wire4022/A VGND VGND VPWR VPWR wire4022/X sky130_fd_sc_hd__dlymetal6s2s_1
Xwire4033 _6405_/A VGND VGND VPWR VPWR _6407_/A sky130_fd_sc_hd__buf_2
XFILLER_123_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire4044 wire4045/X VGND VGND VPWR VPWR wire4044/X sky130_fd_sc_hd__clkbuf_2
Xwire4055 wire4056/A VGND VGND VPWR VPWR wire4055/X sky130_fd_sc_hd__buf_2
Xwire3310 _4630_/A VGND VGND VPWR VPWR _4635_/B sky130_fd_sc_hd__clkbuf_2
Xwire4066 wire4066/A VGND VGND VPWR VPWR wire4066/X sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3321 _4575_/X VGND VGND VPWR VPWR _4814_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_2_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold390 _6765_/Q VGND VGND VPWR VPWR hold390/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire3332 _5105_/A2 VGND VGND VPWR VPWR _5036_/A sky130_fd_sc_hd__clkbuf_1
Xwire4088 wire4088/A VGND VGND VPWR VPWR wire4088/X sky130_fd_sc_hd__clkbuf_1
Xwire3343 wire3344/X VGND VGND VPWR VPWR _4684_/A sky130_fd_sc_hd__clkbuf_2
Xwire3354 _4721_/A VGND VGND VPWR VPWR _5018_/A sky130_fd_sc_hd__buf_2
Xwire4099 wire4100/X VGND VGND VPWR VPWR wire4099/X sky130_fd_sc_hd__clkbuf_1
Xwire2620 _6212_/B1 VGND VGND VPWR VPWR _6173_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire3365 _4369_/X VGND VGND VPWR VPWR _4461_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_77_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2631 _6148_/B VGND VGND VPWR VPWR _6053_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire3387 wire3387/A VGND VGND VPWR VPWR wire3387/X sky130_fd_sc_hd__clkbuf_1
Xwire2642 _6113_/B1 VGND VGND VPWR VPWR _6141_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2653 _6101_/B1 VGND VGND VPWR VPWR _6034_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire2664 _6209_/B1 VGND VGND VPWR VPWR _6086_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire2675 _6173_/A2 VGND VGND VPWR VPWR _6166_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2686 _6017_/X VGND VGND VPWR VPWR _6198_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire1941 wire1942/X VGND VGND VPWR VPWR _3224_/A sky130_fd_sc_hd__clkbuf_1
Xwire2697 _6016_/X VGND VGND VPWR VPWR wire2697/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1952 _5673_/B2 VGND VGND VPWR VPWR _6004_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire1963 _5718_/B2 VGND VGND VPWR VPWR _3709_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire1985 _5786_/A1 VGND VGND VPWR VPWR _3453_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_45_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3580_ _6619_/Q _4153_/A _3720_/B1 _6678_/Q VGND VGND VPWR VPWR _3580_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5250_ _5250_/A _5268_/B VGND VGND VPWR VPWR _5254_/S sky130_fd_sc_hd__and2_1
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4201_ hold392/X _4237_/A0 _4203_/S VGND VGND VPWR VPWR _6657_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5181_ _5123_/X _5180_/X _5160_/X VGND VGND VPWR VPWR _5181_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4132_ hold657/X _6395_/A0 _4134_/S VGND VGND VPWR VPWR _6598_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4063_ hold110/X _4062_/X _4069_/S VGND VGND VPWR VPWR _4063_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4965_ _4965_/A _4965_/B _4816_/X VGND VGND VPWR VPWR _5142_/A sky130_fd_sc_hd__or3b_1
X_6704_ _6705_/CLK _6704_/D wire3959/A VGND VGND VPWR VPWR _6704_/Q sky130_fd_sc_hd__dfrtp_1
Xmax_length4008 wire4007/A VGND VGND VPWR VPWR _7176_/RESET_B sky130_fd_sc_hd__buf_4
X_3916_ _6542_/Q _6545_/Q _3850_/B VGND VGND VPWR VPWR _3917_/B sky130_fd_sc_hd__o21ai_1
X_4896_ _5134_/A _4896_/B _4896_/C _5045_/A VGND VGND VPWR VPWR _4897_/B sky130_fd_sc_hd__or4_1
XFILLER_177_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length3307 _4610_/X VGND VGND VPWR VPWR _4645_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_177_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6635_ _6671_/CLK _6635_/D fanout4028/X VGND VGND VPWR VPWR _6635_/Q sky130_fd_sc_hd__dfrtp_1
X_3847_ _3951_/A1 _6456_/Q _3847_/S VGND VGND VPWR VPWR _6456_/D sky130_fd_sc_hd__mux2_1
XFILLER_149_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6566_ _6973_/CLK _6566_/D wire4069/X VGND VGND VPWR VPWR _6566_/Q sky130_fd_sc_hd__dfrtp_1
X_3778_ _6498_/Q _3287_/Y _5484_/A _5990_/A1 wire743/X VGND VGND VPWR VPWR _3781_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_152_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5517_ _5517_/A0 hold533/X _5517_/S VGND VGND VPWR VPWR _7079_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6497_ _6825_/CLK _6497_/D wire3956/X VGND VGND VPWR VPWR _6497_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_118_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5448_ _5448_/A _5448_/B VGND VGND VPWR VPWR _5448_/Y sky130_fd_sc_hd__nand2_1
XFILLER_160_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5379_ _5442_/A0 hold173/X _5379_/S VGND VGND VPWR VPWR _6956_/D sky130_fd_sc_hd__mux2_1
XFILLER_120_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7118_ _7132_/CLK _7118_/D fanout4077/X VGND VGND VPWR VPWR _7118_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1215 _3314_/Y VGND VGND VPWR VPWR _3425_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1226 _3310_/Y VGND VGND VPWR VPWR _3666_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1237 _3783_/A2 VGND VGND VPWR VPWR _5250_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1248 _3617_/A2 VGND VGND VPWR VPWR wire1248/X sky130_fd_sc_hd__clkbuf_1
X_7049_ _7126_/CLK _7049_/D wire4046/A VGND VGND VPWR VPWR _7049_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1259 _3654_/A2 VGND VGND VPWR VPWR _3522_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_170_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire501 _5310_/S VGND VGND VPWR VPWR _5312_/S sky130_fd_sc_hd__clkbuf_1
Xwire512 wire513/X VGND VGND VPWR VPWR _5269_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_183_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire523 _5012_/X VGND VGND VPWR VPWR _5112_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire534 wire535/X VGND VGND VPWR VPWR _4109_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_10_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire545 wire546/X VGND VGND VPWR VPWR _3688_/B sky130_fd_sc_hd__clkbuf_1
Xwire556 _3604_/X VGND VGND VPWR VPWR wire556/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire567 _3488_/X VGND VGND VPWR VPWR wire567/X sky130_fd_sc_hd__clkbuf_1
Xwire578 wire579/X VGND VGND VPWR VPWR _3371_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_155_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire589 wire590/X VGND VGND VPWR VPWR wire589/X sky130_fd_sc_hd__clkbuf_1
XFILLER_170_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3140 _5656_/X VGND VGND VPWR VPWR _5827_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3151 _5655_/X VGND VGND VPWR VPWR _5824_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3162 _6182_/A2 VGND VGND VPWR VPWR _6214_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_111_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3173 _5152_/B2 VGND VGND VPWR VPWR _4710_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_26_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3184 _4587_/B VGND VGND VPWR VPWR _4677_/B sky130_fd_sc_hd__clkbuf_2
Xwire2450 wire2451/X VGND VGND VPWR VPWR _6391_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire2461 _6306_/B1 VGND VGND VPWR VPWR _6328_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_78_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2472 _6162_/B1 VGND VGND VPWR VPWR _6139_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2483 _6158_/A2 VGND VGND VPWR VPWR _6102_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1760 wire1761/X VGND VGND VPWR VPWR _5739_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire1771 _7015_/Q VGND VGND VPWR VPWR _6150_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire1782 _7011_/Q VGND VGND VPWR VPWR _5723_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire1793 wire1794/X VGND VGND VPWR VPWR _3441_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_46_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4750_ _5002_/A _4754_/B VGND VGND VPWR VPWR _4983_/B sky130_fd_sc_hd__nor2_1
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3701_ _3701_/A _3701_/B _3701_/C _3701_/D VGND VGND VPWR VPWR _3722_/B sky130_fd_sc_hd__or4_1
XFILLER_147_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4681_ _4958_/B1 _5024_/A _5017_/A _5076_/A VGND VGND VPWR VPWR _4681_/X sky130_fd_sc_hd__o22a_1
XFILLER_146_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6420_ _6440_/A _6440_/B VGND VGND VPWR VPWR _6420_/X sky130_fd_sc_hd__and2_1
XFILLER_147_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3632_ _3632_/A _3632_/B _3632_/C _3632_/D VGND VGND VPWR VPWR _3633_/D sky130_fd_sc_hd__or4_1
XFILLER_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6351_ _7191_/Q wire363/X _6353_/S VGND VGND VPWR VPWR _7191_/D sky130_fd_sc_hd__mux2_1
X_3563_ _6668_/Q _3678_/B1 _4198_/A _6658_/Q _3549_/X VGND VGND VPWR VPWR _3563_/X
+ sky130_fd_sc_hd__a221o_1
X_5302_ _5374_/A0 hold310/X _5303_/S VGND VGND VPWR VPWR _6888_/D sky130_fd_sc_hd__mux2_1
X_6282_ _6282_/A1 _6282_/A2 _6282_/B1 _6282_/B2 _6281_/X VGND VGND VPWR VPWR _6292_/B
+ sky130_fd_sc_hd__a221o_1
X_3494_ _3494_/A1 wire971/X _3494_/B1 _3494_/B2 _3493_/X VGND VGND VPWR VPWR _3494_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5233_ _5233_/A0 hold387/X _5240_/S VGND VGND VPWR VPWR _6826_/D sky130_fd_sc_hd__mux2_1
XFILLER_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5164_ _4932_/A _4784_/A _5164_/A3 _4950_/C VGND VGND VPWR VPWR _5165_/C sky130_fd_sc_hd__o31a_1
XFILLER_69_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4115_ _4115_/A0 hold296/X _4115_/S VGND VGND VPWR VPWR _6583_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5095_ _5095_/A _5095_/B _5095_/C _5095_/D VGND VGND VPWR VPWR _5145_/B sky130_fd_sc_hd__or4_1
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4046_ _4046_/A _5210_/B VGND VGND VPWR VPWR _4051_/S sky130_fd_sc_hd__nand2_2
XFILLER_71_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5997_ _6038_/A _6019_/B VGND VGND VPWR VPWR _5997_/Y sky130_fd_sc_hd__nor2_1
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4948_ _4932_/A _4947_/A _4933_/A _4932_/B _4857_/A VGND VGND VPWR VPWR _4950_/B
+ sky130_fd_sc_hd__o41a_1
XFILLER_184_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length3115 wire3119/X VGND VGND VPWR VPWR wire3112/A sky130_fd_sc_hd__clkbuf_1
XFILLER_20_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4879_ _4996_/A _4754_/B _4510_/B VGND VGND VPWR VPWR _5174_/A sky130_fd_sc_hd__o21ai_1
XFILLER_193_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6618_ _7208_/CLK hold59/X wire4026/X VGND VGND VPWR VPWR _6618_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_20_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6549_ _6945_/CLK _6549_/D fanout4078/X VGND VGND VPWR VPWR _6549_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length1724 _7034_/Q VGND VGND VPWR VPWR _5698_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_106_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput270 _6797_/Q VGND VGND VPWR VPWR pll_div[4] sky130_fd_sc_hd__buf_12
Xoutput281 wire2443/X VGND VGND VPWR VPWR pll_trim[15] sky130_fd_sc_hd__buf_12
Xoutput292 _6805_/Q VGND VGND VPWR VPWR pll_trim[25] sky130_fd_sc_hd__buf_12
XFILLER_121_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1012 _5073_/X VGND VGND VPWR VPWR _5155_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_181_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1023 _3711_/Y VGND VGND VPWR VPWR _5200_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_75_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1034 _4330_/A VGND VGND VPWR VPWR _3617_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_181_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1045 _3754_/B1 VGND VGND VPWR VPWR _3625_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_114_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1056 _3706_/B1 VGND VGND VPWR VPWR _3766_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1067 _4216_/A VGND VGND VPWR VPWR _3747_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1078 _3465_/Y VGND VGND VPWR VPWR _4234_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1089 _3454_/Y VGND VGND VPWR VPWR _4240_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire353 _5167_/X VGND VGND VPWR VPWR wire353/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire364 wire365/X VGND VGND VPWR VPWR wire364/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire375 wire376/X VGND VGND VPWR VPWR wire375/X sky130_fd_sc_hd__clkbuf_2
Xwire386 _3633_/X VGND VGND VPWR VPWR _3660_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_109_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire397 wire398/X VGND VGND VPWR VPWR wire397/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length2981 _5781_/B1 VGND VGND VPWR VPWR wire2977/A sky130_fd_sc_hd__clkbuf_1
XFILLER_152_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2280 _6664_/Q VGND VGND VPWR VPWR _6329_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire2291 _6656_/Q VGND VGND VPWR VPWR _6249_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1590 wire1591/X VGND VGND VPWR VPWR wire1590/X sky130_fd_sc_hd__clkbuf_1
X_5920_ _6533_/Q _5920_/A2 _5930_/B1 _6279_/B2 _5919_/X VGND VGND VPWR VPWR _5923_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_74_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5851_ _6203_/B2 _5851_/A2 _5851_/B1 _5850_/X VGND VGND VPWR VPWR _5851_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4802_ _4802_/A _4802_/B _4802_/C _4802_/D VGND VGND VPWR VPWR _4822_/C sky130_fd_sc_hd__nor4_1
X_5782_ _6982_/Q _5782_/A2 _5782_/B1 _5782_/B2 _5781_/X VGND VGND VPWR VPWR _5785_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_9_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4733_ _4656_/Y _4667_/X _5039_/A _4758_/A VGND VGND VPWR VPWR _4761_/A sky130_fd_sc_hd__o22a_1
XFILLER_119_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4664_ _4664_/A _4664_/B VGND VGND VPWR VPWR _4665_/B sky130_fd_sc_hd__or2_1
XFILLER_147_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6403_ _6405_/A _6407_/B VGND VGND VPWR VPWR _6403_/X sky130_fd_sc_hd__and2_1
XFILLER_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3615_ _5736_/A1 _3615_/A2 _3615_/B1 _6956_/Q VGND VGND VPWR VPWR _3615_/X sky130_fd_sc_hd__a22o_1
X_4595_ _4674_/A _4595_/B VGND VGND VPWR VPWR _4595_/Y sky130_fd_sc_hd__nand2_1
XFILLER_162_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6334_ _6334_/A1 _6334_/A2 _6334_/B1 _6334_/B2 _6333_/X VGND VGND VPWR VPWR _6341_/B
+ sky130_fd_sc_hd__a221o_1
X_3546_ _3546_/A _3546_/B VGND VGND VPWR VPWR _3546_/Y sky130_fd_sc_hd__nor2_1
XFILLER_115_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3909 wire3910/X VGND VGND VPWR VPWR _3951_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_143_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6265_ _6265_/A1 _6290_/A2 _6265_/B1 _6707_/Q _6249_/X VGND VGND VPWR VPWR _6266_/D
+ sky130_fd_sc_hd__a221o_1
X_3477_ _3477_/A _3519_/B VGND VGND VPWR VPWR _4216_/A sky130_fd_sc_hd__nor2_1
XFILLER_130_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5216_ _5216_/A0 _5216_/A1 _5220_/S VGND VGND VPWR VPWR _6814_/D sky130_fd_sc_hd__mux2_1
X_6196_ _7181_/Q _5652_/Y _6194_/X _6195_/X VGND VGND VPWR VPWR _7181_/D sky130_fd_sc_hd__a22o_1
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5147_ _5172_/B _5147_/B VGND VGND VPWR VPWR _5147_/X sky130_fd_sc_hd__and2b_1
XFILLER_28_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5078_ _4655_/B _5108_/B _5077_/X VGND VGND VPWR VPWR _5178_/A sky130_fd_sc_hd__o21ai_1
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4029_ hold361/X _5503_/A0 _4032_/S VGND VGND VPWR VPWR _6521_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length2222 hold356/X VGND VGND VPWR VPWR _4263_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_181_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2288 hold489/X VGND VGND VPWR VPWR _4206_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_109_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold208 _7053_/Q VGND VGND VPWR VPWR hold208/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold219 _6971_/Q VGND VGND VPWR VPWR hold219/X sky130_fd_sc_hd__dlygate4sd3_1
X_3400_ _5824_/A1 _5304_/A _3397_/X _3399_/X VGND VGND VPWR VPWR _3409_/C sky130_fd_sc_hd__a211o_1
X_4380_ _4476_/A _4564_/B _4605_/A _4565_/A VGND VGND VPWR VPWR _4380_/X sky130_fd_sc_hd__or4_1
XFILLER_171_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3331_ _3331_/A _3711_/B VGND VGND VPWR VPWR _3331_/Y sky130_fd_sc_hd__nor2_1
XFILLER_152_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ _7136_/Q _6258_/A2 _6258_/B1 _6050_/B2 VGND VGND VPWR VPWR _6050_/X sky130_fd_sc_hd__a22o_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ hold114/X hold81/X _3820_/A VGND VGND VPWR VPWR _3262_/X sky130_fd_sc_hd__mux2_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ _5001_/A _5001_/B _5001_/C VGND VGND VPWR VPWR _5042_/C sky130_fd_sc_hd__and3_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3193_ _6562_/Q VGND VGND VPWR VPWR _5615_/A sky130_fd_sc_hd__inv_2
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6952_ _6973_/CLK _6952_/D _7087_/RESET_B VGND VGND VPWR VPWR _6952_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5903_ _5969_/A1 _7170_/Q wire461/X VGND VGND VPWR VPWR _5903_/X sky130_fd_sc_hd__a21o_1
X_6883_ _7135_/CLK _6883_/D wire4037/X VGND VGND VPWR VPWR _6883_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_179_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5834_ _6992_/Q _5854_/A2 _5834_/B1 _5834_/B2 _5833_/X VGND VGND VPWR VPWR _5834_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5765_ _6098_/A1 _5780_/A2 _5780_/B1 _6113_/A1 VGND VGND VPWR VPWR _5765_/X sky130_fd_sc_hd__a22o_1
X_4716_ _4745_/A _4717_/B VGND VGND VPWR VPWR _5031_/B sky130_fd_sc_hd__nor2_1
XFILLER_148_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5696_ _7152_/Q _5705_/B _5699_/C VGND VGND VPWR VPWR _5696_/X sky130_fd_sc_hd__and3_1
X_4647_ _4647_/A _4647_/B VGND VGND VPWR VPWR _4648_/B sky130_fd_sc_hd__nor2_1
XFILLER_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold720 _6483_/Q VGND VGND VPWR VPWR hold720/X sky130_fd_sc_hd__dlygate4sd3_1
X_4578_ _4588_/A _4588_/B _4621_/B _4935_/A VGND VGND VPWR VPWR _4646_/A sky130_fd_sc_hd__or4b_1
XFILLER_1_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3706 wire3707/X VGND VGND VPWR VPWR _6390_/A1 sky130_fd_sc_hd__clkbuf_1
X_6317_ _6301_/X _6307_/X _6316_/X wire977/X _6317_/B2 VGND VGND VPWR VPWR _6317_/X
+ sky130_fd_sc_hd__o32a_1
X_3529_ _3529_/A1 wire958/X _3528_/Y _6625_/Q wire805/X VGND VGND VPWR VPWR _3541_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3717 _7192_/Q VGND VGND VPWR VPWR wire3717/X sky130_fd_sc_hd__clkbuf_2
Xwire3728 _6780_/Q VGND VGND VPWR VPWR wire3728/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3739 wire3740/X VGND VGND VPWR VPWR _3265_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_39_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6248_ _6248_/A _6248_/B VGND VGND VPWR VPWR _6248_/X sky130_fd_sc_hd__and2_1
XFILLER_130_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6179_ _6179_/A1 _6003_/X _6018_/Y _6896_/Q _6178_/X VGND VGND VPWR VPWR _6180_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length1373 hold70/X VGND VGND VPWR VPWR wire1372/A sky130_fd_sc_hd__clkbuf_1
XFILLER_122_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold80 hold80/A VGND VGND VPWR VPWR hold80/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_36_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold91 hold91/A VGND VGND VPWR VPWR hold91/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3880_ _4337_/C _4337_/D _3880_/C input116/X VGND VGND VPWR VPWR _3887_/B sky130_fd_sc_hd__or4b_1
XFILLER_43_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5550_ _5550_/A0 hold232/X _5550_/S VGND VGND VPWR VPWR _7108_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4501_ _4489_/A _4387_/Y _4393_/X _4500_/X VGND VGND VPWR VPWR _5053_/A sky130_fd_sc_hd__o31ai_2
XFILLER_8_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5481_ _5481_/A0 hold654/X _5482_/S VGND VGND VPWR VPWR _7047_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4432_ _4436_/B _4433_/C VGND VGND VPWR VPWR _4724_/A sky130_fd_sc_hd__nand2_1
XFILLER_144_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7151_ _7180_/CLK _7151_/D wire4014/X VGND VGND VPWR VPWR _7151_/Q sky130_fd_sc_hd__dfrtp_1
X_4363_ _4944_/A _4363_/B _4426_/B VGND VGND VPWR VPWR _4489_/A sky130_fd_sc_hd__or3_2
X_6102_ _6102_/A1 _6102_/A2 _6102_/B1 _6981_/Q _6101_/X VGND VGND VPWR VPWR _6109_/A
+ sky130_fd_sc_hd__a221o_1
X_3314_ _3314_/A _3510_/B VGND VGND VPWR VPWR _3314_/Y sky130_fd_sc_hd__nor2_2
X_7082_ _7083_/CLK _7082_/D wire4037/X VGND VGND VPWR VPWR _7082_/Q sky130_fd_sc_hd__dfstp_1
X_4294_ _4294_/A _5193_/B VGND VGND VPWR VPWR _4299_/S sky130_fd_sc_hd__nand2_2
XFILLER_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6033_ _6033_/A _6040_/B _6040_/C VGND VGND VPWR VPWR _6033_/X sky130_fd_sc_hd__and3_1
X_3245_ wire3726/X _3963_/B VGND VGND VPWR VPWR _3245_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6935_ _7017_/CLK _6935_/D _7047_/RESET_B VGND VGND VPWR VPWR _6935_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6866_ _6939_/CLK _6866_/D _6407_/A VGND VGND VPWR VPWR _6866_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_34_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5817_ _6904_/Q _5817_/A2 _5817_/B1 _6172_/A1 VGND VGND VPWR VPWR _5817_/X sky130_fd_sc_hd__a22o_1
XFILLER_167_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6797_ _6799_/CLK _6797_/D _6743_/SET_B VGND VGND VPWR VPWR _6797_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_10_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire919 wire920/X VGND VGND VPWR VPWR wire919/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5748_ _6956_/Q _5748_/A2 _5748_/B1 _5748_/B2 VGND VGND VPWR VPWR _5748_/X sky130_fd_sc_hd__a22o_1
XFILLER_136_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5679_ _5679_/A1 _5718_/B1 _5727_/B1 _6042_/B2 VGND VGND VPWR VPWR _5679_/X sky130_fd_sc_hd__a22o_1
XFILLER_136_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire4204 wire4205/X VGND VGND VPWR VPWR _3757_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire4215 wire4216/X VGND VGND VPWR VPWR wire4215/X sky130_fd_sc_hd__clkbuf_1
Xwire4226 wire4227/X VGND VGND VPWR VPWR _3959_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_123_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire4237 wire4238/X VGND VGND VPWR VPWR _3540_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_123_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold550 _6769_/Q VGND VGND VPWR VPWR hold550/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 _7076_/Q VGND VGND VPWR VPWR hold561/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire4248 input19/X VGND VGND VPWR VPWR wire4248/X sky130_fd_sc_hd__clkbuf_1
Xwire3514 _5479_/A0 VGND VGND VPWR VPWR _5575_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold572 _6492_/Q VGND VGND VPWR VPWR hold572/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3525 hold49/X VGND VGND VPWR VPWR wire3525/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold583 _6842_/Q VGND VGND VPWR VPWR hold583/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold594 _7140_/Q VGND VGND VPWR VPWR hold594/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire2802 _5990_/A2 VGND VGND VPWR VPWR _6335_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire3547 _4162_/A1 VGND VGND VPWR VPWR _4321_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire3558 _5574_/A0 VGND VGND VPWR VPWR _5487_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_173_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2813 _6161_/A2 VGND VGND VPWR VPWR _6138_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire2824 _5977_/X VGND VGND VPWR VPWR _6198_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire3569 _4273_/A1 VGND VGND VPWR VPWR _4255_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2857 _5889_/A2 VGND VGND VPWR VPWR _5713_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_58_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2879 _5877_/B1 VGND VGND VPWR VPWR _5961_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_181_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout3953 wire4018/A VGND VGND VPWR VPWR wire3956/A sky130_fd_sc_hd__buf_6
Xfanout3964 fanout3964/A VGND VGND VPWR VPWR wire3965/A sky130_fd_sc_hd__buf_6
Xfanout3986 wire3992/A VGND VGND VPWR VPWR fanout3986/X sky130_fd_sc_hd__buf_6
XFILLER_150_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput170 wb_we_i VGND VGND VPWR VPWR _6358_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4981_ _4981_/A _4981_/B _4981_/C VGND VGND VPWR VPWR _4982_/C sky130_fd_sc_hd__nor3_1
XFILLER_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3932_ _3931_/X _3953_/B _6459_/Q VGND VGND VPWR VPWR _3932_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6720_ _6770_/CLK _6720_/D fanout4005/X VGND VGND VPWR VPWR _6720_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_44_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6651_ _7206_/CLK _6651_/D VGND VGND VPWR VPWR _6651_/Q sky130_fd_sc_hd__dfxtp_1
X_3863_ hold47/A hold14/A _3866_/S VGND VGND VPWR VPWR _6449_/D sky130_fd_sc_hd__mux2_1
XFILLER_32_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5602_ _7145_/Q _5595_/Y _5600_/Y _5601_/X VGND VGND VPWR VPWR _7145_/D sky130_fd_sc_hd__a22o_1
X_6582_ _7017_/CLK _6582_/D fanout4078/X VGND VGND VPWR VPWR _6582_/Q sky130_fd_sc_hd__dfrtp_1
X_3794_ _6541_/Q _3794_/B VGND VGND VPWR VPWR _3801_/B sky130_fd_sc_hd__or2_2
XFILLER_192_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5533_ hold676/X _5533_/A1 _5533_/S VGND VGND VPWR VPWR _7093_/D sky130_fd_sc_hd__mux2_1
XFILLER_191_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5464_ _5464_/A0 _5834_/B2 _5464_/S VGND VGND VPWR VPWR _7032_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7203_ _7204_/CLK _7203_/D wire4260/X VGND VGND VPWR VPWR _7203_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_105_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4415_ _4415_/A _4435_/B VGND VGND VPWR VPWR _4444_/B sky130_fd_sc_hd__or2_1
X_5395_ hold416/X _5440_/A0 _5397_/S VGND VGND VPWR VPWR _6970_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7134_ _7134_/CLK _7134_/D _7134_/RESET_B VGND VGND VPWR VPWR _7134_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_160_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4346_ _4544_/B _4359_/B VGND VGND VPWR VPWR _4354_/A sky130_fd_sc_hd__nand2_1
Xwire2109 _6819_/Q VGND VGND VPWR VPWR _5590_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_75_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _7066_/CLK sky130_fd_sc_hd__clkbuf_16
Xwire1408 _6271_/X VGND VGND VPWR VPWR _6281_/C1 sky130_fd_sc_hd__clkbuf_1
XFILLER_101_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7065_ _7079_/CLK _7065_/D wire4049/X VGND VGND VPWR VPWR _7065_/Q sky130_fd_sc_hd__dfrtp_1
X_4277_ _5314_/A0 hold367/X _4281_/S VGND VGND VPWR VPWR _6726_/D sky130_fd_sc_hd__mux2_1
Xwire1419 wire1420/X VGND VGND VPWR VPWR wire1419/X sky130_fd_sc_hd__clkbuf_1
X_6016_ _6039_/A _6039_/C _6020_/C VGND VGND VPWR VPWR _6016_/X sky130_fd_sc_hd__and3_1
X_3228_ _6893_/Q VGND VGND VPWR VPWR _3228_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6918_ _7140_/CLK _6918_/D wire4065/X VGND VGND VPWR VPWR _6918_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_52_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_13_csclk _7059_/CLK VGND VGND VPWR VPWR _6740_/CLK sky130_fd_sc_hd__clkbuf_16
X_6849_ _7109_/CLK _6849_/D wire3999/A VGND VGND VPWR VPWR _6849_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire705 _5258_/S VGND VGND VPWR VPWR _5256_/S sky130_fd_sc_hd__clkbuf_1
Xwire716 _4323_/S VGND VGND VPWR VPWR _4321_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_167_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire727 _4111_/X VGND VGND VPWR VPWR _4119_/S sky130_fd_sc_hd__buf_2
XFILLER_10_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire738 _3783_/X VGND VGND VPWR VPWR wire738/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire749 wire750/X VGND VGND VPWR VPWR wire749/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_28_csclk _7059_/CLK VGND VGND VPWR VPWR _7121_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_163_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4001 wire4001/A VGND VGND VPWR VPWR wire4001/X sky130_fd_sc_hd__buf_2
XFILLER_151_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4034 _6404_/A VGND VGND VPWR VPWR _6405_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire4045 wire4046/X VGND VGND VPWR VPWR wire4045/X sky130_fd_sc_hd__buf_2
XFILLER_123_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3300 _4651_/X VGND VGND VPWR VPWR _4910_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire4056 wire4056/A VGND VGND VPWR VPWR wire4056/X sky130_fd_sc_hd__clkbuf_4
Xwire3311 _4630_/A VGND VGND VPWR VPWR _5089_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3322 _4567_/B VGND VGND VPWR VPWR _5023_/C sky130_fd_sc_hd__clkbuf_2
Xhold380 _6732_/Q VGND VGND VPWR VPWR hold380/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold391 _6764_/Q VGND VGND VPWR VPWR hold391/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3333 _4752_/B VGND VGND VPWR VPWR _4754_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3344 _4465_/X VGND VGND VPWR VPWR wire3344/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3355 _4659_/A VGND VGND VPWR VPWR _4677_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2643 _6215_/B1 VGND VGND VPWR VPWR _6113_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2654 _6154_/B1 VGND VGND VPWR VPWR _6101_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1920 _6932_/Q VGND VGND VPWR VPWR _6081_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2665 _6209_/B1 VGND VGND VPWR VPWR _6158_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire2676 _6200_/B1 VGND VGND VPWR VPWR _6173_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire1931 _3365_/B2 VGND VGND VPWR VPWR _6211_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2687 _6310_/B1 VGND VGND VPWR VPWR _6325_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_65_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1942 _6925_/Q VGND VGND VPWR VPWR wire1942/X sky130_fd_sc_hd__clkbuf_1
Xwire1953 _6922_/Q VGND VGND VPWR VPWR _5673_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_18_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2698 _6024_/C VGND VGND VPWR VPWR _6129_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_58_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1964 _6915_/Q VGND VGND VPWR VPWR _5718_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_93_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1975 _5736_/B2 VGND VGND VPWR VPWR _6090_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire1986 _6902_/Q VGND VGND VPWR VPWR _5786_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_18_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1997 _5787_/A1 VGND VGND VPWR VPWR _6137_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_73_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4200_ hold358/X _4200_/A1 _4203_/S VGND VGND VPWR VPWR _4200_/X sky130_fd_sc_hd__mux2_1
X_5180_ _4939_/C _5066_/C _5180_/C _5180_/D VGND VGND VPWR VPWR _5180_/X sky130_fd_sc_hd__and4bb_1
X_4131_ hold662/X _4131_/A1 _4134_/S VGND VGND VPWR VPWR _6597_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4062_ hold74/X _4116_/A0 _4068_/S VGND VGND VPWR VPWR _4062_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4964_ _4964_/A _5112_/B VGND VGND VPWR VPWR _5103_/A sky130_fd_sc_hd__or2_1
X_6703_ _6705_/CLK _6703_/D wire3959/A VGND VGND VPWR VPWR _6703_/Q sky130_fd_sc_hd__dfstp_1
Xmax_length4009 fanout4005/X VGND VGND VPWR VPWR wire4007/A sky130_fd_sc_hd__buf_2
XFILLER_189_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3915_ _3850_/B _3890_/Y _3834_/B _3850_/A VGND VGND VPWR VPWR _6543_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_20_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4895_ _4742_/A _4742_/C _4741_/C _4741_/X VGND VGND VPWR VPWR _5045_/A sky130_fd_sc_hd__a31o_1
XFILLER_32_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3846_ _6473_/Q _6472_/Q _6471_/Q _6541_/Q VGND VGND VPWR VPWR _3847_/S sky130_fd_sc_hd__or4bb_1
X_6634_ _6671_/CLK _6634_/D wire4029/A VGND VGND VPWR VPWR _6634_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_177_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6565_ _7187_/CLK _6565_/D fanout3986/X VGND VGND VPWR VPWR _6565_/Q sky130_fd_sc_hd__dfrtp_2
X_3777_ input34/X _3777_/A2 _3777_/B1 input20/X VGND VGND VPWR VPWR _3777_/X sky130_fd_sc_hd__a22o_1
X_5516_ _5567_/A0 hold251/X _5516_/S VGND VGND VPWR VPWR _7078_/D sky130_fd_sc_hd__mux2_1
X_6496_ _6825_/CLK _6496_/D wire3956/X VGND VGND VPWR VPWR _6496_/Q sky130_fd_sc_hd__dfstp_1
X_5447_ _5561_/A0 _5447_/A1 _5447_/S VGND VGND VPWR VPWR _7017_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5378_ _5555_/A0 hold476/X _5378_/S VGND VGND VPWR VPWR _6955_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7117_ _7117_/CLK _7117_/D _7141_/RESET_B VGND VGND VPWR VPWR _7117_/Q sky130_fd_sc_hd__dfrtp_1
X_4329_ hold655/X _4329_/A1 _4329_/S VGND VGND VPWR VPWR _6770_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1205 _3625_/A2 VGND VGND VPWR VPWR _5394_/A sky130_fd_sc_hd__clkbuf_2
Xwire1216 wire1217/X VGND VGND VPWR VPWR _3741_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire1227 _3386_/A2 VGND VGND VPWR VPWR _3418_/A2 sky130_fd_sc_hd__clkbuf_1
X_7048_ _7133_/CLK _7048_/D fanout4073/X VGND VGND VPWR VPWR _7048_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1238 wire1238/A VGND VGND VPWR VPWR _3426_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_74_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1249 _3423_/A2 VGND VGND VPWR VPWR _3387_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire502 _5311_/S VGND VGND VPWR VPWR _5310_/S sky130_fd_sc_hd__clkbuf_2
Xmax_length3820 _4611_/A VGND VGND VPWR VPWR _4613_/A sky130_fd_sc_hd__clkbuf_1
Xwire513 _5268_/Y VGND VGND VPWR VPWR wire513/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire524 _4988_/Y VGND VGND VPWR VPWR _4989_/D sky130_fd_sc_hd__clkbuf_1
Xwire535 _4104_/Y VGND VGND VPWR VPWR wire535/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire546 wire547/X VGND VGND VPWR VPWR wire546/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_690 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire557 _3595_/X VGND VGND VPWR VPWR _3600_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_6_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire568 wire569/X VGND VGND VPWR VPWR _3468_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_109_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire579 _3367_/X VGND VGND VPWR VPWR wire579/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire3130 _5963_/A2 VGND VGND VPWR VPWR _5897_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_78_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3141 wire3142/X VGND VGND VPWR VPWR _5953_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire3152 _5650_/Y VGND VGND VPWR VPWR _6047_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_77_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3163 _5642_/X VGND VGND VPWR VPWR _6182_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3174 _4638_/X VGND VGND VPWR VPWR _5152_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2440 wire2441/X VGND VGND VPWR VPWR _3366_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_78_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3185 _4569_/Y VGND VGND VPWR VPWR _4804_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3196 _4535_/B VGND VGND VPWR VPWR _4802_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2451 wire2452/X VGND VGND VPWR VPWR wire2451/X sky130_fd_sc_hd__clkbuf_1
Xwire2462 wire2463/X VGND VGND VPWR VPWR _6306_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_93_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2473 _6213_/B1 VGND VGND VPWR VPWR _6162_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_19_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2484 _6209_/A2 VGND VGND VPWR VPWR _6158_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1750 _7022_/Q VGND VGND VPWR VPWR _3457_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2495 wire2496/X VGND VGND VPWR VPWR _6211_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire1761 wire1762/X VGND VGND VPWR VPWR wire1761/X sky130_fd_sc_hd__clkbuf_1
Xwire1772 _7014_/Q VGND VGND VPWR VPWR _6127_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_18_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1783 _5999_/B2 VGND VGND VPWR VPWR _3787_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_18_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1794 _7007_/Q VGND VGND VPWR VPWR wire1794/X sky130_fd_sc_hd__clkbuf_1
XFILLER_34_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3700_ _3700_/A1 _3700_/A2 wire825/X _6258_/A1 _3699_/X VGND VGND VPWR VPWR _3701_/D
+ sky130_fd_sc_hd__a221o_1
X_4680_ _4680_/A _4680_/B VGND VGND VPWR VPWR _5083_/B sky130_fd_sc_hd__nor2_1
XFILLER_186_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3631_ _6884_/Q wire920/X wire874/X _6081_/A1 _3608_/X VGND VGND VPWR VPWR _3631_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6350_ _7190_/Q wire361/X _6356_/S VGND VGND VPWR VPWR _7190_/D sky130_fd_sc_hd__mux2_1
X_3562_ _6103_/A1 wire929/X _3562_/B1 _6098_/A1 _3548_/X VGND VGND VPWR VPWR _3562_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5301_ _5526_/A0 hold696/X _5303_/S VGND VGND VPWR VPWR _6887_/D sky130_fd_sc_hd__mux2_1
XFILLER_155_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6281_ _6281_/A1 _6308_/A2 _6308_/B1 _6768_/Q _6281_/C1 VGND VGND VPWR VPWR _6281_/X
+ sky130_fd_sc_hd__a221o_1
X_3493_ _5781_/B2 wire912/X _3493_/B1 _3493_/B2 VGND VGND VPWR VPWR _3493_/X sky130_fd_sc_hd__a22o_1
X_5232_ _5232_/A _5571_/B VGND VGND VPWR VPWR _5232_/Y sky130_fd_sc_hd__nand2_1
XFILLER_115_579 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout3591 _5468_/A1 VGND VGND VPWR VPWR _5333_/A0 sky130_fd_sc_hd__clkbuf_1
X_5163_ _5163_/A _5163_/B _5163_/C VGND VGND VPWR VPWR _5163_/X sky130_fd_sc_hd__and3_1
XFILLER_96_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4114_ _4114_/A0 hold554/X _4115_/S VGND VGND VPWR VPWR _6582_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5094_ _5094_/A _5094_/B VGND VGND VPWR VPWR _5095_/D sky130_fd_sc_hd__nor2_1
XFILLER_68_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4045_ _4045_/A0 hold435/X _4045_/S VGND VGND VPWR VPWR _6535_/D sky130_fd_sc_hd__mux2_1
XFILLER_71_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5996_ _6014_/A _6030_/C VGND VGND VPWR VPWR _6019_/B sky130_fd_sc_hd__nand2_1
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4947_ _4947_/A _4947_/B VGND VGND VPWR VPWR _4947_/Y sky130_fd_sc_hd__nor2_1
XFILLER_149_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4878_ _5124_/A _4987_/B VGND VGND VPWR VPWR _4878_/X sky130_fd_sc_hd__or2_1
XFILLER_137_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3127 _5841_/A2 VGND VGND VPWR VPWR wire3123/A sky130_fd_sc_hd__clkbuf_1
Xmax_length3138 _5853_/A2 VGND VGND VPWR VPWR _5761_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_192_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length2404 _6512_/Q VGND VGND VPWR VPWR wire2403/A sky130_fd_sc_hd__clkbuf_1
X_6617_ _7112_/CLK _6617_/D wire4026/X VGND VGND VPWR VPWR _6617_/Q sky130_fd_sc_hd__dfrtp_1
X_3829_ _3252_/B _6541_/Q _6464_/Q VGND VGND VPWR VPWR _3831_/A sky130_fd_sc_hd__o21ai_1
XFILLER_165_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6548_ _6945_/CLK _6548_/D fanout4078/X VGND VGND VPWR VPWR _6548_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_180_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length1736 _7028_/Q VGND VGND VPWR VPWR _3645_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_146_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length1758 _7021_/Q VGND VGND VPWR VPWR wire1757/A sky130_fd_sc_hd__clkbuf_1
X_6479_ _7027_/CLK _6479_/D fanout3976/X VGND VGND VPWR VPWR _6479_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_106_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput260 _3950_/A VGND VGND VPWR VPWR pad_flash_io1_oeb sky130_fd_sc_hd__buf_12
XFILLER_133_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput271 _6791_/Q VGND VGND VPWR VPWR pll_ena sky130_fd_sc_hd__buf_12
Xoutput282 _6474_/Q VGND VGND VPWR VPWR pll_trim[16] sky130_fd_sc_hd__buf_12
XFILLER_160_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput293 _6492_/Q VGND VGND VPWR VPWR pll_trim[2] sky130_fd_sc_hd__buf_12
XFILLER_102_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1002 _5860_/S VGND VGND VPWR VPWR _5970_/S sky130_fd_sc_hd__clkbuf_1
Xwire1013 _5030_/X VGND VGND VPWR VPWR _5032_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_181_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1024 _3674_/Y VGND VGND VPWR VPWR _5184_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1035 hold64/A VGND VGND VPWR VPWR _3532_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_87_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1057 _4016_/A VGND VGND VPWR VPWR _3706_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1068 _4216_/A VGND VGND VPWR VPWR _3567_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1079 _3463_/Y VGND VGND VPWR VPWR _3780_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire354 _5139_/X VGND VGND VPWR VPWR _6780_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire365 _3660_/X VGND VGND VPWR VPWR wire365/X sky130_fd_sc_hd__clkbuf_1
XFILLER_171_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3683 _5688_/A VGND VGND VPWR VPWR _5693_/A sky130_fd_sc_hd__clkbuf_2
Xwire376 wire377/X VGND VGND VPWR VPWR wire376/X sky130_fd_sc_hd__clkbuf_1
Xwire387 wire388/X VGND VGND VPWR VPWR _3601_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire398 _5969_/X VGND VGND VPWR VPWR wire398/X sky130_fd_sc_hd__clkbuf_1
XFILLER_171_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2270 _6673_/Q VGND VGND VPWR VPWR _6311_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2281 _6303_/B2 VGND VGND VPWR VPWR _3597_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2292 _6655_/Q VGND VGND VPWR VPWR _3752_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire1580 _7100_/Q VGND VGND VPWR VPWR wire1580/X sky130_fd_sc_hd__clkbuf_1
Xwire1591 _7096_/Q VGND VGND VPWR VPWR wire1591/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5850_ _6977_/Q _5850_/B VGND VGND VPWR VPWR _5850_/X sky130_fd_sc_hd__or2_1
XFILLER_61_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4801_ _4674_/A _4595_/B _4804_/A2 _4764_/A VGND VGND VPWR VPWR _4813_/B sky130_fd_sc_hd__a31o_1
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5781_ _6130_/A1 _5781_/A2 _5781_/B1 _5781_/B2 VGND VGND VPWR VPWR _5781_/X sky130_fd_sc_hd__a22o_1
X_4732_ _4999_/A _4742_/A _4741_/C VGND VGND VPWR VPWR _5039_/A sky130_fd_sc_hd__and3_1
XFILLER_159_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4663_ _4664_/A _4664_/B VGND VGND VPWR VPWR _4663_/Y sky130_fd_sc_hd__nor2_1
XFILLER_159_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6402_ _6405_/A _6407_/B VGND VGND VPWR VPWR _6402_/X sky130_fd_sc_hd__and2_1
X_3614_ _6868_/Q wire913/X _5286_/A _6075_/B2 VGND VGND VPWR VPWR _3614_/X sky130_fd_sc_hd__a22o_1
X_4594_ _4632_/A _5108_/A VGND VGND VPWR VPWR _4983_/A sky130_fd_sc_hd__nor2_1
X_6333_ _5960_/A _6333_/A2 _6333_/B1 _6333_/B2 VGND VGND VPWR VPWR _6333_/X sky130_fd_sc_hd__a22o_1
X_3545_ _3544_/X _6787_/Q _3791_/B VGND VGND VPWR VPWR _6787_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6264_ _6264_/A1 _6264_/A2 _6264_/B1 _6264_/B2 _6247_/X VGND VGND VPWR VPWR _6266_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3476_ _3476_/A _3607_/B VGND VGND VPWR VPWR _3476_/Y sky130_fd_sc_hd__nor2_1
XFILLER_170_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5215_ _5453_/A0 hold513/X _5220_/S VGND VGND VPWR VPWR _6813_/D sky130_fd_sc_hd__mux2_1
X_6195_ _6219_/S _7180_/Q _6171_/S VGND VGND VPWR VPWR _6195_/X sky130_fd_sc_hd__o21a_1
XFILLER_29_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5146_ _5172_/A _5172_/C _5170_/C VGND VGND VPWR VPWR _5147_/B sky130_fd_sc_hd__or3_1
XFILLER_96_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5077_ _4655_/B _4635_/B _5027_/B _4581_/X _4860_/B VGND VGND VPWR VPWR _5077_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_84_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4028_ _4028_/A _4318_/B VGND VGND VPWR VPWR _4032_/S sky130_fd_sc_hd__and2_1
XFILLER_44_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5979_ _6040_/A _6030_/C VGND VGND VPWR VPWR _6038_/B sky130_fd_sc_hd__nand2_1
XFILLER_100_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length2245 _5900_/A1 VGND VGND VPWR VPWR _6255_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_125_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold209 _6501_/Q VGND VGND VPWR VPWR hold209/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3491 _4298_/A0 VGND VGND VPWR VPWR _5197_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_144_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3330_ _3416_/B hold84/X VGND VGND VPWR VPWR _3342_/B sky130_fd_sc_hd__nand2_1
XFILLER_124_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ _3282_/A hold68/X VGND VGND VPWR VPWR _3303_/A sky130_fd_sc_hd__and2b_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5000_ _4740_/Y _4999_/Y _4453_/A VGND VGND VPWR VPWR _5039_/B sky130_fd_sc_hd__a21oi_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3192_ _6543_/Q VGND VGND VPWR VPWR _3850_/B sky130_fd_sc_hd__inv_2
XFILLER_140_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6951_ _7116_/CLK _6951_/D _7138_/RESET_B VGND VGND VPWR VPWR _6951_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5902_ _6268_/A1 _5902_/A2 _5891_/X _5901_/X _6268_/C1 VGND VGND VPWR VPWR _5902_/X
+ sky130_fd_sc_hd__o221a_1
X_6882_ _6963_/CLK _6882_/D _7042_/SET_B VGND VGND VPWR VPWR _6882_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_179_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5833_ _5833_/A1 _5845_/A2 _5851_/A2 _6912_/Q VGND VGND VPWR VPWR _5833_/X sky130_fd_sc_hd__a22o_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5764_ _5764_/A1 _5764_/A2 _5764_/B1 _6108_/B2 _5763_/X VGND VGND VPWR VPWR _5770_/A
+ sky130_fd_sc_hd__a221o_1
X_4715_ _4478_/Y _4563_/B _4771_/B1 _4714_/X VGND VGND VPWR VPWR _4722_/B sky130_fd_sc_hd__a211o_1
X_5695_ _5990_/B2 _5695_/A2 _5695_/B1 _5995_/B2 _5695_/C1 VGND VGND VPWR VPWR _5708_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_108_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4646_ _4646_/A _4646_/B VGND VGND VPWR VPWR _4646_/X sky130_fd_sc_hd__or2_1
XFILLER_190_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold710 _7034_/Q VGND VGND VPWR VPWR hold710/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold721 _7003_/Q VGND VGND VPWR VPWR hold721/X sky130_fd_sc_hd__dlygate4sd3_1
X_4577_ _4814_/B _5027_/A VGND VGND VPWR VPWR _5115_/A sky130_fd_sc_hd__nor2_1
XFILLER_150_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6316_ _6316_/A _6316_/B _6316_/C VGND VGND VPWR VPWR _6316_/X sky130_fd_sc_hd__or3_1
X_3528_ _3528_/A _3528_/B VGND VGND VPWR VPWR _3528_/Y sky130_fd_sc_hd__nor2_1
XFILLER_115_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3707 wire3708/X VGND VGND VPWR VPWR wire3707/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3718 _7191_/Q VGND VGND VPWR VPWR wire3718/X sky130_fd_sc_hd__clkbuf_2
Xwire3729 _6780_/Q VGND VGND VPWR VPWR _5111_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_103_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6247_ _7091_/Q _6247_/A2 _6247_/B1 _6676_/Q VGND VGND VPWR VPWR _6247_/X sky130_fd_sc_hd__a22o_1
X_3459_ _6950_/Q _3459_/A2 _5439_/A _6127_/B2 VGND VGND VPWR VPWR _3459_/X sky130_fd_sc_hd__a22o_1
XFILLER_39_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6178_ _7101_/Q _6029_/B _6178_/B1 _6984_/Q VGND VGND VPWR VPWR _6178_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5129_ _5123_/X _5128_/X _5160_/A VGND VGND VPWR VPWR _5139_/C sky130_fd_sc_hd__a21oi_1
XFILLER_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold70 hold70/A VGND VGND VPWR VPWR hold70/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold81 hold81/A VGND VGND VPWR VPWR hold81/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 hold92/A VGND VGND VPWR VPWR hold92/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4500_ _4351_/A _4351_/B _4497_/A _4981_/A _4391_/Y VGND VGND VPWR VPWR _4500_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_172_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5480_ _5480_/A0 hold129/X _5480_/S VGND VGND VPWR VPWR _7046_/D sky130_fd_sc_hd__mux2_1
XFILLER_8_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1 _3444_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4431_ _4846_/C _4459_/B VGND VGND VPWR VPWR _4491_/B sky130_fd_sc_hd__nand2_1
XFILLER_172_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4362_ _4363_/B _4426_/B VGND VGND VPWR VPWR _4362_/Y sky130_fd_sc_hd__nor2_1
X_7150_ _7180_/CLK _7150_/D wire3996/X VGND VGND VPWR VPWR _7150_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3313_ _3416_/A _3313_/B VGND VGND VPWR VPWR hold70/A sky130_fd_sc_hd__nand2_1
X_6101_ _6101_/A1 _6161_/A2 _6101_/B1 _6101_/B2 VGND VGND VPWR VPWR _6101_/X sky130_fd_sc_hd__a22o_1
X_7081_ _7081_/CLK _7081_/D fanout3986/X VGND VGND VPWR VPWR _7081_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4293_ _4305_/A0 hold234/X _4293_/S VGND VGND VPWR VPWR _6740_/D sky130_fd_sc_hd__mux2_1
X_3244_ _3244_/A _3820_/A VGND VGND VPWR VPWR _3244_/X sky130_fd_sc_hd__and2_1
XFILLER_113_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6032_ _7111_/Q _6032_/A2 _6032_/B1 _6032_/B2 _6031_/X VGND VGND VPWR VPWR _6044_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_140_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6934_ _7130_/CLK _6934_/D wire4061/X VGND VGND VPWR VPWR _6934_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6865_ _7064_/CLK _6865_/D wire4045/X VGND VGND VPWR VPWR _6865_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_179_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5816_ _7167_/Q _5815_/X _5838_/S VGND VGND VPWR VPWR _7167_/D sky130_fd_sc_hd__mux2_1
X_6796_ _6799_/CLK _6796_/D wire3935/A VGND VGND VPWR VPWR _6796_/Q sky130_fd_sc_hd__dfrtp_1
Xwire909 wire910/X VGND VGND VPWR VPWR _5277_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_148_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5747_ _5747_/A1 _5775_/B1 _5747_/B1 _6916_/Q _5747_/C1 VGND VGND VPWR VPWR _5750_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_136_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5678_ _7152_/Q _5705_/B _5706_/C VGND VGND VPWR VPWR _5678_/X sky130_fd_sc_hd__and3_1
XFILLER_108_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4629_ _4629_/A _4680_/A VGND VGND VPWR VPWR _5017_/A sky130_fd_sc_hd__or2_1
XFILLER_135_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire4205 wire4206/X VGND VGND VPWR VPWR wire4205/X sky130_fd_sc_hd__clkbuf_1
Xwire4216 input39/X VGND VGND VPWR VPWR wire4216/X sky130_fd_sc_hd__clkbuf_1
Xwire4227 wire4228/X VGND VGND VPWR VPWR wire4227/X sky130_fd_sc_hd__clkbuf_1
Xhold540 _7208_/Q VGND VGND VPWR VPWR hold540/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold551 _6506_/Q VGND VGND VPWR VPWR hold551/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire4238 input30/X VGND VGND VPWR VPWR wire4238/X sky130_fd_sc_hd__clkbuf_1
Xwire4249 wire4250/X VGND VGND VPWR VPWR _3407_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire3504 _5452_/A0 VGND VGND VPWR VPWR _5216_/A0 sky130_fd_sc_hd__clkbuf_1
Xwire3515 _5479_/A0 VGND VGND VPWR VPWR _5398_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold562 _6493_/Q VGND VGND VPWR VPWR hold562/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 _6960_/Q VGND VGND VPWR VPWR hold573/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 _7081_/Q VGND VGND VPWR VPWR hold584/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 _7056_/Q VGND VGND VPWR VPWR hold595/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire2803 _5988_/X VGND VGND VPWR VPWR _5990_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire2814 _6212_/A2 VGND VGND VPWR VPWR _6161_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire3559 _4114_/A0 VGND VGND VPWR VPWR _5244_/A0 sky130_fd_sc_hd__clkbuf_1
Xwire2836 wire2836/A VGND VGND VPWR VPWR _5941_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire2847 _5952_/B1 VGND VGND VPWR VPWR _5893_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire2858 _5958_/A2 VGND VGND VPWR VPWR _5930_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire2869 _5701_/B1 VGND VGND VPWR VPWR _5931_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_66_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout3976 wire3985/A VGND VGND VPWR VPWR fanout3976/X sky130_fd_sc_hd__buf_8
XFILLER_122_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout3998 wire4013/X VGND VGND VPWR VPWR wire4001/A sky130_fd_sc_hd__buf_6
XFILLER_122_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput160 wb_dat_i[6] VGND VGND VPWR VPWR _6382_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4980_ _5059_/A _5130_/A _5158_/B VGND VGND VPWR VPWR _4980_/X sky130_fd_sc_hd__or3_1
XFILLER_63_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3931_ _3930_/X _3931_/A1 _6461_/Q VGND VGND VPWR VPWR _3931_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6650_ _7206_/CLK _6650_/D VGND VGND VPWR VPWR _6650_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3862_ hold14/A _6450_/Q _3866_/S VGND VGND VPWR VPWR _6450_/D sky130_fd_sc_hd__mux2_1
XFILLER_31_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5601_ _7144_/Q _7145_/Q _6565_/Q _5593_/B _5592_/Y VGND VGND VPWR VPWR _5601_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_149_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6581_ _6945_/CLK _6581_/D fanout4078/X VGND VGND VPWR VPWR _6581_/Q sky130_fd_sc_hd__dfrtp_1
X_3793_ _3850_/A _6543_/Q VGND VGND VPWR VPWR _3794_/B sky130_fd_sc_hd__or2_1
XFILLER_164_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5532_ hold556/X _5532_/A1 _5533_/S VGND VGND VPWR VPWR _7092_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_9_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _7067_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_172_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5463_ _5463_/A0 hold178/X _5463_/S VGND VGND VPWR VPWR _5463_/X sky130_fd_sc_hd__mux2_1
X_7202_ _7204_/CLK _7202_/D wire4260/X VGND VGND VPWR VPWR _7202_/Q sky130_fd_sc_hd__dfrtp_1
X_4414_ _4544_/B _4538_/B _4402_/A VGND VGND VPWR VPWR _4435_/B sky130_fd_sc_hd__a21oi_1
XFILLER_172_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5394_ _5394_/A _5562_/B VGND VGND VPWR VPWR _5402_/S sky130_fd_sc_hd__and2_1
X_7133_ _7133_/CLK hold53/X fanout4077/X VGND VGND VPWR VPWR hold52/A sky130_fd_sc_hd__dfrtp_1
X_4345_ _4570_/A _4570_/B _4570_/C _4570_/D VGND VGND VPWR VPWR _4781_/A sky130_fd_sc_hd__o211a_1
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4276_ _4276_/A _4276_/B VGND VGND VPWR VPWR _4281_/S sky130_fd_sc_hd__nand2_2
X_7064_ _7064_/CLK _7064_/D wire4049/X VGND VGND VPWR VPWR _7064_/Q sky130_fd_sc_hd__dfrtp_1
Xwire1409 wire1410/X VGND VGND VPWR VPWR _6233_/C1 sky130_fd_sc_hd__clkbuf_1
XFILLER_101_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6015_ _6039_/C _6020_/C _6040_/C VGND VGND VPWR VPWR _6015_/X sky130_fd_sc_hd__and3_1
X_3227_ _3227_/A VGND VGND VPWR VPWR _3227_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6917_ _6921_/CLK _6917_/D wire4046/X VGND VGND VPWR VPWR _6917_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6848_ _7072_/CLK _6848_/D wire3995/X VGND VGND VPWR VPWR _6848_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire706 _5254_/S VGND VGND VPWR VPWR _5258_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_183_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire717 _4317_/S VGND VGND VPWR VPWR _4316_/S sky130_fd_sc_hd__clkbuf_2
X_6779_ _7196_/CLK _6779_/D _6780_/RESET_B VGND VGND VPWR VPWR _6779_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_183_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire728 _4032_/S VGND VGND VPWR VPWR _4033_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_183_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire739 wire740/X VGND VGND VPWR VPWR wire739/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire4013 wire4015/X VGND VGND VPWR VPWR wire4013/X sky130_fd_sc_hd__dlymetal6s2s_1
Xwire4046 wire4046/A VGND VGND VPWR VPWR wire4046/X sky130_fd_sc_hd__clkbuf_2
Xwire3301 _4651_/X VGND VGND VPWR VPWR _4707_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_117_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold370 _4161_/X VGND VGND VPWR VPWR _6622_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 _6733_/Q VGND VGND VPWR VPWR hold381/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3323 _4680_/A VGND VGND VPWR VPWR _4693_/C sky130_fd_sc_hd__clkbuf_1
Xwire3334 _5105_/A2 VGND VGND VPWR VPWR _4752_/B sky130_fd_sc_hd__clkbuf_2
Xwire2600 _4671_/Y VGND VGND VPWR VPWR _4897_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold392 _6657_/Q VGND VGND VPWR VPWR hold392/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3345 _4738_/A VGND VGND VPWR VPWR _4527_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire2611 _4393_/X VGND VGND VPWR VPWR _4932_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_77_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3356 _5023_/A VGND VGND VPWR VPWR _4659_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3367 _4397_/A VGND VGND VPWR VPWR _4931_/A sky130_fd_sc_hd__clkbuf_1
Xwire2622 wire2623/X VGND VGND VPWR VPWR _6212_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire3378 _3991_/A1 VGND VGND VPWR VPWR _4000_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2633 _6207_/A2 VGND VGND VPWR VPWR _6148_/B sky130_fd_sc_hd__clkbuf_2
Xwire2644 _6181_/B1 VGND VGND VPWR VPWR _6215_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire2655 _6205_/B1 VGND VGND VPWR VPWR _6154_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire1921 _6931_/Q VGND VGND VPWR VPWR _3695_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2666 wire2667/X VGND VGND VPWR VPWR _6209_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire1932 hold79/A VGND VGND VPWR VPWR _3365_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire2688 wire2689/X VGND VGND VPWR VPWR _6310_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_46_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1943 _5764_/A1 VGND VGND VPWR VPWR _6114_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2699 _6303_/B1 VGND VGND VPWR VPWR _6329_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1965 _6914_/Q VGND VGND VPWR VPWR _5679_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_92_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1976 wire1977/X VGND VGND VPWR VPWR _5736_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_133_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1987 _6901_/Q VGND VGND VPWR VPWR _3227_/A sky130_fd_sc_hd__clkbuf_1
Xwire1998 wire1999/X VGND VGND VPWR VPWR _5787_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_73_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length893 wire894/X VGND VGND VPWR VPWR _5571_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_181_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__1134_ clkbuf_0__1134_/X VGND VGND VPWR VPWR _4194_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_96_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4130_ hold619/X _4130_/A1 _4134_/S VGND VGND VPWR VPWR _6596_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3890 input89/X VGND VGND VPWR VPWR wire3890/X sky130_fd_sc_hd__clkbuf_1
X_4061_ hold388/X _4060_/X _4061_/S VGND VGND VPWR VPWR _6549_/D sky130_fd_sc_hd__mux2_1
XFILLER_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4963_ _4963_/A _4963_/B VGND VGND VPWR VPWR _5112_/B sky130_fd_sc_hd__or2_1
X_6702_ _6702_/CLK _6702_/D fanout3964/A VGND VGND VPWR VPWR _6702_/Q sky130_fd_sc_hd__dfrtp_1
X_3914_ _6444_/Q _6445_/Q _3835_/S _3834_/B _3190_/Y VGND VGND VPWR VPWR _6544_/D
+ sky130_fd_sc_hd__o32ai_1
XFILLER_51_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4894_ _4894_/A _4894_/B _4894_/C _4490_/X VGND VGND VPWR VPWR _4896_/C sky130_fd_sc_hd__or4b_1
XFILLER_149_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6633_ _7196_/CLK _6633_/D VGND VGND VPWR VPWR _6633_/Q sky130_fd_sc_hd__dfxtp_1
X_3845_ _3859_/A1 _6457_/Q _3845_/S VGND VGND VPWR VPWR _6457_/D sky130_fd_sc_hd__mux2_1
XFILLER_165_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6564_ _7180_/CLK _6564_/D _6562_/SET_B VGND VGND VPWR VPWR _6564_/Q sky130_fd_sc_hd__dfrtp_4
X_3776_ _3776_/A1 _3776_/A2 _3776_/B1 _7207_/Q _3775_/X VGND VGND VPWR VPWR _3781_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_138_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5515_ _5515_/A0 hold687/X _5515_/S VGND VGND VPWR VPWR _7077_/D sky130_fd_sc_hd__mux2_1
X_6495_ _6825_/CLK _6495_/D _6495_/SET_B VGND VGND VPWR VPWR _6495_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_173_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5446_ _5587_/A0 hold686/X _5446_/S VGND VGND VPWR VPWR _7016_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5377_ _5563_/A0 _5377_/A1 _5378_/S VGND VGND VPWR VPWR _6954_/D sky130_fd_sc_hd__mux2_1
X_7116_ _7116_/CLK _7116_/D _7138_/RESET_B VGND VGND VPWR VPWR _7116_/Q sky130_fd_sc_hd__dfrtp_1
X_4328_ hold550/X _5539_/A1 _4328_/S VGND VGND VPWR VPWR _6769_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1206 wire1206/A VGND VGND VPWR VPWR _3625_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire1217 _3311_/Y VGND VGND VPWR VPWR wire1217/X sky130_fd_sc_hd__clkbuf_1
X_7047_ _7133_/CLK _7047_/D _7047_/RESET_B VGND VGND VPWR VPWR _7047_/Q sky130_fd_sc_hd__dfrtp_1
Xwire1228 _3568_/A2 VGND VGND VPWR VPWR _3386_/A2 sky130_fd_sc_hd__clkbuf_2
X_4259_ hold497/X _4259_/A1 _4263_/S VGND VGND VPWR VPWR _6711_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire503 _5304_/Y VGND VGND VPWR VPWR _5311_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire514 _5275_/S VGND VGND VPWR VPWR _5276_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire525 _4269_/S VGND VGND VPWR VPWR _4268_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_7_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire536 wire536/A VGND VGND VPWR VPWR wire536/X sky130_fd_sc_hd__clkbuf_1
Xwire547 wire548/X VGND VGND VPWR VPWR wire547/X sky130_fd_sc_hd__clkbuf_1
Xwire558 _3580_/X VGND VGND VPWR VPWR wire558/X sky130_fd_sc_hd__clkbuf_1
Xwire569 _3461_/X VGND VGND VPWR VPWR wire569/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3120 _5661_/X VGND VGND VPWR VPWR wire3120/X sky130_fd_sc_hd__clkbuf_1
Xwire3131 _5928_/A2 VGND VGND VPWR VPWR _5963_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire3142 wire3142/A VGND VGND VPWR VPWR wire3142/X sky130_fd_sc_hd__clkbuf_1
Xwire3153 wire3153/A VGND VGND VPWR VPWR _6298_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_151_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3164 _4675_/B VGND VGND VPWR VPWR _4680_/B sky130_fd_sc_hd__clkbuf_2
Xwire2430 wire2431/X VGND VGND VPWR VPWR _5732_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_78_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3175 _4689_/B VGND VGND VPWR VPWR _4831_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire2441 wire2442/X VGND VGND VPWR VPWR wire2441/X sky130_fd_sc_hd__clkbuf_1
Xwire3186 _4567_/X VGND VGND VPWR VPWR _4632_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_78_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3197 _4816_/A2 VGND VGND VPWR VPWR _4805_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2452 wire2453/X VGND VGND VPWR VPWR wire2452/X sky130_fd_sc_hd__clkbuf_1
Xwire2463 _6038_/Y VGND VGND VPWR VPWR wire2463/X sky130_fd_sc_hd__clkbuf_1
XFILLER_120_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2474 wire2474/A VGND VGND VPWR VPWR _6213_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire1740 _7027_/Q VGND VGND VPWR VPWR wire1740/X sky130_fd_sc_hd__clkbuf_1
Xwire2485 _6189_/B1 VGND VGND VPWR VPWR _6209_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire1751 wire1751/A VGND VGND VPWR VPWR _6130_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire2496 _6018_/Y VGND VGND VPWR VPWR wire2496/X sky130_fd_sc_hd__clkbuf_1
Xwire1762 _7020_/Q VGND VGND VPWR VPWR wire1762/X sky130_fd_sc_hd__clkbuf_1
Xwire1773 wire1774/X VGND VGND VPWR VPWR _3596_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire1784 wire1785/X VGND VGND VPWR VPWR _5999_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire1795 _3533_/A1 VGND VGND VPWR VPWR _5788_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_523 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_74_csclk _7117_/CLK VGND VGND VPWR VPWR _7068_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_147_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3630_ _6636_/Q wire836/X _3489_/Y _3630_/B2 _3610_/X VGND VGND VPWR VPWR _3632_/C
+ sky130_fd_sc_hd__a221o_1
X_3561_ _3561_/A1 _3561_/A2 _4028_/A _6524_/Q VGND VGND VPWR VPWR _3561_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5300_ _5489_/A0 hold454/X _5303_/S VGND VGND VPWR VPWR _6886_/D sky130_fd_sc_hd__mux2_1
XFILLER_6_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3492_ _3525_/A _3492_/B VGND VGND VPWR VPWR _4016_/A sky130_fd_sc_hd__nor2_1
X_6280_ _6280_/A _6280_/B _6280_/C _6280_/D VGND VGND VPWR VPWR _6280_/X sky130_fd_sc_hd__or4_1
XFILLER_154_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5231_ _5231_/A0 hold344/X _5231_/S VGND VGND VPWR VPWR _6825_/D sky130_fd_sc_hd__mux2_1
XFILLER_170_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_580 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5162_ _5162_/A _5162_/B _5162_/C _5162_/D VGND VGND VPWR VPWR _5163_/C sky130_fd_sc_hd__nor4_1
XFILLER_111_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_12_csclk _7059_/CLK VGND VGND VPWR VPWR _6979_/CLK sky130_fd_sc_hd__clkbuf_16
X_4113_ _4113_/A0 hold102/X _4115_/S VGND VGND VPWR VPWR _6581_/D sky130_fd_sc_hd__mux2_1
X_5093_ _4425_/B _4728_/B _5083_/A _4785_/X VGND VGND VPWR VPWR _5114_/C sky130_fd_sc_hd__a211o_1
XFILLER_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4044_ _6396_/A0 hold430/X _4045_/S VGND VGND VPWR VPWR _6534_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_27_csclk _7059_/CLK VGND VGND VPWR VPWR _7104_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_25_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5995_ _6498_/Q _5995_/A2 _5995_/B1 _5995_/B2 VGND VGND VPWR VPWR _5995_/X sky130_fd_sc_hd__a22o_1
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4946_ _5064_/B _5126_/C _5053_/B _4945_/X VGND VGND VPWR VPWR _4960_/A sky130_fd_sc_hd__or4b_1
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4877_ _4485_/B _4524_/B _4983_/B VGND VGND VPWR VPWR _5049_/C sky130_fd_sc_hd__a21o_1
XFILLER_177_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6616_ _7112_/CLK _6616_/D wire4026/X VGND VGND VPWR VPWR _6616_/Q sky130_fd_sc_hd__dfrtp_1
X_3828_ _3827_/X hold66/A _3828_/S VGND VGND VPWR VPWR _6465_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length2427 _6501_/Q VGND VGND VPWR VPWR _3203_/A sky130_fd_sc_hd__clkbuf_1
X_6547_ _6945_/CLK _6547_/D fanout4078/X VGND VGND VPWR VPWR _6547_/Q sky130_fd_sc_hd__dfrtp_1
Xmax_length2438 _6495_/Q VGND VGND VPWR VPWR wire2437/A sky130_fd_sc_hd__clkbuf_1
Xmax_length2449 _6481_/Q VGND VGND VPWR VPWR wire2448/A sky130_fd_sc_hd__clkbuf_1
Xmax_length1704 _5777_/A1 VGND VGND VPWR VPWR wire1703/A sky130_fd_sc_hd__clkbuf_1
X_3759_ _7119_/Q wire889/X wire871/X _5986_/B2 wire538/X VGND VGND VPWR VPWR _3760_/D
+ sky130_fd_sc_hd__a221o_1
X_6478_ _6824_/CLK _6478_/D _6483_/SET_B VGND VGND VPWR VPWR _6478_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_145_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5429_ _5429_/A0 hold507/X _5429_/S VGND VGND VPWR VPWR _7001_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput250 _3927_/X VGND VGND VPWR VPWR mgmt_gpio_out[9] sky130_fd_sc_hd__clkbuf_1
XFILLER_160_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput261 _6801_/Q VGND VGND VPWR VPWR pll90_sel[0] sky130_fd_sc_hd__buf_12
XFILLER_160_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput272 _6798_/Q VGND VGND VPWR VPWR pll_sel[0] sky130_fd_sc_hd__buf_12
XFILLER_133_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput283 _6475_/Q VGND VGND VPWR VPWR pll_trim[17] sky130_fd_sc_hd__buf_12
XFILLER_160_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput294 _6493_/Q VGND VGND VPWR VPWR pll_trim[3] sky130_fd_sc_hd__buf_12
XFILLER_58_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1014 _4983_/Y VGND VGND VPWR VPWR _4989_/C sky130_fd_sc_hd__clkbuf_1
Xwire1025 wire1026/X VGND VGND VPWR VPWR _5225_/A sky130_fd_sc_hd__clkbuf_2
Xwire1036 hold64/X VGND VGND VPWR VPWR _4270_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1047 _3767_/A2 VGND VGND VPWR VPWR _3665_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1058 _4258_/A VGND VGND VPWR VPWR _3579_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire1069 _3480_/B1 VGND VGND VPWR VPWR _3667_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire355 _5104_/X VGND VGND VPWR VPWR _6779_/D sky130_fd_sc_hd__clkbuf_1
Xwire366 wire367/X VGND VGND VPWR VPWR wire366/X sky130_fd_sc_hd__dlymetal6s2s_1
Xwire377 _3410_/X VGND VGND VPWR VPWR wire377/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire388 _3583_/X VGND VGND VPWR VPWR wire388/X sky130_fd_sc_hd__clkbuf_1
XFILLER_99_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire399 _5859_/X VGND VGND VPWR VPWR wire399/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_1_wb_clk_i clkbuf_1_1_1_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire2260 _6679_/Q VGND VGND VPWR VPWR _6327_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2271 _6672_/Q VGND VGND VPWR VPWR _5922_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2282 _6663_/Q VGND VGND VPWR VPWR _6303_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2293 _4199_/A0 VGND VGND VPWR VPWR _6224_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_65_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1570 wire1571/X VGND VGND VPWR VPWR wire1570/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1581 wire1581/A VGND VGND VPWR VPWR _6134_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4800_ _4804_/A2 _4800_/A2 _4753_/Y VGND VGND VPWR VPWR _5090_/A sky130_fd_sc_hd__a21o_1
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5780_ _6958_/Q _5780_/A2 _5780_/B1 _5780_/B2 _5779_/X VGND VGND VPWR VPWR _5780_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4731_ _4484_/B _4731_/B _4731_/C VGND VGND VPWR VPWR _4731_/X sky130_fd_sc_hd__and3b_1
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4662_ _4931_/A _4662_/B VGND VGND VPWR VPWR _4662_/Y sky130_fd_sc_hd__nand2_1
X_6401_ _6401_/A _6407_/B VGND VGND VPWR VPWR _6401_/X sky130_fd_sc_hd__and2_1
X_3613_ _5735_/B2 _5367_/A _3613_/B1 hold91/A VGND VGND VPWR VPWR _3613_/X sky130_fd_sc_hd__a22o_1
X_4593_ _4661_/B _4707_/A VGND VGND VPWR VPWR _4620_/A sky130_fd_sc_hd__or2_1
X_6332_ _6332_/A _6332_/B _6332_/C VGND VGND VPWR VPWR _6332_/X sky130_fd_sc_hd__or3_1
X_3544_ _4194_/A1 _6786_/Q _3791_/A VGND VGND VPWR VPWR _3544_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6263_ _6607_/Q _6286_/A2 _6286_/B1 _6622_/Q _6262_/X VGND VGND VPWR VPWR _6266_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3475_ _3475_/A1 _3475_/A2 _4264_/A _6720_/Q _3473_/X VGND VGND VPWR VPWR _3484_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_170_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5214_ _5214_/A _5511_/B VGND VGND VPWR VPWR _5220_/S sky130_fd_sc_hd__nand2_2
X_6194_ _6194_/A1 wire992/X _6193_/X _6194_/C1 VGND VGND VPWR VPWR _6194_/X sky130_fd_sc_hd__a211o_1
XFILLER_69_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5145_ _5145_/A _5145_/B _5144_/X VGND VGND VPWR VPWR _5145_/X sky130_fd_sc_hd__or3b_1
XFILLER_57_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5076_ _5076_/A _5076_/B VGND VGND VPWR VPWR _5108_/B sky130_fd_sc_hd__and2_2
X_4027_ hold329/X _4209_/A1 _4027_/S VGND VGND VPWR VPWR _6520_/D sky130_fd_sc_hd__mux2_1
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5978_ _7156_/Q _7155_/Q VGND VGND VPWR VPWR _6030_/C sky130_fd_sc_hd__nor2_2
XFILLER_80_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4929_ _4929_/A1 _5034_/B1 _4825_/X _4928_/X VGND VGND VPWR VPWR _6777_/D sky130_fd_sc_hd__o22a_1
XFILLER_100_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length1556 _7122_/Q VGND VGND VPWR VPWR wire1555/A sky130_fd_sc_hd__clkbuf_1
XFILLER_69_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length3492 _4286_/A0 VGND VGND VPWR VPWR _4298_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ hold67/X _3260_/A1 _3265_/S VGND VGND VPWR VPWR hold68/A sky130_fd_sc_hd__mux2_1
XFILLER_98_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3191_ _6697_/Q VGND VGND VPWR VPWR _3191_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2090 _6850_/Q VGND VGND VPWR VPWR _5981_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_26_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6950_ _7139_/CLK _6950_/D wire4065/X VGND VGND VPWR VPWR _6950_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5901_ _5901_/A _5901_/B _5901_/C _5901_/D VGND VGND VPWR VPWR _5901_/X sky130_fd_sc_hd__or4_1
X_6881_ _7134_/CLK _6881_/D _7134_/RESET_B VGND VGND VPWR VPWR _6881_/Q sky130_fd_sc_hd__dfrtp_1
X_5832_ _6952_/Q _5832_/A2 _5832_/B1 _6172_/B2 _5831_/X VGND VGND VPWR VPWR _5832_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5763_ _5763_/A1 _5763_/A2 _5763_/B1 _5763_/B2 VGND VGND VPWR VPWR _5763_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4714_ _4714_/A _4714_/B _4822_/A _4686_/X VGND VGND VPWR VPWR _4714_/X sky130_fd_sc_hd__or4b_1
XFILLER_187_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5694_ _7152_/Q _5706_/C _5703_/C VGND VGND VPWR VPWR _5694_/X sky130_fd_sc_hd__and3_1
XFILLER_147_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4645_ _5013_/B _4645_/B VGND VGND VPWR VPWR _4645_/X sky130_fd_sc_hd__or2_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold700 _6486_/Q VGND VGND VPWR VPWR hold700/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold711 _6478_/Q VGND VGND VPWR VPWR hold711/X sky130_fd_sc_hd__dlygate4sd3_1
X_4576_ _4814_/A _4704_/A VGND VGND VPWR VPWR _5027_/A sky130_fd_sc_hd__or2_4
XFILLER_146_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold722 _7200_/Q VGND VGND VPWR VPWR hold722/X sky130_fd_sc_hd__dlygate4sd3_1
X_6315_ _6315_/A _6315_/B _6315_/C _6315_/D VGND VGND VPWR VPWR _6315_/X sky130_fd_sc_hd__or4_1
XFILLER_190_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3527_ _6540_/Q _4046_/A _5187_/A _6797_/Q VGND VGND VPWR VPWR _3527_/X sky130_fd_sc_hd__a22o_1
Xwire3708 wire3709/X VGND VGND VPWR VPWR wire3708/X sky130_fd_sc_hd__clkbuf_1
Xwire3719 _7188_/Q VGND VGND VPWR VPWR wire3719/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6246_ _6727_/Q _6296_/A2 _6296_/B1 _6246_/B2 VGND VGND VPWR VPWR _6246_/X sky130_fd_sc_hd__a22o_1
X_3458_ _6337_/A1 _3454_/Y _3771_/B1 _6336_/B2 wire831/X VGND VGND VPWR VPWR _3458_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6177_ _6177_/A1 _6006_/Y _6176_/X VGND VGND VPWR VPWR _6180_/C sky130_fd_sc_hd__a21o_1
X_3389_ _3389_/A1 _5340_/A _5358_/A _6172_/B2 VGND VGND VPWR VPWR _3389_/X sky130_fd_sc_hd__a22o_1
X_5128_ _5160_/B _5128_/B _5128_/C _5159_/B VGND VGND VPWR VPWR _5128_/X sky130_fd_sc_hd__and4b_1
XFILLER_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5059_ _5059_/A _5059_/B _5059_/C VGND VGND VPWR VPWR _5059_/Y sky130_fd_sc_hd__nor3_1
XFILLER_57_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length2054 _6869_/Q VGND VGND VPWR VPWR _5281_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_181_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length2087 hold51/X VGND VGND VPWR VPWR _5263_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_107_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold60 hold60/A VGND VGND VPWR VPWR hold60/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 hold71/A VGND VGND VPWR VPWR hold71/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_36_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold82 hold82/A VGND VGND VPWR VPWR hold82/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 hold93/A VGND VGND VPWR VPWR hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_35_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4430_ _4495_/A _4738_/A VGND VGND VPWR VPWR _4931_/B sky130_fd_sc_hd__nor2_2
XANTENNA_2 _5828_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4361_ _4412_/A1 _4359_/B _4360_/B _4591_/A VGND VGND VPWR VPWR _4426_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6100_ _6100_/A1 _6197_/A2 _6197_/B1 _6100_/B2 _6099_/X VGND VGND VPWR VPWR _6110_/A
+ sky130_fd_sc_hd__a221o_1
X_3312_ _3324_/A _3466_/A VGND VGND VPWR VPWR _3312_/Y sky130_fd_sc_hd__nor2_1
X_7080_ _7080_/CLK _7080_/D fanout3986/X VGND VGND VPWR VPWR _7080_/Q sky130_fd_sc_hd__dfrtp_1
X_4292_ _4304_/A0 hold127/X _4293_/S VGND VGND VPWR VPWR _4292_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6031_ _6031_/A1 _6054_/B1 _6031_/B1 _6031_/B2 VGND VGND VPWR VPWR _6031_/X sky130_fd_sc_hd__a22o_1
X_3243_ hold60/X _3820_/A hold158/X VGND VGND VPWR VPWR _3243_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_86_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6933_ _7031_/CLK _6933_/D wire4044/X VGND VGND VPWR VPWR _6933_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6864_ _7109_/CLK _6864_/D wire3999/A VGND VGND VPWR VPWR _6864_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_179_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5815_ _5859_/A1 _7166_/Q wire463/X VGND VGND VPWR VPWR _5815_/X sky130_fd_sc_hd__a21o_1
XFILLER_179_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6795_ _6799_/CLK _6795_/D wire3935/A VGND VGND VPWR VPWR _6795_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_50_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5746_ _6075_/B2 _5784_/A2 _5746_/B1 _6081_/A1 VGND VGND VPWR VPWR _5746_/X sky130_fd_sc_hd__a22o_1
XFILLER_182_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5677_ _5693_/A _5703_/C _5699_/C VGND VGND VPWR VPWR _5677_/X sky130_fd_sc_hd__and3_1
XFILLER_157_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4628_ _4675_/A _4646_/B VGND VGND VPWR VPWR _5083_/A sky130_fd_sc_hd__nor2_1
XFILLER_135_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire4206 input43/X VGND VGND VPWR VPWR wire4206/X sky130_fd_sc_hd__clkbuf_1
Xwire4217 wire4218/X VGND VGND VPWR VPWR _3931_/A1 sky130_fd_sc_hd__clkbuf_1
Xhold530 _6895_/Q VGND VGND VPWR VPWR hold530/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire4228 _3751_/B2 VGND VGND VPWR VPWR wire4228/X sky130_fd_sc_hd__clkbuf_1
XFILLER_151_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4559_ _4560_/A _4573_/B VGND VGND VPWR VPWR _4797_/A sky130_fd_sc_hd__and2_1
Xhold541 _6893_/Q VGND VGND VPWR VPWR hold541/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4239 wire4240/X VGND VGND VPWR VPWR _3406_/A1 sky130_fd_sc_hd__clkbuf_1
Xhold552 _7211_/Q VGND VGND VPWR VPWR hold552/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3505 _5539_/A1 VGND VGND VPWR VPWR _5452_/A0 sky130_fd_sc_hd__clkbuf_2
Xhold563 _6497_/Q VGND VGND VPWR VPWR hold563/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 _7109_/Q VGND VGND VPWR VPWR hold574/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3527 _4304_/A0 VGND VGND VPWR VPWR _4274_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3538 _5532_/A1 VGND VGND VPWR VPWR _6395_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold585 _6996_/Q VGND VGND VPWR VPWR hold585/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 _7027_/Q VGND VGND VPWR VPWR hold596/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire2804 _6172_/A2 VGND VGND VPWR VPWR _6124_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3549 _5514_/A0 VGND VGND VPWR VPWR _5469_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2815 wire2816/X VGND VGND VPWR VPWR _6212_/A2 sky130_fd_sc_hd__clkbuf_2
X_6229_ _6229_/A1 _6304_/A2 _6304_/B1 _6756_/Q _6228_/X VGND VGND VPWR VPWR _6232_/C
+ sky130_fd_sc_hd__a221o_1
Xwire2826 _5943_/B1 VGND VGND VPWR VPWR _5958_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2837 _5921_/B1 VGND VGND VPWR VPWR _5955_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2848 _5912_/B1 VGND VGND VPWR VPWR _5952_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout3944 wire3948/X VGND VGND VPWR VPWR fanout3944/X sky130_fd_sc_hd__buf_6
XFILLER_49_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout3977 wire3985/X VGND VGND VPWR VPWR wire3981/A sky130_fd_sc_hd__buf_6
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput150 wb_dat_i[26] VGND VGND VPWR VPWR _6370_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput161 wb_dat_i[7] VGND VGND VPWR VPWR _6385_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3930_ _6555_/Q _6790_/Q _6432_/B VGND VGND VPWR VPWR _3930_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3861_ _6450_/Q hold42/A _3866_/S VGND VGND VPWR VPWR _6451_/D sky130_fd_sc_hd__mux2_1
XFILLER_149_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5600_ _7144_/Q _7145_/Q VGND VGND VPWR VPWR _5600_/Y sky130_fd_sc_hd__nand2_1
XFILLER_176_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6580_ _6945_/CLK _6580_/D fanout4078/X VGND VGND VPWR VPWR _6580_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_32_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3792_ _6783_/Q _3791_/B wire358/X _3791_/Y VGND VGND VPWR VPWR _6783_/D sky130_fd_sc_hd__a22o_1
XFILLER_192_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5531_ hold693/X _5531_/A1 _5534_/S VGND VGND VPWR VPWR _7091_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5462_ _5462_/A0 hold593/X _5462_/S VGND VGND VPWR VPWR _7030_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7201_ _7204_/CLK _7201_/D wire4260/X VGND VGND VPWR VPWR _7201_/Q sky130_fd_sc_hd__dfrtp_1
X_4413_ _4544_/B _4538_/B _4435_/A VGND VGND VPWR VPWR _4434_/B sky130_fd_sc_hd__a21boi_1
XFILLER_133_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5393_ _5528_/A0 hold134/X _5393_/S VGND VGND VPWR VPWR _6969_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7132_ _7132_/CLK _7132_/D fanout4077/X VGND VGND VPWR VPWR _7132_/Q sky130_fd_sc_hd__dfrtp_1
X_4344_ _4419_/B _4450_/A VGND VGND VPWR VPWR _4596_/B sky130_fd_sc_hd__or2_1
XFILLER_99_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7063_ _7133_/CLK _7063_/D fanout4073/X VGND VGND VPWR VPWR _7063_/Q sky130_fd_sc_hd__dfrtp_1
X_4275_ hold223/X _4305_/A0 _4275_/S VGND VGND VPWR VPWR _6725_/D sky130_fd_sc_hd__mux2_1
XFILLER_98_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6014_ _6014_/A _6039_/A _6020_/C VGND VGND VPWR VPWR _6014_/X sky130_fd_sc_hd__and3_1
X_3226_ _3226_/A VGND VGND VPWR VPWR _3226_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6916_ _7142_/CLK _6916_/D wire4039/X VGND VGND VPWR VPWR _6916_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6847_ _6921_/CLK _6847_/D wire4046/X VGND VGND VPWR VPWR _6847_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6778_ _7204_/CLK _6778_/D wire4261/X VGND VGND VPWR VPWR _6778_/Q sky130_fd_sc_hd__dfrtp_1
Xwire707 _5255_/S VGND VGND VPWR VPWR _5253_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire718 _4139_/S VGND VGND VPWR VPWR _4140_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire729 _4014_/S VGND VGND VPWR VPWR _4015_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_148_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5729_ _6070_/A1 _5729_/A2 _5719_/X wire996/X _5729_/C1 VGND VGND VPWR VPWR _5729_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_6_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4014 wire4015/X VGND VGND VPWR VPWR wire4014/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3313 _5074_/A2 VGND VGND VPWR VPWR _4613_/B sky130_fd_sc_hd__clkbuf_2
Xhold360 _6755_/Q VGND VGND VPWR VPWR hold360/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire4058 wire4058/A VGND VGND VPWR VPWR wire4058/X sky130_fd_sc_hd__buf_2
Xhold371 _6729_/Q VGND VGND VPWR VPWR hold371/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 _6775_/Q VGND VGND VPWR VPWR hold382/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4069 wire4069/A VGND VGND VPWR VPWR wire4069/X sky130_fd_sc_hd__clkbuf_4
Xhold393 _7132_/Q VGND VGND VPWR VPWR hold393/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3335 _4609_/A VGND VGND VPWR VPWR _5105_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire2601 _4670_/Y VGND VGND VPWR VPWR _4771_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire3346 _4739_/A VGND VGND VPWR VPWR _4520_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3357 _4689_/A VGND VGND VPWR VPWR _5023_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2612 _4362_/Y VGND VGND VPWR VPWR _4957_/A sky130_fd_sc_hd__clkbuf_1
Xwire3368 _4363_/B VGND VGND VPWR VPWR _4428_/B sky130_fd_sc_hd__clkbuf_1
Xwire2623 _6040_/X VGND VGND VPWR VPWR wire2623/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3379 _5519_/A0 VGND VGND VPWR VPWR _3991_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2634 _6186_/B1 VGND VGND VPWR VPWR _6207_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1900 _6945_/Q VGND VGND VPWR VPWR wire1900/X sky130_fd_sc_hd__clkbuf_1
Xwire2645 _6036_/X VGND VGND VPWR VPWR _6181_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire1911 _6939_/Q VGND VGND VPWR VPWR _6061_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire2667 _6191_/B1 VGND VGND VPWR VPWR wire2667/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1922 wire1923/X VGND VGND VPWR VPWR _6048_/B2 sky130_fd_sc_hd__clkbuf_2
Xwire2678 wire2679/X VGND VGND VPWR VPWR _6200_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire1933 wire1934/X VGND VGND VPWR VPWR _6179_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1944 _5344_/A1 VGND VGND VPWR VPWR _5764_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire2689 _6024_/D VGND VGND VPWR VPWR wire2689/X sky130_fd_sc_hd__clkbuf_1
XFILLER_133_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1955 wire1956/X VGND VGND VPWR VPWR _3442_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_46_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1966 _6913_/Q VGND VGND VPWR VPWR _6203_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1977 _6908_/Q VGND VGND VPWR VPWR wire1977/X sky130_fd_sc_hd__clkbuf_1
Xwire1988 _6901_/Q VGND VGND VPWR VPWR _6103_/A1 sky130_fd_sc_hd__clkbuf_2
Xwire1999 _3529_/A1 VGND VGND VPWR VPWR wire1999/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3880 wire3881/X VGND VGND VPWR VPWR wire3880/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4060_ hold296/X _4115_/A0 _4060_/S VGND VGND VPWR VPWR _4060_/X sky130_fd_sc_hd__mux2_1
Xwire3891 wire3892/X VGND VGND VPWR VPWR _3949_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_95_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4962_ _5068_/B _4962_/B VGND VGND VPWR VPWR _4962_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3913_ _6445_/Q _6541_/Q _3834_/B _6545_/Q VGND VGND VPWR VPWR _6545_/D sky130_fd_sc_hd__a31o_1
X_6701_ _6701_/CLK _6701_/D wire3959/A VGND VGND VPWR VPWR _6701_/Q sky130_fd_sc_hd__dfrtp_1
X_4893_ _4524_/B _4871_/Y _4892_/X VGND VGND VPWR VPWR _4894_/B sky130_fd_sc_hd__a21o_1
X_6632_ _7196_/CLK _6632_/D VGND VGND VPWR VPWR _6632_/Q sky130_fd_sc_hd__dfxtp_1
X_3844_ _6473_/Q _6472_/Q _6471_/Q _6541_/Q VGND VGND VPWR VPWR _3845_/S sky130_fd_sc_hd__or4b_1
XFILLER_192_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6563_ _7180_/CLK _6563_/D _6562_/SET_B VGND VGND VPWR VPWR _6563_/Q sky130_fd_sc_hd__dfrtp_1
X_3775_ _6798_/Q _3417_/Y _5529_/A _7090_/Q VGND VGND VPWR VPWR _3775_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5514_ _5514_/A0 hold561/X _5514_/S VGND VGND VPWR VPWR _7076_/D sky130_fd_sc_hd__mux2_1
XFILLER_192_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6494_ _6825_/CLK _6494_/D _6495_/SET_B VGND VGND VPWR VPWR _6494_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_173_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5445_ _5481_/A0 hold645/X _5447_/S VGND VGND VPWR VPWR _7015_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5376_ _5376_/A _5553_/B VGND VGND VPWR VPWR _5376_/Y sky130_fd_sc_hd__nand2_1
XFILLER_154_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7115_ _7115_/CLK _7115_/D _7185_/RESET_B VGND VGND VPWR VPWR _7115_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4327_ hold549/X _4327_/A1 _4328_/S VGND VGND VPWR VPWR _6768_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1218 _3548_/A2 VGND VGND VPWR VPWR _5349_/A sky130_fd_sc_hd__clkbuf_1
X_7046_ _7046_/CLK _7046_/D wire4037/X VGND VGND VPWR VPWR _7046_/Q sky130_fd_sc_hd__dfrtp_1
X_4258_ _4258_/A _5223_/B VGND VGND VPWR VPWR _4263_/S sky130_fd_sc_hd__and2_2
Xwire1229 _3310_/Y VGND VGND VPWR VPWR _3568_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
X_3209_ hold95/A VGND VGND VPWR VPWR _3209_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4189_ _6694_/Q _4189_/B VGND VGND VPWR VPWR _4197_/S sky130_fd_sc_hd__and2_1
XFILLER_28_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire504 _5298_/S VGND VGND VPWR VPWR _5303_/S sky130_fd_sc_hd__buf_2
XFILLER_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire548 _3683_/X VGND VGND VPWR VPWR wire548/X sky130_fd_sc_hd__clkbuf_1
Xwire559 _3575_/X VGND VGND VPWR VPWR _3582_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_578 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3110 _5966_/A2 VGND VGND VPWR VPWR _5936_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_151_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3121 _5906_/A2 VGND VGND VPWR VPWR _5953_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire3132 wire3133/X VGND VGND VPWR VPWR _5928_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_151_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold190 _6746_/Q VGND VGND VPWR VPWR hold190/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3143 _5758_/A2 VGND VGND VPWR VPWR _5787_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_120_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3154 _6323_/A2 VGND VGND VPWR VPWR _6247_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire2420 _3523_/A1 VGND VGND VPWR VPWR _5782_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire3165 _4692_/B VGND VGND VPWR VPWR _4675_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2431 _6500_/Q VGND VGND VPWR VPWR wire2431/X sky130_fd_sc_hd__clkbuf_1
Xwire2442 _6489_/Q VGND VGND VPWR VPWR wire2442/X sky130_fd_sc_hd__clkbuf_1
XFILLER_120_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire3187 _4688_/B VGND VGND VPWR VPWR _5016_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2453 _6390_/X VGND VGND VPWR VPWR wire2453/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2464 _6178_/B1 VGND VGND VPWR VPWR _6132_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire1730 _6151_/A1 VGND VGND VPWR VPWR _3423_/B2 sky130_fd_sc_hd__clkbuf_1
Xwire2486 _6025_/C VGND VGND VPWR VPWR _6189_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1741 wire1742/X VGND VGND VPWR VPWR _6005_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire2497 _6278_/B1 VGND VGND VPWR VPWR _6304_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1763 _7019_/Q VGND VGND VPWR VPWR _6055_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1774 _5762_/B2 VGND VGND VPWR VPWR wire1774/X sky130_fd_sc_hd__clkbuf_1
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1785 wire1786/X VGND VGND VPWR VPWR wire1785/X sky130_fd_sc_hd__clkbuf_1
Xwire1796 _6128_/B2 VGND VGND VPWR VPWR _3533_/A1 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_8_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _7211_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_160_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3560_ _3560_/A1 _3617_/A2 _3786_/B1 _6764_/Q VGND VGND VPWR VPWR _3560_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3491_ _6715_/Q _4258_/A wire820/A _3491_/B2 wire566/X VGND VGND VPWR VPWR _3491_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_142_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5230_ _5212_/C hold335/X _5231_/S VGND VGND VPWR VPWR _6824_/D sky130_fd_sc_hd__mux2_1
XFILLER_154_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5161_ _4614_/A _5161_/A2 _4490_/X VGND VGND VPWR VPWR _5162_/D sky130_fd_sc_hd__o21ai_1
XFILLER_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4112_ _5242_/A0 hold341/X _4115_/S VGND VGND VPWR VPWR _6580_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5092_ _5119_/A _5119_/B _5092_/C _5092_/D VGND VGND VPWR VPWR _5102_/A sky130_fd_sc_hd__or4_1
XFILLER_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4043_ _4285_/A0 hold439/X _4045_/S VGND VGND VPWR VPWR _6533_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5994_ _6040_/A _6039_/A _6040_/B VGND VGND VPWR VPWR _5994_/X sky130_fd_sc_hd__and3_1
X_4945_ _4419_/B _4483_/A _4944_/X _4839_/A _4847_/A VGND VGND VPWR VPWR _4945_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_178_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4876_ _4876_/A _4876_/B VGND VGND VPWR VPWR _4887_/D sky130_fd_sc_hd__nand2_1
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length3107 _5781_/A2 VGND VGND VPWR VPWR wire3102/A sky130_fd_sc_hd__clkbuf_1
Xmax_length3118 wire3119/X VGND VGND VPWR VPWR _5756_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_138_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6615_ _6702_/CLK _6615_/D wire3958/X VGND VGND VPWR VPWR _6615_/Q sky130_fd_sc_hd__dfrtp_1
X_3827_ _3807_/B _3820_/A _3820_/Y _3826_/X VGND VGND VPWR VPWR _3827_/X sky130_fd_sc_hd__a22o_1
XFILLER_137_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6546_ _6945_/CLK _6546_/D fanout4078/X VGND VGND VPWR VPWR _6546_/Q sky130_fd_sc_hd__dfrtp_1
X_3758_ _6031_/A1 wire858/X wire820/X _3758_/B2 _3728_/X VGND VGND VPWR VPWR _3760_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_192_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6477_ _6824_/CLK _6477_/D fanout3973/X VGND VGND VPWR VPWR _6477_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_106_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3689_ _3689_/A _3689_/B VGND VGND VPWR VPWR _3723_/B sky130_fd_sc_hd__or2_1
XFILLER_160_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5428_ _5491_/A0 hold505/X _5429_/S VGND VGND VPWR VPWR _7000_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput240 _6576_/Q VGND VGND VPWR VPWR mgmt_gpio_out[34] sky130_fd_sc_hd__buf_12
Xoutput251 _3945_/X VGND VGND VPWR VPWR pad_flash_clk sky130_fd_sc_hd__clkbuf_1
Xoutput262 _6802_/Q VGND VGND VPWR VPWR pll90_sel[1] sky130_fd_sc_hd__buf_12
Xoutput273 _6799_/Q VGND VGND VPWR VPWR pll_sel[1] sky130_fd_sc_hd__buf_12
X_5359_ _5359_/A0 hold325/X _5361_/S VGND VGND VPWR VPWR _6938_/D sky130_fd_sc_hd__mux2_1
Xoutput284 _6476_/Q VGND VGND VPWR VPWR pll_trim[18] sky130_fd_sc_hd__buf_12
Xoutput295 _6494_/Q VGND VGND VPWR VPWR pll_trim[4] sky130_fd_sc_hd__buf_12
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1004 _6319_/S VGND VGND VPWR VPWR _6171_/S sky130_fd_sc_hd__buf_2
XFILLER_87_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1015 _4947_/Y VGND VGND VPWR VPWR _5064_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1026 _3783_/B1 VGND VGND VPWR VPWR wire1026/X sky130_fd_sc_hd__clkbuf_1
XFILLER_102_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1037 _3526_/Y VGND VGND VPWR VPWR _5187_/A sky130_fd_sc_hd__clkbuf_2
X_7029_ _7130_/CLK _7029_/D wire4058/A VGND VGND VPWR VPWR hold92/A sky130_fd_sc_hd__dfrtp_1
XFILLER_74_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1059 _3489_/Y VGND VGND VPWR VPWR _4258_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire356 _3375_/X VGND VGND VPWR VPWR wire356/X sky130_fd_sc_hd__clkbuf_1
XFILLER_99_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire367 wire368/X VGND VGND VPWR VPWR wire367/X sky130_fd_sc_hd__clkbuf_2
Xwire378 wire379/X VGND VGND VPWR VPWR wire378/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire389 wire390/X VGND VGND VPWR VPWR _3447_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire2250 _5915_/A1 VGND VGND VPWR VPWR wire2250/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2272 _6671_/Q VGND VGND VPWR VPWR _6261_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2283 wire2284/X VGND VGND VPWR VPWR _3629_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_93_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1560 wire1561/X VGND VGND VPWR VPWR _6135_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire1571 wire1572/X VGND VGND VPWR VPWR wire1571/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1593 _7094_/Q VGND VGND VPWR VPWR _6323_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4730_ _4753_/A _5002_/A VGND VGND VPWR VPWR _4815_/A sky130_fd_sc_hd__nor2_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4661_ _4677_/A _4661_/B VGND VGND VPWR VPWR _4704_/B sky130_fd_sc_hd__or2_1
XFILLER_147_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6400_ _6433_/A _6433_/B VGND VGND VPWR VPWR _6400_/X sky130_fd_sc_hd__and2_1
X_3612_ _5738_/B2 _3612_/A2 wire825/X _3612_/B2 VGND VGND VPWR VPWR _3612_/X sky130_fd_sc_hd__a22o_1
X_4592_ _4592_/A VGND VGND VPWR VPWR _4592_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6331_ _6331_/A _6331_/B _6331_/C _6331_/D VGND VGND VPWR VPWR _6332_/C sky130_fd_sc_hd__or4_1
X_3543_ _3543_/A _3543_/B _3543_/C VGND VGND VPWR VPWR _3543_/X sky130_fd_sc_hd__or3_2
X_6262_ _6262_/A1 _6262_/A2 _6262_/B1 _6262_/B2 VGND VGND VPWR VPWR _6262_/X sky130_fd_sc_hd__a22o_1
X_3474_ _3546_/A _3528_/B VGND VGND VPWR VPWR _3474_/Y sky130_fd_sc_hd__nor2_1
XFILLER_143_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5213_ hold350/X _3727_/Y _5229_/B _5212_/X VGND VGND VPWR VPWR _6812_/D sky130_fd_sc_hd__o211a_1
X_6193_ _6193_/A _6193_/B _6193_/C VGND VGND VPWR VPWR _6193_/X sky130_fd_sc_hd__or3_1
XFILLER_142_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5144_ _4794_/A _5143_/Y _4810_/C _5144_/C1 VGND VGND VPWR VPWR _5144_/X sky130_fd_sc_hd__o211a_1
XFILLER_97_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5075_ _5018_/A _5074_/X _5028_/X _5013_/X _4911_/X VGND VGND VPWR VPWR _5156_/B
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_111_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4026_ hold322/X _4139_/A1 _4027_/S VGND VGND VPWR VPWR _4026_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5977_ _6014_/A _6039_/A _6040_/B VGND VGND VPWR VPWR _5977_/X sky130_fd_sc_hd__and3_1
X_4928_ _6362_/A _4928_/B _4928_/C _4928_/D VGND VGND VPWR VPWR _4928_/X sky130_fd_sc_hd__or4_1
XFILLER_33_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4859_ _4660_/B _4581_/X _4858_/X _4504_/A VGND VGND VPWR VPWR _4860_/D sky130_fd_sc_hd__o211a_1
XFILLER_166_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length1502 _3414_/Y VGND VGND VPWR VPWR _3415_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_119_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6529_ _6811_/CLK _6529_/D wire3935/X VGND VGND VPWR VPWR _6529_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_length1546 hold196/X VGND VGND VPWR VPWR _3198_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_134_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_730 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_73_csclk _7117_/CLK VGND VGND VPWR VPWR _6770_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_102_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_11_csclk _7059_/CLK VGND VGND VPWR VPWR _7112_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_11_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3460 _5558_/A0 VGND VGND VPWR VPWR _5462_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_109_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_26_csclk _7059_/CLK VGND VGND VPWR VPWR _7136_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_125_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3190_ _3850_/A VGND VGND VPWR VPWR _3190_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2080 wire2081/X VGND VGND VPWR VPWR wire2080/X sky130_fd_sc_hd__clkbuf_1
Xwire2091 _6849_/Q VGND VGND VPWR VPWR _6218_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1390 _3285_/Y VGND VGND VPWR VPWR _3714_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_19_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5900_ _5900_/A1 _5906_/A2 _5965_/B1 _5900_/B2 _5899_/X VGND VGND VPWR VPWR _5901_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6880_ _7140_/CLK _6880_/D _7138_/RESET_B VGND VGND VPWR VPWR _6880_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5831_ _5831_/A1 _5831_/A2 _5831_/B1 _6173_/B2 VGND VGND VPWR VPWR _5831_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5762_ _6104_/A1 _5853_/B1 _5762_/B1 _5762_/B2 _5761_/X VGND VGND VPWR VPWR _5771_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4713_ _4713_/A _4713_/B _4713_/C _4713_/D VGND VGND VPWR VPWR _4713_/Y sky130_fd_sc_hd__nand4_1
X_5693_ _5693_/A _5706_/B _5700_/C VGND VGND VPWR VPWR _5693_/X sky130_fd_sc_hd__and3_1
XFILLER_147_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4644_ _5059_/A _4644_/B _4644_/C _4643_/X VGND VGND VPWR VPWR _4647_/B sky130_fd_sc_hd__or4b_1
XFILLER_163_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold701 _6807_/Q VGND VGND VPWR VPWR hold701/X sky130_fd_sc_hd__dlygate4sd3_1
X_4575_ _4591_/A _4575_/B _4621_/C VGND VGND VPWR VPWR _4575_/X sky130_fd_sc_hd__or3_1
XFILLER_162_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold712 _6477_/Q VGND VGND VPWR VPWR hold712/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold723 _6781_/Q VGND VGND VPWR VPWR hold723/X sky130_fd_sc_hd__dlygate4sd3_1
X_3526_ _3526_/A _3714_/B VGND VGND VPWR VPWR _3526_/Y sky130_fd_sc_hd__nor2_1
X_6314_ _6314_/A1 _6314_/A2 _6314_/B1 _6314_/B2 _6298_/X VGND VGND VPWR VPWR _6315_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3709 wire3709/A VGND VGND VPWR VPWR wire3709/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6245_ _7183_/Q _6319_/S wire448/X _6244_/X VGND VGND VPWR VPWR _7183_/D sky130_fd_sc_hd__o22a_1
X_3457_ _3457_/A1 _3327_/Y _4282_/A _6735_/Q VGND VGND VPWR VPWR _3457_/X sky130_fd_sc_hd__a22o_1
XFILLER_103_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6176_ _7141_/Q _6023_/B _6176_/B1 _6176_/B2 VGND VGND VPWR VPWR _6176_/X sky130_fd_sc_hd__a22o_1
XFILLER_162_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3388_ _5834_/B2 _3557_/A2 wire877/X _3388_/B2 _3387_/X VGND VGND VPWR VPWR _3392_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_57_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5127_ _5127_/A _5127_/B _5127_/C VGND VGND VPWR VPWR _5159_/B sky130_fd_sc_hd__nor3_1
XFILLER_69_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5058_ _4397_/A _4951_/B _4846_/D VGND VGND VPWR VPWR _5059_/C sky130_fd_sc_hd__o21a_1
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4009_ _5429_/A0 hold529/X _4009_/S VGND VGND VPWR VPWR _6505_/D sky130_fd_sc_hd__mux2_1
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length1343 _4488_/B VGND VGND VPWR VPWR _5133_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_4_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_length1398 hold244/X VGND VGND VPWR VPWR wire1394/A sky130_fd_sc_hd__clkbuf_1
XFILLER_161_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold50 hold50/A VGND VGND VPWR VPWR hold50/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold61 hold61/A VGND VGND VPWR VPWR hold61/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold72 hold72/A VGND VGND VPWR VPWR hold72/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold83/A VGND VGND VPWR VPWR hold83/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 hold94/A VGND VGND VPWR VPWR hold94/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_mgmt_gpio_in[4] clkbuf_2_3_0_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR _3487_/B2
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_189_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_3 mgmt_gpio_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4360_ _4360_/A _4360_/B VGND VGND VPWR VPWR _4462_/B sky130_fd_sc_hd__or2_1
X_3311_ hold85/A _3511_/B VGND VGND VPWR VPWR _3311_/Y sky130_fd_sc_hd__nor2_1
XFILLER_98_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4291_ hold22/X _6738_/Q _4293_/S VGND VGND VPWR VPWR hold23/A sky130_fd_sc_hd__mux2_1
XFILLER_140_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6030_ _6033_/A _6040_/B _6030_/C VGND VGND VPWR VPWR _6030_/X sky130_fd_sc_hd__and3_1
X_3242_ _3242_/A _3252_/B VGND VGND VPWR VPWR _3242_/X sky130_fd_sc_hd__and2_1
XFILLER_67_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6932_ _7131_/CLK _6932_/D wire4061/A VGND VGND VPWR VPWR _6932_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6863_ _7017_/CLK _6863_/D wire4081/X VGND VGND VPWR VPWR _6863_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5814_ _6169_/A1 _5814_/A2 _5804_/X wire993/X _6169_/C1 VGND VGND VPWR VPWR _5814_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6794_ _6811_/CLK _6794_/D wire3935/A VGND VGND VPWR VPWR _6794_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5745_ _6074_/B2 _5745_/A2 _5745_/B1 _6900_/Q _5744_/X VGND VGND VPWR VPWR _5750_/B
+ sky130_fd_sc_hd__a221o_1
Xmax_length509 _5273_/S VGND VGND VPWR VPWR wire508/A sky130_fd_sc_hd__clkbuf_1
X_5676_ _7152_/Q _5703_/C _5699_/C VGND VGND VPWR VPWR _5676_/X sky130_fd_sc_hd__and3_1
XFILLER_148_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4627_ _4986_/A _5115_/B _4627_/C _5177_/A VGND VGND VPWR VPWR _4634_/A sky130_fd_sc_hd__or4_1
XFILLER_135_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4207 wire4208/X VGND VGND VPWR VPWR _3350_/B2 sky130_fd_sc_hd__clkbuf_1
Xhold520 _6959_/Q VGND VGND VPWR VPWR hold520/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4558_ _4802_/B _4609_/B VGND VGND VPWR VPWR _4778_/B sky130_fd_sc_hd__nor2_1
Xwire4218 wire4219/X VGND VGND VPWR VPWR wire4218/X sky130_fd_sc_hd__clkbuf_1
Xhold531 _6991_/Q VGND VGND VPWR VPWR hold531/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire4229 wire4230/X VGND VGND VPWR VPWR _3751_/B2 sky130_fd_sc_hd__clkbuf_2
Xhold542 _7072_/Q VGND VGND VPWR VPWR hold542/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold553 _6576_/Q VGND VGND VPWR VPWR hold553/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3506 _5254_/A1 VGND VGND VPWR VPWR _5539_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold564 _6495_/Q VGND VGND VPWR VPWR hold564/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 _7080_/Q VGND VGND VPWR VPWR hold575/X sky130_fd_sc_hd__dlygate4sd3_1
X_3509_ _7099_/Q _3605_/A2 _3509_/B1 _3509_/B2 wire810/X VGND VGND VPWR VPWR _3515_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3528 _5281_/A0 VGND VGND VPWR VPWR _4304_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold586 _7090_/Q VGND VGND VPWR VPWR hold586/X sky130_fd_sc_hd__dlygate4sd3_1
X_4489_ _4489_/A _4932_/A _4942_/B VGND VGND VPWR VPWR _4489_/X sky130_fd_sc_hd__or3_1
Xwire3539 wire3539/A VGND VGND VPWR VPWR _4327_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_104_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold597 _6967_/Q VGND VGND VPWR VPWR hold597/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire2805 _6199_/A2 VGND VGND VPWR VPWR _6172_/A2 sky130_fd_sc_hd__clkbuf_2
Xwire2816 _5982_/X VGND VGND VPWR VPWR wire2816/X sky130_fd_sc_hd__clkbuf_1
X_6228_ _6228_/A1 _6277_/A2 _6303_/B1 _6228_/B2 VGND VGND VPWR VPWR _6228_/X sky130_fd_sc_hd__a22o_1
Xwire2827 _5707_/B1 VGND VGND VPWR VPWR _5943_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire2838 _5738_/B1 VGND VGND VPWR VPWR _5921_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire2849 wire2850/X VGND VGND VPWR VPWR _5912_/B1 sky130_fd_sc_hd__clkbuf_2
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ _6919_/Q _6159_/A2 _6159_/B1 _6943_/Q VGND VGND VPWR VPWR _6159_/X sky130_fd_sc_hd__a22o_1
XFILLER_57_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length1140 _5493_/A VGND VGND VPWR VPWR _3522_/B1 sky130_fd_sc_hd__clkbuf_1
Xfanout3934 _3946_/B VGND VGND VPWR VPWR wire3935/A sky130_fd_sc_hd__buf_6
XFILLER_107_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout3967 wire4022/X VGND VGND VPWR VPWR wire3970/A sky130_fd_sc_hd__clkbuf_1
XFILLER_68_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput140 wb_dat_i[17] VGND VGND VPWR VPWR _6367_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput151 wb_dat_i[27] VGND VGND VPWR VPWR _6373_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput162 wb_dat_i[8] VGND VGND VPWR VPWR _6364_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3860_ hold42/A hold1/A _3866_/S VGND VGND VPWR VPWR _6452_/D sky130_fd_sc_hd__mux2_1
XFILLER_32_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3791_ _3791_/A _3791_/B VGND VGND VPWR VPWR _3791_/Y sky130_fd_sc_hd__nor2_1
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5530_ hold586/X _5530_/A1 _5533_/S VGND VGND VPWR VPWR _7090_/D sky130_fd_sc_hd__mux2_1
XFILLER_75_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5461_ _5479_/A0 hold92/X _5461_/S VGND VGND VPWR VPWR _7029_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7200_ _7204_/CLK _7200_/D wire4260/X VGND VGND VPWR VPWR _7200_/Q sky130_fd_sc_hd__dfrtp_1
X_4412_ _4412_/A1 _4538_/B _4379_/A VGND VGND VPWR VPWR _4435_/A sky130_fd_sc_hd__a21o_1
XFILLER_172_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5392_ _5392_/A0 hold429/X _5393_/S VGND VGND VPWR VPWR _6968_/D sky130_fd_sc_hd__mux2_1
X_7131_ _7131_/CLK _7131_/D wire4058/A VGND VGND VPWR VPWR _7131_/Q sky130_fd_sc_hd__dfrtp_1
X_4343_ _4846_/B _4398_/C VGND VGND VPWR VPWR _4596_/A sky130_fd_sc_hd__nand2_2
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7062_ _7075_/CLK _7062_/D _7075_/SET_B VGND VGND VPWR VPWR _7062_/Q sky130_fd_sc_hd__dfrtp_1
X_4274_ hold253/X _4274_/A1 _4275_/S VGND VGND VPWR VPWR _6724_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6013_ _6040_/A _6020_/C _6040_/C VGND VGND VPWR VPWR _6027_/C sky130_fd_sc_hd__and3_1
XFILLER_113_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3225_ _6917_/Q VGND VGND VPWR VPWR _3225_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6915_ _6939_/CLK _6915_/D _7042_/SET_B VGND VGND VPWR VPWR _6915_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_23_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6846_ _7102_/CLK _6846_/D _7176_/RESET_B VGND VGND VPWR VPWR _6846_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6777_ _7204_/CLK _6777_/D wire4261/X VGND VGND VPWR VPWR _6777_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3989_ hold708/X _5436_/A0 _3991_/S VGND VGND VPWR VPWR _6487_/D sky130_fd_sc_hd__mux2_1
XFILLER_139_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire719 wire720/X VGND VGND VPWR VPWR _4127_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_109_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5728_ _5728_/A _5728_/B _5728_/C _5728_/D VGND VGND VPWR VPWR _5728_/X sky130_fd_sc_hd__or4_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5659_ _5688_/A _5699_/B _5706_/C VGND VGND VPWR VPWR _5659_/X sky130_fd_sc_hd__and3_1
XFILLER_191_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4004 wire4004/A VGND VGND VPWR VPWR wire4004/X sky130_fd_sc_hd__clkbuf_2
XFILLER_151_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4015 wire4016/X VGND VGND VPWR VPWR wire4015/X sky130_fd_sc_hd__clkbuf_2
XFILLER_123_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4026 wire4026/A VGND VGND VPWR VPWR wire4026/X sky130_fd_sc_hd__clkbuf_4
Xhold350 _6812_/Q VGND VGND VPWR VPWR hold350/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire4037 _6401_/A VGND VGND VPWR VPWR wire4037/X sky130_fd_sc_hd__buf_2
Xhold361 _6521_/Q VGND VGND VPWR VPWR hold361/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire4048 wire4049/X VGND VGND VPWR VPWR wire4048/X sky130_fd_sc_hd__buf_2
Xwire3303 _4621_/X VGND VGND VPWR VPWR _4639_/B sky130_fd_sc_hd__buf_2
XFILLER_116_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3314 _4592_/A VGND VGND VPWR VPWR _4707_/A sky130_fd_sc_hd__clkbuf_2
Xwire3325 _4565_/X VGND VGND VPWR VPWR _4784_/A sky130_fd_sc_hd__clkbuf_2
Xhold372 _6721_/Q VGND VGND VPWR VPWR hold372/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3336 _4538_/Y VGND VGND VPWR VPWR _4609_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold383 _7070_/Q VGND VGND VPWR VPWR hold383/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 _6667_/Q VGND VGND VPWR VPWR hold394/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire2602 wire2603/X VGND VGND VPWR VPWR wire2602/X sky130_fd_sc_hd__clkbuf_1
XFILLER_117_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3347 _4662_/B VGND VGND VPWR VPWR _4674_/A sky130_fd_sc_hd__clkbuf_2
Xwire3358 _4492_/A VGND VGND VPWR VPWR _4689_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2613 _3833_/S VGND VGND VPWR VPWR _3828_/S sky130_fd_sc_hd__buf_2
Xwire3369 _4197_/S VGND VGND VPWR VPWR _4196_/S sky130_fd_sc_hd__buf_2
Xwire2635 _6039_/X VGND VGND VPWR VPWR _6186_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire1901 _6944_/Q VGND VGND VPWR VPWR _6172_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2646 _6326_/B1 VGND VGND VPWR VPWR _6255_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire1912 wire1913/X VGND VGND VPWR VPWR _5707_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_58_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2657 _6188_/B1 VGND VGND VPWR VPWR _6205_/B1 sky130_fd_sc_hd__clkbuf_2
Xwire2668 _6030_/X VGND VGND VPWR VPWR _6191_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1923 _6931_/Q VGND VGND VPWR VPWR wire1923/X sky130_fd_sc_hd__clkbuf_1
Xwire2679 _6020_/X VGND VGND VPWR VPWR wire2679/X sky130_fd_sc_hd__clkbuf_1
Xwire1934 wire1935/X VGND VGND VPWR VPWR wire1934/X sky130_fd_sc_hd__clkbuf_1
Xwire1945 hold203/X VGND VGND VPWR VPWR _5344_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire1956 wire1957/X VGND VGND VPWR VPWR wire1956/X sky130_fd_sc_hd__clkbuf_1
Xwire1967 _6912_/Q VGND VGND VPWR VPWR _6184_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1978 _6054_/B2 VGND VGND VPWR VPWR _3707_/A1 sky130_fd_sc_hd__clkbuf_1
Xwire1989 _6899_/Q VGND VGND VPWR VPWR _3691_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length873 _3339_/Y VGND VGND VPWR VPWR _3361_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_142_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3870 wire3871/X VGND VGND VPWR VPWR wire3870/X sky130_fd_sc_hd__clkbuf_1
Xwire3881 _3785_/A1 VGND VGND VPWR VPWR wire3881/X sky130_fd_sc_hd__clkbuf_1
Xwire3892 wire3893/X VGND VGND VPWR VPWR wire3892/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4961_ _4961_/A _4961_/B VGND VGND VPWR VPWR _4961_/Y sky130_fd_sc_hd__nor2_1
X_6700_ _7193_/CLK _6700_/D _6780_/RESET_B VGND VGND VPWR VPWR _6700_/Q sky130_fd_sc_hd__dfrtp_1
X_3912_ _6444_/Q _3868_/A _6541_/Q _3834_/B _6542_/Q VGND VGND VPWR VPWR _6542_/D
+ sky130_fd_sc_hd__a41o_1
XFILLER_51_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4892_ _4454_/Y _4871_/Y _5049_/C _4878_/X _4891_/X VGND VGND VPWR VPWR _4892_/X
+ sky130_fd_sc_hd__a2111o_1
X_6631_ _7196_/CLK _6631_/D VGND VGND VPWR VPWR _6631_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3843_ _3794_/B _3890_/A _3842_/Y _6541_/Q VGND VGND VPWR VPWR _6458_/D sky130_fd_sc_hd__a211oi_1
XFILLER_20_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3774_ _6243_/A1 _3496_/Y _3774_/B1 _6756_/Q _3773_/X VGND VGND VPWR VPWR _3781_/A
+ sky130_fd_sc_hd__a221o_1
X_6562_ _7187_/CLK _6562_/D _6562_/SET_B VGND VGND VPWR VPWR _6562_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_158_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5513_ _5513_/A0 hold229/X _5515_/S VGND VGND VPWR VPWR _7075_/D sky130_fd_sc_hd__mux2_1
XFILLER_185_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6493_ _6825_/CLK _6493_/D _6495_/SET_B VGND VGND VPWR VPWR _6493_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5444_ _5585_/A0 hold280/X _5444_/S VGND VGND VPWR VPWR _7014_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5375_ _5375_/A0 hold343/X _5375_/S VGND VGND VPWR VPWR _6953_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7114_ _7130_/CLK _7114_/D fanout4077/X VGND VGND VPWR VPWR _7114_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4326_ hold582/X _4326_/A1 _4329_/S VGND VGND VPWR VPWR _6767_/D sky130_fd_sc_hd__mux2_1
X_7045_ _7134_/CLK _7045_/D wire4058/A VGND VGND VPWR VPWR hold95/A sky130_fd_sc_hd__dfrtp_1
Xwire1208 _3596_/A2 VGND VGND VPWR VPWR _3383_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_59_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4257_ hold357/X _4263_/A1 _4257_/S VGND VGND VPWR VPWR _6710_/D sky130_fd_sc_hd__mux2_1
Xwire1219 _3615_/A2 VGND VGND VPWR VPWR _3548_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_101_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3208_ _7053_/Q VGND VGND VPWR VPWR _3208_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4188_ _6646_/Q wire378/X _4188_/S VGND VGND VPWR VPWR _6646_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6829_ _7130_/CLK _6829_/D _6833_/RESET_B VGND VGND VPWR VPWR _6829_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire505 _5291_/S VGND VGND VPWR VPWR _5294_/S sky130_fd_sc_hd__clkbuf_2
Xwire516 _5264_/S VGND VGND VPWR VPWR _5263_/S sky130_fd_sc_hd__clkbuf_2
Xwire527 _4104_/Y VGND VGND VPWR VPWR _4107_/S sky130_fd_sc_hd__clkbuf_1
Xmax_length3834 _6432_/B VGND VGND VPWR VPWR _6433_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_149_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire538 wire539/X VGND VGND VPWR VPWR wire538/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire549 _3673_/X VGND VGND VPWR VPWR _3679_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_183_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3100 _5663_/X VGND VGND VPWR VPWR _5843_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3111 _5922_/A2 VGND VGND VPWR VPWR _5966_/A2 sky130_fd_sc_hd__clkbuf_1
Xhold180 _7083_/Q VGND VGND VPWR VPWR hold180/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3122 _5748_/A2 VGND VGND VPWR VPWR _5906_/A2 sky130_fd_sc_hd__clkbuf_2
Xhold191 _7085_/Q VGND VGND VPWR VPWR hold191/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire3133 _5656_/X VGND VGND VPWR VPWR wire3133/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire3144 _5739_/A2 VGND VGND VPWR VPWR _5898_/A2 sky130_fd_sc_hd__clkbuf_1
Xwire2410 _6509_/Q VGND VGND VPWR VPWR _6302_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3155 wire3156/X VGND VGND VPWR VPWR _6323_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2421 _6502_/Q VGND VGND VPWR VPWR _3523_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2432 _6499_/Q VGND VGND VPWR VPWR _5711_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3177 _4611_/X VGND VGND VPWR VPWR _5024_/A sky130_fd_sc_hd__clkbuf_2
Xwire3188 _4688_/B VGND VGND VPWR VPWR _4721_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2443 _6489_/Q VGND VGND VPWR VPWR wire2443/X sky130_fd_sc_hd__clkbuf_2
Xwire3199 _4535_/B VGND VGND VPWR VPWR _4734_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2454 _6155_/B1 VGND VGND VPWR VPWR _6102_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire2465 _6038_/Y VGND VGND VPWR VPWR _6178_/B1 sky130_fd_sc_hd__clkbuf_1
Xwire1720 wire1721/X VGND VGND VPWR VPWR wire1720/X sky130_fd_sc_hd__clkbuf_1
XFILLER_144_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1731 _7031_/Q VGND VGND VPWR VPWR _6151_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2476 _6027_/D VGND VGND VPWR VPWR _6182_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2487 _6337_/B1 VGND VGND VPWR VPWR _6284_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1742 wire1743/X VGND VGND VPWR VPWR wire1742/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire1753 _5767_/A1 VGND VGND VPWR VPWR _3212_/A sky130_fd_sc_hd__clkbuf_1
Xwire2498 _6025_/B VGND VGND VPWR VPWR _6278_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_58_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1764 wire1765/X VGND VGND VPWR VPWR _6004_/A1 sky130_fd_sc_hd__clkbuf_2
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1775 _6108_/A1 VGND VGND VPWR VPWR _5762_/B2 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1786 wire1787/X VGND VGND VPWR VPWR wire1786/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire1797 _7006_/Q VGND VGND VPWR VPWR _6128_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_18_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3490_ _3490_/A _3519_/B VGND VGND VPWR VPWR hold30/A sky130_fd_sc_hd__nor2_1
XFILLER_115_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length681 _5381_/S VGND VGND VPWR VPWR wire679/A sky130_fd_sc_hd__clkbuf_1
XFILLER_154_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5160_ _5160_/A _5160_/B _5160_/C VGND VGND VPWR VPWR _5160_/X sky130_fd_sc_hd__or3_1
XFILLER_170_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout3583 wire3617/X VGND VGND VPWR VPWR _4200_/A1 sky130_fd_sc_hd__buf_6
X_4111_ _5241_/A _4111_/B _5241_/C _5241_/D VGND VGND VPWR VPWR _4111_/X sky130_fd_sc_hd__or4_1
XFILLER_68_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5091_ _4516_/B _4729_/Y _4988_/B _4627_/C _4635_/Y VGND VGND VPWR VPWR _5091_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4042_ _4131_/A1 hold442/X _4045_/S VGND VGND VPWR VPWR _6532_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5993_ _7095_/Q _6338_/B1 _5993_/B1 _5993_/B2 _5990_/X VGND VGND VPWR VPWR _5993_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_178_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4944_ _4944_/A _4944_/B VGND VGND VPWR VPWR _4944_/X sky130_fd_sc_hd__or2_1
X_4875_ _4964_/A _4875_/B VGND VGND VPWR VPWR _4875_/X sky130_fd_sc_hd__or2_1
XFILLER_177_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6614_ _6705_/CLK _6614_/D wire3958/X VGND VGND VPWR VPWR _6614_/Q sky130_fd_sc_hd__dfstp_1
X_3826_ _3807_/B hold81/A hold66/A VGND VGND VPWR VPWR _3826_/X sky130_fd_sc_hd__a21o_1
XFILLER_193_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6545_ _6545_/CLK _6545_/D _6433_/X VGND VGND VPWR VPWR _6545_/Q sky130_fd_sc_hd__dfrtp_1
X_3757_ _3757_/A1 wire944/X _3757_/B1 _3757_/B2 _3740_/X VGND VGND VPWR VPWR _3757_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6476_ _6824_/CLK _6476_/D fanout3973/X VGND VGND VPWR VPWR _6476_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_161_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3688_ _3688_/A _3688_/B _3688_/C _3688_/D VGND VGND VPWR VPWR _3689_/B sky130_fd_sc_hd__or4_1
XFILLER_106_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput230 _6827_/Q VGND VGND VPWR VPWR mgmt_gpio_out[25] sky130_fd_sc_hd__buf_12
X_5427_ _5427_/A0 hold508/X _5429_/S VGND VGND VPWR VPWR _6999_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput241 wire1463/X VGND VGND VPWR VPWR mgmt_gpio_out[35] sky130_fd_sc_hd__buf_12
XFILLER_133_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput252 _3946_/Y VGND VGND VPWR VPWR pad_flash_clk_oeb sky130_fd_sc_hd__buf_12
Xoutput263 _6803_/Q VGND VGND VPWR VPWR pll90_sel[2] sky130_fd_sc_hd__buf_12
Xoutput274 _6800_/Q VGND VGND VPWR VPWR pll_sel[2] sky130_fd_sc_hd__buf_12
X_5358_ _5358_/A _5571_/B VGND VGND VPWR VPWR _5363_/S sky130_fd_sc_hd__nand2_1
Xoutput285 _6477_/Q VGND VGND VPWR VPWR pll_trim[19] sky130_fd_sc_hd__buf_12
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput296 _6495_/Q VGND VGND VPWR VPWR pll_trim[5] sky130_fd_sc_hd__buf_12
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4309_ _4309_/A0 hold362/X _4311_/S VGND VGND VPWR VPWR _6753_/D sky130_fd_sc_hd__mux2_1
Xwire1005 _5860_/S VGND VGND VPWR VPWR _6319_/S sky130_fd_sc_hd__buf_2
X_5289_ _5487_/A0 _6075_/B2 _5291_/S VGND VGND VPWR VPWR _6876_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1016 _4734_/Y VGND VGND VPWR VPWR _4770_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1027 _3607_/Y VGND VGND VPWR VPWR _3783_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_75_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7028_ _7056_/CLK _7028_/D fanout3976/X VGND VGND VPWR VPWR _7028_/Q sky130_fd_sc_hd__dfrtp_1
Xwire1049 _3686_/B1 VGND VGND VPWR VPWR _4034_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3653 wire3652/A VGND VGND VPWR VPWR _5572_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_23_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire357 _4710_/X VGND VGND VPWR VPWR wire357/X sky130_fd_sc_hd__clkbuf_1
Xwire368 _3601_/X VGND VGND VPWR VPWR wire368/X sky130_fd_sc_hd__clkbuf_1
Xwire379 wire380/X VGND VGND VPWR VPWR wire379/X sky130_fd_sc_hd__clkbuf_2
XFILLER_137_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length2963 _5839_/B1 VGND VGND VPWR VPWR wire2959/A sky130_fd_sc_hd__clkbuf_1
XFILLER_136_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length2996 _5920_/A2 VGND VGND VPWR VPWR _5928_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_152_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2240 _6706_/Q VGND VGND VPWR VPWR wire2240/X sky130_fd_sc_hd__clkbuf_1
XFILLER_78_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2251 _6688_/Q VGND VGND VPWR VPWR _5915_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_66_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2262 _4226_/A1 VGND VGND VPWR VPWR _6298_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_78_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2273 _6670_/Q VGND VGND VPWR VPWR _3747_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2284 _6277_/B2 VGND VGND VPWR VPWR wire2284/X sky130_fd_sc_hd__clkbuf_1
Xwire1550 _7127_/Q VGND VGND VPWR VPWR _5986_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2295 _6337_/B2 VGND VGND VPWR VPWR _3452_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_65_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1561 wire1562/X VGND VGND VPWR VPWR wire1561/X sky130_fd_sc_hd__clkbuf_1
Xwire1572 _7107_/Q VGND VGND VPWR VPWR wire1572/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1583 wire1584/X VGND VGND VPWR VPWR _3202_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1594 _7093_/Q VGND VGND VPWR VPWR _3594_/B2 sky130_fd_sc_hd__clkbuf_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4660_ _4677_/A _4660_/B VGND VGND VPWR VPWR _4660_/X sky130_fd_sc_hd__and2_1
XFILLER_30_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3611_ _3611_/A1 _3324_/Y _3465_/Y _5921_/B2 VGND VGND VPWR VPWR _3611_/X sky130_fd_sc_hd__a22o_1
X_4591_ _4591_/A _4621_/B _4621_/C VGND VGND VPWR VPWR _4592_/A sky130_fd_sc_hd__or3_2
X_6330_ _6330_/A1 _6330_/A2 _6330_/B1 _6625_/Q _6329_/X VGND VGND VPWR VPWR _6331_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire880 wire881/X VGND VGND VPWR VPWR _4083_/S sky130_fd_sc_hd__clkbuf_2
X_3542_ _3542_/A _3542_/B _3542_/C _3542_/D VGND VGND VPWR VPWR _3543_/C sky130_fd_sc_hd__or4_2
XFILLER_128_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire891 wire892/X VGND VGND VPWR VPWR _5562_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_155_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3473_ _6765_/Q _4318_/A _3472_/Y _3473_/C1 VGND VGND VPWR VPWR _3473_/X sky130_fd_sc_hd__a211o_1
X_6261_ _6261_/A1 _6284_/A2 _6284_/B1 _6261_/B2 _6260_/X VGND VGND VPWR VPWR _6266_/A
+ sky130_fd_sc_hd__a221o_1
Xfanout4070 wire4082/X VGND VGND VPWR VPWR wire4071/A sky130_fd_sc_hd__buf_6
X_5212_ _5212_/A _5212_/B _5212_/C VGND VGND VPWR VPWR _5212_/X sky130_fd_sc_hd__or3_1
XFILLER_115_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6192_ _6192_/A _6192_/B _6192_/C _6192_/D VGND VGND VPWR VPWR _6193_/C sky130_fd_sc_hd__or4_1
X_5143_ _4664_/B _4610_/X _4795_/Y _4494_/Y VGND VGND VPWR VPWR _5143_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_97_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5074_ _4380_/X _5074_/A2 _4665_/B VGND VGND VPWR VPWR _5074_/X sky130_fd_sc_hd__o21a_1
XFILLER_84_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4025_ hold338/X _5532_/A1 _4027_/S VGND VGND VPWR VPWR _6518_/D sky130_fd_sc_hd__mux2_1
XFILLER_37_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5976_ _6006_/B _6021_/A VGND VGND VPWR VPWR _6022_/A sky130_fd_sc_hd__nor2_1
XFILLER_12_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4927_ _5130_/B wire401/X _4650_/Y VGND VGND VPWR VPWR _4928_/D sky130_fd_sc_hd__o21a_1
XFILLER_166_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4858_ _4858_/A1 _4506_/B _4694_/X wire714/X VGND VGND VPWR VPWR _4858_/X sky130_fd_sc_hd__o211a_1
XFILLER_21_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3809_ hold60/A _6468_/Q _6467_/Q _3821_/S VGND VGND VPWR VPWR _3811_/S sky130_fd_sc_hd__nand4_1
XFILLER_20_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length2226 _6714_/Q VGND VGND VPWR VPWR wire2223/A sky130_fd_sc_hd__clkbuf_1
X_4789_ _4958_/A1 _4816_/A2 _4590_/A _5108_/A VGND VGND VPWR VPWR _4983_/C sky130_fd_sc_hd__o22ai_1
X_6528_ _6799_/CLK _6528_/D wire3935/X VGND VGND VPWR VPWR _6528_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_4_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_7_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _7094_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_106_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6459_ _6545_/CLK _6459_/D _6414_/X VGND VGND VPWR VPWR _6459_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_69_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length4151 _3859_/A1 VGND VGND VPWR VPWR _3951_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_12_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2070 _6859_/Q VGND VGND VPWR VPWR _6064_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire2081 _3575_/A1 VGND VGND VPWR VPWR wire2081/X sky130_fd_sc_hd__clkbuf_1
Xwire2092 _6848_/Q VGND VGND VPWR VPWR _6194_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1380 _3711_/A VGND VGND VPWR VPWR _3714_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_53_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire1391 wire1391/A VGND VGND VPWR VPWR _5241_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_19_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5830_ _7072_/Q _5830_/A2 _5830_/B1 _6185_/A1 _5829_/X VGND VGND VPWR VPWR _5835_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_179_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5761_ _5761_/A1 _5761_/A2 _5761_/B1 _5761_/B2 VGND VGND VPWR VPWR _5761_/X sky130_fd_sc_hd__a22o_1
XFILLER_91_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4712_ _5018_/A _4712_/B _5018_/C VGND VGND VPWR VPWR _4713_/D sky130_fd_sc_hd__or3_1
XFILLER_148_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5692_ _6858_/Q _5788_/B1 _5783_/A2 _5692_/B2 _5783_/C1 VGND VGND VPWR VPWR _5692_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_30_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4643_ _4562_/X _4976_/B1 _4643_/B1 _4847_/A _4530_/B VGND VGND VPWR VPWR _4643_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_147_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4574_ _4609_/A _4609_/B _4981_/C VGND VGND VPWR VPWR _4574_/Y sky130_fd_sc_hd__nor3_1
Xhold702 _6808_/Q VGND VGND VPWR VPWR hold702/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 _6476_/Q VGND VGND VPWR VPWR hold713/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold724 _6447_/Q VGND VGND VPWR VPWR hold20/A sky130_fd_sc_hd__dlygate4sd3_1
X_6313_ _6313_/A1 _6326_/A2 _6313_/B1 _6624_/Q _6312_/X VGND VGND VPWR VPWR _6315_/C
+ sky130_fd_sc_hd__a221o_1
X_3525_ _3525_/A _3525_/B VGND VGND VPWR VPWR _4046_/A sky130_fd_sc_hd__nor2_1
XFILLER_171_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6244_ _7182_/Q _6343_/A2 _5650_/Y VGND VGND VPWR VPWR _6244_/X sky130_fd_sc_hd__o21ba_1
XFILLER_115_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3456_ _3534_/A _3456_/B VGND VGND VPWR VPWR _4282_/A sky130_fd_sc_hd__nor2_2
XFILLER_170_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3387_ _6992_/Q _3387_/A2 _5475_/A _3387_/B2 VGND VGND VPWR VPWR _3387_/X sky130_fd_sc_hd__a22o_1
X_6175_ _6992_/Q _6175_/A2 _6175_/B1 _7125_/Q _6174_/X VGND VGND VPWR VPWR _6175_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_97_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5126_ _5126_/A _5126_/B _5126_/C _4945_/X VGND VGND VPWR VPWR _5160_/B sky130_fd_sc_hd__or4b_1
XFILLER_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5057_ _4932_/A _4942_/B _4675_/A _5056_/X _4503_/C VGND VGND VPWR VPWR _5123_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_55_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4008_ _5518_/A0 hold532/X _4009_/S VGND VGND VPWR VPWR _6504_/D sky130_fd_sc_hd__mux2_1
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5959_ _6620_/Q _5959_/A2 _5959_/B1 _5959_/B2 _5958_/X VGND VGND VPWR VPWR _5967_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_187_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length1344 _5060_/A VGND VGND VPWR VPWR _4488_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length1399 _3314_/A VGND VGND VPWR VPWR _5212_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_121_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold40 hold40/A VGND VGND VPWR VPWR hold40/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A VGND VGND VPWR VPWR hold51/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold62 hold62/A VGND VGND VPWR VPWR hold62/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hold73/A VGND VGND VPWR VPWR hold73/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold84 hold84/A VGND VGND VPWR VPWR hold84/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 hold95/A VGND VGND VPWR VPWR hold95/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_4 mgmt_gpio_in[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmax_length2590 _5836_/A2 VGND VGND VPWR VPWR _5858_/A2 sky130_fd_sc_hd__clkbuf_2
X_3310_ _3318_/B _3511_/B VGND VGND VPWR VPWR _3310_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4290_ _5555_/A0 hold473/X _4293_/S VGND VGND VPWR VPWR _6737_/D sky130_fd_sc_hd__mux2_1
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3241_ _6473_/Q _6472_/Q _6471_/Q VGND VGND VPWR VPWR _3241_/X sky130_fd_sc_hd__or3_1
XFILLER_3_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6931_ _7088_/CLK _6931_/D wire4069/A VGND VGND VPWR VPWR _6931_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6862_ _7127_/CLK hold19/X fanout4054/A VGND VGND VPWR VPWR hold18/A sky130_fd_sc_hd__dfrtp_1
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5813_ _5813_/A _5813_/B _5813_/C _5813_/D VGND VGND VPWR VPWR _5813_/X sky130_fd_sc_hd__or4_1
XFILLER_50_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6793_ _6799_/CLK _6793_/D _6743_/SET_B VGND VGND VPWR VPWR _6793_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5744_ _5744_/A1 _5783_/B1 _5743_/X _5744_/B2 VGND VGND VPWR VPWR _5744_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5675_ _5683_/A _5706_/B _5706_/C VGND VGND VPWR VPWR _5675_/X sky130_fd_sc_hd__and3_1
XFILLER_136_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_72_csclk _7117_/CLK VGND VGND VPWR VPWR _7141_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4626_ _5177_/A VGND VGND VPWR VPWR _4626_/Y sky130_fd_sc_hd__inv_2
XFILLER_163_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold510 _7125_/Q VGND VGND VPWR VPWR hold510/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire4208 wire4209/X VGND VGND VPWR VPWR wire4208/X sky130_fd_sc_hd__clkbuf_1
XFILLER_144_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4557_ _4605_/A _4793_/B _4802_/C VGND VGND VPWR VPWR _4609_/B sky130_fd_sc_hd__or3_1
Xhold521 _6814_/Q VGND VGND VPWR VPWR hold521/X sky130_fd_sc_hd__dlygate4sd3_1
Xwire4219 _3549_/A1 VGND VGND VPWR VPWR wire4219/X sky130_fd_sc_hd__clkbuf_1
Xhold532 _6504_/Q VGND VGND VPWR VPWR hold532/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold543 _7066_/Q VGND VGND VPWR VPWR hold543/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold554 _6582_/Q VGND VGND VPWR VPWR hold554/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 _6494_/Q VGND VGND VPWR VPWR hold565/X sky130_fd_sc_hd__dlygate4sd3_1
X_3508_ _6486_/Q _3735_/A2 _3686_/B1 _3508_/B2 VGND VGND VPWR VPWR _3508_/X sky130_fd_sc_hd__a22o_1
Xwire3507 _5506_/A0 VGND VGND VPWR VPWR _5254_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_104_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire3518 _5515_/A0 VGND VGND VPWR VPWR _5566_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
X_4488_ _4488_/A _4488_/B VGND VGND VPWR VPWR _4847_/A sky130_fd_sc_hd__nand2_2
XFILLER_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold576 _6933_/Q VGND VGND VPWR VPWR hold576/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 _6994_/Q VGND VGND VPWR VPWR hold587/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 _6903_/Q VGND VGND VPWR VPWR hold598/X sky130_fd_sc_hd__dlygate4sd3_1
X_6227_ _6227_/A1 _6302_/A2 _6302_/B1 _6227_/B2 _6222_/X VGND VGND VPWR VPWR _6232_/B
+ sky130_fd_sc_hd__a221o_1
Xwire2806 wire2807/X VGND VGND VPWR VPWR _6199_/A2 sky130_fd_sc_hd__clkbuf_2
X_3439_ input8/X _3439_/A2 _3682_/B1 input25/X VGND VGND VPWR VPWR _3439_/X sky130_fd_sc_hd__a22o_1
Xwire2828 _5707_/B1 VGND VGND VPWR VPWR _5782_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2839 _5707_/A2 VGND VGND VPWR VPWR _5738_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_131_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6158_ _6158_/A1 _6158_/A2 _6158_/B1 _6158_/B2 _6157_/X VGND VGND VPWR VPWR _6168_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5109_ _5109_/A _5109_/B _5109_/C _5109_/D VGND VGND VPWR VPWR _5110_/C sky130_fd_sc_hd__or4_1
XFILLER_73_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6089_ _6089_/A1 _6089_/A2 _6089_/B1 _6089_/B2 _6088_/X VGND VGND VPWR VPWR _6094_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_45_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length1163 _3326_/Y VGND VGND VPWR VPWR _3645_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_134_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length1196 _3321_/Y VGND VGND VPWR VPWR _3736_/A2 sky130_fd_sc_hd__clkbuf_2
Xfanout3957 wire3963/A VGND VGND VPWR VPWR wire3959/A sky130_fd_sc_hd__buf_6
XFILLER_122_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput130 wb_adr_i[9] VGND VGND VPWR VPWR _4339_/A sky130_fd_sc_hd__clkbuf_1
Xinput141 wb_dat_i[18] VGND VGND VPWR VPWR _6369_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput152 wb_dat_i[28] VGND VGND VPWR VPWR _6376_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput163 wb_dat_i[9] VGND VGND VPWR VPWR _6366_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3790_ _3790_/A _3790_/B _3790_/C _3790_/D VGND VGND VPWR VPWR _3790_/X sky130_fd_sc_hd__or4_1
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5460_ _5514_/A0 hold566/X _5462_/S VGND VGND VPWR VPWR _7028_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4411_ _4758_/A _5001_/A VGND VGND VPWR VPWR _4445_/A sky130_fd_sc_hd__nand2_1
X_5391_ _5586_/A0 hold597/X _5391_/S VGND VGND VPWR VPWR _6967_/D sky130_fd_sc_hd__mux2_1
X_7130_ _7130_/CLK _7130_/D wire4061/X VGND VGND VPWR VPWR _7130_/Q sky130_fd_sc_hd__dfrtp_1
X_4342_ _4476_/A _4342_/B _4342_/C VGND VGND VPWR VPWR _4819_/C sky130_fd_sc_hd__and3_1
XFILLER_141_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7061_ _7134_/CLK _7061_/D fanout4057/X VGND VGND VPWR VPWR _7061_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_140_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4273_ _6723_/Q _4273_/A1 _4275_/S VGND VGND VPWR VPWR hold65/A sky130_fd_sc_hd__mux2_1
XFILLER_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6012_ _6012_/A _6012_/B _6012_/C _6012_/D VGND VGND VPWR VPWR _6045_/B sky130_fd_sc_hd__or4_1
X_3224_ _3224_/A VGND VGND VPWR VPWR _3224_/Y sky130_fd_sc_hd__inv_2
.ends

