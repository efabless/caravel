magic
tech sky130A
magscale 1 2
timestamp 1638030917
<< viali >>
rect 8493 765 8527 799
<< metal1 >>
rect 0 1114 19964 1136
rect 0 1062 4174 1114
rect 4226 1062 12174 1114
rect 12226 1062 19964 1114
rect 0 1040 19964 1062
rect 8478 796 8484 808
rect 8439 768 8484 796
rect 8478 756 8484 768
rect 8536 756 8542 808
rect 0 570 19964 592
rect 0 518 174 570
rect 226 518 8174 570
rect 8226 518 16174 570
rect 16226 518 19964 570
rect 0 496 19964 518
rect 0 26 19964 48
rect 0 -26 4174 26
rect 4226 -26 12174 26
rect 12226 -26 19964 26
rect 0 -48 19964 -26
<< via1 >>
rect 4174 1062 4226 1114
rect 12174 1062 12226 1114
rect 8484 799 8536 808
rect 8484 765 8493 799
rect 8493 765 8527 799
rect 8527 765 8536 799
rect 8484 756 8536 765
rect 174 518 226 570
rect 8174 518 8226 570
rect 16174 518 16226 570
rect 4174 -26 4226 26
rect 12174 -26 12226 26
<< metal2 >>
rect 170 570 230 1136
rect 170 518 174 570
rect 226 518 230 570
rect 170 380 230 518
rect 170 324 172 380
rect 228 324 230 380
rect 170 -48 230 324
rect 4170 1114 4230 1136
rect 4170 1062 4174 1114
rect 4226 1062 4230 1114
rect 4170 960 4230 1062
rect 4170 904 4172 960
rect 4228 904 4230 960
rect 4170 26 4230 904
rect 4170 -26 4174 26
rect 4226 -26 4230 26
rect 4170 -48 4230 -26
rect 8170 570 8230 1136
rect 12170 1114 12230 1136
rect 12170 1062 12174 1114
rect 12226 1062 12230 1114
rect 12170 960 12230 1062
rect 12170 904 12172 960
rect 12228 904 12230 960
rect 8484 808 8536 814
rect 8482 776 8484 785
rect 8536 776 8538 785
rect 8482 711 8538 720
rect 8170 518 8174 570
rect 8226 518 8230 570
rect 8170 380 8230 518
rect 8170 324 8172 380
rect 8228 324 8230 380
rect 8170 -48 8230 324
rect 12170 26 12230 904
rect 12170 -26 12174 26
rect 12226 -26 12230 26
rect 12170 -48 12230 -26
rect 16170 570 16230 1136
rect 16170 518 16174 570
rect 16226 518 16230 570
rect 16170 380 16230 518
rect 16170 324 16172 380
rect 16228 324 16230 380
rect 16170 -48 16230 324
<< via2 >>
rect 172 324 228 380
rect 4172 904 4228 960
rect 12172 904 12228 960
rect 8482 756 8484 776
rect 8484 756 8536 776
rect 8536 756 8538 776
rect 8482 720 8538 756
rect 8172 324 8228 380
rect 16172 324 16228 380
<< metal3 >>
rect 0 960 19964 982
rect 0 904 4172 960
rect 4228 904 12172 960
rect 12228 904 19964 960
rect 0 882 19964 904
rect 0 778 800 808
rect 8477 778 8543 781
rect 0 776 8543 778
rect 0 720 8482 776
rect 8538 720 8543 776
rect 0 718 8543 720
rect 0 688 800 718
rect 8477 715 8543 718
rect 0 380 19964 402
rect 0 324 172 380
rect 228 324 8172 380
rect 8228 324 16172 380
rect 16228 324 19964 380
rect 0 302 19964 324
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 0 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1638025753
transform 1 0 0 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 276 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1638025753
transform 1 0 276 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1638025753
transform 1 0 1380 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1638025753
transform 1 0 1380 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 2484 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 1638025753
transform 1 0 2484 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_29
timestamp 1638025753
transform 1 0 2668 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29
timestamp 1638025753
transform 1 0 2668 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 2576 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_11
timestamp 1638025753
transform 1 0 2576 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_41
timestamp 1638025753
transform 1 0 3772 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_41
timestamp 1638025753
transform 1 0 3772 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_53
timestamp 1638025753
transform 1 0 4876 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1638025753
transform 1 0 4876 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1638025753
transform 1 0 5244 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_57
timestamp 1638025753
transform 1 0 5244 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_5
timestamp 1638025753
transform 1 0 5152 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_12
timestamp 1638025753
transform 1 0 5152 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_69
timestamp 1638025753
transform 1 0 6348 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_69
timestamp 1638025753
transform 1 0 6348 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_81
timestamp 1638025753
transform 1 0 7452 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1638025753
transform 1 0 7452 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_85
timestamp 1638025753
transform 1 0 7820 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_6
timestamp 1638025753
transform 1 0 7728 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_13
timestamp 1638025753
transform 1 0 7728 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 7820 0 -1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_91
timestamp 1638025753
transform 1 0 8372 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_95
timestamp 1638025753
transform 1 0 8740 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_97
timestamp 1638025753
transform 1 0 8924 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  inst $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 8464 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1638025753
transform 1 0 10212 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_107 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1638025753
transform 1 0 9844 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1638025753
transform 1 0 10028 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_113
timestamp 1638025753
transform 1 0 10396 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113
timestamp 1638025753
transform 1 0 10396 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_7
timestamp 1638025753
transform 1 0 10304 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_14
timestamp 1638025753
transform 1 0 10304 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_125
timestamp 1638025753
transform 1 0 11500 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1638025753
transform 1 0 11500 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_137
timestamp 1638025753
transform 1 0 12604 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1638025753
transform 1 0 12604 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_141
timestamp 1638025753
transform 1 0 12972 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1638025753
transform 1 0 12972 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_8
timestamp 1638025753
transform 1 0 12880 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_15
timestamp 1638025753
transform 1 0 12880 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_153
timestamp 1638025753
transform 1 0 14076 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_153
timestamp 1638025753
transform 1 0 14076 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp 1638025753
transform 1 0 15180 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1638025753
transform 1 0 15180 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_169
timestamp 1638025753
transform 1 0 15548 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_169
timestamp 1638025753
transform 1 0 15548 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_9
timestamp 1638025753
transform 1 0 15456 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_16
timestamp 1638025753
transform 1 0 15456 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_181
timestamp 1638025753
transform 1 0 16652 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_181
timestamp 1638025753
transform 1 0 16652 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_193
timestamp 1638025753
transform 1 0 17756 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1638025753
transform 1 0 17756 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_197
timestamp 1638025753
transform 1 0 18124 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_197
timestamp 1638025753
transform 1 0 18124 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_17
timestamp 1638025753
transform 1 0 18032 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_10
timestamp 1638025753
transform 1 0 18032 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_213
timestamp 1638025753
transform 1 0 19596 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_213
timestamp 1638025753
transform 1 0 19596 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_209
timestamp 1638025753
transform 1 0 19228 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_209
timestamp 1638025753
transform 1 0 19228 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1638025753
transform -1 0 19964 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1638025753
transform -1 0 19964 0 1 0
box -38 -48 314 592
<< labels >>
rlabel metal3 s 0 688 800 808 6 HI
port 0 nsew signal tristate
rlabel metal3 s 0 302 19964 402 6 vccd2
port 1 nsew power input
rlabel metal2 s 170 -48 230 1136 6 vccd2
port 1 nsew power input
rlabel metal2 s 8170 -48 8230 1136 6 vccd2
port 1 nsew power input
rlabel metal2 s 16170 -48 16230 1136 6 vccd2
port 1 nsew power input
rlabel metal3 s 0 882 19964 982 6 vssd2
port 2 nsew ground input
rlabel metal2 s 4170 -48 4230 1136 6 vssd2
port 2 nsew ground input
rlabel metal2 s 12170 -48 12230 1136 6 vssd2
port 2 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 20000 1400
<< end >>
