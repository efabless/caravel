magic
tech sky130A
magscale 1 2
timestamp 1638030917
<< checkpaint >>
rect 7506 3785 11790 4559
rect 5010 325 11790 3785
rect 12594 325 15726 3785
rect 26802 325 31278 4559
<< isosubstrate >>
rect 6116 1496 7106 2652
rect 13698 1476 14528 2638
<< viali >>
rect 8959 2610 8993 2644
rect 28255 2610 28289 2644
rect 6655 2240 6689 2274
rect 28831 1944 28865 1978
rect 14047 1870 14081 1904
rect 9535 1796 9569 1830
<< metal1 >>
rect 8578 3282 29952 3307
rect 8578 3230 10934 3282
rect 10986 3230 26934 3282
rect 26986 3230 29952 3282
rect 8578 3205 29952 3230
rect 6640 2601 6646 2653
rect 6698 2641 6704 2653
rect 8947 2644 9005 2650
rect 8947 2641 8959 2644
rect 6698 2613 8959 2641
rect 6698 2601 6704 2613
rect 8947 2610 8959 2613
rect 8993 2610 9005 2644
rect 28240 2641 28246 2653
rect 28201 2613 28246 2641
rect 8947 2604 9005 2610
rect 28240 2601 28246 2613
rect 28298 2601 28304 2653
rect 5442 2468 8042 2493
rect 5442 2416 5800 2468
rect 5852 2416 8042 2468
rect 5442 2391 8042 2416
rect 8760 2468 10540 2493
rect 8760 2416 9974 2468
rect 10026 2416 10540 2468
rect 8760 2391 10540 2416
rect 13362 2468 15306 2493
rect 13362 2416 14664 2468
rect 14716 2416 15306 2468
rect 13362 2391 15306 2416
rect 15766 2468 27494 2493
rect 15766 2416 18934 2468
rect 18986 2416 27494 2468
rect 15766 2391 27494 2416
rect 28056 2468 29952 2493
rect 28056 2416 29190 2468
rect 29242 2416 29952 2468
rect 28056 2391 29952 2416
rect 10113 2286 28290 2289
rect 6640 2271 6646 2283
rect 6601 2243 6646 2271
rect 6640 2231 6646 2243
rect 6698 2231 6704 2283
rect 10113 2234 18927 2286
rect 18979 2234 28290 2286
rect 10113 2232 28290 2234
rect 784 1935 790 1987
rect 842 1975 848 1987
rect 28819 1978 28877 1984
rect 28819 1975 28831 1978
rect 842 1947 28831 1975
rect 842 1935 848 1947
rect 28819 1944 28831 1947
rect 28865 1944 28877 1978
rect 28819 1938 28877 1944
rect 14035 1904 14093 1910
rect 14035 1870 14047 1904
rect 14081 1901 14093 1904
rect 28240 1901 28246 1913
rect 14081 1873 28246 1901
rect 14081 1870 14093 1873
rect 14035 1864 14093 1870
rect 28240 1861 28246 1873
rect 28298 1861 28304 1913
rect 784 1787 790 1839
rect 842 1827 848 1839
rect 9523 1830 9581 1836
rect 9523 1827 9535 1830
rect 842 1799 9535 1827
rect 842 1787 848 1799
rect 9523 1796 9535 1799
rect 9569 1796 9581 1830
rect 9523 1790 9581 1796
rect 5406 1654 8010 1679
rect 5406 1602 7460 1654
rect 7512 1602 8010 1654
rect 5406 1577 8010 1602
rect 8510 1654 12920 1679
rect 8510 1602 10934 1654
rect 10986 1602 12920 1654
rect 8510 1577 12920 1602
rect 13380 1654 15310 1679
rect 13380 1602 13488 1654
rect 13540 1602 15310 1654
rect 13380 1577 15310 1602
rect 15770 1654 29952 1679
rect 15770 1602 26934 1654
rect 26986 1602 29952 1654
rect 15770 1577 29952 1602
rect 8510 840 29952 865
rect 8510 788 18934 840
rect 18986 788 29952 840
rect 8510 763 29952 788
<< via1 >>
rect 10934 3230 10986 3282
rect 26934 3230 26986 3282
rect 6646 2601 6698 2653
rect 28246 2644 28298 2653
rect 28246 2610 28255 2644
rect 28255 2610 28289 2644
rect 28289 2610 28298 2644
rect 28246 2601 28298 2610
rect 5800 2416 5852 2468
rect 9974 2416 10026 2468
rect 14664 2416 14716 2468
rect 18934 2416 18986 2468
rect 29190 2416 29242 2468
rect 6646 2274 6698 2283
rect 6646 2240 6655 2274
rect 6655 2240 6689 2274
rect 6689 2240 6698 2274
rect 6646 2231 6698 2240
rect 18927 2234 18979 2286
rect 790 1935 842 1987
rect 28246 1861 28298 1913
rect 790 1787 842 1839
rect 7460 1602 7512 1654
rect 10934 1602 10986 1654
rect 13488 1602 13540 1654
rect 26934 1602 26986 1654
rect 18934 788 18986 840
<< metal2 >>
rect 10930 3282 10990 3307
rect 10930 3230 10934 3282
rect 10986 3230 10990 3282
rect 7412 2930 7612 2971
rect 788 2914 844 2923
rect 788 2849 844 2858
rect 802 1993 830 2849
rect 7412 2794 7444 2930
rect 7580 2794 7612 2930
rect 6646 2653 6698 2659
rect 6646 2595 6698 2601
rect 5775 2494 5877 2499
rect 5744 2468 5904 2494
rect 5744 2416 5800 2468
rect 5852 2416 5904 2468
rect 790 1987 842 1993
rect 790 1929 842 1935
rect 5744 1900 5904 2416
rect 6658 2289 6686 2595
rect 6646 2283 6698 2289
rect 6646 2225 6698 2231
rect 790 1839 842 1845
rect 790 1781 842 1787
rect 802 999 830 1781
rect 5744 1764 5756 1900
rect 5892 1764 5904 1900
rect 5744 1743 5904 1764
rect 7412 1654 7612 2794
rect 9886 2468 10096 2566
rect 9886 2416 9974 2468
rect 10026 2416 10096 2468
rect 9886 1864 10096 2416
rect 9886 1728 9923 1864
rect 10059 1728 10096 1864
rect 9886 1682 10096 1728
rect 10930 2071 10990 3230
rect 10930 2015 10932 2071
rect 10988 2015 10990 2071
rect 7412 1602 7460 1654
rect 7512 1602 7612 1654
rect 7412 1576 7612 1602
rect 10930 1654 10990 2015
rect 10930 1602 10934 1654
rect 10986 1602 10990 1654
rect 7435 1571 7537 1576
rect 788 990 844 999
rect 788 925 844 934
rect 10930 763 10990 1602
rect 11330 2522 11390 3256
rect 11330 2466 11332 2522
rect 11388 2466 11390 2522
rect 11330 814 11390 2466
rect 11730 2922 11790 3256
rect 11730 2866 11732 2922
rect 11788 2866 11790 2922
rect 11730 814 11790 2866
rect 18930 3151 18990 3307
rect 26930 3282 26990 3307
rect 18930 3095 18932 3151
rect 18988 3095 18990 3151
rect 13420 2538 13614 2576
rect 13420 2402 13449 2538
rect 13585 2402 13614 2538
rect 14639 2484 14741 2499
rect 13420 1654 13614 2402
rect 13420 1602 13488 1654
rect 13540 1602 13614 1654
rect 13420 1574 13614 1602
rect 14618 2468 14818 2484
rect 14618 2416 14664 2468
rect 14716 2416 14818 2468
rect 13463 1571 13565 1574
rect 14618 1506 14818 2416
rect 18930 2468 18990 3095
rect 18930 2416 18934 2468
rect 18986 2416 18990 2468
rect 18930 2295 18990 2416
rect 18925 2286 18990 2295
rect 18925 2234 18927 2286
rect 18979 2234 18990 2286
rect 18925 2226 18990 2234
rect 14618 1370 14650 1506
rect 14786 1370 14818 1506
rect 14618 1329 14818 1370
rect 18930 991 18990 2226
rect 18930 935 18932 991
rect 18988 935 18990 991
rect 18930 840 18990 935
rect 18930 788 18934 840
rect 18986 788 18990 840
rect 19330 1442 19390 3256
rect 19330 1386 19332 1442
rect 19388 1386 19390 1442
rect 19330 814 19390 1386
rect 19730 1842 19790 3256
rect 19730 1786 19732 1842
rect 19788 1786 19790 1842
rect 19730 814 19790 1786
rect 26930 3230 26934 3282
rect 26986 3230 26990 3282
rect 26930 2071 26990 3230
rect 26930 2015 26932 2071
rect 26988 2015 26990 2071
rect 26930 1654 26990 2015
rect 26930 1602 26934 1654
rect 26986 1602 26990 1654
rect 18930 763 18990 788
rect 26930 763 26990 1602
rect 27330 2522 27390 3256
rect 27330 2466 27332 2522
rect 27388 2466 27390 2522
rect 27330 814 27390 2466
rect 27730 2922 27790 3256
rect 27730 2866 27732 2922
rect 27788 2866 27790 2922
rect 27730 814 27790 2866
rect 28246 2653 28298 2659
rect 28246 2595 28298 2601
rect 28258 1919 28286 2595
rect 29132 2468 29312 2562
rect 29132 2416 29190 2468
rect 29242 2416 29312 2468
rect 28246 1913 28298 1919
rect 28246 1855 28298 1861
rect 29132 1502 29312 2416
rect 29132 1366 29154 1502
rect 29290 1366 29312 1502
rect 29132 1335 29312 1366
<< via2 >>
rect 788 2858 844 2914
rect 7444 2794 7580 2930
rect 5756 1764 5892 1900
rect 9923 1728 10059 1864
rect 10932 2015 10988 2071
rect 788 934 844 990
rect 11332 2466 11388 2522
rect 11732 2866 11788 2922
rect 18932 3095 18988 3151
rect 13449 2402 13585 2538
rect 14650 1370 14786 1506
rect 18932 935 18988 991
rect 19332 1386 19388 1442
rect 19732 1786 19788 1842
rect 26932 2015 26988 2071
rect 27332 2466 27388 2522
rect 27732 2866 27788 2922
rect 29154 1366 29290 1502
<< metal3 >>
rect 18927 3153 18993 3156
rect 960 3151 29952 3153
rect 960 3095 18932 3151
rect 18988 3095 29952 3151
rect 960 3093 29952 3095
rect 18927 3090 18993 3093
rect 0 2919 800 2946
rect 7407 2930 7617 2967
rect 7407 2924 7444 2930
rect 0 2914 849 2919
rect 0 2858 788 2914
rect 844 2858 849 2914
rect 960 2864 7444 2924
rect 0 2853 849 2858
rect 0 2826 800 2853
rect 7407 2794 7444 2864
rect 7580 2924 7617 2930
rect 11727 2924 11793 2927
rect 27727 2924 27793 2927
rect 7580 2922 29952 2924
rect 7580 2866 11732 2922
rect 11788 2866 27732 2922
rect 27788 2866 29952 2922
rect 7580 2864 29952 2866
rect 7580 2794 7617 2864
rect 11727 2861 11793 2864
rect 27727 2861 27793 2864
rect 7407 2757 7617 2794
rect 13415 2538 13619 2572
rect 11327 2524 11393 2527
rect 13415 2524 13449 2538
rect 960 2522 13449 2524
rect 960 2466 11332 2522
rect 11388 2466 13449 2522
rect 960 2464 13449 2466
rect 11327 2461 11393 2464
rect 13415 2402 13449 2464
rect 13585 2524 13619 2538
rect 27327 2524 27393 2527
rect 13585 2522 29952 2524
rect 13585 2466 27332 2522
rect 27388 2466 29952 2522
rect 13585 2464 29952 2466
rect 13585 2402 13619 2464
rect 27327 2461 27393 2464
rect 13415 2368 13619 2402
rect 10927 2073 10993 2076
rect 26927 2073 26993 2076
rect 960 2071 29952 2073
rect 960 2015 10932 2071
rect 10988 2015 26932 2071
rect 26988 2015 29952 2071
rect 960 2013 29952 2015
rect 10927 2010 10993 2013
rect 26927 2010 26993 2013
rect 5739 1900 5909 1917
rect 5739 1844 5756 1900
rect 960 1784 5756 1844
rect 5739 1764 5756 1784
rect 5892 1844 5909 1900
rect 9881 1864 10101 1906
rect 9881 1844 9923 1864
rect 5892 1784 9923 1844
rect 5892 1764 5909 1784
rect 5739 1747 5909 1764
rect 9881 1728 9923 1784
rect 10059 1844 10101 1864
rect 19727 1844 19793 1847
rect 10059 1842 29952 1844
rect 10059 1786 19732 1842
rect 19788 1786 29952 1842
rect 10059 1784 29952 1786
rect 10059 1728 10101 1784
rect 19727 1781 19793 1784
rect 9881 1686 10101 1728
rect 14613 1506 14823 1543
rect 14613 1444 14650 1506
rect 960 1384 14650 1444
rect 14613 1370 14650 1384
rect 14786 1444 14823 1506
rect 29127 1502 29317 1529
rect 19327 1444 19393 1447
rect 29127 1444 29154 1502
rect 14786 1442 29154 1444
rect 14786 1386 19332 1442
rect 19388 1386 29154 1442
rect 14786 1384 29154 1386
rect 14786 1370 14823 1384
rect 19327 1381 19393 1384
rect 14613 1333 14823 1370
rect 29127 1366 29154 1384
rect 29290 1444 29317 1502
rect 29290 1384 29952 1444
rect 29290 1366 29317 1384
rect 29127 1339 29317 1366
rect 0 995 800 1022
rect 0 990 849 995
rect 18927 993 18993 996
rect 0 934 788 990
rect 844 934 849 990
rect 0 929 849 934
rect 960 991 29952 993
rect 960 935 18932 991
rect 18988 935 29952 991
rect 960 933 29952 935
rect 18927 930 18993 933
rect 0 902 800 929
use sky130_fd_sc_hvl__fill_2  FILLER_2_300 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1638906210
transform 1 0 29760 0 -1 3256
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  FILLER_1_300
timestamp 1638906210
transform 1 0 29760 0 1 1628
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_1  FILLER_1_56 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1638906210
transform 1 0 6336 0 1 1628
box -66 -43 162 897
use sky130_fd_sc_hvl__lsbufhv2lv_1  mprj2_logic_high_lv $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1638906210
transform 1 0 8832 0 1 1628
box -66 -43 1698 1671
use sky130_fd_sc_hvl__lsbufhv2lv_1  mprj_logic_high_lv
timestamp 1638906210
transform 1 0 28128 0 1 1628
box -66 -43 1698 1671
use sky130_fd_sc_hvl__conb_1  mprj_logic_high_hvl $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1638906210
transform 1 0 13920 0 1 1628
box -66 -43 546 897
use sky130_fd_sc_hvl__conb_1  mprj2_logic_high_hvl
timestamp 1638906210
transform 1 0 6432 0 1 1628
box -66 -43 546 897
<< labels >>
rlabel metal3 s 0 902 800 1022 4 mprj2_vdd_logic1
rlabel metal3 s 0 2826 800 2946 4 mprj_vdd_logic1
rlabel metal3 s 960 3093 29952 3153 4 vccd
rlabel metal3 s 960 933 29952 993 4 vccd
rlabel metal3 s 960 2013 29952 2073 4 vssd
rlabel metal3 s 960 1384 29952 1444 4 vdda1
rlabel metal3 s 960 2464 29952 2524 4 vssa1
rlabel metal3 s 960 1784 29952 1844 4 vdda2
rlabel metal3 s 960 2864 29952 2924 4 vssa2
rlabel metal2 s 18930 763 18990 3307 4 vccd
rlabel metal2 s 26930 763 26990 3307 4 vssd
rlabel metal2 s 10930 763 10990 3307 4 vssd
rlabel metal2 s 19330 814 19390 3256 4 vdda1
rlabel metal2 s 27330 814 27390 3256 4 vssa1
rlabel metal2 s 11330 814 11390 3256 4 vssa1
rlabel metal2 s 19730 814 19790 3256 4 vdda2
rlabel metal2 s 27730 814 27790 3256 4 vssa2
rlabel metal2 s 11730 814 11790 3256 4 vssa2
rlabel metal2 s 18960 2035 18960 2035 4 vccd
port 1 nsew
rlabel metal2 s 26960 2035 26960 2035 4 vssd
port 2 nsew
rlabel metal2 s 10960 2035 10960 2035 4 vssd
port 2 nsew
rlabel metal2 s 19360 2035 19360 2035 4 vdda1
port 3 nsew
rlabel metal2 s 27360 2035 27360 2035 4 vssa1
port 4 nsew
rlabel metal2 s 11360 2035 11360 2035 4 vssa1
port 4 nsew
rlabel metal2 s 19760 2035 19760 2035 4 vdda2
port 5 nsew
rlabel metal2 s 27760 2035 27760 2035 4 vssa2
port 6 nsew
rlabel metal2 s 11760 2035 11760 2035 4 vssa2
port 6 nsew
rlabel metal3 s 400 962 400 962 4 mprj2_vdd_logic1
port 7 nsew
rlabel metal3 s 400 2886 400 2886 4 mprj_vdd_logic1
port 8 nsew
rlabel metal3 s 15456 3123 15456 3123 4 vccd
port 1 nsew
rlabel metal3 s 15456 963 15456 963 4 vccd
port 1 nsew
rlabel metal3 s 15456 2043 15456 2043 4 vssd
port 2 nsew
rlabel metal3 s 15456 1414 15456 1414 4 vdda1
port 3 nsew
rlabel metal3 s 15456 2494 15456 2494 4 vssa1
port 4 nsew
rlabel metal3 s 15456 1814 15456 1814 4 vdda2
port 5 nsew
rlabel metal3 s 15456 2894 15456 2894 4 vssa2
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 30000 4000
<< end >>
